module NRISC_InstructionDecoder (CORE_InstructionIN, CORE_ctrl, CORE_ULA_flags, clk, rst, CORE_InstructionToULAMux, CORE_Status_ctrl, CORE_ULA_ctrl, CORE_ULAMux_inc_dec, CORE_REG_RF1, CORE_REG_RF2, CORE_REG_RD, CORE_REG_write, CORE_DATA_write, CORE_DATA_load, CORE_DATA_ctrl, CORE_DATA_ADDR_mux, CORE_DATA_REGMux, CORE_STACK_ctrl, CORE_PC_ctrl, CORE_PC_clk, CORE_INT_CHA, CORE_INT_ctrl);

input clk;
input rst;
output CORE_ULAMux_inc_dec;
output CORE_REG_write;
output CORE_DATA_write;
output CORE_DATA_load;
output CORE_DATA_ADDR_mux;
output CORE_DATA_REGMux;
output CORE_PC_clk;
input [15:0] CORE_InstructionIN;
input [2:0] CORE_ctrl;
input [2:0] CORE_ULA_flags;
output [1:0] CORE_InstructionToULAMux;
output [4:0] CORE_Status_ctrl;
output [3:0] CORE_ULA_ctrl;
output [3:0] CORE_REG_RF1;
output [3:0] CORE_REG_RF2;
output [3:0] CORE_REG_RD;
output [2:0] CORE_DATA_ctrl;
output [1:0] CORE_STACK_ctrl;
output [1:0] CORE_PC_ctrl;
output [7:0] CORE_INT_CHA;
output [1:0] CORE_INT_ctrl;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(_16_), .Y(_16__bF_buf3) );
BUFX4 BUFX4_2 ( .A(_16_), .Y(_16__bF_buf2) );
BUFX4 BUFX4_3 ( .A(_16_), .Y(_16__bF_buf1) );
BUFX4 BUFX4_4 ( .A(_16_), .Y(_16__bF_buf0) );
BUFX4 BUFX4_5 ( .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_6 ( .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_7 ( .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_8 ( .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_9 ( .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_10 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_11 ( .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf3) );
BUFX4 BUFX4_12 ( .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf2) );
BUFX4 BUFX4_13 ( .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf1) );
BUFX4 BUFX4_14 ( .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf0) );
INVX8 INVX8_1 ( .A(CORE_InstructionIN_15_bF_buf3), .Y(_16_) );
INVX8 INVX8_2 ( .A(CORE_InstructionIN[11]), .Y(_17_) );
INVX4 INVX4_1 ( .A(CORE_InstructionIN[13]), .Y(_18_) );
NOR2X1 NOR2X1_1 ( .A(CORE_InstructionIN[14]), .B(CORE_InstructionIN[12]), .Y(_19_) );
AND2X2 AND2X2_1 ( .A(_19_), .B(_18_), .Y(_20_) );
NAND3X1 NAND3X1_1 ( .A(_16__bF_buf3), .B(_17_), .C(_20_), .Y(_21_) );
NAND3X1 NAND3X1_2 ( .A(_216__0_), .B(CORE_InstructionIN[14]), .C(_16__bF_buf2), .Y(_22_) );
INVX2 INVX2_1 ( .A(CORE_InstructionIN[10]), .Y(_23_) );
NAND2X1 NAND2X1_1 ( .A(CORE_InstructionIN[9]), .B(_23_), .Y(_24_) );
NOR2X1 NOR2X1_2 ( .A(CORE_InstructionIN[8]), .B(_24_), .Y(_25_) );
AOI21X1 AOI21X1_1 ( .A(_216__0_), .B(CORE_InstructionIN[10]), .C(_25_), .Y(_26_) );
OAI21X1 OAI21X1_1 ( .A(_26_), .B(_21_), .C(_22_), .Y(_6__0_) );
INVX4 INVX4_2 ( .A(CORE_InstructionIN[14]), .Y(_27_) );
NOR2X1 NOR2X1_3 ( .A(CORE_InstructionIN_15_bF_buf2), .B(_27_), .Y(_28_) );
NAND2X1 NAND2X1_2 ( .A(_216__1_), .B(_28_), .Y(_29_) );
AOI21X1 AOI21X1_2 ( .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[9]), .C(CORE_InstructionIN[10]), .Y(_30_) );
INVX2 INVX2_2 ( .A(_30_), .Y(_31_) );
OAI21X1 OAI21X1_2 ( .A(_23_), .B(_216__1_), .C(_31_), .Y(_32_) );
OAI21X1 OAI21X1_3 ( .A(_21_), .B(_32_), .C(_29_), .Y(_6__1_) );
INVX1 INVX1_1 ( .A(_215__0_), .Y(_33_) );
INVX2 INVX2_3 ( .A(CORE_InstructionIN[0]), .Y(_34_) );
NOR2X1 NOR2X1_4 ( .A(_24_), .B(_21_), .Y(_35_) );
MUX2X1 MUX2X1_1 ( .A(_34_), .B(_33_), .S(_35_), .Y(_5__0_) );
INVX1 INVX1_2 ( .A(_215__1_), .Y(_36_) );
INVX4 INVX4_3 ( .A(CORE_InstructionIN[1]), .Y(_37_) );
MUX2X1 MUX2X1_2 ( .A(_37_), .B(_36_), .S(_35_), .Y(_5__1_) );
INVX1 INVX1_3 ( .A(_215__2_), .Y(_38_) );
INVX2 INVX2_4 ( .A(CORE_InstructionIN[2]), .Y(_39_) );
MUX2X1 MUX2X1_3 ( .A(_39_), .B(_38_), .S(_35_), .Y(_5__2_) );
INVX1 INVX1_4 ( .A(_215__3_), .Y(_40_) );
INVX2 INVX2_5 ( .A(CORE_InstructionIN[3]), .Y(_41_) );
MUX2X1 MUX2X1_4 ( .A(_41_), .B(_40_), .S(_35_), .Y(_5__3_) );
INVX1 INVX1_5 ( .A(_215__4_), .Y(_42_) );
INVX1 INVX1_6 ( .A(CORE_InstructionIN[4]), .Y(_43_) );
MUX2X1 MUX2X1_5 ( .A(_43_), .B(_42_), .S(_35_), .Y(_5__4_) );
INVX1 INVX1_7 ( .A(_215__5_), .Y(_44_) );
INVX1 INVX1_8 ( .A(CORE_InstructionIN[5]), .Y(_45_) );
MUX2X1 MUX2X1_6 ( .A(_45_), .B(_44_), .S(_35_), .Y(_5__5_) );
INVX1 INVX1_9 ( .A(_215__6_), .Y(_46_) );
INVX1 INVX1_10 ( .A(CORE_InstructionIN[6]), .Y(_47_) );
MUX2X1 MUX2X1_7 ( .A(_47_), .B(_46_), .S(_35_), .Y(_5__6_) );
INVX1 INVX1_11 ( .A(_215__7_), .Y(_48_) );
INVX1 INVX1_12 ( .A(CORE_InstructionIN[7]), .Y(_49_) );
MUX2X1 MUX2X1_8 ( .A(_49_), .B(_48_), .S(_35_), .Y(_5__7_) );
INVX4 INVX4_4 ( .A(CORE_InstructionIN[9]), .Y(_50_) );
NAND3X1 NAND3X1_3 ( .A(CORE_InstructionIN[8]), .B(CORE_ULA_flags[1]), .C(_50_), .Y(_51_) );
NAND3X1 NAND3X1_4 ( .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[9]), .C(CORE_ULA_flags[0]), .Y(_52_) );
INVX2 INVX2_6 ( .A(CORE_InstructionIN[8]), .Y(_53_) );
OAI21X1 OAI21X1_4 ( .A(_50_), .B(CORE_ULA_flags[2]), .C(_53_), .Y(_54_) );
NAND3X1 NAND3X1_5 ( .A(_52_), .B(_51_), .C(_54_), .Y(_55_) );
NAND2X1 NAND2X1_3 ( .A(CORE_InstructionIN[12]), .B(_27_), .Y(_56_) );
OR2X2 OR2X2_1 ( .A(_56_), .B(CORE_InstructionIN[13]), .Y(_57_) );
NOR2X1 NOR2X1_5 ( .A(_218__0_), .B(_17_), .Y(_58_) );
NOR2X1 NOR2X1_6 ( .A(_58_), .B(_57_), .Y(_59_) );
OAI21X1 OAI21X1_5 ( .A(_55_), .B(CORE_InstructionIN[11]), .C(_59_), .Y(_60_) );
NAND2X1 NAND2X1_4 ( .A(_18_), .B(_19_), .Y(_61_) );
NOR2X1 NOR2X1_7 ( .A(_17_), .B(_61_), .Y(_62_) );
OAI21X1 OAI21X1_6 ( .A(_23_), .B(_50_), .C(_218__0_), .Y(_63_) );
NAND2X1 NAND2X1_5 ( .A(_31_), .B(_63_), .Y(_64_) );
AOI22X1 AOI22X1_1 ( .A(CORE_InstructionIN[14]), .B(_218__0_), .C(_62_), .D(_64_), .Y(_65_) );
AOI21X1 AOI21X1_3 ( .A(_65_), .B(_60_), .C(CORE_InstructionIN_15_bF_buf1), .Y(_8__0_) );
INVX1 INVX1_13 ( .A(_218__1_), .Y(_66_) );
NAND2X1 NAND2X1_6 ( .A(CORE_InstructionIN[10]), .B(CORE_InstructionIN[9]), .Y(_67_) );
AOI21X1 AOI21X1_4 ( .A(_66_), .B(_67_), .C(_30_), .Y(_68_) );
NOR2X1 NOR2X1_8 ( .A(_66_), .B(_57_), .Y(_69_) );
AOI22X1 AOI22X1_2 ( .A(_62_), .B(_68_), .C(_69_), .D(CORE_InstructionIN[11]), .Y(_70_) );
NAND2X1 NAND2X1_7 ( .A(CORE_InstructionIN[14]), .B(_218__1_), .Y(_71_) );
AOI21X1 AOI21X1_5 ( .A(_71_), .B(_70_), .C(CORE_InstructionIN_15_bF_buf0), .Y(_8__1_) );
NAND2X1 NAND2X1_8 ( .A(CORE_InstructionIN[11]), .B(_20_), .Y(_72_) );
NAND2X1 NAND2X1_9 ( .A(CORE_InstructionIN[14]), .B(_223__0_), .Y(_73_) );
AOI21X1 AOI21X1_6 ( .A(_223__0_), .B(_67_), .C(_30_), .Y(_74_) );
OAI21X1 OAI21X1_7 ( .A(_72_), .B(_74_), .C(_73_), .Y(_75_) );
AND2X2 AND2X2_2 ( .A(_75_), .B(_16__bF_buf1), .Y(_13__0_) );
NOR2X1 NOR2X1_9 ( .A(_67_), .B(_72_), .Y(_76_) );
NOR2X1 NOR2X1_10 ( .A(_223__1_), .B(_76_), .Y(_77_) );
OAI21X1 OAI21X1_8 ( .A(_72_), .B(_30_), .C(_27_), .Y(_78_) );
NAND2X1 NAND2X1_10 ( .A(_16__bF_buf0), .B(_78_), .Y(_79_) );
NOR2X1 NOR2X1_11 ( .A(_77_), .B(_79_), .Y(_13__1_) );
NAND3X1 NAND3X1_6 ( .A(CORE_InstructionIN[2]), .B(_37_), .C(_41_), .Y(_80_) );
NOR2X1 NOR2X1_12 ( .A(CORE_InstructionIN[0]), .B(CORE_InstructionIN[1]), .Y(_81_) );
OR2X2 OR2X2_2 ( .A(CORE_InstructionIN[2]), .B(CORE_InstructionIN[3]), .Y(_82_) );
OAI21X1 OAI21X1_9 ( .A(_81_), .B(_82_), .C(_80_), .Y(_83_) );
NOR2X1 NOR2X1_13 ( .A(CORE_InstructionIN[2]), .B(CORE_InstructionIN[3]), .Y(_84_) );
NAND2X1 NAND2X1_11 ( .A(_81_), .B(_84_), .Y(_85_) );
AOI21X1 AOI21X1_7 ( .A(_211_), .B(_85_), .C(_83_), .Y(_86_) );
NOR3X1 NOR3X1_1 ( .A(CORE_InstructionIN[14]), .B(CORE_InstructionIN[12]), .C(_18_), .Y(_87_) );
NAND2X1 NAND2X1_12 ( .A(_16__bF_buf3), .B(_87_), .Y(_88_) );
NAND2X1 NAND2X1_13 ( .A(_211_), .B(_28_), .Y(_89_) );
OAI21X1 OAI21X1_10 ( .A(_86_), .B(_88_), .C(_89_), .Y(_1_) );
NOR2X1 NOR2X1_14 ( .A(CORE_InstructionIN[14]), .B(_18_), .Y(_90_) );
INVX2 INVX2_7 ( .A(_90_), .Y(_91_) );
OAI21X1 OAI21X1_11 ( .A(_91_), .B(CORE_InstructionIN_15_bF_buf3), .C(_212__0_), .Y(_92_) );
INVX1 INVX1_14 ( .A(_212__0_), .Y(_93_) );
OAI21X1 OAI21X1_12 ( .A(CORE_InstructionIN[0]), .B(CORE_InstructionIN[1]), .C(_84_), .Y(_94_) );
NAND3X1 NAND3X1_7 ( .A(_93_), .B(_80_), .C(_94_), .Y(_95_) );
NOR3X1 NOR3X1_2 ( .A(CORE_InstructionIN[1]), .B(CORE_InstructionIN[3]), .C(_39_), .Y(_96_) );
NAND2X1 NAND2X1_14 ( .A(CORE_InstructionIN[0]), .B(_37_), .Y(_97_) );
NOR2X1 NOR2X1_15 ( .A(_82_), .B(_97_), .Y(_98_) );
NAND2X1 NAND2X1_15 ( .A(CORE_InstructionIN[13]), .B(_19_), .Y(_99_) );
NOR3X1 NOR3X1_3 ( .A(_96_), .B(_99_), .C(_98_), .Y(_100_) );
OR2X2 OR2X2_3 ( .A(_56_), .B(_18_), .Y(_101_) );
NAND2X1 NAND2X1_16 ( .A(CORE_InstructionIN[10]), .B(CORE_InstructionIN[11]), .Y(_102_) );
OAI22X1 OAI22X1_1 ( .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[11]), .C(_102_), .D(_212__0_), .Y(_103_) );
NOR2X1 NOR2X1_16 ( .A(_103_), .B(_101_), .Y(_104_) );
AOI21X1 AOI21X1_8 ( .A(_95_), .B(_100_), .C(_104_), .Y(_105_) );
OAI21X1 OAI21X1_13 ( .A(_105_), .B(CORE_InstructionIN_15_bF_buf2), .C(_92_), .Y(_2__0_) );
INVX1 INVX1_15 ( .A(_212__1_), .Y(_106_) );
NOR2X1 NOR2X1_17 ( .A(CORE_InstructionIN_15_bF_buf1), .B(_91_), .Y(_107_) );
INVX1 INVX1_16 ( .A(_101_), .Y(_108_) );
NOR2X1 NOR2X1_18 ( .A(_212__1_), .B(_102_), .Y(_109_) );
AOI21X1 AOI21X1_9 ( .A(_17_), .B(_24_), .C(_109_), .Y(_110_) );
AOI21X1 AOI21X1_10 ( .A(_106_), .B(_80_), .C(_99_), .Y(_111_) );
AOI22X1 AOI22X1_3 ( .A(_94_), .B(_111_), .C(_108_), .D(_110_), .Y(_112_) );
OAI22X1 OAI22X1_2 ( .A(_106_), .B(_107_), .C(_112_), .D(CORE_InstructionIN_15_bF_buf0), .Y(_2__1_) );
OAI21X1 OAI21X1_14 ( .A(_91_), .B(CORE_InstructionIN_15_bF_buf3), .C(_212__2_), .Y(_113_) );
INVX1 INVX1_17 ( .A(_212__2_), .Y(_114_) );
NAND3X1 NAND3X1_8 ( .A(_114_), .B(_80_), .C(_94_), .Y(_115_) );
NAND2X1 NAND2X1_17 ( .A(CORE_InstructionIN[2]), .B(_41_), .Y(_116_) );
NOR2X1 NOR2X1_19 ( .A(_116_), .B(_97_), .Y(_117_) );
NAND2X1 NAND2X1_18 ( .A(CORE_InstructionIN[0]), .B(_84_), .Y(_118_) );
NAND2X1 NAND2X1_19 ( .A(_118_), .B(_87_), .Y(_119_) );
NOR2X1 NOR2X1_20 ( .A(_117_), .B(_119_), .Y(_120_) );
NOR2X1 NOR2X1_21 ( .A(CORE_InstructionIN[10]), .B(CORE_InstructionIN[11]), .Y(_121_) );
INVX1 INVX1_18 ( .A(_121_), .Y(_122_) );
OAI21X1 OAI21X1_15 ( .A(_212__2_), .B(_102_), .C(_122_), .Y(_123_) );
NOR2X1 NOR2X1_22 ( .A(_123_), .B(_101_), .Y(_124_) );
AOI21X1 AOI21X1_11 ( .A(_115_), .B(_120_), .C(_124_), .Y(_125_) );
OAI21X1 OAI21X1_16 ( .A(_125_), .B(CORE_InstructionIN_15_bF_buf2), .C(_113_), .Y(_2__2_) );
AOI21X1 AOI21X1_12 ( .A(CORE_InstructionIN[13]), .B(CORE_InstructionIN[12]), .C(CORE_InstructionIN[14]), .Y(_126_) );
OAI21X1 OAI21X1_17 ( .A(_27_), .B(_210_), .C(_16__bF_buf2), .Y(_127_) );
NOR2X1 NOR2X1_23 ( .A(_126_), .B(_127_), .Y(_0_) );
INVX1 INVX1_19 ( .A(_83_), .Y(_128_) );
INVX1 INVX1_20 ( .A(_85_), .Y(_129_) );
NOR2X1 NOR2X1_24 ( .A(_129_), .B(_88_), .Y(_130_) );
OAI21X1 OAI21X1_18 ( .A(_130_), .B(_28_), .C(_213_), .Y(_131_) );
OAI21X1 OAI21X1_19 ( .A(_128_), .B(_88_), .C(_131_), .Y(_3_) );
OAI21X1 OAI21X1_20 ( .A(_27_), .B(_214_), .C(_16__bF_buf1), .Y(_132_) );
NOR2X1 NOR2X1_25 ( .A(_126_), .B(_132_), .Y(_4_) );
INVX1 INVX1_21 ( .A(CORE_InstructionIN[12]), .Y(_133_) );
OAI21X1 OAI21X1_21 ( .A(_133_), .B(CORE_InstructionIN[14]), .C(_16__bF_buf0), .Y(_134_) );
AOI21X1 AOI21X1_13 ( .A(_30_), .B(_62_), .C(_134_), .Y(_135_) );
NAND2X1 NAND2X1_20 ( .A(CORE_InstructionIN[11]), .B(_30_), .Y(_136_) );
AOI21X1 AOI21X1_14 ( .A(_136_), .B(_20_), .C(CORE_InstructionIN[14]), .Y(_137_) );
NAND2X1 NAND2X1_21 ( .A(_221__0_), .B(_16__bF_buf3), .Y(_138_) );
OAI22X1 OAI22X1_3 ( .A(_137_), .B(_138_), .C(_135_), .D(_34_), .Y(_11__0_) );
NAND2X1 NAND2X1_22 ( .A(_221__1_), .B(_16__bF_buf2), .Y(_139_) );
OAI22X1 OAI22X1_4 ( .A(_137_), .B(_139_), .C(_135_), .D(_37_), .Y(_11__1_) );
NAND2X1 NAND2X1_23 ( .A(_221__2_), .B(_16__bF_buf1), .Y(_140_) );
OAI22X1 OAI22X1_5 ( .A(_137_), .B(_140_), .C(_135_), .D(_39_), .Y(_11__2_) );
NAND2X1 NAND2X1_24 ( .A(_221__3_), .B(_16__bF_buf0), .Y(_141_) );
OAI22X1 OAI22X1_6 ( .A(_137_), .B(_141_), .C(_135_), .D(_41_), .Y(_11__3_) );
NOR2X1 NOR2X1_26 ( .A(_53_), .B(_17_), .Y(_142_) );
AOI21X1 AOI21X1_15 ( .A(_30_), .B(_142_), .C(CORE_InstructionIN_15_bF_buf1), .Y(_143_) );
INVX1 INVX1_22 ( .A(_220__0_), .Y(_144_) );
AOI21X1 AOI21X1_16 ( .A(_144_), .B(_136_), .C(_61_), .Y(_145_) );
OAI21X1 OAI21X1_22 ( .A(_143_), .B(CORE_InstructionIN[4]), .C(_145_), .Y(_146_) );
OAI21X1 OAI21X1_23 ( .A(_90_), .B(CORE_InstructionIN_15_bF_buf0), .C(CORE_InstructionIN[4]), .Y(_147_) );
AOI21X1 AOI21X1_17 ( .A(CORE_InstructionIN[11]), .B(_144_), .C(_57_), .Y(_148_) );
OAI21X1 OAI21X1_24 ( .A(_121_), .B(CORE_InstructionIN_15_bF_buf3), .C(_43_), .Y(_149_) );
AOI22X1 AOI22X1_4 ( .A(_220__0_), .B(_28_), .C(_148_), .D(_149_), .Y(_150_) );
NAND3X1 NAND3X1_9 ( .A(_146_), .B(_147_), .C(_150_), .Y(_10__0_) );
NOR2X1 NOR2X1_27 ( .A(_17_), .B(_57_), .Y(_151_) );
OAI21X1 OAI21X1_25 ( .A(_17_), .B(_31_), .C(_20_), .Y(_152_) );
NAND2X1 NAND2X1_25 ( .A(_27_), .B(_152_), .Y(_153_) );
NOR2X1 NOR2X1_28 ( .A(_151_), .B(_153_), .Y(_154_) );
NAND2X1 NAND2X1_26 ( .A(_220__1_), .B(_16__bF_buf3), .Y(_155_) );
NAND2X1 NAND2X1_27 ( .A(CORE_InstructionIN[8]), .B(_30_), .Y(_156_) );
NOR2X1 NOR2X1_29 ( .A(_156_), .B(_72_), .Y(_157_) );
OAI21X1 OAI21X1_26 ( .A(_18_), .B(CORE_InstructionIN[14]), .C(_16__bF_buf2), .Y(_158_) );
INVX1 INVX1_23 ( .A(_158_), .Y(_159_) );
OAI21X1 OAI21X1_27 ( .A(_57_), .B(_122_), .C(_159_), .Y(_160_) );
OAI21X1 OAI21X1_28 ( .A(_157_), .B(_160_), .C(CORE_InstructionIN[5]), .Y(_161_) );
OAI21X1 OAI21X1_29 ( .A(_154_), .B(_155_), .C(_161_), .Y(_10__1_) );
NAND2X1 NAND2X1_28 ( .A(_220__2_), .B(_16__bF_buf1), .Y(_162_) );
OAI21X1 OAI21X1_30 ( .A(_157_), .B(_160_), .C(CORE_InstructionIN[6]), .Y(_163_) );
OAI21X1 OAI21X1_31 ( .A(_154_), .B(_162_), .C(_163_), .Y(_10__2_) );
NAND2X1 NAND2X1_29 ( .A(_220__3_), .B(_16__bF_buf0), .Y(_164_) );
OAI21X1 OAI21X1_32 ( .A(_157_), .B(_160_), .C(CORE_InstructionIN[7]), .Y(_165_) );
OAI21X1 OAI21X1_33 ( .A(_154_), .B(_164_), .C(_165_), .Y(_10__3_) );
NOR2X1 NOR2X1_30 ( .A(_219__0_), .B(_158_), .Y(_166_) );
AOI21X1 AOI21X1_18 ( .A(_53_), .B(_158_), .C(_166_), .Y(_9__0_) );
NOR2X1 NOR2X1_31 ( .A(_219__1_), .B(_158_), .Y(_167_) );
AOI21X1 AOI21X1_19 ( .A(_50_), .B(_158_), .C(_167_), .Y(_9__1_) );
NOR2X1 NOR2X1_32 ( .A(_219__2_), .B(_158_), .Y(_168_) );
AOI21X1 AOI21X1_20 ( .A(_23_), .B(_158_), .C(_168_), .Y(_9__2_) );
NOR2X1 NOR2X1_33 ( .A(_219__3_), .B(_158_), .Y(_169_) );
AOI21X1 AOI21X1_21 ( .A(_17_), .B(_107_), .C(_169_), .Y(_9__3_) );
NAND2X1 NAND2X1_30 ( .A(_126_), .B(_152_), .Y(_170_) );
NAND2X1 NAND2X1_31 ( .A(_225__0_), .B(_170_), .Y(_171_) );
OAI21X1 OAI21X1_34 ( .A(_99_), .B(_17_), .C(_57_), .Y(_172_) );
NAND2X1 NAND2X1_32 ( .A(CORE_InstructionIN_15_bF_buf2), .B(_172_), .Y(_173_) );
OAI21X1 OAI21X1_35 ( .A(_171_), .B(CORE_InstructionIN_15_bF_buf1), .C(_173_), .Y(_15__0_) );
OAI21X1 OAI21X1_36 ( .A(_27_), .B(_133_), .C(_99_), .Y(_174_) );
AOI21X1 AOI21X1_22 ( .A(CORE_InstructionIN[11]), .B(_108_), .C(_174_), .Y(_175_) );
NAND3X1 NAND3X1_10 ( .A(_16__bF_buf3), .B(_225__1_), .C(_170_), .Y(_176_) );
OAI21X1 OAI21X1_37 ( .A(_16__bF_buf2), .B(_175_), .C(_176_), .Y(_15__1_) );
OAI21X1 OAI21X1_38 ( .A(CORE_InstructionIN[14]), .B(CORE_InstructionIN[12]), .C(CORE_InstructionIN[13]), .Y(_177_) );
NAND3X1 NAND3X1_11 ( .A(_16__bF_buf1), .B(_225__2_), .C(_170_), .Y(_178_) );
OAI21X1 OAI21X1_39 ( .A(_16__bF_buf0), .B(_177_), .C(_178_), .Y(_15__2_) );
NAND3X1 NAND3X1_12 ( .A(_16__bF_buf3), .B(_225__3_), .C(_170_), .Y(_179_) );
OAI21X1 OAI21X1_40 ( .A(_16__bF_buf2), .B(_27_), .C(_179_), .Y(_15__3_) );
NOR2X1 NOR2X1_34 ( .A(CORE_InstructionIN_15_bF_buf0), .B(_61_), .Y(_180_) );
AOI22X1 AOI22X1_5 ( .A(CORE_InstructionIN_15_bF_buf3), .B(_91_), .C(_180_), .D(_25_), .Y(_181_) );
AND2X2 AND2X2_3 ( .A(_16__bF_buf1), .B(_217__0_), .Y(_182_) );
OAI21X1 OAI21X1_41 ( .A(_170_), .B(_151_), .C(_182_), .Y(_183_) );
OAI21X1 OAI21X1_42 ( .A(_17_), .B(_181_), .C(_183_), .Y(_7__0_) );
INVX1 INVX1_24 ( .A(_217__1_), .Y(_184_) );
OR2X2 OR2X2_4 ( .A(_126_), .B(_184_), .Y(_185_) );
OAI21X1 OAI21X1_43 ( .A(_136_), .B(_61_), .C(_184_), .Y(_186_) );
OAI21X1 OAI21X1_44 ( .A(_151_), .B(_20_), .C(_186_), .Y(_187_) );
AOI21X1 AOI21X1_23 ( .A(_185_), .B(_187_), .C(CORE_InstructionIN_15_bF_buf2), .Y(_7__1_) );
NOR2X1 NOR2X1_35 ( .A(CORE_InstructionIN[4]), .B(CORE_InstructionIN[5]), .Y(_188_) );
NOR2X1 NOR2X1_36 ( .A(CORE_InstructionIN[6]), .B(CORE_InstructionIN[7]), .Y(_189_) );
NAND2X1 NAND2X1_33 ( .A(_188_), .B(_189_), .Y(_190_) );
NOR2X1 NOR2X1_37 ( .A(_190_), .B(_156_), .Y(_191_) );
NAND2X1 NAND2X1_34 ( .A(_98_), .B(_191_), .Y(_192_) );
OAI21X1 OAI21X1_45 ( .A(_192_), .B(_21_), .C(_224__0_), .Y(_193_) );
NAND2X1 NAND2X1_35 ( .A(_129_), .B(_191_), .Y(_194_) );
OAI21X1 OAI21X1_46 ( .A(_21_), .B(_194_), .C(_193_), .Y(_14__0_) );
INVX1 INVX1_25 ( .A(_94_), .Y(_195_) );
OAI21X1 OAI21X1_47 ( .A(_34_), .B(_37_), .C(_195_), .Y(_196_) );
INVX1 INVX1_26 ( .A(_190_), .Y(_197_) );
NAND3X1 NAND3X1_13 ( .A(_53_), .B(_50_), .C(_121_), .Y(_198_) );
INVX1 INVX1_27 ( .A(_198_), .Y(_199_) );
NAND3X1 NAND3X1_14 ( .A(_197_), .B(_199_), .C(_180_), .Y(_200_) );
NAND2X1 NAND2X1_36 ( .A(_199_), .B(_180_), .Y(_201_) );
NOR2X1 NOR2X1_38 ( .A(_34_), .B(_37_), .Y(_202_) );
NAND3X1 NAND3X1_15 ( .A(_84_), .B(_202_), .C(_197_), .Y(_203_) );
OAI21X1 OAI21X1_48 ( .A(_201_), .B(_203_), .C(_224__1_), .Y(_204_) );
OAI21X1 OAI21X1_49 ( .A(_196_), .B(_200_), .C(_204_), .Y(_14__1_) );
OAI21X1 OAI21X1_50 ( .A(_200_), .B(_196_), .C(_224__2_), .Y(_205_) );
OAI21X1 OAI21X1_51 ( .A(_118_), .B(_200_), .C(_205_), .Y(_14__2_) );
INVX1 INVX1_28 ( .A(_224__3_), .Y(_206_) );
NAND2X1 NAND2X1_37 ( .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[9]), .Y(_207_) );
NOR2X1 NOR2X1_39 ( .A(_207_), .B(_102_), .Y(_208_) );
AOI21X1 AOI21X1_24 ( .A(_208_), .B(_180_), .C(_206_), .Y(_14__3_) );
NAND2X1 NAND2X1_38 ( .A(_222_), .B(_78_), .Y(_209_) );
NAND3X1 NAND3X1_16 ( .A(_16__bF_buf0), .B(_99_), .C(_209_), .Y(_12_) );
BUFX2 BUFX2_1 ( .A(_210_), .Y(CORE_DATA_ADDR_mux) );
BUFX2 BUFX2_2 ( .A(_211_), .Y(CORE_DATA_REGMux) );
BUFX2 BUFX2_3 ( .A(_212__0_), .Y(CORE_DATA_ctrl[0]) );
BUFX2 BUFX2_4 ( .A(_212__1_), .Y(CORE_DATA_ctrl[1]) );
BUFX2 BUFX2_5 ( .A(_212__2_), .Y(CORE_DATA_ctrl[2]) );
BUFX2 BUFX2_6 ( .A(_213_), .Y(CORE_DATA_load) );
BUFX2 BUFX2_7 ( .A(_214_), .Y(CORE_DATA_write) );
BUFX2 BUFX2_8 ( .A(_215__0_), .Y(CORE_INT_CHA[0]) );
BUFX2 BUFX2_9 ( .A(_215__1_), .Y(CORE_INT_CHA[1]) );
BUFX2 BUFX2_10 ( .A(_215__2_), .Y(CORE_INT_CHA[2]) );
BUFX2 BUFX2_11 ( .A(_215__3_), .Y(CORE_INT_CHA[3]) );
BUFX2 BUFX2_12 ( .A(_215__4_), .Y(CORE_INT_CHA[4]) );
BUFX2 BUFX2_13 ( .A(_215__5_), .Y(CORE_INT_CHA[5]) );
BUFX2 BUFX2_14 ( .A(_215__6_), .Y(CORE_INT_CHA[6]) );
BUFX2 BUFX2_15 ( .A(_215__7_), .Y(CORE_INT_CHA[7]) );
BUFX2 BUFX2_16 ( .A(_216__0_), .Y(CORE_INT_ctrl[0]) );
BUFX2 BUFX2_17 ( .A(_216__1_), .Y(CORE_INT_ctrl[1]) );
BUFX2 BUFX2_18 ( .A(_217__0_), .Y(CORE_InstructionToULAMux[0]) );
BUFX2 BUFX2_19 ( .A(_217__1_), .Y(CORE_InstructionToULAMux[1]) );
BUFX2 BUFX2_20 ( .A(_undef), .Y(CORE_PC_clk) );
BUFX2 BUFX2_21 ( .A(_218__0_), .Y(CORE_PC_ctrl[0]) );
BUFX2 BUFX2_22 ( .A(_218__1_), .Y(CORE_PC_ctrl[1]) );
BUFX2 BUFX2_23 ( .A(_219__0_), .Y(CORE_REG_RD[0]) );
BUFX2 BUFX2_24 ( .A(_219__1_), .Y(CORE_REG_RD[1]) );
BUFX2 BUFX2_25 ( .A(_219__2_), .Y(CORE_REG_RD[2]) );
BUFX2 BUFX2_26 ( .A(_219__3_), .Y(CORE_REG_RD[3]) );
BUFX2 BUFX2_27 ( .A(_220__0_), .Y(CORE_REG_RF1[0]) );
BUFX2 BUFX2_28 ( .A(_220__1_), .Y(CORE_REG_RF1[1]) );
BUFX2 BUFX2_29 ( .A(_220__2_), .Y(CORE_REG_RF1[2]) );
BUFX2 BUFX2_30 ( .A(_220__3_), .Y(CORE_REG_RF1[3]) );
BUFX2 BUFX2_31 ( .A(_221__0_), .Y(CORE_REG_RF2[0]) );
BUFX2 BUFX2_32 ( .A(_221__1_), .Y(CORE_REG_RF2[1]) );
BUFX2 BUFX2_33 ( .A(_221__2_), .Y(CORE_REG_RF2[2]) );
BUFX2 BUFX2_34 ( .A(_221__3_), .Y(CORE_REG_RF2[3]) );
BUFX2 BUFX2_35 ( .A(_222_), .Y(CORE_REG_write) );
BUFX2 BUFX2_36 ( .A(_223__0_), .Y(CORE_STACK_ctrl[0]) );
BUFX2 BUFX2_37 ( .A(_223__1_), .Y(CORE_STACK_ctrl[1]) );
BUFX2 BUFX2_38 ( .A(_224__0_), .Y(CORE_Status_ctrl[0]) );
BUFX2 BUFX2_39 ( .A(_224__1_), .Y(CORE_Status_ctrl[1]) );
BUFX2 BUFX2_40 ( .A(_224__2_), .Y(CORE_Status_ctrl[2]) );
BUFX2 BUFX2_41 ( .A(_224__3_), .Y(CORE_Status_ctrl[3]) );
BUFX2 BUFX2_42 ( .A(_undef), .Y(CORE_Status_ctrl[4]) );
BUFX2 BUFX2_43 ( .A(_undef), .Y(CORE_ULAMux_inc_dec) );
BUFX2 BUFX2_44 ( .A(_225__0_), .Y(CORE_ULA_ctrl[0]) );
BUFX2 BUFX2_45 ( .A(_225__1_), .Y(CORE_ULA_ctrl[1]) );
BUFX2 BUFX2_46 ( .A(_225__2_), .Y(CORE_ULA_ctrl[2]) );
BUFX2 BUFX2_47 ( .A(_225__3_), .Y(CORE_ULA_ctrl[3]) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf5), .D(_14__0_), .Q(_224__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf4), .D(_14__1_), .Q(_224__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf3), .D(_14__2_), .Q(_224__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf2), .D(_14__3_), .Q(_224__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf1), .D(_7__0_), .Q(_217__0_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf0), .D(_7__1_), .Q(_217__1_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf5), .D(_15__0_), .Q(_225__0_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf4), .D(_15__1_), .Q(_225__1_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf3), .D(_15__2_), .Q(_225__2_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf2), .D(_15__3_), .Q(_225__3_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf1), .D(_9__0_), .Q(_219__0_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf0), .D(_9__1_), .Q(_219__1_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf5), .D(_9__2_), .Q(_219__2_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf4), .D(_9__3_), .Q(_219__3_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf3), .D(_10__0_), .Q(_220__0_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf2), .D(_10__1_), .Q(_220__1_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf1), .D(_10__2_), .Q(_220__2_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf0), .D(_10__3_), .Q(_220__3_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf5), .D(_11__0_), .Q(_221__0_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf4), .D(_11__1_), .Q(_221__1_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf3), .D(_11__2_), .Q(_221__2_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf2), .D(_11__3_), .Q(_221__3_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf1), .D(_12_), .Q(_222_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf0), .D(_4_), .Q(_214_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf5), .D(_3_), .Q(_213_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf4), .D(_0_), .Q(_210_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf3), .D(_2__0_), .Q(_212__0_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf2), .D(_2__1_), .Q(_212__1_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf1), .D(_2__2_), .Q(_212__2_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf0), .D(_1_), .Q(_211_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf5), .D(_13__0_), .Q(_223__0_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf4), .D(_13__1_), .Q(_223__1_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf3), .D(_8__0_), .Q(_218__0_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf2), .D(_8__1_), .Q(_218__1_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf1), .D(_5__0_), .Q(_215__0_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf0), .D(_5__1_), .Q(_215__1_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf5), .D(_5__2_), .Q(_215__2_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf4), .D(_5__3_), .Q(_215__3_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf3), .D(_5__4_), .Q(_215__4_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf2), .D(_5__5_), .Q(_215__5_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf1), .D(_5__6_), .Q(_215__6_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf0), .D(_5__7_), .Q(_215__7_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf5), .D(_6__0_), .Q(_216__0_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf4), .D(_6__1_), .Q(_216__1_) );
endmodule
