magic
tech scmos
magscale 1 4
timestamp 1515852544
<< metal1 >>
rect 1928 4777 1955 4783
rect 3309 4737 3336 4743
rect 4877 4717 4888 4723
rect 4909 4717 4931 4723
rect 93 4697 131 4703
rect 829 4697 851 4703
rect 845 4683 851 4697
rect 1000 4697 1011 4703
rect 2044 4703 2052 4706
rect 2029 4697 2052 4703
rect 4012 4703 4020 4708
rect 3981 4697 4020 4703
rect 4141 4697 4168 4703
rect 4252 4703 4260 4706
rect 4252 4697 4275 4703
rect 4396 4703 4404 4708
rect 4396 4697 4435 4703
rect 4829 4697 4840 4703
rect 4909 4703 4915 4717
rect 4861 4697 4915 4703
rect 5080 4697 5107 4703
rect 5868 4703 5876 4706
rect 5868 4697 5896 4703
rect 5981 4697 6008 4703
rect 845 4677 883 4683
rect 3688 4677 3699 4683
rect 3960 4677 3971 4683
rect 4712 4677 4723 4683
rect 4776 4677 4787 4683
rect 5661 4677 5700 4683
rect 152 4657 163 4663
rect 205 4657 227 4663
rect 381 4657 403 4663
rect 669 4657 691 4663
rect 957 4657 979 4663
rect 6717 4657 6739 4663
rect 93 4517 116 4523
rect 108 4514 116 4517
rect 1165 4517 1203 4523
rect 1197 4497 1203 4517
rect 1309 4523 1315 4543
rect 1805 4537 1816 4543
rect 3272 4537 3283 4543
rect 3720 4537 3731 4543
rect 4344 4537 4355 4543
rect 4648 4537 4659 4543
rect 1288 4517 1315 4523
rect 1341 4517 1379 4523
rect 1469 4517 1508 4523
rect 1500 4512 1508 4517
rect 1629 4517 1667 4523
rect 1677 4517 1688 4523
rect 1741 4517 1779 4523
rect 1741 4497 1747 4517
rect 1816 4517 1875 4523
rect 1885 4517 1923 4523
rect 1917 4497 1923 4517
rect 2173 4517 2211 4523
rect 2509 4517 2547 4523
rect 1933 4497 1971 4503
rect 2541 4497 2547 4517
rect 2717 4517 2755 4523
rect 2861 4517 2899 4523
rect 2632 4497 2643 4503
rect 2861 4503 2867 4517
rect 3037 4517 3075 4523
rect 2829 4497 2867 4503
rect 3037 4497 3043 4517
rect 3197 4517 3235 4523
rect 3256 4517 3267 4523
rect 3373 4517 3411 4523
rect 3373 4497 3379 4517
rect 3597 4517 3635 4523
rect 3629 4497 3635 4517
rect 3848 4517 3859 4523
rect 3917 4517 3987 4523
rect 4157 4517 4195 4523
rect 4408 4517 4419 4523
rect 4536 4517 4547 4523
rect 4557 4517 4595 4523
rect 3837 4497 3843 4512
rect 3944 4497 3971 4503
rect 4445 4497 4456 4503
rect 4552 4496 4556 4504
rect 4589 4497 4595 4517
rect 4733 4523 4739 4543
rect 5821 4537 5843 4543
rect 6109 4537 6147 4543
rect 4728 4517 4739 4523
rect 4925 4517 4968 4523
rect 5160 4517 5187 4523
rect 5309 4517 5347 4523
rect 5341 4497 5347 4517
rect 5805 4517 5816 4523
rect 6696 4517 6707 4523
rect 5384 4497 5395 4503
rect 5501 4497 5523 4503
rect 2328 4476 2330 4484
rect 2605 4477 2632 4483
rect 6342 4476 6344 4484
rect 6632 4476 6634 4484
rect 2508 4337 2520 4343
rect 2508 4332 2516 4337
rect 6781 4337 6808 4343
rect 541 4317 579 4323
rect 733 4317 744 4323
rect 1064 4316 1068 4324
rect 125 4297 163 4303
rect 253 4297 280 4303
rect 696 4297 707 4303
rect 760 4297 771 4303
rect 781 4297 824 4303
rect 984 4297 995 4303
rect 1837 4297 1880 4303
rect 2077 4303 2083 4323
rect 2045 4297 2083 4303
rect 2173 4303 2179 4323
rect 2829 4317 2840 4323
rect 2968 4316 2972 4324
rect 3144 4317 3155 4323
rect 3229 4317 3267 4323
rect 3805 4317 3816 4323
rect 3853 4317 3880 4323
rect 2173 4297 2195 4303
rect 2253 4297 2291 4303
rect 2461 4297 2472 4303
rect 2524 4303 2532 4308
rect 2493 4297 2532 4303
rect 2637 4297 2648 4303
rect 2952 4297 2963 4303
rect 3000 4297 3011 4303
rect 3309 4297 3320 4303
rect 4061 4303 4067 4323
rect 4061 4297 4099 4303
rect 4109 4297 4147 4303
rect 1112 4277 1123 4283
rect 2445 4277 2456 4283
rect 4141 4283 4147 4297
rect 4200 4297 4211 4303
rect 4333 4303 4339 4323
rect 4408 4316 4412 4324
rect 4301 4297 4339 4303
rect 4477 4297 4515 4303
rect 4856 4297 4867 4303
rect 4141 4277 4163 4283
rect 4989 4277 4995 4292
rect 5373 4303 5379 4323
rect 5565 4317 5587 4323
rect 5341 4297 5379 4303
rect 6424 4297 6435 4303
rect 5037 4277 5059 4283
rect 5421 4277 5427 4292
rect 5624 4277 5635 4283
rect 5816 4277 5827 4283
rect 5853 4277 5891 4283
rect 5832 4256 5836 4264
rect 3373 4157 3384 4163
rect 188 4137 212 4143
rect 536 4137 547 4143
rect 781 4137 824 4143
rect 1133 4137 1144 4143
rect 1693 4137 1720 4143
rect 1773 4137 1784 4143
rect 1880 4137 1896 4143
rect 2152 4137 2163 4143
rect 2189 4137 2200 4143
rect 2840 4137 2851 4143
rect 2904 4137 2947 4143
rect 3341 4137 3363 4143
rect 3597 4137 3608 4143
rect 3656 4137 3667 4143
rect 3736 4137 3747 4143
rect 3773 4137 3784 4143
rect 3880 4137 3912 4143
rect 4701 4143 4707 4163
rect 4637 4137 4675 4143
rect 4701 4137 4739 4143
rect 4749 4137 4787 4143
rect 5085 4137 5096 4143
rect 5165 4137 5176 4143
rect 5309 4137 5347 4143
rect 6136 4137 6147 4143
rect 269 4117 296 4123
rect 472 4117 483 4123
rect 493 4117 531 4123
rect 637 4117 664 4123
rect 525 4097 531 4117
rect 1048 4117 1075 4123
rect 1149 4117 1187 4123
rect 797 4097 824 4103
rect 1037 4097 1048 4103
rect 1149 4097 1155 4117
rect 1645 4117 1656 4123
rect 1789 4117 1800 4123
rect 1933 4117 1971 4123
rect 1373 4097 1384 4103
rect 1933 4097 1939 4117
rect 2088 4117 2099 4123
rect 2109 4117 2147 4123
rect 2621 4117 2659 4123
rect 2221 4088 2227 4103
rect 2308 4096 2312 4104
rect 2509 4097 2520 4103
rect 2653 4097 2659 4117
rect 2797 4117 2835 4123
rect 2893 4117 2904 4123
rect 2973 4117 3011 4123
rect 3005 4097 3011 4117
rect 3149 4117 3187 4123
rect 3101 4097 3139 4103
rect 3149 4097 3155 4117
rect 3384 4117 3395 4123
rect 3693 4117 3731 4123
rect 3789 4117 3800 4123
rect 3837 4117 3864 4123
rect 3965 4117 4003 4123
rect 4013 4117 4024 4123
rect 4397 4117 4424 4123
rect 4461 4117 4499 4123
rect 4493 4097 4499 4117
rect 4856 4117 4899 4123
rect 4909 4117 4979 4123
rect 4760 4097 4771 4103
rect 4973 4097 4979 4117
rect 5245 4117 5256 4123
rect 5533 4117 5544 4123
rect 5576 4117 5587 4123
rect 5933 4117 5992 4123
rect 6429 4117 6440 4123
rect 5773 4097 5795 4103
rect 6088 4096 6092 4104
rect 5789 4077 5800 4083
rect 4168 3937 4196 3943
rect 4908 3937 4936 3943
rect 4188 3932 4196 3937
rect 5736 3936 5738 3944
rect 6765 3937 6808 3943
rect 108 3903 116 3906
rect 93 3897 116 3903
rect 200 3897 227 3903
rect 653 3903 659 3923
rect 541 3897 579 3903
rect 637 3897 659 3903
rect 925 3903 931 3923
rect 856 3897 883 3903
rect 893 3897 931 3903
rect 1005 3897 1043 3903
rect 1117 3903 1123 3923
rect 1112 3897 1123 3903
rect 1373 3897 1384 3903
rect 1864 3897 1891 3903
rect 1917 3903 1923 3923
rect 1917 3897 1944 3903
rect 2061 3903 2067 3923
rect 2861 3917 2899 3923
rect 2061 3897 2099 3903
rect 2861 3903 2867 3917
rect 2808 3897 2819 3903
rect 2829 3897 2867 3903
rect 3069 3897 3107 3903
rect 3117 3897 3128 3903
rect 3352 3897 3379 3903
rect 3501 3897 3512 3903
rect 3741 3903 3747 3923
rect 3741 3897 3779 3903
rect 3912 3897 3923 3903
rect 3981 3897 4019 3903
rect 4172 3903 4180 3908
rect 4269 3903 4275 3923
rect 4408 3917 4419 3923
rect 4493 3917 4504 3923
rect 4797 3917 4808 3923
rect 4172 3897 4211 3903
rect 4269 3897 4307 3903
rect 4781 3897 4792 3903
rect 4952 3897 4979 3903
rect 5325 3903 5331 3923
rect 5272 3897 5283 3903
rect 5293 3897 5331 3903
rect 5784 3897 5811 3903
rect 6680 3897 6691 3903
rect 648 3877 659 3883
rect 1981 3877 1992 3883
rect 4573 3877 4611 3883
rect 3224 3856 3228 3864
rect 4573 3857 4579 3877
rect 4696 3877 4723 3883
rect 5005 3877 5043 3883
rect 5229 3877 5267 3883
rect 5373 3877 5384 3883
rect 5464 3877 5475 3883
rect 5501 3877 5512 3883
rect 6077 3877 6104 3883
rect 6396 3868 6404 3872
rect 5549 3857 5571 3863
rect 5976 3857 5987 3863
rect 861 3777 888 3783
rect 1764 3756 1768 3764
rect 2477 3757 2488 3763
rect 2861 3757 2888 3763
rect 3788 3757 3816 3763
rect 3788 3748 3796 3757
rect 6541 3757 6563 3763
rect 6653 3757 6675 3763
rect 541 3737 552 3743
rect 1340 3743 1348 3748
rect 1340 3737 1363 3743
rect 1624 3737 1635 3743
rect 1960 3737 1971 3743
rect 2397 3737 2424 3743
rect 2637 3737 2648 3743
rect 2749 3737 2771 3743
rect 3437 3737 3464 3743
rect 4285 3737 4296 3743
rect 5096 3737 5123 3743
rect 5229 3737 5256 3743
rect 6365 3737 6376 3743
rect 6781 3737 6808 3743
rect 349 3717 387 3723
rect 349 3697 355 3717
rect 605 3717 616 3723
rect 749 3717 776 3723
rect 1229 3717 1240 3723
rect 1485 3717 1528 3723
rect 1672 3717 1699 3723
rect 1917 3717 1955 3723
rect 2776 3717 2787 3723
rect 2941 3717 2979 3723
rect 2941 3697 2947 3717
rect 3496 3717 3507 3723
rect 3613 3717 3651 3723
rect 3645 3697 3651 3717
rect 4381 3717 4392 3723
rect 4685 3717 4723 3723
rect 3661 3697 3699 3703
rect 4685 3697 4691 3717
rect 4744 3717 4755 3723
rect 5149 3717 5160 3723
rect 5656 3717 5683 3723
rect 6077 3717 6088 3723
rect 6184 3717 6195 3723
rect 6696 3717 6707 3723
rect 5357 3697 5379 3703
rect 6093 3697 6115 3703
rect 6509 3697 6520 3703
rect 3224 3537 3235 3543
rect 3848 3537 3859 3543
rect 4888 3537 4915 3543
rect 5741 3537 5752 3543
rect 5864 3537 5907 3543
rect 301 3517 339 3523
rect 493 3517 504 3523
rect 77 3497 104 3503
rect 541 3497 552 3503
rect 605 3497 632 3503
rect 669 3503 675 3523
rect 781 3517 819 3523
rect 669 3497 707 3503
rect 813 3503 819 3517
rect 1709 3517 1731 3523
rect 2061 3517 2083 3523
rect 2189 3517 2227 3523
rect 2664 3517 2675 3523
rect 813 3497 851 3503
rect 1052 3503 1060 3508
rect 1052 3497 1091 3503
rect 1208 3497 1235 3503
rect 1437 3497 1464 3503
rect 1613 3497 1640 3503
rect 1292 3477 1331 3483
rect 1613 3477 1619 3497
rect 1928 3497 1939 3503
rect 2024 3497 2035 3503
rect 2124 3497 2147 3503
rect 2124 3492 2132 3497
rect 2376 3497 2387 3503
rect 2397 3497 2435 3503
rect 3245 3503 3251 3523
rect 3869 3517 3907 3523
rect 3245 3497 3283 3503
rect 3389 3497 3427 3503
rect 3772 3503 3780 3508
rect 3741 3497 3780 3503
rect 3901 3503 3907 3517
rect 3901 3497 3939 3503
rect 4205 3503 4211 3523
rect 4205 3497 4243 3503
rect 4253 3497 4264 3503
rect 5213 3503 5219 3523
rect 5213 3497 5251 3503
rect 5496 3497 5523 3503
rect 5656 3497 5667 3503
rect 5832 3497 5843 3503
rect 5944 3497 5971 3503
rect 6109 3497 6120 3503
rect 6237 3503 6243 3523
rect 6237 3497 6275 3503
rect 6285 3497 6296 3503
rect 6392 3497 6403 3503
rect 2984 3477 2995 3483
rect 1852 3463 1860 3472
rect 1852 3457 1880 3463
rect 2989 3457 2995 3477
rect 3336 3477 3347 3483
rect 4552 3477 4563 3483
rect 5272 3477 5299 3483
rect 5976 3477 5987 3483
rect 6013 3477 6024 3483
rect 6093 3477 6131 3483
rect 6680 3477 6691 3483
rect 6701 3477 6739 3483
rect 6588 3463 6596 3472
rect 6568 3457 6596 3463
rect 5912 3356 5916 3364
rect 6008 3357 6019 3363
rect 6093 3357 6104 3363
rect 6125 3357 6147 3363
rect 701 3337 723 3343
rect 221 3317 232 3323
rect 381 3317 392 3323
rect 717 3323 723 3337
rect 781 3337 792 3343
rect 1053 3337 1064 3343
rect 1144 3337 1155 3343
rect 1789 3337 1800 3343
rect 2285 3337 2296 3343
rect 4317 3337 4328 3343
rect 717 3317 755 3323
rect 1325 3317 1336 3323
rect 1612 3323 1620 3328
rect 1612 3317 1624 3323
rect 1704 3317 1715 3323
rect 1773 3317 1827 3323
rect 1837 3317 1864 3323
rect 1997 3317 2036 3323
rect 2028 3312 2036 3317
rect 2200 3317 2227 3323
rect 2493 3317 2536 3323
rect 2797 3317 2808 3323
rect 2909 3317 2920 3323
rect 3213 3317 3224 3323
rect 3277 3317 3288 3323
rect 212 3296 216 3304
rect 781 3297 792 3303
rect 856 3296 860 3304
rect 2440 3297 2451 3303
rect 3277 3297 3283 3317
rect 3357 3317 3395 3323
rect 3725 3317 3763 3323
rect 3757 3297 3763 3317
rect 3880 3317 3923 3323
rect 3981 3317 3992 3323
rect 4077 3317 4104 3323
rect 4333 3317 4371 3323
rect 4445 3317 4483 3323
rect 3773 3297 3811 3303
rect 4445 3297 4451 3317
rect 4765 3317 4776 3323
rect 4861 3317 4920 3323
rect 4989 3323 4995 3343
rect 5064 3337 5075 3343
rect 5245 3337 5256 3343
rect 5821 3337 5832 3343
rect 6040 3337 6051 3343
rect 6253 3337 6291 3343
rect 4968 3317 4995 3323
rect 5325 3317 5336 3323
rect 5992 3317 6003 3323
rect 6445 3323 6451 3343
rect 6573 3337 6611 3343
rect 6445 3317 6467 3323
rect 6728 3317 6739 3323
rect 4548 3296 4552 3304
rect 4589 3288 4595 3303
rect 4792 3297 4803 3303
rect 6360 3296 6364 3304
rect 4221 3277 4232 3283
rect 4616 3277 4627 3283
rect 1837 3177 1864 3183
rect 797 3137 808 3143
rect 941 3137 1011 3143
rect 2909 3137 2936 3143
rect 5256 3137 5299 3143
rect 237 3103 243 3123
rect 237 3097 275 3103
rect 349 3103 355 3123
rect 349 3097 387 3103
rect 685 3097 696 3103
rect 728 3097 739 3103
rect 824 3097 851 3103
rect 1069 3103 1075 3123
rect 2221 3117 2232 3123
rect 2941 3117 2979 3123
rect 1069 3097 1107 3103
rect 1272 3097 1299 3103
rect 1533 3097 1560 3103
rect 2013 3097 2072 3103
rect 2157 3097 2211 3103
rect 2749 3097 2787 3103
rect 2989 3103 2995 3123
rect 2989 3097 3027 3103
rect 3053 3097 3064 3103
rect 3053 3088 3059 3097
rect 3101 3103 3107 3123
rect 3272 3116 3276 3124
rect 5752 3117 5763 3123
rect 3101 3097 3139 3103
rect 3149 3097 3176 3103
rect 3341 3097 3352 3103
rect 3405 3097 3443 3103
rect 3661 3097 3672 3103
rect 4221 3097 4248 3103
rect 4504 3097 4520 3103
rect 4872 3097 4952 3103
rect 5453 3097 5475 3103
rect 1629 3077 1640 3083
rect 2040 3077 2083 3083
rect 2317 3077 2376 3083
rect 2632 3077 2659 3083
rect 3544 3077 3571 3083
rect 3645 3077 3656 3083
rect 3773 3077 3784 3083
rect 5469 3077 5475 3097
rect 5528 3097 5539 3103
rect 5560 3097 5571 3103
rect 5693 3097 5704 3103
rect 5837 3097 5875 3103
rect 6044 3103 6052 3108
rect 6044 3097 6083 3103
rect 6700 3106 6708 3112
rect 6141 3077 6152 3083
rect 1357 3057 1379 3063
rect 1389 3057 1400 3063
rect 2024 3057 2035 3063
rect 2664 3056 2668 3064
rect 4893 3057 4904 3063
rect 4952 3057 4963 3063
rect 5037 3057 5059 3063
rect 5229 3037 5240 3043
rect 4909 2977 4920 2983
rect 1140 2956 1144 2964
rect 1853 2957 1880 2963
rect 2860 2948 2868 2952
rect 232 2937 243 2943
rect 1149 2937 1160 2943
rect 2109 2937 2120 2943
rect 2173 2937 2184 2943
rect 2285 2937 2312 2943
rect 3160 2937 3171 2943
rect 4120 2937 4147 2943
rect 4364 2937 4376 2943
rect 4637 2937 4648 2943
rect 4968 2937 4979 2943
rect 5229 2937 5251 2943
rect 5656 2937 5667 2943
rect 5949 2937 6003 2943
rect 6024 2937 6051 2943
rect 77 2917 104 2923
rect 477 2917 515 2923
rect 477 2897 483 2917
rect 829 2917 856 2923
rect 1309 2917 1320 2923
rect 1548 2923 1556 2928
rect 1548 2917 1560 2923
rect 1581 2917 1620 2923
rect 1612 2912 1620 2917
rect 2301 2917 2312 2923
rect 2461 2917 2499 2923
rect 516 2896 520 2904
rect 2493 2897 2499 2917
rect 2573 2917 2611 2923
rect 2605 2897 2611 2917
rect 3224 2917 3251 2923
rect 3288 2917 3315 2923
rect 4253 2917 4264 2923
rect 4509 2917 4520 2923
rect 4920 2917 4963 2923
rect 5565 2917 5603 2923
rect 2621 2897 2659 2903
rect 3256 2896 3260 2904
rect 3341 2897 3379 2903
rect 4548 2896 4552 2904
rect 4909 2897 4920 2903
rect 5597 2897 5603 2917
rect 5709 2917 5747 2923
rect 5757 2917 5795 2923
rect 5869 2917 5907 2923
rect 5757 2897 5763 2917
rect 5901 2897 5907 2917
rect 6093 2917 6131 2923
rect 6157 2923 6163 2943
rect 6781 2937 6808 2943
rect 6157 2917 6196 2923
rect 6188 2916 6196 2917
rect 6264 2917 6275 2923
rect 6301 2917 6339 2923
rect 6301 2897 6307 2917
rect 6461 2917 6499 2923
rect 6493 2897 6499 2917
rect 6568 2917 6579 2923
rect 2893 2837 2904 2843
rect 5976 2837 6003 2843
rect 5389 2737 5400 2743
rect 6312 2736 6314 2744
rect 348 2703 356 2706
rect 348 2697 371 2703
rect 429 2697 467 2703
rect 573 2697 584 2703
rect 765 2703 771 2723
rect 781 2717 851 2723
rect 733 2697 771 2703
rect 973 2697 1011 2703
rect 1021 2697 1032 2703
rect 1085 2703 1091 2723
rect 1085 2697 1123 2703
rect 1197 2703 1203 2723
rect 1197 2697 1235 2703
rect 1384 2697 1411 2703
rect 1432 2697 1459 2703
rect 957 2677 968 2683
rect 1453 2677 1459 2697
rect 1485 2697 1523 2703
rect 1725 2703 1731 2723
rect 1672 2697 1683 2703
rect 1693 2697 1731 2703
rect 1848 2697 1891 2703
rect 1917 2703 1923 2723
rect 4552 2717 4563 2723
rect 1912 2697 1923 2703
rect 2408 2697 2419 2703
rect 2600 2697 2659 2703
rect 2712 2697 2723 2703
rect 2776 2697 2787 2703
rect 1864 2677 1875 2683
rect 2445 2677 2472 2683
rect 2605 2677 2616 2683
rect 2669 2677 2680 2683
rect 2797 2683 2803 2703
rect 2824 2697 2835 2703
rect 2888 2697 2931 2703
rect 3224 2697 3235 2703
rect 3661 2697 3672 2703
rect 3725 2697 3736 2703
rect 4093 2697 4131 2703
rect 4189 2697 4200 2703
rect 4264 2697 4275 2703
rect 4749 2697 4760 2703
rect 4984 2697 4995 2703
rect 5005 2697 5043 2703
rect 5149 2703 5155 2723
rect 5325 2717 5336 2723
rect 5149 2697 5187 2703
rect 6008 2697 6019 2703
rect 2797 2677 2808 2683
rect 3197 2677 3208 2683
rect 3240 2677 3251 2683
rect 3677 2677 3699 2683
rect 3965 2677 3976 2683
rect 4136 2677 4147 2683
rect 6573 2697 6595 2703
rect 4605 2677 4616 2683
rect 4968 2677 4979 2683
rect 5085 2677 5096 2683
rect 5448 2677 5459 2683
rect 5517 2677 5555 2683
rect 5992 2677 6003 2683
rect 6589 2677 6595 2697
rect 6621 2697 6659 2703
rect 6664 2677 6675 2683
rect 2349 2657 2360 2663
rect 2493 2657 2536 2663
rect 5757 2657 5779 2663
rect 2861 2637 2888 2643
rect 2296 2576 2302 2584
rect 2237 2557 2264 2563
rect 2920 2556 2924 2564
rect 5101 2557 5112 2563
rect 589 2537 627 2543
rect 877 2537 915 2543
rect 1901 2537 1912 2543
rect 2189 2537 2200 2543
rect 2333 2537 2360 2543
rect 2845 2537 2856 2543
rect 2941 2537 2952 2543
rect 3085 2537 3096 2543
rect 3544 2537 3555 2543
rect 4013 2537 4024 2543
rect 93 2517 131 2523
rect 93 2497 99 2517
rect 301 2517 312 2523
rect 344 2517 355 2523
rect 536 2517 547 2523
rect 541 2497 547 2517
rect 765 2517 835 2523
rect 829 2497 835 2517
rect 1373 2517 1400 2523
rect 1549 2517 1560 2523
rect 1549 2497 1555 2517
rect 1741 2517 1779 2523
rect 1832 2517 1859 2523
rect 1917 2517 1939 2523
rect 1581 2497 1619 2503
rect 1933 2497 1939 2517
rect 2317 2517 2328 2523
rect 2461 2517 2500 2523
rect 2492 2512 2500 2517
rect 2701 2517 2712 2523
rect 2856 2517 2899 2523
rect 3032 2517 3043 2523
rect 3101 2517 3139 2523
rect 3277 2517 3315 2523
rect 2653 2497 2664 2503
rect 3277 2497 3283 2517
rect 3912 2517 3939 2523
rect 4077 2517 4115 2523
rect 3672 2497 3683 2503
rect 3784 2497 3795 2503
rect 4077 2497 4083 2517
rect 4157 2523 4163 2543
rect 4605 2537 4643 2543
rect 4136 2517 4163 2523
rect 4317 2517 4344 2523
rect 4429 2517 4440 2523
rect 4637 2517 4643 2537
rect 4760 2537 4771 2543
rect 5197 2537 5224 2543
rect 5992 2537 6019 2543
rect 6189 2537 6200 2543
rect 6408 2537 6419 2543
rect 6525 2537 6563 2543
rect 4893 2517 4947 2523
rect 4248 2496 4252 2504
rect 4861 2497 4872 2503
rect 4941 2503 4947 2517
rect 5053 2517 5091 2523
rect 5629 2517 5656 2523
rect 5901 2517 5912 2523
rect 5933 2517 5992 2523
rect 6317 2517 6355 2523
rect 6381 2517 6392 2523
rect 4941 2497 4963 2503
rect 6349 2497 6355 2517
rect 6621 2523 6627 2543
rect 6605 2517 6627 2523
rect 6669 2517 6707 2523
rect 6669 2497 6675 2517
rect 6728 2517 6739 2523
rect 1640 2477 1651 2483
rect 2568 2477 2579 2483
rect 3197 2477 3267 2483
rect 3868 2483 3876 2488
rect 3868 2477 3896 2483
rect 6540 2483 6548 2488
rect 6540 2477 6552 2483
rect 2397 2337 2451 2343
rect 3816 2337 3827 2343
rect 109 2317 147 2323
rect 404 2316 408 2324
rect 232 2297 243 2303
rect 301 2297 339 2303
rect 413 2297 440 2303
rect 477 2297 488 2303
rect 605 2297 643 2303
rect 701 2297 712 2303
rect 813 2297 824 2303
rect 973 2297 1011 2303
rect 1597 2303 1603 2323
rect 1917 2317 1928 2323
rect 1565 2297 1603 2303
rect 1741 2297 1779 2303
rect 2732 2306 2740 2312
rect 2872 2297 2883 2303
rect 3325 2303 3331 2323
rect 3293 2297 3331 2303
rect 3501 2297 3528 2303
rect 3693 2303 3699 2323
rect 3709 2317 3747 2323
rect 3661 2297 3699 2303
rect 3837 2303 3843 2323
rect 3837 2297 3875 2303
rect 4653 2303 4659 2323
rect 5384 2317 5395 2323
rect 5412 2316 5416 2324
rect 5992 2317 6003 2323
rect 4621 2297 4659 2303
rect 4957 2297 4968 2303
rect 5117 2297 5144 2303
rect 5277 2297 5288 2303
rect 5448 2297 5475 2303
rect 5677 2297 5688 2303
rect 5976 2297 6019 2303
rect 6029 2297 6040 2303
rect 6157 2297 6168 2303
rect 6493 2303 6499 2323
rect 6461 2297 6499 2303
rect 285 2277 296 2283
rect 696 2277 712 2283
rect 829 2277 840 2283
rect 872 2277 899 2283
rect 1053 2277 1064 2283
rect 1821 2277 1875 2283
rect 1949 2277 1971 2283
rect 2925 2277 2936 2283
rect 4237 2277 4248 2283
rect 4728 2277 4739 2283
rect 4765 2277 4792 2283
rect 5261 2277 5299 2283
rect 5341 2277 5363 2283
rect 5565 2277 5603 2283
rect 5709 2277 5715 2292
rect 5757 2277 5795 2283
rect 5949 2277 5960 2283
rect 1224 2256 1228 2264
rect 2525 2257 2556 2263
rect 6637 2157 6659 2163
rect 349 2137 371 2143
rect 1528 2137 1539 2143
rect 1965 2137 1976 2143
rect 2109 2137 2120 2143
rect 2429 2137 2451 2143
rect 2472 2137 2499 2143
rect 2904 2137 2915 2143
rect 3197 2137 3208 2143
rect 3885 2137 3928 2143
rect 4349 2137 4360 2143
rect 5356 2143 5364 2148
rect 5341 2137 5364 2143
rect 5532 2137 5556 2143
rect 5724 2143 5732 2148
rect 5724 2137 5747 2143
rect 6152 2137 6163 2143
rect 6333 2137 6344 2143
rect 477 2117 515 2123
rect 477 2097 483 2117
rect 648 2117 680 2123
rect 701 2117 739 2123
rect 733 2097 739 2117
rect 1736 2117 1747 2123
rect 1912 2117 1923 2123
rect 2029 2117 2067 2123
rect 2061 2097 2067 2117
rect 2317 2117 2328 2123
rect 2349 2117 2387 2123
rect 2765 2117 2792 2123
rect 2829 2117 2899 2123
rect 3069 2117 3107 2123
rect 2184 2097 2195 2103
rect 3069 2097 3075 2117
rect 3160 2117 3171 2123
rect 3181 2117 3192 2123
rect 3437 2117 3475 2123
rect 3501 2117 3512 2123
rect 3469 2097 3475 2117
rect 3544 2117 3555 2123
rect 3677 2117 3688 2123
rect 3725 2117 3763 2123
rect 3832 2117 3843 2123
rect 3837 2097 3843 2117
rect 4216 2117 4259 2123
rect 4269 2117 4307 2123
rect 4365 2117 4376 2123
rect 4477 2117 4515 2123
rect 4509 2097 4515 2117
rect 4760 2117 4787 2123
rect 5133 2117 5144 2123
rect 5165 2117 5203 2123
rect 5292 2117 5331 2123
rect 5292 2112 5300 2117
rect 5448 2117 5475 2123
rect 5757 2117 5795 2123
rect 4525 2097 4563 2103
rect 5789 2097 5795 2117
rect 5949 2117 6019 2123
rect 5949 2097 5955 2117
rect 6397 2117 6424 2123
rect 2989 2077 3059 2083
rect 5686 2076 5688 2084
rect 6120 2077 6131 2083
rect 189 1937 200 1943
rect 1302 1936 1304 1944
rect 2280 1937 2323 1943
rect 3494 1936 3496 1944
rect 477 1917 488 1923
rect 1464 1917 1475 1923
rect 1645 1917 1667 1923
rect 2280 1917 2291 1923
rect 2669 1917 2680 1923
rect 77 1897 104 1903
rect 252 1903 260 1908
rect 221 1897 260 1903
rect 381 1897 392 1903
rect 440 1897 451 1903
rect 525 1897 536 1903
rect 696 1897 707 1903
rect 925 1897 963 1903
rect 1229 1897 1256 1903
rect 1672 1897 1683 1903
rect 1880 1897 1923 1903
rect 2365 1897 2403 1903
rect 2653 1897 2664 1903
rect 2717 1903 2723 1923
rect 2717 1897 2755 1903
rect 2776 1897 2803 1903
rect 968 1877 979 1883
rect 1608 1877 1619 1883
rect 1853 1877 1880 1883
rect 2184 1877 2211 1883
rect 2445 1877 2467 1883
rect 2797 1877 2803 1897
rect 2989 1903 2995 1923
rect 2872 1897 2915 1903
rect 2989 1897 3027 1903
rect 3192 1897 3203 1903
rect 3272 1897 3283 1903
rect 3708 1903 3716 1906
rect 3704 1897 3716 1903
rect 4157 1897 4168 1903
rect 4221 1897 4232 1903
rect 4296 1897 4323 1903
rect 4621 1897 4659 1903
rect 4797 1903 4803 1923
rect 4984 1917 4995 1923
rect 4765 1897 4803 1903
rect 5085 1903 5091 1923
rect 5085 1897 5096 1903
rect 5261 1897 5299 1903
rect 5405 1903 5411 1923
rect 5757 1917 5779 1923
rect 5917 1917 5928 1923
rect 5405 1897 5443 1903
rect 5741 1897 5752 1903
rect 5965 1903 5971 1923
rect 5901 1897 5971 1903
rect 6093 1897 6104 1903
rect 6141 1897 6152 1903
rect 6264 1897 6291 1903
rect 3245 1877 3256 1883
rect 3884 1877 3944 1883
rect 4664 1877 4675 1883
rect 4957 1877 4984 1883
rect 5176 1877 5187 1883
rect 6077 1877 6088 1883
rect 6493 1877 6531 1883
rect 6685 1877 6739 1883
rect 6749 1877 6808 1883
rect 984 1856 988 1864
rect 6669 1757 6691 1763
rect 77 1717 104 1723
rect 301 1717 339 1723
rect 504 1717 515 1723
rect 525 1717 563 1723
rect 557 1697 563 1717
rect 600 1717 627 1723
rect 701 1717 739 1723
rect 733 1697 739 1717
rect 813 1717 851 1723
rect 845 1703 851 1717
rect 989 1717 1027 1723
rect 1053 1717 1064 1723
rect 845 1697 883 1703
rect 984 1696 988 1704
rect 1021 1697 1027 1717
rect 1213 1717 1224 1723
rect 1357 1723 1363 1743
rect 1389 1737 1416 1743
rect 1901 1737 1912 1743
rect 3101 1737 3112 1743
rect 3256 1737 3267 1743
rect 4376 1737 4387 1743
rect 1357 1717 1368 1723
rect 1485 1717 1496 1723
rect 1581 1723 1587 1732
rect 1576 1717 1587 1723
rect 1613 1717 1651 1723
rect 1645 1697 1651 1717
rect 1917 1717 1955 1723
rect 2344 1717 2355 1723
rect 2813 1717 2824 1723
rect 3037 1717 3075 1723
rect 3149 1717 3187 1723
rect 3245 1717 3256 1723
rect 3293 1717 3331 1723
rect 3325 1697 3331 1717
rect 3436 1717 3475 1723
rect 3436 1712 3444 1717
rect 3592 1717 3619 1723
rect 3725 1717 3763 1723
rect 4152 1717 4179 1723
rect 4205 1717 4216 1723
rect 3956 1696 3960 1704
rect 4173 1697 4179 1717
rect 4269 1717 4296 1723
rect 4333 1717 4371 1723
rect 4728 1717 4739 1723
rect 5005 1723 5011 1743
rect 5005 1717 5016 1723
rect 5581 1723 5587 1743
rect 6397 1737 6408 1743
rect 6717 1737 6755 1743
rect 5581 1717 5603 1723
rect 5789 1717 5800 1723
rect 5917 1717 5971 1723
rect 5965 1703 5971 1717
rect 6264 1717 6291 1723
rect 5965 1697 5987 1703
rect 2157 1677 2168 1683
rect 2925 1677 2952 1683
rect 3452 1683 3460 1688
rect 3432 1677 3460 1683
rect 3544 1676 3546 1684
rect 5960 1677 6019 1683
rect 2861 1637 2872 1643
rect 2941 1577 2968 1583
rect 221 1537 232 1543
rect 392 1537 403 1543
rect 2056 1536 2058 1544
rect 2968 1537 3011 1543
rect 253 1517 291 1523
rect 301 1503 307 1523
rect 301 1497 339 1503
rect 413 1503 419 1523
rect 413 1497 451 1503
rect 824 1497 856 1503
rect 909 1503 915 1523
rect 877 1497 915 1503
rect 1005 1503 1011 1523
rect 1005 1497 1043 1503
rect 1064 1497 1091 1503
rect 669 1477 680 1483
rect 840 1477 851 1483
rect 1085 1477 1091 1497
rect 1149 1503 1155 1523
rect 1117 1497 1155 1503
rect 1501 1497 1539 1503
rect 1645 1503 1651 1523
rect 1900 1517 1955 1523
rect 1900 1512 1908 1517
rect 1645 1497 1683 1503
rect 2333 1503 2339 1523
rect 2301 1497 2339 1503
rect 2376 1497 2403 1503
rect 2829 1497 2856 1503
rect 3021 1503 3027 1523
rect 3021 1497 3059 1503
rect 3069 1497 3112 1503
rect 3165 1503 3171 1523
rect 3261 1517 3299 1523
rect 4413 1517 4451 1523
rect 5405 1517 5443 1523
rect 3133 1497 3171 1503
rect 3224 1497 3235 1503
rect 3245 1497 3272 1503
rect 4541 1497 4579 1503
rect 4696 1497 4707 1503
rect 4877 1497 4904 1503
rect 5016 1497 5043 1503
rect 5149 1497 5160 1503
rect 5277 1497 5315 1503
rect 5644 1503 5652 1504
rect 5533 1497 5571 1503
rect 5644 1497 5683 1503
rect 5789 1497 5800 1503
rect 5885 1497 5955 1503
rect 6061 1497 6099 1503
rect 6120 1497 6131 1503
rect 6173 1497 6184 1503
rect 6444 1503 6452 1508
rect 6444 1497 6483 1503
rect 1229 1477 1256 1483
rect 1400 1477 1411 1483
rect 2648 1477 2659 1483
rect 3384 1477 3395 1483
rect 3485 1477 3523 1483
rect 3624 1477 3635 1483
rect 4333 1477 4344 1483
rect 4808 1477 4820 1483
rect 5016 1477 5059 1483
rect 5357 1477 5368 1483
rect 6136 1477 6147 1483
rect 6652 1463 6660 1472
rect 6632 1457 6660 1463
rect 4381 1437 4392 1443
rect 4989 1437 5000 1443
rect 1816 1377 1843 1383
rect 6781 1377 6792 1383
rect 4968 1357 4995 1363
rect 152 1337 163 1343
rect 2216 1337 2227 1343
rect 4412 1337 4436 1343
rect 5400 1337 5427 1343
rect 6237 1337 6275 1343
rect 93 1317 131 1323
rect 141 1317 152 1323
rect 493 1317 520 1323
rect 1021 1317 1059 1323
rect 1021 1297 1027 1317
rect 1165 1317 1192 1323
rect 1725 1317 1736 1323
rect 1928 1317 1955 1323
rect 2093 1317 2104 1323
rect 2616 1317 2643 1323
rect 2749 1317 2787 1323
rect 2797 1317 2808 1323
rect 1421 1297 1432 1303
rect 2781 1297 2787 1317
rect 2861 1317 2931 1323
rect 3101 1317 3139 1323
rect 3101 1297 3107 1317
rect 3421 1317 3432 1323
rect 3421 1297 3427 1317
rect 3496 1317 3507 1323
rect 3613 1317 3651 1323
rect 3645 1297 3651 1317
rect 3704 1317 3715 1323
rect 3773 1317 3796 1323
rect 3788 1314 3796 1317
rect 3992 1317 4035 1323
rect 4120 1317 4131 1323
rect 4157 1317 4195 1323
rect 4157 1297 4163 1317
rect 4328 1317 4355 1323
rect 4829 1317 4840 1323
rect 5069 1317 5107 1323
rect 5069 1297 5075 1317
rect 5160 1317 5171 1323
rect 5197 1317 5235 1323
rect 5176 1296 5180 1304
rect 5197 1297 5203 1317
rect 5645 1317 5683 1323
rect 5645 1297 5651 1317
rect 5800 1317 5827 1323
rect 5917 1317 5987 1323
rect 5981 1297 5987 1317
rect 6333 1323 6339 1343
rect 6381 1337 6392 1343
rect 6317 1317 6339 1323
rect 6381 1317 6419 1323
rect 6381 1297 6387 1317
rect 6541 1317 6579 1323
rect 6573 1297 6579 1317
rect 342 1276 344 1284
rect 941 1277 952 1283
rect 1389 1277 1459 1283
rect 1880 1276 1882 1284
rect 3080 1277 3091 1283
rect 3832 1276 3834 1284
rect 4989 1277 5000 1283
rect 4941 1237 4968 1243
rect 29 1137 40 1143
rect 328 1097 355 1103
rect 413 1097 424 1103
rect 557 1097 568 1103
rect 669 1103 675 1123
rect 1228 1117 1251 1123
rect 1228 1112 1236 1117
rect 1517 1117 1528 1123
rect 669 1097 707 1103
rect 717 1097 728 1103
rect 877 1097 915 1103
rect 1277 1097 1304 1103
rect 1480 1097 1491 1103
rect 1576 1097 1603 1103
rect 152 1077 163 1083
rect 504 1077 531 1083
rect 584 1077 595 1083
rect 781 1077 851 1083
rect 920 1077 931 1083
rect 957 1077 968 1083
rect 1597 1083 1603 1097
rect 2013 1097 2024 1103
rect 2424 1097 2435 1103
rect 2557 1097 2568 1103
rect 2621 1097 2632 1103
rect 2685 1103 2691 1123
rect 2653 1097 2691 1103
rect 2813 1097 2840 1103
rect 2872 1097 2899 1103
rect 3304 1097 3331 1103
rect 3709 1103 3715 1123
rect 4348 1123 4356 1128
rect 4344 1117 4356 1123
rect 4968 1117 4979 1123
rect 3677 1097 3715 1103
rect 3880 1097 3923 1103
rect 4077 1097 4120 1103
rect 4189 1097 4227 1103
rect 4316 1103 4324 1108
rect 4285 1097 4324 1103
rect 4749 1097 4760 1103
rect 5005 1097 5043 1103
rect 5116 1103 5124 1108
rect 5116 1097 5155 1103
rect 5581 1103 5587 1123
rect 5992 1117 6003 1123
rect 5581 1097 5619 1103
rect 5896 1097 5907 1103
rect 6301 1097 6328 1103
rect 6604 1106 6612 1112
rect 6680 1097 6691 1103
rect 1597 1077 1619 1083
rect 2680 1077 2691 1083
rect 2733 1077 2771 1083
rect 3789 1077 3800 1083
rect 4104 1077 4115 1083
rect 4909 1077 4952 1083
rect 5304 1077 5315 1083
rect 5517 1077 5528 1083
rect 5672 1077 5683 1083
rect 6141 1077 6163 1083
rect 6349 1077 6387 1083
rect 4157 1057 4168 1063
rect 4524 1063 4532 1072
rect 4504 1057 4532 1063
rect 4909 977 4936 983
rect 2333 957 2344 963
rect 2696 957 2724 963
rect 2716 948 2724 957
rect 829 937 840 943
rect 856 937 872 943
rect 333 917 371 923
rect 477 917 504 923
rect 701 917 739 923
rect 701 897 707 917
rect 845 917 915 923
rect 941 923 947 943
rect 1912 937 1924 943
rect 3112 937 3123 943
rect 3576 937 3587 943
rect 4301 937 4312 943
rect 4429 937 4451 943
rect 4813 937 4835 943
rect 4936 937 4963 943
rect 5101 937 5139 943
rect 5192 937 5203 943
rect 5245 937 5283 943
rect 941 917 968 923
rect 1053 917 1064 923
rect 1096 917 1107 923
rect 1485 917 1523 923
rect 1005 897 1016 903
rect 1517 897 1523 917
rect 1629 917 1667 923
rect 2060 908 2068 914
rect 2301 917 2339 923
rect 2397 917 2435 923
rect 2508 917 2547 923
rect 2508 912 2516 917
rect 2861 917 2920 923
rect 2957 917 2995 923
rect 2989 897 2995 917
rect 3069 917 3107 923
rect 3213 917 3251 923
rect 3213 897 3219 917
rect 3416 917 3427 923
rect 3992 917 4003 923
rect 4040 917 4051 923
rect 4349 917 4387 923
rect 3453 897 3491 903
rect 4381 897 4387 917
rect 5176 917 5192 923
rect 5453 923 5459 943
rect 5768 937 5795 943
rect 5901 937 5928 943
rect 6365 937 6376 943
rect 6424 937 6435 943
rect 5437 917 5459 923
rect 5640 917 5667 923
rect 5677 917 5715 923
rect 5709 897 5715 917
rect 5752 917 5779 923
rect 5837 917 5848 923
rect 6024 917 6035 923
rect 6061 917 6099 923
rect 6173 917 6184 923
rect 6061 897 6067 917
rect 6285 917 6323 923
rect 6349 917 6360 923
rect 6317 897 6323 917
rect 6397 917 6424 923
rect 6488 917 6499 923
rect 6696 917 6723 923
rect 621 877 691 883
rect 2710 876 2712 884
rect 3894 876 3896 884
rect 1960 737 1987 743
rect 2344 737 2355 743
rect 3276 737 3288 743
rect 396 717 419 723
rect 396 712 404 717
rect 93 697 131 703
rect 509 703 515 723
rect 509 697 547 703
rect 557 697 568 703
rect 621 703 627 723
rect 1869 717 1907 723
rect 1917 717 1955 723
rect 621 697 659 703
rect 765 697 792 703
rect 1020 703 1028 708
rect 1020 697 1059 703
rect 1149 697 1160 703
rect 1613 697 1624 703
rect 1869 703 1875 717
rect 1837 697 1875 703
rect 2077 703 2083 723
rect 2024 697 2035 703
rect 2045 697 2083 703
rect 2413 703 2419 723
rect 2792 717 2803 723
rect 2413 697 2451 703
rect 2637 697 2675 703
rect 2941 703 2947 723
rect 3256 716 3260 724
rect 3805 717 3827 723
rect 4648 717 4659 723
rect 4952 717 4979 723
rect 5389 717 5400 723
rect 2909 697 2947 703
rect 3176 697 3187 703
rect 3240 697 3251 703
rect 3405 697 3416 703
rect 3501 697 3528 703
rect 3981 697 4008 703
rect 4536 697 4547 703
rect 4696 697 4723 703
rect 4936 697 4995 703
rect 5021 697 5043 703
rect 1133 677 1144 683
rect 1661 677 1672 683
rect 2152 677 2163 683
rect 2349 677 2371 683
rect 2989 677 3027 683
rect 3688 677 3699 683
rect 3853 677 3880 683
rect 3912 677 3924 683
rect 4092 677 4104 683
rect 4092 672 4100 677
rect 4205 677 4227 683
rect 4813 677 4851 683
rect 5021 677 5027 697
rect 5133 697 5144 703
rect 5517 703 5523 723
rect 5480 697 5491 703
rect 5517 697 5555 703
rect 5656 697 5667 703
rect 5821 697 5843 703
rect 5224 677 5235 683
rect 5837 677 5843 697
rect 6152 697 6179 703
rect 6408 697 6435 703
rect 6685 703 6691 723
rect 6685 697 6723 703
rect 5949 677 6019 683
rect 2168 656 2172 664
rect 3277 657 3299 663
rect 2893 577 2904 583
rect 5928 577 5939 583
rect 1900 557 1928 563
rect 1900 554 1908 557
rect 2093 557 2115 563
rect 2972 557 3000 563
rect 2972 548 2980 557
rect 3565 557 3587 563
rect 3597 557 3619 563
rect 6765 557 6808 563
rect 813 537 840 543
rect 1277 537 1288 543
rect 2221 537 2232 543
rect 125 517 163 523
rect 221 517 259 523
rect 253 497 259 517
rect 429 517 467 523
rect 504 517 531 523
rect 637 517 664 523
rect 748 517 771 523
rect 829 517 856 523
rect 748 514 756 517
rect 1032 517 1059 523
rect 1096 517 1123 523
rect 1341 517 1352 523
rect 1453 517 1491 523
rect 269 497 307 503
rect 1085 497 1096 503
rect 1453 497 1459 517
rect 1624 517 1651 523
rect 1789 517 1816 523
rect 2045 517 2083 523
rect 2237 517 2275 523
rect 2557 523 2563 543
rect 2541 517 2563 523
rect 3261 523 3267 543
rect 3565 537 3576 543
rect 3880 537 3923 543
rect 4029 537 4040 543
rect 4200 537 4211 543
rect 4280 537 4291 543
rect 5181 537 5192 543
rect 5704 537 5715 543
rect 5784 537 5795 543
rect 5832 537 5843 543
rect 6365 537 6403 543
rect 6440 537 6451 543
rect 6461 537 6499 543
rect 3245 517 3267 523
rect 3389 517 3416 523
rect 3800 517 3827 523
rect 4184 517 4195 523
rect 4893 517 4904 523
rect 5341 517 5352 523
rect 5565 517 5603 523
rect 5629 517 5656 523
rect 2132 496 2136 504
rect 3133 497 3144 503
rect 5597 497 5603 517
rect 6024 517 6051 523
rect 6157 517 6195 523
rect 5620 496 5624 504
rect 6189 497 6195 517
rect 6248 517 6275 523
rect 710 476 712 484
rect 893 477 963 483
rect 2008 477 2020 483
rect 1421 337 1491 343
rect 4198 336 4200 344
rect 4733 337 4744 343
rect 4876 337 4904 343
rect 6029 337 6052 343
rect 6044 332 6052 337
rect 6184 337 6195 343
rect 461 297 472 303
rect 600 297 627 303
rect 637 297 648 303
rect 728 297 739 303
rect 765 303 771 323
rect 765 297 803 303
rect 941 303 947 323
rect 909 297 947 303
rect 1021 297 1059 303
rect 1133 303 1139 323
rect 1128 297 1139 303
rect 1229 297 1267 303
rect 1405 303 1411 323
rect 1448 317 1459 323
rect 1352 297 1363 303
rect 1373 297 1411 303
rect 2045 297 2067 303
rect 829 277 856 283
rect 1272 277 1283 283
rect 1336 277 1347 283
rect 1884 277 1928 283
rect 2045 277 2051 297
rect 2381 297 2424 303
rect 2637 288 2643 303
rect 2973 303 2979 323
rect 3720 316 3724 324
rect 2941 297 2979 303
rect 3005 297 3016 303
rect 3453 297 3480 303
rect 4413 297 4440 303
rect 4605 303 4611 323
rect 4717 317 4739 323
rect 4573 297 4611 303
rect 4776 297 4787 303
rect 5112 297 5123 303
rect 5261 303 5267 323
rect 5229 297 5267 303
rect 5533 303 5539 323
rect 5556 316 5560 324
rect 5501 297 5539 303
rect 5565 297 5576 303
rect 5741 303 5747 323
rect 5741 297 5763 303
rect 2205 277 2216 283
rect 2648 277 2675 283
rect 3112 277 3128 283
rect 3197 283 3203 292
rect 3197 277 3219 283
rect 3325 277 3363 283
rect 3533 277 3571 283
rect 3768 277 3779 283
rect 3885 277 3939 283
rect 5336 277 5347 283
rect 5384 277 5427 283
rect 5757 277 5763 297
rect 5912 297 5939 303
rect 6280 297 6307 303
rect 6573 297 6611 303
rect 5832 277 5843 283
rect 6077 277 6104 283
rect 6125 277 6136 283
rect 6364 277 6387 283
rect 2141 257 2163 263
rect 2301 257 2323 263
rect 2525 257 2547 263
rect 3165 257 3187 263
rect 6381 257 6387 277
rect 6397 257 6419 263
rect 5960 177 5987 183
rect 152 157 163 163
rect 221 157 243 163
rect 2904 157 2931 163
rect 4397 157 4419 163
rect 6221 157 6243 163
rect 2156 148 2164 152
rect 1085 137 1096 143
rect 2188 143 2196 148
rect 2188 137 2211 143
rect 2605 137 2616 143
rect 2877 137 2947 143
rect 3901 137 3939 143
rect 93 117 131 123
rect 264 117 275 123
rect 1277 128 1283 132
rect 1101 117 1139 123
rect 1213 117 1251 123
rect 493 97 531 103
rect 1213 97 1219 117
rect 1789 117 1828 123
rect 1820 116 1828 117
rect 2077 117 2104 123
rect 2221 117 2260 123
rect 2252 112 2260 117
rect 2477 117 2515 123
rect 1373 97 1411 103
rect 2509 97 2515 117
rect 2568 117 2579 123
rect 3021 117 3032 123
rect 3144 117 3171 123
rect 3389 117 3400 123
rect 3933 123 3939 137
rect 4461 137 4472 143
rect 4904 137 4947 143
rect 3933 117 3955 123
rect 4445 117 4456 123
rect 4584 117 4595 123
rect 3341 97 3363 103
rect 3380 96 3384 104
rect 4045 97 4067 103
rect 4589 97 4595 117
rect 5640 117 5651 123
rect 5720 117 5747 123
rect 5501 97 5523 103
rect 461 77 488 83
rect 6088 77 6099 83
rect 1896 37 1923 43
<< m2contact >>
rect 797 4802 833 4818
rect 2861 4802 2897 4818
rect 4909 4802 4945 4818
rect 344 4772 360 4788
rect 520 4772 536 4788
rect 568 4772 584 4788
rect 792 4772 808 4788
rect 1080 4772 1096 4788
rect 1672 4772 1688 4788
rect 1912 4772 1928 4788
rect 2424 4772 2440 4788
rect 3080 4772 3096 4788
rect 5432 4772 5448 4788
rect 5608 4772 5624 4788
rect 6296 4772 6312 4788
rect 6472 4772 6488 4788
rect 6568 4772 6600 4788
rect 4024 4752 4040 4768
rect 8 4732 24 4748
rect 248 4732 264 4748
rect 424 4732 440 4748
rect 632 4732 648 4748
rect 920 4732 936 4748
rect 1112 4732 1128 4748
rect 1160 4732 1176 4748
rect 2232 4732 2248 4748
rect 2728 4732 2744 4748
rect 2776 4732 2792 4748
rect 3336 4732 3352 4748
rect 3624 4732 3640 4748
rect 4040 4732 4056 4748
rect 4360 4732 4376 4748
rect 4952 4732 4968 4748
rect 4984 4732 5000 4748
rect 6280 4732 6296 4748
rect 6680 4732 6696 4748
rect 1128 4712 1144 4728
rect 1192 4712 1208 4728
rect 2744 4712 2760 4728
rect 2808 4712 2824 4728
rect 3336 4712 3352 4728
rect 3608 4712 3624 4728
rect 3656 4712 3672 4728
rect 3992 4712 4008 4728
rect 4312 4712 4328 4728
rect 4408 4712 4424 4728
rect 4744 4712 4760 4728
rect 4888 4712 4904 4728
rect 40 4692 56 4708
rect 136 4692 152 4708
rect 248 4692 280 4708
rect 312 4692 328 4708
rect 424 4692 456 4708
rect 488 4692 504 4708
rect 536 4692 552 4708
rect 616 4692 648 4708
rect 56 4672 72 4688
rect 296 4672 312 4688
rect 472 4672 488 4688
rect 584 4672 600 4688
rect 776 4672 792 4688
rect 904 4692 936 4708
rect 984 4692 1000 4708
rect 1048 4692 1064 4708
rect 1144 4692 1160 4708
rect 1176 4692 1192 4708
rect 1256 4690 1272 4706
rect 1320 4692 1336 4708
rect 1464 4692 1480 4708
rect 1512 4692 1528 4708
rect 1592 4692 1608 4708
rect 1640 4692 1656 4708
rect 1832 4692 1848 4708
rect 1976 4692 1992 4708
rect 2168 4690 2184 4706
rect 2360 4690 2376 4706
rect 2456 4692 2472 4708
rect 2504 4692 2520 4708
rect 2568 4690 2584 4706
rect 2632 4692 2648 4708
rect 2760 4692 2776 4708
rect 2792 4692 2808 4708
rect 2904 4690 2920 4706
rect 2968 4692 2984 4708
rect 3048 4692 3064 4708
rect 3224 4690 3240 4706
rect 3288 4692 3320 4708
rect 3400 4692 3416 4708
rect 3544 4690 3560 4706
rect 3640 4692 3656 4708
rect 3720 4692 3736 4708
rect 3864 4690 3880 4706
rect 4024 4692 4040 4708
rect 4168 4692 4200 4708
rect 4328 4692 4360 4708
rect 4376 4692 4392 4708
rect 4584 4690 4600 4706
rect 4760 4692 4776 4708
rect 4792 4692 4808 4708
rect 4840 4692 4856 4708
rect 4936 4692 4952 4708
rect 4968 4692 4984 4708
rect 5064 4692 5080 4708
rect 5176 4692 5192 4708
rect 5304 4692 5320 4708
rect 5352 4692 5368 4708
rect 5464 4692 5480 4708
rect 5512 4692 5544 4708
rect 5576 4692 5592 4708
rect 5624 4692 5640 4708
rect 5736 4690 5752 4706
rect 5896 4692 5912 4708
rect 6008 4692 6024 4708
rect 6152 4690 6168 4706
rect 6328 4692 6344 4708
rect 6376 4692 6408 4708
rect 6440 4692 6456 4708
rect 6488 4692 6504 4708
rect 6536 4692 6552 4708
rect 6616 4692 6632 4708
rect 6664 4692 6696 4708
rect 1032 4672 1048 4688
rect 1096 4672 1112 4688
rect 1624 4672 1640 4688
rect 1704 4672 1720 4688
rect 1880 4672 1896 4688
rect 1992 4672 2008 4688
rect 2200 4672 2216 4688
rect 2392 4672 2408 4688
rect 2472 4672 2488 4688
rect 2712 4672 2728 4688
rect 3256 4672 3272 4688
rect 3576 4672 3592 4688
rect 3672 4672 3688 4688
rect 3896 4672 3912 4688
rect 3944 4672 3960 4688
rect 4280 4672 4296 4688
rect 4312 4672 4328 4688
rect 4440 4672 4456 4688
rect 4616 4672 4632 4688
rect 4696 4672 4712 4688
rect 4760 4672 4776 4688
rect 4808 4672 4824 4688
rect 4840 4672 4856 4688
rect 5048 4672 5064 4688
rect 5144 4672 5160 4688
rect 5208 4672 5224 4688
rect 5480 4672 5496 4688
rect 5560 4672 5576 4688
rect 5800 4672 5816 4688
rect 5928 4672 5944 4688
rect 6120 4672 6136 4688
rect 6216 4672 6232 4688
rect 6344 4672 6360 4688
rect 6424 4672 6440 4688
rect 6520 4672 6536 4688
rect 6632 4672 6648 4688
rect 104 4652 120 4668
rect 136 4652 152 4668
rect 168 4652 200 4668
rect 360 4652 376 4668
rect 696 4652 712 4668
rect 984 4652 1000 4668
rect 1256 4652 1272 4668
rect 3368 4652 3384 4668
rect 4648 4652 4664 4668
rect 4696 4652 4712 4668
rect 6744 4652 6760 4668
rect 728 4632 744 4648
rect 1384 4632 1416 4648
rect 1688 4632 1704 4648
rect 1720 4632 1736 4648
rect 2696 4632 2712 4648
rect 3032 4632 3048 4648
rect 3096 4632 3112 4648
rect 3416 4632 3432 4648
rect 3736 4632 3752 4648
rect 4248 4632 4264 4648
rect 4456 4632 4472 4648
rect 4664 4632 4696 4648
rect 4728 4632 4744 4648
rect 5240 4632 5256 4648
rect 6088 4632 6104 4648
rect 1837 4602 1873 4618
rect 3885 4602 3921 4618
rect 5933 4602 5969 4618
rect 488 4572 504 4588
rect 632 4572 648 4588
rect 936 4572 952 4588
rect 1192 4572 1208 4588
rect 1240 4572 1256 4588
rect 1384 4572 1400 4588
rect 1528 4572 1544 4588
rect 1592 4572 1608 4588
rect 1992 4572 2008 4588
rect 2216 4572 2232 4588
rect 2280 4572 2296 4588
rect 2936 4572 2952 4588
rect 3016 4572 3032 4588
rect 3304 4572 3320 4588
rect 3352 4572 3368 4588
rect 3512 4572 3528 4588
rect 3624 4572 3640 4588
rect 3688 4572 3704 4588
rect 3880 4572 3896 4588
rect 4024 4572 4040 4588
rect 4120 4572 4136 4588
rect 4296 4572 4312 4588
rect 4360 4572 4376 4588
rect 4584 4572 4600 4588
rect 4776 4572 4792 4588
rect 4888 4572 4904 4588
rect 5336 4572 5352 4588
rect 5384 4572 5400 4588
rect 6040 4572 6056 4588
rect 6392 4572 6408 4588
rect 6584 4572 6600 4588
rect 3112 4552 3128 4568
rect 3240 4552 3256 4568
rect 4456 4552 4472 4568
rect 5560 4552 5576 4568
rect 8 4532 24 4548
rect 56 4532 72 4548
rect 264 4532 280 4548
rect 456 4532 472 4548
rect 536 4532 552 4548
rect 584 4532 600 4548
rect 920 4532 936 4548
rect 1128 4532 1144 4548
rect 1224 4532 1240 4548
rect 1288 4532 1304 4548
rect 40 4512 56 4528
rect 232 4514 248 4530
rect 360 4512 376 4528
rect 424 4514 440 4530
rect 520 4512 536 4528
rect 568 4512 584 4528
rect 696 4512 712 4528
rect 744 4512 760 4528
rect 1000 4512 1016 4528
rect 1064 4514 1080 4530
rect 1144 4512 1160 4528
rect 1176 4492 1192 4508
rect 1272 4512 1288 4528
rect 1384 4532 1400 4548
rect 1416 4532 1432 4548
rect 1448 4532 1464 4548
rect 1576 4532 1592 4548
rect 1608 4532 1624 4548
rect 1688 4532 1720 4548
rect 1816 4532 1832 4548
rect 1848 4532 1864 4548
rect 1944 4532 1960 4548
rect 2024 4532 2040 4548
rect 2072 4532 2088 4548
rect 2136 4532 2152 4548
rect 2216 4532 2232 4548
rect 2248 4532 2264 4548
rect 2440 4532 2456 4548
rect 2472 4532 2488 4548
rect 2568 4532 2584 4548
rect 2664 4532 2712 4548
rect 2776 4532 2824 4548
rect 2920 4532 2936 4548
rect 2984 4532 3016 4548
rect 3096 4532 3112 4548
rect 3144 4532 3160 4548
rect 3208 4532 3224 4548
rect 3256 4532 3272 4548
rect 3304 4532 3320 4548
rect 3336 4532 3352 4548
rect 3432 4532 3448 4548
rect 3496 4532 3512 4548
rect 3544 4532 3576 4548
rect 3656 4532 3688 4548
rect 3704 4532 3720 4548
rect 3784 4532 3800 4548
rect 3864 4532 3880 4548
rect 3896 4532 3912 4548
rect 4008 4532 4024 4548
rect 4072 4532 4088 4548
rect 4104 4532 4120 4548
rect 4136 4532 4152 4548
rect 4216 4532 4232 4548
rect 4248 4532 4264 4548
rect 4280 4532 4296 4548
rect 4328 4532 4344 4548
rect 4392 4532 4408 4548
rect 4504 4532 4536 4548
rect 4632 4532 4648 4548
rect 4712 4532 4728 4548
rect 1320 4512 1336 4528
rect 1432 4512 1448 4528
rect 1512 4512 1528 4528
rect 1560 4512 1576 4528
rect 1688 4512 1704 4528
rect 1240 4492 1256 4508
rect 1352 4492 1368 4508
rect 1640 4492 1656 4508
rect 1720 4492 1736 4508
rect 1784 4512 1816 4528
rect 1752 4492 1768 4508
rect 1896 4492 1912 4508
rect 1976 4512 1992 4528
rect 2088 4512 2120 4528
rect 2152 4512 2168 4528
rect 2264 4512 2280 4528
rect 2392 4512 2408 4528
rect 2488 4512 2504 4528
rect 2120 4492 2136 4508
rect 2184 4492 2200 4508
rect 2520 4492 2536 4508
rect 2552 4512 2568 4528
rect 2584 4512 2600 4528
rect 2616 4512 2632 4528
rect 2648 4512 2664 4528
rect 2760 4512 2776 4528
rect 2616 4492 2632 4508
rect 2728 4492 2744 4508
rect 2904 4512 2920 4528
rect 2968 4512 2984 4528
rect 2872 4492 2888 4508
rect 2936 4492 2952 4508
rect 3080 4512 3096 4528
rect 3128 4512 3144 4528
rect 3160 4512 3176 4528
rect 3240 4512 3256 4528
rect 3320 4512 3336 4528
rect 3048 4492 3064 4508
rect 3416 4512 3432 4528
rect 3480 4512 3496 4528
rect 3576 4512 3592 4528
rect 3384 4492 3400 4508
rect 3448 4492 3464 4508
rect 3468 4492 3484 4508
rect 3512 4492 3528 4508
rect 3608 4492 3624 4508
rect 3736 4512 3768 4528
rect 3800 4512 3848 4528
rect 3992 4512 4008 4528
rect 4056 4512 4072 4528
rect 4088 4512 4104 4528
rect 4200 4512 4216 4528
rect 4264 4512 4280 4528
rect 4392 4512 4408 4528
rect 4488 4512 4504 4528
rect 4520 4512 4536 4528
rect 3768 4492 3784 4508
rect 3928 4492 3944 4508
rect 4024 4492 4040 4508
rect 4168 4492 4184 4508
rect 4232 4492 4248 4508
rect 4296 4492 4312 4508
rect 4376 4492 4392 4508
rect 4420 4492 4436 4508
rect 4456 4492 4472 4508
rect 4536 4492 4552 4508
rect 4568 4492 4584 4508
rect 4616 4512 4632 4528
rect 4664 4512 4680 4528
rect 4696 4512 4728 4528
rect 4872 4532 4888 4548
rect 4904 4532 4920 4548
rect 4968 4532 4984 4548
rect 5032 4532 5048 4548
rect 5064 4532 5080 4548
rect 5144 4532 5160 4548
rect 5192 4532 5224 4548
rect 5240 4532 5256 4548
rect 5272 4532 5288 4548
rect 5368 4532 5384 4548
rect 5432 4532 5464 4548
rect 5480 4532 5496 4548
rect 5544 4532 5560 4548
rect 5768 4532 5784 4548
rect 5880 4532 5896 4548
rect 5912 4532 5928 4548
rect 5944 4532 5960 4548
rect 5992 4532 6008 4548
rect 6072 4532 6088 4548
rect 6184 4532 6200 4548
rect 6216 4532 6232 4548
rect 4744 4512 4760 4528
rect 4808 4512 4824 4528
rect 4856 4512 4872 4528
rect 4968 4512 5016 4528
rect 5048 4512 5064 4528
rect 5112 4512 5160 4528
rect 5224 4512 5240 4528
rect 5288 4512 5304 4528
rect 4776 4492 4808 4508
rect 5016 4492 5032 4508
rect 5080 4492 5112 4508
rect 5160 4492 5176 4508
rect 5256 4492 5272 4508
rect 5320 4492 5336 4508
rect 5416 4512 5432 4528
rect 5464 4512 5480 4528
rect 5640 4512 5656 4528
rect 5704 4514 5720 4530
rect 5816 4512 5832 4528
rect 5864 4512 5880 4528
rect 5928 4512 5944 4528
rect 6008 4512 6024 4528
rect 6056 4512 6072 4528
rect 6088 4512 6104 4528
rect 6120 4512 6136 4528
rect 6168 4512 6184 4528
rect 6248 4514 6264 4530
rect 6376 4512 6392 4528
rect 6456 4512 6472 4528
rect 6504 4512 6520 4528
rect 6648 4512 6664 4528
rect 6680 4512 6696 4528
rect 5368 4492 5384 4508
rect 5768 4492 5784 4508
rect 5896 4492 5912 4508
rect 6040 4492 6056 4508
rect 6136 4492 6152 4508
rect 296 4472 312 4488
rect 616 4472 632 4488
rect 1480 4472 1496 4488
rect 1528 4472 1544 4488
rect 1992 4472 2008 4488
rect 2040 4472 2072 4488
rect 2312 4472 2328 4488
rect 2632 4472 2648 4488
rect 3704 4472 3720 4488
rect 4824 4472 4840 4488
rect 5832 4472 5848 4488
rect 6344 4472 6360 4488
rect 6616 4472 6632 4488
rect 4808 4452 4824 4468
rect 600 4432 616 4448
rect 872 4432 888 4448
rect 2280 4432 2296 4448
rect 3176 4432 3192 4448
rect 4680 4432 4696 4448
rect 5576 4432 5592 4448
rect 797 4402 833 4418
rect 2861 4402 2897 4418
rect 4909 4402 4945 4418
rect 1448 4372 1464 4388
rect 1736 4372 1752 4388
rect 1800 4372 1816 4388
rect 1912 4372 1928 4388
rect 1960 4372 1976 4388
rect 2136 4372 2152 4388
rect 2232 4372 2248 4388
rect 2568 4372 2584 4388
rect 2600 4372 2616 4388
rect 3768 4372 3784 4388
rect 3896 4372 3912 4388
rect 4152 4372 4168 4388
rect 4344 4372 4360 4388
rect 4856 4372 4872 4388
rect 5480 4372 5496 4388
rect 5528 4372 5544 4388
rect 5656 4372 5672 4388
rect 5992 4372 6008 4388
rect 6680 4372 6696 4388
rect 936 4352 952 4368
rect 3336 4352 3352 4368
rect 40 4332 56 4348
rect 504 4332 520 4348
rect 584 4332 600 4348
rect 1192 4332 1208 4348
rect 1752 4332 1768 4348
rect 2168 4332 2184 4348
rect 2520 4332 2536 4348
rect 2552 4332 2568 4348
rect 2792 4332 2808 4348
rect 3288 4332 3304 4348
rect 3320 4332 3336 4348
rect 3912 4332 3928 4348
rect 4616 4332 4632 4348
rect 6808 4332 6824 4348
rect 408 4312 424 4328
rect 452 4312 468 4328
rect 472 4312 488 4328
rect 708 4312 724 4328
rect 744 4312 760 4328
rect 840 4312 856 4328
rect 904 4312 920 4328
rect 996 4312 1012 4328
rect 1016 4312 1032 4328
rect 1048 4312 1064 4328
rect 1080 4312 1096 4328
rect 1144 4312 1160 4328
rect 1224 4312 1240 4328
rect 1480 4312 1496 4328
rect 1720 4312 1736 4328
rect 1992 4312 2008 4328
rect 2056 4312 2072 4328
rect 72 4292 88 4308
rect 168 4292 184 4308
rect 280 4292 296 4308
rect 440 4292 456 4308
rect 488 4292 504 4308
rect 520 4292 536 4308
rect 600 4292 616 4308
rect 632 4292 648 4308
rect 664 4292 696 4308
rect 744 4292 760 4308
rect 824 4292 840 4308
rect 856 4292 888 4308
rect 936 4292 952 4308
rect 968 4292 984 4308
rect 1048 4292 1064 4308
rect 1096 4292 1112 4308
rect 1160 4292 1176 4308
rect 1208 4292 1224 4308
rect 1288 4290 1304 4306
rect 1352 4292 1368 4308
rect 1448 4292 1464 4308
rect 1656 4290 1672 4306
rect 1752 4292 1768 4308
rect 1880 4292 1896 4308
rect 1960 4292 1976 4308
rect 2024 4292 2040 4308
rect 2136 4292 2152 4308
rect 2264 4312 2280 4328
rect 2440 4312 2456 4328
rect 2740 4312 2756 4328
rect 2760 4312 2776 4328
rect 2840 4312 2856 4328
rect 2920 4312 2936 4328
rect 2952 4312 2968 4328
rect 2984 4312 3000 4328
rect 3128 4312 3144 4328
rect 3164 4312 3180 4328
rect 3208 4312 3224 4328
rect 3816 4312 3848 4328
rect 3880 4312 3896 4328
rect 3944 4312 3976 4328
rect 2296 4292 2312 4308
rect 2376 4292 2408 4308
rect 2472 4292 2488 4308
rect 2536 4292 2552 4308
rect 2648 4292 2664 4308
rect 2728 4292 2744 4308
rect 2792 4292 2808 4308
rect 2888 4292 2904 4308
rect 2936 4292 2952 4308
rect 2984 4292 3000 4308
rect 3032 4292 3048 4308
rect 3064 4292 3080 4308
rect 3096 4292 3112 4308
rect 3176 4292 3192 4308
rect 3272 4292 3288 4308
rect 3320 4292 3336 4308
rect 3416 4290 3432 4306
rect 3480 4292 3496 4308
rect 3672 4292 3688 4308
rect 3768 4292 3784 4308
rect 3928 4292 3944 4308
rect 3976 4292 4008 4308
rect 4072 4312 4088 4328
rect 4312 4312 4328 4328
rect 88 4272 104 4288
rect 248 4272 264 4288
rect 376 4272 392 4288
rect 424 4272 440 4288
rect 552 4272 568 4288
rect 616 4272 632 4288
rect 648 4272 664 4288
rect 680 4272 696 4288
rect 792 4272 808 4288
rect 888 4272 904 4288
rect 952 4272 984 4288
rect 1032 4272 1048 4288
rect 1096 4272 1112 4288
rect 1144 4272 1160 4288
rect 1256 4272 1272 4288
rect 1432 4272 1448 4288
rect 1496 4272 1512 4288
rect 1944 4272 1960 4288
rect 2008 4272 2024 4288
rect 2104 4272 2136 4288
rect 2200 4272 2216 4288
rect 2232 4272 2248 4288
rect 2312 4272 2328 4288
rect 2408 4272 2424 4288
rect 2456 4272 2488 4288
rect 2712 4272 2728 4288
rect 2776 4272 2792 4288
rect 2872 4272 2888 4288
rect 2920 4272 2952 4288
rect 3016 4272 3032 4288
rect 3048 4272 3064 4288
rect 3080 4272 3096 4288
rect 3128 4272 3144 4288
rect 3192 4272 3208 4288
rect 3240 4272 3256 4288
rect 3352 4272 3368 4288
rect 3720 4272 3736 4288
rect 3752 4272 3768 4288
rect 3816 4272 3832 4288
rect 4008 4272 4040 4288
rect 4120 4272 4136 4288
rect 4184 4292 4200 4308
rect 4280 4292 4296 4308
rect 4392 4312 4408 4328
rect 4424 4312 4440 4328
rect 4488 4312 4504 4328
rect 4584 4312 4600 4328
rect 4632 4312 4648 4328
rect 4888 4312 4904 4328
rect 4952 4312 4984 4328
rect 5032 4312 5048 4328
rect 5096 4312 5112 4328
rect 5352 4312 5368 4328
rect 4392 4292 4408 4308
rect 4456 4292 4472 4308
rect 4536 4292 4552 4308
rect 4568 4292 4584 4308
rect 4600 4292 4616 4308
rect 4696 4290 4712 4306
rect 4840 4292 4856 4308
rect 4984 4292 5016 4308
rect 5064 4292 5096 4308
rect 4232 4272 4248 4288
rect 4264 4272 4280 4288
rect 4360 4272 4392 4288
rect 4440 4272 4456 4288
rect 4520 4272 4536 4288
rect 4552 4272 4568 4288
rect 4664 4272 4680 4288
rect 4840 4272 4856 4288
rect 4936 4272 4952 4288
rect 5160 4290 5176 4306
rect 5320 4292 5336 4308
rect 5700 4312 5716 4328
rect 5720 4312 5736 4328
rect 5784 4312 5800 4328
rect 5880 4312 5896 4328
rect 6024 4312 6040 4328
rect 5400 4292 5448 4308
rect 5496 4292 5512 4308
rect 5528 4292 5544 4308
rect 5688 4292 5704 4308
rect 5752 4292 5784 4308
rect 5800 4292 5816 4308
rect 5864 4292 5880 4308
rect 5912 4292 5928 4308
rect 5992 4292 6008 4308
rect 6232 4292 6248 4308
rect 6408 4292 6424 4308
rect 5304 4272 5320 4288
rect 5384 4272 5400 4288
rect 6552 4290 6568 4306
rect 6616 4292 6632 4308
rect 6696 4292 6712 4308
rect 6744 4292 6760 4308
rect 5448 4272 5464 4288
rect 5480 4272 5496 4288
rect 5512 4272 5528 4288
rect 5608 4272 5624 4288
rect 5672 4272 5688 4288
rect 5736 4272 5752 4288
rect 5800 4272 5816 4288
rect 5928 4272 5944 4288
rect 5976 4272 5992 4288
rect 6056 4272 6072 4288
rect 6104 4272 6120 4288
rect 6280 4272 6296 4288
rect 6424 4272 6440 4288
rect 6728 4272 6744 4288
rect 8 4252 40 4268
rect 136 4252 152 4268
rect 1192 4252 1208 4268
rect 1656 4252 1672 4268
rect 5160 4252 5176 4268
rect 5592 4252 5624 4268
rect 5816 4252 5832 4268
rect 360 4232 376 4248
rect 392 4232 408 4248
rect 1416 4232 1432 4248
rect 1512 4232 1544 4248
rect 2088 4232 2104 4248
rect 2344 4232 2360 4248
rect 2680 4232 2696 4248
rect 3544 4232 3576 4248
rect 4040 4232 4056 4248
rect 4824 4232 4840 4248
rect 5288 4232 5304 4248
rect 5576 4232 5592 4248
rect 6120 4232 6136 4248
rect 6312 4232 6328 4248
rect 1837 4202 1873 4218
rect 3885 4202 3921 4218
rect 5933 4202 5969 4218
rect 744 4172 760 4188
rect 1240 4172 1256 4188
rect 1288 4172 1304 4188
rect 1448 4172 1464 4188
rect 1752 4172 1768 4188
rect 1912 4172 1928 4188
rect 2280 4172 2296 4188
rect 2504 4172 2536 4188
rect 2712 4172 2728 4188
rect 3448 4172 3464 4188
rect 3928 4172 3944 4188
rect 4200 4172 4216 4188
rect 4504 4172 4520 4188
rect 4680 4172 4696 4188
rect 5144 4172 5160 4188
rect 5640 4172 5656 4188
rect 5704 4172 5720 4188
rect 5832 4172 5848 4188
rect 6232 4172 6248 4188
rect 6728 4172 6744 4188
rect 248 4152 264 4168
rect 1368 4152 1384 4168
rect 1576 4152 1592 4168
rect 3384 4152 3400 4168
rect 3416 4152 3432 4168
rect 3640 4152 3656 4168
rect 4536 4152 4552 4168
rect 456 4132 472 4148
rect 520 4132 536 4148
rect 552 4132 568 4148
rect 760 4132 776 4148
rect 824 4132 840 4148
rect 920 4132 968 4148
rect 984 4132 1000 4148
rect 1096 4132 1128 4148
rect 1144 4132 1160 4148
rect 1208 4132 1240 4148
rect 1272 4132 1288 4148
rect 1320 4132 1336 4148
rect 1384 4132 1400 4148
rect 1432 4132 1448 4148
rect 1496 4132 1512 4148
rect 1528 4132 1544 4148
rect 1560 4132 1576 4148
rect 1656 4132 1688 4148
rect 1720 4132 1752 4148
rect 1784 4132 1816 4148
rect 1864 4132 1880 4148
rect 1896 4132 1912 4148
rect 1992 4132 2008 4148
rect 2072 4132 2088 4148
rect 2136 4132 2152 4148
rect 2200 4132 2216 4148
rect 2328 4132 2344 4148
rect 2392 4132 2408 4148
rect 2440 4132 2472 4148
rect 2568 4132 2600 4148
rect 2696 4132 2712 4148
rect 2744 4132 2776 4148
rect 2824 4132 2840 4148
rect 2872 4132 2904 4148
rect 3032 4132 3048 4148
rect 3112 4132 3128 4148
rect 3208 4132 3224 4148
rect 3272 4132 3288 4148
rect 3608 4132 3624 4148
rect 3640 4132 3656 4148
rect 3720 4132 3736 4148
rect 3784 4132 3816 4148
rect 3864 4132 3880 4148
rect 3912 4132 3928 4148
rect 3944 4132 3976 4148
rect 4024 4132 4040 4148
rect 4088 4132 4104 4148
rect 4136 4132 4152 4148
rect 4296 4132 4312 4148
rect 4360 4132 4376 4148
rect 4424 4132 4440 4148
rect 4520 4132 4536 4148
rect 4584 4132 4600 4148
rect 5240 4152 5256 4168
rect 5512 4152 5528 4168
rect 5800 4152 5832 4168
rect 6200 4152 6216 4168
rect 4792 4132 4808 4148
rect 4856 4132 4888 4148
rect 5016 4132 5032 4148
rect 5048 4132 5064 4148
rect 5096 4132 5112 4148
rect 5128 4132 5144 4148
rect 5176 4132 5192 4148
rect 5208 4132 5224 4148
rect 5256 4132 5272 4148
rect 5368 4132 5384 4148
rect 5400 4132 5416 4148
rect 5656 4132 5672 4148
rect 5720 4132 5736 4148
rect 5848 4132 5864 4148
rect 5880 4132 5896 4148
rect 5944 4132 5960 4148
rect 5992 4132 6008 4148
rect 6040 4132 6072 4148
rect 6120 4132 6136 4148
rect 6168 4132 6184 4148
rect 6280 4132 6312 4148
rect 6328 4132 6344 4148
rect 6616 4132 6632 4148
rect 136 4114 152 4130
rect 296 4112 328 4128
rect 408 4112 424 4128
rect 456 4112 472 4128
rect 392 4092 408 4108
rect 504 4092 520 4108
rect 664 4112 696 4128
rect 872 4112 888 4128
rect 904 4112 920 4128
rect 968 4112 984 4128
rect 1000 4112 1016 4128
rect 1032 4112 1048 4128
rect 1080 4112 1096 4128
rect 824 4092 840 4108
rect 888 4092 904 4108
rect 1012 4092 1028 4108
rect 1048 4092 1064 4108
rect 1192 4112 1208 4128
rect 1336 4112 1352 4128
rect 1416 4112 1432 4128
rect 1480 4112 1496 4128
rect 1544 4112 1560 4128
rect 1656 4112 1672 4128
rect 1704 4112 1736 4128
rect 1800 4112 1832 4128
rect 1160 4092 1176 4108
rect 1256 4092 1272 4108
rect 1304 4092 1320 4108
rect 1384 4092 1400 4108
rect 1448 4092 1464 4108
rect 1512 4092 1528 4108
rect 1608 4092 1624 4108
rect 1828 4092 1844 4108
rect 1848 4092 1864 4108
rect 1976 4112 1992 4128
rect 2056 4112 2088 4128
rect 2168 4112 2184 4128
rect 2200 4112 2216 4128
rect 2232 4112 2248 4128
rect 2312 4112 2328 4128
rect 2376 4112 2392 4128
rect 2472 4112 2488 4128
rect 2552 4112 2568 4128
rect 2600 4112 2616 4128
rect 1944 4092 1960 4108
rect 2024 4092 2040 4108
rect 2120 4092 2136 4108
rect 2280 4092 2296 4108
rect 2312 4092 2328 4108
rect 2344 4092 2360 4108
rect 2364 4092 2380 4108
rect 2408 4092 2440 4108
rect 2520 4092 2536 4108
rect 2632 4092 2648 4108
rect 2680 4112 2696 4128
rect 2776 4112 2792 4128
rect 2856 4112 2872 4128
rect 2904 4112 2920 4128
rect 2952 4112 2968 4128
rect 2668 4092 2684 4108
rect 2808 4092 2824 4108
rect 2984 4092 3000 4108
rect 3080 4112 3096 4128
rect 3192 4112 3208 4128
rect 3256 4112 3272 4128
rect 3320 4112 3336 4128
rect 3368 4112 3384 4128
rect 3480 4112 3512 4128
rect 3560 4112 3576 4128
rect 3672 4112 3688 4128
rect 3800 4112 3832 4128
rect 3864 4112 3880 4128
rect 3896 4112 3912 4128
rect 4024 4112 4040 4128
rect 4072 4112 4088 4128
rect 4104 4112 4120 4128
rect 4168 4112 4184 4128
rect 4232 4112 4248 4128
rect 4312 4112 4328 4128
rect 4376 4112 4392 4128
rect 4424 4112 4456 4128
rect 3160 4092 3176 4108
rect 3224 4092 3240 4108
rect 3288 4092 3304 4108
rect 3308 4092 3324 4108
rect 3704 4092 3720 4108
rect 3848 4092 3864 4108
rect 3976 4092 3992 4108
rect 4040 4092 4056 4108
rect 4264 4092 4280 4108
rect 4344 4092 4360 4108
rect 4408 4092 4424 4108
rect 4472 4092 4488 4108
rect 4568 4112 4584 4128
rect 4600 4112 4616 4128
rect 4632 4112 4664 4128
rect 4840 4112 4856 4128
rect 4632 4092 4648 4108
rect 4712 4092 4728 4108
rect 4744 4092 4760 4108
rect 4792 4092 4824 4108
rect 4920 4092 4936 4108
rect 5000 4112 5016 4128
rect 5032 4112 5048 4128
rect 5096 4112 5128 4128
rect 5176 4112 5208 4128
rect 5256 4112 5288 4128
rect 5320 4112 5336 4128
rect 5384 4112 5400 4128
rect 5416 4112 5432 4128
rect 5544 4112 5576 4128
rect 5672 4112 5688 4128
rect 5736 4112 5752 4128
rect 5864 4112 5880 4128
rect 5896 4112 5912 4128
rect 5992 4112 6024 4128
rect 6072 4112 6088 4128
rect 6120 4112 6136 4128
rect 6152 4112 6168 4128
rect 6184 4112 6200 4128
rect 6264 4112 6280 4128
rect 6312 4112 6328 4128
rect 6440 4112 6456 4128
rect 6472 4112 6488 4128
rect 6600 4114 6616 4130
rect 6744 4112 6760 4128
rect 4988 4092 5004 4108
rect 5304 4092 5320 4108
rect 5428 4092 5444 4108
rect 5448 4092 5464 4108
rect 5704 4092 5720 4108
rect 6040 4092 6056 4108
rect 6072 4092 6088 4108
rect 6104 4092 6120 4108
rect 6232 4092 6248 4108
rect 6344 4092 6360 4108
rect 6536 4092 6552 4108
rect 424 4072 440 4088
rect 840 4072 872 4088
rect 1640 4072 1656 4088
rect 1704 4072 1720 4088
rect 2216 4072 2232 4088
rect 2248 4072 2264 4088
rect 2712 4072 2728 4088
rect 3064 4072 3080 4088
rect 4072 4072 4088 4088
rect 5080 4072 5096 4088
rect 5736 4072 5752 4088
rect 5800 4072 5816 4088
rect 408 4052 424 4068
rect 2600 4052 2616 4068
rect 3016 4052 3032 4068
rect 3256 4052 3272 4068
rect 4840 4052 4856 4068
rect 6216 4052 6232 4068
rect 8 4032 24 4048
rect 376 4032 392 4048
rect 1592 4032 1608 4048
rect 2264 4032 2280 4048
rect 3080 4032 3096 4048
rect 3384 4032 3400 4048
rect 3528 4032 3544 4048
rect 3624 4032 3640 4048
rect 3736 4032 3752 4048
rect 4312 4032 4328 4048
rect 4568 4032 4584 4048
rect 5336 4032 5352 4048
rect 5912 4032 5928 4048
rect 6776 4032 6792 4048
rect 797 4002 833 4018
rect 2861 4002 2897 4018
rect 4909 4002 4945 4018
rect 312 3972 328 3988
rect 584 3972 600 3988
rect 1272 3972 1288 3988
rect 1416 3972 1432 3988
rect 1608 3972 1624 3988
rect 2152 3972 2168 3988
rect 2520 3972 2536 3988
rect 2744 3972 2760 3988
rect 3256 3972 3272 3988
rect 3656 3972 3672 3988
rect 3848 3972 3864 3988
rect 5224 3972 5240 3988
rect 5912 3972 5928 3988
rect 5976 3972 5992 3988
rect 2536 3952 2552 3968
rect 8 3932 24 3948
rect 328 3932 344 3948
rect 648 3932 664 3948
rect 2952 3932 2968 3948
rect 3048 3932 3064 3948
rect 3208 3932 3224 3948
rect 4136 3932 4168 3948
rect 4936 3932 4952 3948
rect 5688 3932 5704 3948
rect 5720 3932 5736 3948
rect 6360 3932 6376 3948
rect 6808 3932 6824 3948
rect 296 3912 312 3928
rect 440 3912 456 3928
rect 552 3912 568 3928
rect 40 3892 56 3908
rect 168 3892 200 3908
rect 312 3892 328 3908
rect 360 3892 376 3908
rect 392 3892 408 3908
rect 424 3892 440 3908
rect 472 3892 488 3908
rect 520 3892 536 3908
rect 744 3912 760 3928
rect 808 3912 824 3928
rect 904 3912 920 3928
rect 680 3892 696 3908
rect 776 3892 808 3908
rect 840 3892 856 3908
rect 1016 3912 1032 3928
rect 984 3892 1000 3908
rect 1096 3892 1112 3908
rect 1132 3912 1148 3928
rect 1304 3912 1320 3928
rect 1656 3912 1672 3928
rect 1704 3912 1720 3928
rect 1144 3892 1160 3908
rect 1176 3892 1192 3908
rect 1240 3892 1256 3908
rect 1272 3892 1288 3908
rect 1384 3892 1400 3908
rect 1496 3892 1528 3908
rect 1544 3892 1560 3908
rect 1576 3892 1592 3908
rect 1640 3892 1656 3908
rect 1736 3892 1752 3908
rect 1816 3892 1832 3908
rect 1848 3892 1864 3908
rect 1896 3892 1912 3908
rect 1928 3912 1944 3928
rect 1944 3892 1976 3908
rect 2072 3912 2088 3928
rect 2776 3912 2792 3928
rect 2840 3912 2856 3928
rect 2104 3892 2120 3908
rect 2184 3892 2216 3908
rect 2264 3892 2280 3908
rect 2296 3892 2312 3908
rect 2392 3890 2408 3906
rect 2456 3892 2472 3908
rect 2600 3892 2616 3908
rect 2648 3892 2664 3908
rect 2744 3892 2760 3908
rect 2792 3892 2808 3908
rect 2936 3912 2952 3928
rect 2984 3912 3000 3928
rect 3080 3912 3096 3928
rect 3144 3912 3160 3928
rect 3164 3912 3180 3928
rect 2968 3892 2984 3908
rect 3000 3892 3016 3908
rect 3128 3892 3144 3908
rect 3176 3892 3192 3908
rect 3336 3892 3352 3908
rect 3512 3892 3528 3908
rect 3560 3892 3576 3908
rect 3688 3892 3704 3908
rect 3752 3912 3768 3928
rect 3816 3912 3832 3928
rect 3992 3912 4008 3928
rect 4056 3912 4072 3928
rect 3784 3892 3800 3908
rect 3848 3892 3864 3908
rect 3896 3892 3912 3908
rect 3944 3892 3960 3908
rect 4024 3892 4040 3908
rect 4088 3892 4104 3908
rect 4120 3892 4136 3908
rect 4152 3892 4168 3908
rect 4280 3912 4296 3928
rect 4392 3912 4408 3928
rect 4472 3912 4488 3928
rect 4504 3912 4520 3928
rect 4584 3912 4600 3928
rect 4744 3912 4760 3928
rect 4808 3912 4824 3928
rect 4840 3912 4856 3928
rect 5000 3912 5016 3928
rect 5080 3912 5096 3928
rect 5144 3912 5160 3928
rect 5304 3912 5320 3928
rect 4312 3892 4328 3908
rect 4360 3892 4392 3908
rect 4440 3892 4456 3908
rect 4520 3892 4536 3908
rect 4632 3892 4648 3908
rect 4696 3892 4712 3908
rect 4792 3892 4808 3908
rect 4872 3892 4888 3908
rect 4936 3892 4952 3908
rect 5016 3892 5032 3908
rect 5096 3892 5128 3908
rect 5192 3892 5208 3908
rect 5256 3892 5272 3908
rect 5400 3912 5416 3928
rect 5672 3912 5688 3928
rect 6552 3912 6568 3928
rect 6616 3912 6632 3928
rect 6636 3912 6652 3928
rect 5352 3892 5368 3908
rect 5432 3892 5464 3908
rect 5512 3892 5528 3908
rect 5608 3892 5624 3908
rect 5640 3892 5656 3908
rect 5752 3892 5784 3908
rect 5880 3892 5896 3908
rect 6024 3892 6040 3908
rect 6088 3892 6104 3908
rect 6152 3892 6168 3908
rect 6232 3892 6248 3908
rect 6280 3892 6296 3908
rect 6424 3892 6440 3908
rect 6488 3890 6504 3906
rect 6568 3892 6600 3908
rect 6648 3892 6680 3908
rect 6728 3892 6744 3908
rect 56 3872 72 3888
rect 264 3872 280 3888
rect 376 3872 392 3888
rect 408 3872 424 3888
rect 456 3872 472 3888
rect 488 3872 520 3888
rect 584 3872 600 3888
rect 616 3872 648 3888
rect 696 3872 728 3888
rect 760 3872 776 3888
rect 856 3872 872 3888
rect 952 3872 984 3888
rect 1048 3872 1064 3888
rect 1080 3872 1096 3888
rect 1160 3872 1176 3888
rect 1192 3872 1208 3888
rect 1224 3872 1240 3888
rect 1256 3872 1272 3888
rect 1528 3872 1544 3888
rect 1560 3872 1576 3888
rect 1688 3872 1704 3888
rect 1720 3872 1736 3888
rect 1752 3872 1768 3888
rect 1800 3872 1816 3888
rect 1864 3872 1880 3888
rect 1992 3872 2008 3888
rect 2024 3872 2040 3888
rect 2120 3872 2136 3888
rect 2216 3872 2232 3888
rect 2248 3872 2264 3888
rect 2280 3872 2296 3888
rect 2552 3872 2568 3888
rect 2728 3872 2744 3888
rect 2792 3872 2808 3888
rect 2920 3872 2936 3888
rect 3016 3872 3032 3888
rect 3048 3872 3064 3888
rect 3128 3872 3144 3888
rect 3192 3872 3208 3888
rect 3240 3872 3256 3888
rect 3416 3872 3432 3888
rect 3464 3872 3480 3888
rect 3544 3872 3560 3888
rect 3704 3872 3720 3888
rect 3800 3872 3816 3888
rect 3864 3872 3880 3888
rect 3912 3872 3944 3888
rect 3960 3872 3976 3888
rect 4040 3872 4056 3888
rect 4104 3872 4120 3888
rect 4216 3872 4248 3888
rect 4328 3872 4360 3888
rect 4424 3872 4440 3888
rect 4456 3872 4472 3888
rect 4504 3872 4520 3888
rect 4536 3872 4552 3888
rect 1336 3852 1352 3868
rect 1768 3852 1784 3868
rect 1992 3852 2008 3868
rect 2232 3852 2248 3868
rect 2904 3852 2920 3868
rect 3208 3852 3224 3868
rect 3528 3852 3544 3868
rect 3656 3852 3672 3868
rect 4248 3852 4264 3868
rect 4616 3872 4632 3888
rect 4648 3872 4664 3888
rect 4680 3872 4696 3888
rect 4760 3872 4776 3888
rect 4808 3872 4824 3888
rect 4856 3872 4872 3888
rect 4888 3872 4904 3888
rect 4952 3872 4968 3888
rect 5128 3872 5144 3888
rect 5176 3872 5192 3888
rect 5336 3872 5352 3888
rect 5384 3872 5400 3888
rect 5448 3872 5464 3888
rect 5512 3872 5528 3888
rect 5576 3872 5608 3888
rect 5624 3872 5640 3888
rect 5672 3872 5688 3888
rect 5848 3872 5864 3888
rect 6008 3872 6024 3888
rect 6104 3872 6120 3888
rect 6136 3872 6152 3888
rect 6600 3872 6616 3888
rect 6664 3872 6680 3888
rect 6712 3872 6728 3888
rect 5064 3852 5080 3868
rect 5528 3852 5544 3868
rect 5960 3852 5976 3868
rect 6040 3852 6056 3868
rect 6104 3852 6120 3868
rect 6392 3852 6408 3868
rect 6488 3852 6504 3868
rect 744 3832 760 3848
rect 936 3832 952 3848
rect 1064 3832 1080 3848
rect 1208 3832 1224 3848
rect 1464 3832 1480 3848
rect 1656 3832 1672 3848
rect 1784 3832 1800 3848
rect 2008 3832 2024 3848
rect 2056 3832 2072 3848
rect 2328 3832 2344 3848
rect 2520 3832 2536 3848
rect 3544 3832 3560 3848
rect 3720 3832 3736 3848
rect 4056 3832 4072 3848
rect 4552 3832 4568 3848
rect 4664 3832 4680 3848
rect 4728 3832 4744 3848
rect 4840 3832 4856 3848
rect 5048 3832 5064 3848
rect 5144 3832 5160 3848
rect 5480 3832 5496 3848
rect 6056 3832 6072 3848
rect 6120 3832 6136 3848
rect 6344 3832 6376 3848
rect 1837 3802 1873 3818
rect 3885 3802 3921 3818
rect 5933 3802 5969 3818
rect 184 3772 200 3788
rect 232 3772 248 3788
rect 328 3772 344 3788
rect 424 3772 440 3788
rect 568 3772 584 3788
rect 648 3772 664 3788
rect 888 3772 904 3788
rect 984 3772 1000 3788
rect 1064 3772 1080 3788
rect 2088 3772 2104 3788
rect 3032 3772 3048 3788
rect 3112 3772 3128 3788
rect 3240 3772 3256 3788
rect 3304 3772 3320 3788
rect 4152 3772 4168 3788
rect 4312 3772 4328 3788
rect 4520 3772 4536 3788
rect 4776 3772 4792 3788
rect 4808 3772 4824 3788
rect 4872 3772 4888 3788
rect 5528 3772 5544 3788
rect 5560 3772 5576 3788
rect 6216 3772 6232 3788
rect 6408 3772 6424 3788
rect 6568 3772 6584 3788
rect 1608 3752 1624 3768
rect 1720 3752 1736 3768
rect 1768 3752 1784 3768
rect 2424 3752 2472 3768
rect 2488 3752 2520 3768
rect 2552 3752 2568 3768
rect 2728 3752 2744 3768
rect 2888 3752 2904 3768
rect 3464 3752 3480 3768
rect 3816 3752 3832 3768
rect 5304 3752 5320 3768
rect 5368 3752 5384 3768
rect 6152 3752 6168 3768
rect 6504 3752 6536 3768
rect 6680 3752 6696 3768
rect 56 3732 72 3748
rect 200 3732 216 3748
rect 248 3732 264 3748
rect 312 3732 328 3748
rect 408 3732 424 3748
rect 472 3732 488 3748
rect 552 3732 568 3748
rect 1176 3732 1192 3748
rect 1448 3732 1480 3748
rect 1512 3732 1528 3748
rect 1608 3732 1624 3748
rect 1672 3732 1688 3748
rect 1736 3732 1752 3748
rect 1784 3732 1800 3748
rect 1880 3732 1896 3748
rect 1944 3732 1960 3748
rect 1992 3732 2008 3748
rect 2136 3732 2152 3748
rect 2232 3732 2248 3748
rect 2360 3732 2376 3748
rect 2424 3732 2440 3748
rect 2520 3732 2536 3748
rect 2568 3732 2584 3748
rect 2648 3732 2680 3748
rect 2696 3732 2712 3748
rect 2824 3732 2840 3748
rect 2904 3732 2920 3748
rect 3000 3732 3016 3748
rect 3464 3732 3496 3748
rect 3512 3732 3528 3748
rect 3576 3732 3592 3748
rect 3672 3732 3688 3748
rect 3848 3732 3864 3748
rect 3992 3732 4008 3748
rect 4024 3732 4040 3748
rect 4296 3732 4312 3748
rect 4616 3732 4648 3748
rect 4664 3732 4680 3748
rect 4728 3732 4744 3748
rect 4840 3732 4856 3748
rect 4872 3732 4888 3748
rect 4904 3732 4920 3748
rect 4984 3732 5000 3748
rect 5016 3732 5032 3748
rect 5080 3732 5096 3748
rect 5176 3732 5192 3748
rect 5256 3732 5272 3748
rect 5320 3732 5336 3748
rect 5416 3732 5448 3748
rect 5720 3732 5736 3748
rect 5848 3732 5864 3748
rect 6040 3732 6056 3748
rect 6136 3732 6152 3748
rect 6168 3732 6184 3748
rect 6248 3732 6264 3748
rect 6280 3732 6296 3748
rect 6312 3732 6328 3748
rect 6376 3732 6408 3748
rect 6424 3732 6440 3748
rect 6456 3732 6472 3748
rect 6584 3732 6600 3748
rect 6728 3732 6744 3748
rect 6808 3732 6824 3748
rect 72 3712 88 3728
rect 264 3712 296 3728
rect 232 3692 248 3708
rect 296 3692 312 3708
rect 392 3712 408 3728
rect 456 3712 472 3728
rect 520 3712 552 3728
rect 616 3712 632 3728
rect 776 3712 808 3728
rect 920 3712 936 3728
rect 1016 3712 1048 3728
rect 1144 3712 1160 3728
rect 1240 3712 1256 3728
rect 1384 3712 1400 3728
rect 1528 3712 1544 3728
rect 1576 3712 1592 3728
rect 1656 3712 1672 3728
rect 1800 3712 1832 3728
rect 1896 3712 1912 3728
rect 2008 3712 2024 3728
rect 2040 3712 2056 3728
rect 2072 3712 2088 3728
rect 2120 3712 2136 3728
rect 2200 3714 2216 3730
rect 2344 3712 2360 3728
rect 2408 3712 2424 3728
rect 2488 3712 2504 3728
rect 2584 3712 2600 3728
rect 2616 3712 2632 3728
rect 2648 3712 2664 3728
rect 2712 3712 2728 3728
rect 2760 3712 2776 3728
rect 2808 3712 2824 3728
rect 2840 3712 2856 3728
rect 360 3692 376 3708
rect 424 3692 440 3708
rect 488 3692 504 3708
rect 508 3692 524 3708
rect 904 3692 920 3708
rect 1496 3692 1512 3708
rect 1560 3692 1576 3708
rect 1624 3692 1640 3708
rect 1768 3692 1784 3708
rect 1832 3692 1848 3708
rect 1928 3692 1944 3708
rect 2024 3692 2040 3708
rect 2088 3692 2104 3708
rect 2984 3712 3000 3728
rect 3064 3712 3096 3728
rect 3144 3712 3160 3728
rect 3208 3712 3224 3728
rect 3272 3712 3288 3728
rect 3384 3712 3400 3728
rect 3480 3712 3496 3728
rect 3592 3712 3608 3728
rect 2952 3692 2968 3708
rect 3400 3692 3416 3708
rect 3624 3692 3640 3708
rect 3704 3712 3720 3728
rect 3864 3712 3880 3728
rect 3976 3712 3992 3728
rect 4040 3712 4056 3728
rect 4072 3712 4088 3728
rect 4120 3712 4136 3728
rect 4184 3712 4200 3728
rect 4248 3712 4264 3728
rect 4392 3712 4408 3728
rect 4440 3714 4456 3730
rect 4552 3712 4568 3728
rect 4584 3712 4616 3728
rect 4648 3712 4664 3728
rect 4056 3692 4072 3708
rect 4568 3692 4584 3708
rect 4728 3712 4744 3728
rect 4856 3712 4872 3728
rect 4920 3712 4936 3728
rect 5000 3712 5016 3728
rect 5032 3712 5048 3728
rect 5160 3712 5176 3728
rect 5288 3712 5304 3728
rect 5400 3712 5416 3728
rect 5448 3712 5480 3728
rect 5496 3712 5512 3728
rect 5640 3712 5656 3728
rect 5880 3714 5896 3730
rect 5976 3712 5992 3728
rect 6056 3712 6072 3728
rect 6088 3712 6104 3728
rect 6168 3712 6184 3728
rect 6232 3712 6248 3728
rect 6264 3712 6280 3728
rect 6296 3712 6312 3728
rect 6328 3712 6344 3728
rect 6376 3712 6392 3728
rect 6440 3712 6456 3728
rect 6472 3712 6488 3728
rect 6600 3712 6648 3728
rect 6680 3712 6696 3728
rect 6744 3712 6760 3728
rect 4696 3692 4712 3708
rect 4808 3692 4824 3708
rect 4968 3692 4984 3708
rect 5480 3692 5496 3708
rect 6216 3692 6232 3708
rect 6360 3692 6376 3708
rect 6520 3692 6536 3708
rect 936 3672 952 3688
rect 1960 3672 1976 3688
rect 2056 3672 2072 3688
rect 2328 3672 2344 3688
rect 3720 3672 3736 3688
rect 4024 3672 4040 3688
rect 4088 3672 4104 3688
rect 5064 3672 5080 3688
rect 920 3652 936 3668
rect 5208 3652 5224 3668
rect 648 3632 664 3648
rect 1112 3632 1128 3648
rect 1336 3632 1352 3648
rect 1528 3632 1544 3648
rect 1576 3632 1592 3648
rect 1688 3632 1704 3648
rect 2392 3632 2408 3648
rect 2536 3632 2552 3648
rect 2600 3632 2616 3648
rect 2664 3632 2680 3648
rect 2792 3632 2808 3648
rect 2920 3632 2936 3648
rect 3176 3632 3192 3648
rect 3352 3632 3368 3648
rect 3416 3632 3432 3648
rect 3736 3632 3768 3648
rect 4072 3632 4088 3648
rect 4216 3632 4232 3648
rect 5752 3632 5768 3648
rect 6008 3632 6024 3648
rect 797 3602 833 3618
rect 2861 3602 2897 3618
rect 4909 3602 4945 3618
rect 2312 3572 2328 3588
rect 2680 3572 2696 3588
rect 2744 3572 2760 3588
rect 3032 3572 3048 3588
rect 3096 3572 3112 3588
rect 4152 3572 4168 3588
rect 5608 3572 5624 3588
rect 5688 3572 5704 3588
rect 5880 3572 5896 3588
rect 6344 3572 6360 3588
rect 6392 3572 6408 3588
rect 184 3552 200 3568
rect 1112 3552 1128 3568
rect 3784 3552 3800 3568
rect 216 3532 232 3548
rect 264 3532 280 3548
rect 1016 3532 1032 3548
rect 2152 3532 2168 3548
rect 2280 3532 2296 3548
rect 2728 3532 2744 3548
rect 3016 3532 3032 3548
rect 3176 3532 3192 3548
rect 3208 3532 3224 3548
rect 3752 3532 3768 3548
rect 3800 3532 3816 3548
rect 3832 3532 3848 3548
rect 4872 3532 4888 3548
rect 5752 3532 5768 3548
rect 5848 3532 5864 3548
rect 232 3512 264 3528
rect 344 3512 360 3528
rect 504 3512 520 3528
rect 568 3512 584 3528
rect 104 3492 120 3508
rect 280 3492 296 3508
rect 360 3492 376 3508
rect 392 3492 408 3508
rect 424 3492 440 3508
rect 456 3492 488 3508
rect 552 3492 568 3508
rect 632 3492 648 3508
rect 680 3512 696 3528
rect 712 3492 728 3508
rect 824 3512 840 3528
rect 1000 3512 1016 3528
rect 1064 3512 1080 3528
rect 1560 3512 1576 3528
rect 2232 3512 2248 3528
rect 2360 3512 2376 3528
rect 2648 3512 2664 3528
rect 2760 3512 2776 3528
rect 2936 3512 2952 3528
rect 3048 3512 3064 3528
rect 3080 3512 3096 3528
rect 3144 3512 3160 3528
rect 856 3492 872 3508
rect 920 3492 936 3508
rect 984 3492 1000 3508
rect 1032 3492 1048 3508
rect 1176 3492 1208 3508
rect 1352 3492 1368 3508
rect 1464 3492 1496 3508
rect 1592 3492 1608 3508
rect 200 3472 216 3488
rect 312 3472 328 3488
rect 376 3472 392 3488
rect 408 3472 456 3488
rect 504 3472 520 3488
rect 552 3472 568 3488
rect 616 3472 648 3488
rect 728 3472 776 3488
rect 872 3472 888 3488
rect 936 3472 984 3488
rect 1096 3472 1112 3488
rect 1384 3472 1400 3488
rect 1640 3492 1656 3508
rect 1672 3492 1688 3508
rect 1752 3492 1768 3508
rect 1912 3492 1928 3508
rect 2008 3492 2024 3508
rect 2040 3492 2056 3508
rect 2104 3492 2120 3508
rect 2168 3492 2184 3508
rect 2280 3492 2296 3508
rect 2344 3492 2376 3508
rect 2472 3492 2488 3508
rect 2504 3492 2552 3508
rect 2568 3492 2600 3508
rect 2744 3492 2760 3508
rect 2824 3492 2840 3508
rect 2920 3492 2936 3508
rect 2952 3492 2968 3508
rect 3016 3492 3032 3508
rect 3064 3492 3080 3508
rect 3128 3492 3144 3508
rect 3160 3492 3176 3508
rect 3256 3512 3272 3528
rect 3400 3512 3416 3528
rect 3684 3512 3700 3528
rect 3704 3512 3720 3528
rect 3288 3492 3304 3508
rect 3320 3492 3336 3508
rect 3352 3492 3368 3508
rect 3432 3492 3448 3508
rect 3528 3492 3544 3508
rect 3576 3492 3592 3508
rect 3672 3492 3688 3508
rect 3784 3492 3800 3508
rect 3912 3512 3928 3528
rect 3944 3492 3960 3508
rect 4040 3492 4056 3508
rect 4216 3512 4232 3528
rect 4328 3512 4344 3528
rect 5096 3512 5112 3528
rect 4264 3492 4280 3508
rect 4296 3492 4312 3508
rect 4408 3492 4424 3508
rect 4584 3492 4600 3508
rect 4632 3492 4680 3508
rect 4728 3492 4744 3508
rect 4792 3492 4824 3508
rect 5032 3490 5048 3506
rect 5112 3492 5144 3508
rect 5176 3492 5192 3508
rect 5224 3512 5240 3528
rect 5720 3512 5736 3528
rect 5816 3512 5832 3528
rect 5864 3512 5880 3528
rect 6120 3512 6136 3528
rect 6212 3512 6228 3528
rect 5320 3492 5352 3508
rect 5464 3492 5496 3508
rect 5640 3492 5656 3508
rect 5784 3492 5800 3508
rect 5816 3492 5832 3508
rect 5880 3492 5896 3508
rect 5928 3492 5944 3508
rect 5992 3492 6008 3508
rect 6024 3492 6056 3508
rect 6120 3492 6136 3508
rect 6152 3492 6168 3508
rect 6200 3492 6216 3508
rect 6248 3512 6264 3528
rect 6424 3512 6440 3528
rect 6632 3512 6648 3528
rect 6712 3512 6728 3528
rect 6296 3492 6328 3508
rect 6376 3492 6392 3508
rect 6504 3492 6520 3508
rect 1624 3472 1640 3488
rect 1656 3472 1672 3488
rect 1720 3472 1736 3488
rect 1768 3472 1784 3488
rect 1976 3472 1992 3488
rect 2008 3472 2024 3488
rect 2200 3472 2216 3488
rect 2408 3472 2424 3488
rect 2456 3472 2472 3488
rect 2488 3472 2504 3488
rect 2552 3472 2568 3488
rect 2616 3472 2632 3488
rect 2696 3472 2712 3488
rect 2968 3472 2984 3488
rect 56 3452 72 3468
rect 568 3452 584 3468
rect 904 3452 920 3468
rect 1880 3452 1896 3468
rect 2248 3452 2264 3468
rect 2424 3452 2440 3468
rect 2600 3452 2616 3468
rect 3208 3472 3224 3488
rect 3304 3472 3336 3488
rect 3368 3472 3384 3488
rect 3448 3472 3464 3488
rect 3656 3472 3672 3488
rect 3720 3472 3736 3488
rect 3832 3472 3848 3488
rect 3960 3472 3976 3488
rect 3992 3472 4008 3488
rect 4168 3472 4184 3488
rect 4264 3472 4296 3488
rect 4312 3472 4328 3488
rect 4360 3472 4376 3488
rect 4536 3472 4552 3488
rect 4744 3472 4792 3488
rect 5064 3472 5080 3488
rect 5144 3472 5176 3488
rect 5192 3472 5208 3488
rect 5256 3472 5272 3488
rect 5752 3472 5784 3488
rect 5816 3472 5832 3488
rect 5960 3472 5976 3488
rect 6024 3472 6040 3488
rect 6056 3472 6072 3488
rect 6168 3472 6200 3488
rect 6296 3472 6312 3488
rect 6376 3472 6392 3488
rect 6456 3472 6472 3488
rect 6488 3472 6504 3488
rect 6664 3472 6680 3488
rect 6744 3476 6760 3492
rect 4184 3452 4200 3468
rect 4840 3452 4856 3468
rect 5848 3452 5864 3468
rect 6552 3452 6568 3468
rect 648 3432 664 3448
rect 888 3432 904 3448
rect 1544 3432 1576 3448
rect 1816 3432 1832 3448
rect 2648 3432 2664 3448
rect 2792 3432 2808 3448
rect 2888 3432 2904 3448
rect 3176 3432 3192 3448
rect 3464 3432 3480 3448
rect 4520 3432 4536 3448
rect 4600 3432 4616 3448
rect 4696 3432 4712 3448
rect 5368 3432 5384 3448
rect 5400 3432 5416 3448
rect 5608 3432 5624 3448
rect 6072 3432 6088 3448
rect 6632 3432 6648 3448
rect 6776 3432 6792 3448
rect 1837 3402 1873 3418
rect 3885 3402 3921 3418
rect 5933 3402 5969 3418
rect 248 3372 264 3388
rect 936 3372 952 3388
rect 968 3372 984 3388
rect 1000 3372 1016 3388
rect 1080 3372 1096 3388
rect 1208 3372 1224 3388
rect 1496 3372 1512 3388
rect 1704 3372 1720 3388
rect 1736 3372 1752 3388
rect 1944 3372 1960 3388
rect 2056 3372 2072 3388
rect 2088 3372 2104 3388
rect 2408 3372 2424 3388
rect 3080 3372 3096 3388
rect 3336 3372 3352 3388
rect 3832 3372 3848 3388
rect 4184 3372 4200 3388
rect 4920 3372 4936 3388
rect 5032 3372 5048 3388
rect 5176 3372 5192 3388
rect 5224 3372 5240 3388
rect 5288 3372 5304 3388
rect 5768 3372 5800 3388
rect 5864 3372 5880 3388
rect 6152 3372 6168 3388
rect 6392 3372 6408 3388
rect 6696 3372 6712 3388
rect 104 3352 120 3368
rect 152 3352 184 3368
rect 520 3352 536 3368
rect 1544 3352 1560 3368
rect 1800 3352 1816 3368
rect 1880 3352 1896 3368
rect 2200 3352 2216 3368
rect 2328 3352 2344 3368
rect 2520 3352 2536 3368
rect 3464 3352 3480 3368
rect 4808 3352 4824 3368
rect 5528 3352 5544 3368
rect 5704 3352 5720 3368
rect 5896 3352 5912 3368
rect 5992 3352 6008 3368
rect 6024 3352 6040 3368
rect 6104 3352 6120 3368
rect 6312 3352 6328 3368
rect 6376 3352 6392 3368
rect 6632 3352 6648 3368
rect 4696 3348 4712 3350
rect 88 3332 104 3348
rect 120 3332 136 3348
rect 232 3332 248 3348
rect 296 3332 312 3348
rect 328 3332 344 3348
rect 360 3332 376 3348
rect 392 3332 408 3348
rect 568 3332 600 3348
rect 648 3332 664 3348
rect 40 3312 56 3328
rect 72 3312 88 3328
rect 136 3312 152 3328
rect 232 3312 248 3328
rect 280 3312 296 3328
rect 312 3312 328 3328
rect 392 3312 424 3328
rect 488 3312 504 3328
rect 552 3312 568 3328
rect 600 3312 616 3328
rect 632 3312 648 3328
rect 664 3312 680 3328
rect 728 3332 744 3348
rect 792 3332 808 3348
rect 824 3332 840 3348
rect 888 3332 904 3348
rect 984 3332 1000 3348
rect 1064 3332 1080 3348
rect 1128 3332 1144 3348
rect 1448 3332 1464 3348
rect 1528 3332 1544 3348
rect 1640 3332 1656 3348
rect 1672 3332 1688 3348
rect 1720 3332 1736 3348
rect 1800 3332 1816 3348
rect 1960 3332 1976 3348
rect 2008 3332 2024 3348
rect 2120 3332 2152 3348
rect 2168 3332 2184 3348
rect 2296 3332 2312 3348
rect 2376 3332 2392 3348
rect 2504 3332 2520 3348
rect 2712 3332 2728 3348
rect 2760 3332 2776 3348
rect 2856 3332 2872 3348
rect 2904 3332 2920 3348
rect 3032 3332 3048 3348
rect 3144 3332 3160 3348
rect 3224 3332 3240 3348
rect 3272 3332 3288 3348
rect 3304 3332 3320 3348
rect 3336 3332 3352 3348
rect 3416 3332 3432 3348
rect 3496 3332 3512 3348
rect 3560 3332 3576 3348
rect 3592 3332 3608 3348
rect 3624 3332 3640 3348
rect 3688 3332 3704 3348
rect 3784 3332 3800 3348
rect 3944 3332 3976 3348
rect 4280 3332 4296 3348
rect 4328 3332 4344 3348
rect 4392 3332 4440 3348
rect 4504 3332 4520 3348
rect 4568 3332 4584 3348
rect 4648 3332 4664 3348
rect 4696 3334 4744 3348
rect 4712 3332 4744 3334
rect 4824 3332 4840 3348
rect 4968 3332 4984 3348
rect 840 3312 856 3328
rect 904 3312 920 3328
rect 1032 3312 1048 3328
rect 1112 3312 1128 3328
rect 1176 3312 1192 3328
rect 1240 3312 1256 3328
rect 1336 3312 1352 3328
rect 1368 3312 1384 3328
rect 1592 3312 1608 3328
rect 1624 3312 1640 3328
rect 1656 3312 1672 3328
rect 1688 3312 1704 3328
rect 1864 3312 1880 3328
rect 1912 3312 1928 3328
rect 2040 3312 2056 3328
rect 2152 3312 2168 3328
rect 2184 3312 2200 3328
rect 2232 3312 2264 3328
rect 2344 3312 2360 3328
rect 2536 3312 2552 3328
rect 2680 3314 2696 3330
rect 2808 3312 2824 3328
rect 2920 3312 2936 3328
rect 3048 3312 3064 3328
rect 3112 3312 3144 3328
rect 3224 3312 3256 3328
rect 56 3292 72 3308
rect 184 3292 200 3308
rect 216 3292 232 3308
rect 248 3292 264 3308
rect 360 3292 376 3308
rect 440 3292 456 3308
rect 504 3292 536 3308
rect 792 3292 808 3308
rect 840 3292 856 3308
rect 872 3292 888 3308
rect 936 3292 968 3308
rect 1000 3292 1016 3308
rect 1480 3292 1496 3308
rect 1560 3292 1576 3308
rect 1624 3292 1640 3308
rect 1736 3292 1752 3308
rect 1896 3292 1912 3308
rect 2088 3292 2104 3308
rect 2184 3292 2200 3308
rect 2360 3292 2376 3308
rect 2408 3292 2440 3308
rect 3080 3292 3112 3308
rect 3288 3312 3304 3328
rect 3400 3312 3416 3328
rect 3432 3312 3448 3328
rect 3544 3312 3560 3328
rect 3608 3312 3624 3328
rect 3640 3312 3672 3328
rect 3704 3312 3720 3328
rect 3368 3292 3384 3308
rect 3528 3292 3544 3308
rect 3592 3292 3608 3308
rect 3672 3292 3688 3308
rect 3736 3292 3752 3308
rect 3816 3312 3832 3328
rect 3864 3312 3880 3328
rect 3928 3312 3944 3328
rect 3992 3312 4008 3328
rect 4104 3312 4136 3328
rect 4200 3312 4216 3328
rect 4232 3312 4248 3328
rect 4264 3312 4280 3328
rect 4296 3312 4312 3328
rect 4376 3312 4392 3328
rect 3896 3292 3912 3308
rect 4248 3292 4264 3308
rect 4344 3292 4360 3308
rect 4488 3312 4504 3328
rect 4552 3312 4568 3328
rect 4616 3312 4632 3328
rect 4664 3312 4680 3328
rect 4696 3312 4712 3328
rect 4744 3312 4760 3328
rect 4776 3312 4792 3328
rect 4840 3312 4856 3328
rect 4920 3312 4936 3328
rect 4952 3312 4968 3328
rect 5048 3332 5064 3348
rect 5096 3332 5112 3348
rect 5128 3332 5144 3348
rect 5208 3332 5224 3348
rect 5256 3332 5272 3348
rect 5560 3332 5576 3348
rect 5656 3332 5672 3348
rect 5720 3332 5736 3348
rect 5832 3332 5848 3348
rect 5896 3332 5912 3348
rect 5928 3332 5944 3348
rect 6024 3332 6040 3348
rect 6168 3332 6184 3348
rect 6200 3332 6216 3348
rect 6328 3332 6344 3348
rect 5000 3312 5016 3328
rect 5048 3312 5064 3328
rect 5080 3312 5096 3328
rect 5112 3312 5128 3328
rect 5144 3312 5160 3328
rect 5192 3312 5208 3328
rect 5256 3312 5272 3328
rect 5336 3312 5352 3328
rect 5384 3312 5400 3328
rect 5448 3312 5480 3328
rect 5544 3312 5560 3328
rect 5576 3312 5592 3328
rect 5624 3312 5640 3328
rect 5672 3312 5688 3328
rect 5736 3312 5752 3328
rect 5880 3312 5896 3328
rect 5944 3312 5960 3328
rect 5976 3312 5992 3328
rect 6056 3312 6072 3328
rect 6184 3312 6200 3328
rect 6216 3312 6232 3328
rect 6264 3312 6280 3328
rect 6344 3312 6360 3328
rect 6424 3312 6440 3328
rect 6504 3332 6536 3348
rect 6648 3332 6664 3348
rect 6712 3332 6728 3348
rect 6744 3332 6760 3348
rect 6488 3312 6504 3328
rect 6536 3312 6552 3328
rect 6584 3312 6600 3328
rect 6664 3312 6680 3328
rect 6712 3312 6728 3328
rect 4456 3292 4472 3308
rect 4520 3292 4536 3308
rect 4552 3292 4568 3308
rect 4776 3292 4792 3308
rect 4872 3292 4888 3308
rect 4920 3292 4936 3308
rect 5032 3292 5048 3308
rect 5176 3292 5192 3308
rect 5496 3292 5512 3308
rect 5640 3292 5656 3308
rect 5704 3292 5720 3308
rect 5784 3292 5800 3308
rect 5864 3292 5880 3308
rect 6088 3292 6104 3308
rect 6248 3292 6264 3308
rect 6344 3292 6360 3308
rect 6376 3292 6408 3308
rect 6568 3292 6584 3308
rect 6696 3292 6712 3308
rect 6760 3292 6776 3308
rect 24 3272 40 3288
rect 408 3272 424 3288
rect 472 3272 488 3288
rect 2056 3272 2072 3288
rect 2232 3272 2248 3288
rect 2328 3272 2344 3288
rect 3832 3272 3848 3288
rect 3992 3272 4008 3288
rect 4232 3272 4248 3288
rect 4584 3272 4616 3288
rect 5608 3272 5624 3288
rect 696 3252 712 3268
rect 40 3232 56 3248
rect 488 3232 504 3248
rect 616 3232 632 3248
rect 1432 3232 1448 3248
rect 1464 3232 1480 3248
rect 1992 3232 2008 3248
rect 2552 3232 2568 3248
rect 3016 3232 3032 3248
rect 3176 3232 3192 3248
rect 3512 3232 3528 3248
rect 4600 3232 4616 3248
rect 5352 3232 5368 3248
rect 5416 3232 5432 3248
rect 5592 3232 5608 3248
rect 6008 3232 6024 3248
rect 6312 3232 6328 3248
rect 6632 3232 6648 3248
rect 797 3202 833 3218
rect 2861 3202 2897 3218
rect 4909 3202 4945 3218
rect 184 3172 200 3188
rect 216 3172 232 3188
rect 328 3172 344 3188
rect 1496 3172 1512 3188
rect 1864 3172 1880 3188
rect 2200 3172 2216 3188
rect 2920 3172 2936 3188
rect 3688 3172 3704 3188
rect 3928 3172 3944 3188
rect 4376 3172 4392 3188
rect 4968 3172 4984 3188
rect 5288 3172 5304 3188
rect 5336 3172 5352 3188
rect 5720 3172 5736 3188
rect 5768 3172 5784 3188
rect 6024 3172 6040 3188
rect 6760 3172 6776 3188
rect 920 3152 936 3168
rect 4488 3152 4504 3168
rect 600 3132 616 3148
rect 808 3132 824 3148
rect 1896 3132 1912 3148
rect 2936 3132 2952 3148
rect 3512 3132 3528 3148
rect 5224 3132 5256 3148
rect 56 3090 72 3106
rect 120 3092 136 3108
rect 248 3112 264 3128
rect 280 3092 296 3108
rect 360 3112 376 3128
rect 888 3112 904 3128
rect 968 3112 984 3128
rect 1016 3112 1032 3128
rect 392 3092 408 3108
rect 488 3092 504 3108
rect 536 3092 552 3108
rect 696 3092 728 3108
rect 808 3092 824 3108
rect 904 3092 920 3108
rect 936 3092 952 3108
rect 1080 3112 1096 3128
rect 1144 3112 1160 3128
rect 1208 3112 1224 3128
rect 1272 3112 1288 3128
rect 1928 3112 1944 3128
rect 2104 3112 2136 3128
rect 2232 3112 2248 3128
rect 2760 3112 2776 3128
rect 1112 3092 1128 3108
rect 1176 3092 1192 3108
rect 1224 3092 1272 3108
rect 1304 3092 1320 3108
rect 1400 3092 1416 3108
rect 1560 3092 1576 3108
rect 1608 3092 1624 3108
rect 1672 3092 1688 3108
rect 1752 3092 1768 3108
rect 1832 3092 1848 3108
rect 1912 3092 1928 3108
rect 2072 3092 2088 3108
rect 2296 3092 2312 3108
rect 2424 3092 2440 3108
rect 2504 3092 2520 3108
rect 2536 3092 2552 3108
rect 2600 3092 2616 3108
rect 2632 3092 2648 3108
rect 2696 3092 2712 3108
rect 2728 3092 2744 3108
rect 2808 3092 2824 3108
rect 2840 3092 2856 3108
rect 2920 3092 2936 3108
rect 3000 3112 3016 3128
rect 3032 3092 3048 3108
rect 3064 3092 3080 3108
rect 3112 3112 3128 3128
rect 3224 3112 3240 3128
rect 3256 3112 3272 3128
rect 3288 3112 3304 3128
rect 3352 3112 3368 3128
rect 3416 3112 3432 3128
rect 4008 3112 4024 3128
rect 4056 3112 4072 3128
rect 4456 3112 4472 3128
rect 4520 3112 4536 3128
rect 4696 3112 4712 3128
rect 4728 3112 4744 3128
rect 5048 3112 5064 3128
rect 5256 3112 5272 3128
rect 5384 3112 5400 3128
rect 5512 3112 5528 3128
rect 5736 3112 5752 3128
rect 5800 3112 5816 3128
rect 5944 3112 5960 3128
rect 6008 3112 6024 3128
rect 6056 3112 6072 3128
rect 6280 3112 6296 3128
rect 6536 3112 6552 3128
rect 6696 3112 6712 3128
rect 6744 3112 6760 3128
rect 3176 3092 3208 3108
rect 3256 3092 3272 3108
rect 3320 3092 3336 3108
rect 3352 3092 3368 3108
rect 3384 3092 3400 3108
rect 3496 3092 3512 3108
rect 3592 3092 3608 3108
rect 3672 3092 3688 3108
rect 3720 3092 3752 3108
rect 3800 3092 3816 3108
rect 3896 3092 3912 3108
rect 3976 3092 4008 3108
rect 4024 3092 4040 3108
rect 4088 3092 4104 3108
rect 4248 3092 4280 3108
rect 4344 3092 4360 3108
rect 4440 3092 4456 3108
rect 4488 3092 4504 3108
rect 4520 3092 4568 3108
rect 4616 3092 4632 3108
rect 4648 3092 4664 3108
rect 4712 3092 4728 3108
rect 4760 3092 4776 3108
rect 4856 3092 4872 3108
rect 4952 3092 4968 3108
rect 4984 3092 5000 3108
rect 5032 3092 5048 3108
rect 5080 3092 5096 3108
rect 5160 3092 5192 3108
rect 5240 3092 5256 3108
rect 5336 3092 5352 3108
rect 5416 3092 5432 3108
rect 88 3072 104 3088
rect 200 3072 216 3088
rect 296 3072 328 3088
rect 408 3072 424 3088
rect 440 3072 456 3088
rect 632 3072 648 3088
rect 856 3072 872 3088
rect 888 3072 904 3088
rect 984 3072 1000 3088
rect 1032 3072 1048 3088
rect 1128 3072 1144 3088
rect 1192 3072 1208 3088
rect 1256 3072 1272 3088
rect 1320 3072 1336 3088
rect 1432 3072 1448 3088
rect 1640 3072 1656 3088
rect 1704 3072 1720 3088
rect 1736 3072 1752 3088
rect 2024 3072 2040 3088
rect 2088 3072 2104 3088
rect 2168 3072 2200 3088
rect 2376 3072 2392 3088
rect 2440 3072 2456 3088
rect 2488 3072 2504 3088
rect 2520 3072 2536 3088
rect 2552 3072 2568 3088
rect 2616 3072 2632 3088
rect 2680 3072 2696 3088
rect 2712 3072 2728 3088
rect 2792 3072 2808 3088
rect 2824 3072 2840 3088
rect 2952 3072 2968 3088
rect 3048 3072 3080 3088
rect 3160 3072 3192 3088
rect 3240 3072 3256 3088
rect 3304 3072 3320 3088
rect 3368 3072 3384 3088
rect 3448 3072 3464 3088
rect 3480 3072 3496 3088
rect 3528 3072 3544 3088
rect 3656 3072 3672 3088
rect 3784 3072 3800 3088
rect 3960 3072 3976 3088
rect 4168 3072 4184 3088
rect 4504 3072 4520 3088
rect 4568 3072 4584 3088
rect 4632 3072 4648 3088
rect 4664 3072 4680 3088
rect 4696 3072 4712 3088
rect 4728 3072 4744 3088
rect 4776 3072 4792 3088
rect 4872 3072 4888 3088
rect 5000 3072 5016 3088
rect 5096 3072 5112 3088
rect 5192 3072 5208 3088
rect 5352 3072 5368 3088
rect 5400 3072 5416 3088
rect 5480 3092 5496 3108
rect 5512 3092 5528 3108
rect 5544 3092 5560 3108
rect 5624 3092 5640 3108
rect 5656 3092 5672 3108
rect 5704 3092 5720 3108
rect 5816 3092 5832 3108
rect 5912 3092 5928 3108
rect 6024 3092 6040 3108
rect 6104 3092 6120 3108
rect 6168 3092 6184 3108
rect 6248 3092 6264 3108
rect 6360 3092 6376 3108
rect 6504 3092 6536 3108
rect 6600 3090 6616 3106
rect 5560 3072 5592 3088
rect 5608 3072 5624 3088
rect 5640 3072 5656 3088
rect 5704 3072 5720 3088
rect 5784 3072 5800 3088
rect 5848 3072 5864 3088
rect 5896 3072 5912 3088
rect 6088 3072 6104 3088
rect 6152 3072 6168 3088
rect 6232 3072 6248 3088
rect 6280 3072 6296 3088
rect 6312 3072 6328 3088
rect 6408 3072 6424 3088
rect 6488 3072 6504 3088
rect 6568 3072 6584 3088
rect 6776 3072 6792 3088
rect 1336 3052 1352 3068
rect 1400 3052 1432 3068
rect 1624 3052 1640 3068
rect 1800 3052 1816 3068
rect 2008 3052 2024 3068
rect 2328 3052 2344 3068
rect 2456 3052 2472 3068
rect 2568 3052 2600 3068
rect 2616 3052 2632 3068
rect 2648 3052 2664 3068
rect 3528 3052 3544 3068
rect 3608 3052 3624 3068
rect 4408 3052 4440 3068
rect 4904 3052 4920 3068
rect 4936 3052 4952 3068
rect 5272 3052 5288 3068
rect 5304 3052 5320 3068
rect 5544 3052 5560 3068
rect 5880 3052 5896 3068
rect 5944 3052 5960 3068
rect 1048 3032 1064 3048
rect 1144 3032 1160 3048
rect 1464 3032 1480 3048
rect 1624 3032 1640 3048
rect 1784 3032 1800 3048
rect 1896 3032 1912 3048
rect 2024 3032 2040 3048
rect 2120 3032 2136 3048
rect 2280 3032 2296 3048
rect 2408 3032 2424 3048
rect 3080 3032 3096 3048
rect 3224 3032 3240 3048
rect 3480 3032 3496 3048
rect 3624 3032 3640 3048
rect 3832 3032 3848 3048
rect 4120 3032 4136 3048
rect 4328 3032 4344 3048
rect 4584 3032 4600 3048
rect 4872 3032 4888 3048
rect 5128 3032 5144 3048
rect 5240 3032 5256 3048
rect 5384 3032 5400 3048
rect 5512 3032 5528 3048
rect 5592 3032 5608 3048
rect 6200 3032 6216 3048
rect 6472 3032 6488 3048
rect 6728 3032 6744 3048
rect 1837 3002 1873 3018
rect 3885 3002 3921 3018
rect 5933 3002 5969 3018
rect 264 2972 280 2988
rect 616 2972 632 2988
rect 968 2972 984 2988
rect 1496 2972 1512 2988
rect 1576 2972 1592 2988
rect 2152 2972 2168 2988
rect 2200 2972 2216 2988
rect 2344 2972 2360 2988
rect 2376 2972 2392 2988
rect 3048 2972 3064 2988
rect 3464 2972 3480 2988
rect 4168 2972 4184 2988
rect 4392 2972 4408 2988
rect 4616 2972 4632 2988
rect 4664 2972 4680 2988
rect 4808 2972 4824 2988
rect 4920 2972 4936 2988
rect 5144 2972 5160 2988
rect 5288 2972 5304 2988
rect 5816 2972 5832 2988
rect 6040 2972 6056 2988
rect 6392 2972 6408 2988
rect 6488 2972 6504 2988
rect 216 2952 232 2968
rect 1144 2952 1160 2968
rect 1192 2952 1208 2968
rect 1336 2952 1352 2968
rect 1720 2952 1736 2968
rect 1880 2952 1896 2968
rect 1992 2952 2008 2968
rect 2120 2952 2136 2968
rect 2264 2952 2280 2968
rect 2760 2952 2776 2968
rect 2856 2952 2872 2968
rect 3032 2952 3048 2968
rect 3064 2952 3080 2968
rect 3352 2952 3368 2968
rect 4088 2952 4136 2968
rect 4440 2952 4456 2968
rect 4472 2952 4488 2968
rect 5000 2952 5032 2968
rect 5608 2952 5624 2968
rect 5832 2952 5848 2968
rect 6008 2952 6024 2968
rect 216 2932 232 2948
rect 296 2932 312 2948
rect 328 2932 344 2948
rect 424 2932 440 2948
rect 456 2932 472 2948
rect 536 2932 552 2948
rect 568 2932 584 2948
rect 600 2932 616 2948
rect 648 2932 664 2948
rect 776 2932 792 2948
rect 1032 2932 1048 2948
rect 1064 2932 1080 2948
rect 1112 2932 1128 2948
rect 1160 2932 1176 2948
rect 1288 2932 1304 2948
rect 1320 2932 1336 2948
rect 1544 2932 1560 2948
rect 1592 2932 1608 2948
rect 1704 2932 1720 2948
rect 2120 2932 2136 2948
rect 2184 2932 2200 2948
rect 2216 2932 2232 2948
rect 2248 2932 2264 2948
rect 2312 2932 2328 2948
rect 2424 2932 2440 2948
rect 2520 2932 2552 2948
rect 2632 2932 2648 2948
rect 2792 2932 2808 2948
rect 2936 2932 2952 2948
rect 3000 2932 3016 2948
rect 3096 2932 3112 2948
rect 3128 2932 3160 2948
rect 3208 2932 3240 2948
rect 3288 2932 3304 2948
rect 3400 2932 3416 2948
rect 3432 2932 3448 2948
rect 3560 2932 3576 2948
rect 3816 2932 3832 2948
rect 4104 2932 4120 2948
rect 4376 2932 4392 2948
rect 4568 2932 4584 2948
rect 4600 2932 4616 2948
rect 4648 2932 4664 2948
rect 4712 2932 4744 2948
rect 4856 2932 4872 2948
rect 4952 2932 4968 2948
rect 5176 2932 5192 2948
rect 5368 2932 5384 2948
rect 5544 2932 5560 2948
rect 5624 2932 5656 2948
rect 5688 2932 5704 2948
rect 5720 2932 5736 2948
rect 5800 2932 5816 2948
rect 5848 2932 5864 2948
rect 5912 2932 5928 2948
rect 6008 2932 6024 2948
rect 6072 2932 6088 2948
rect 104 2912 136 2928
rect 280 2912 296 2928
rect 344 2912 360 2928
rect 392 2912 408 2928
rect 440 2912 456 2928
rect 264 2892 280 2908
rect 328 2892 344 2908
rect 408 2892 424 2908
rect 520 2912 552 2928
rect 584 2912 600 2928
rect 712 2912 728 2928
rect 856 2912 872 2928
rect 1000 2912 1032 2928
rect 1080 2912 1112 2928
rect 1160 2912 1176 2928
rect 1224 2912 1240 2928
rect 1320 2912 1336 2928
rect 1368 2912 1384 2928
rect 1448 2912 1464 2928
rect 1528 2912 1544 2928
rect 1560 2912 1576 2928
rect 1624 2912 1640 2928
rect 1784 2912 1800 2928
rect 1816 2912 1832 2928
rect 1928 2912 1944 2928
rect 1960 2912 1976 2928
rect 2040 2912 2056 2928
rect 2216 2912 2248 2928
rect 2312 2912 2328 2928
rect 2392 2912 2408 2928
rect 2440 2912 2456 2928
rect 488 2892 504 2908
rect 520 2892 536 2908
rect 552 2892 568 2908
rect 616 2892 632 2908
rect 680 2892 696 2908
rect 1064 2892 1080 2908
rect 1432 2892 1448 2908
rect 1672 2892 1688 2908
rect 1768 2892 1784 2908
rect 1800 2892 1816 2908
rect 1832 2892 1848 2908
rect 1912 2892 1928 2908
rect 1944 2892 1960 2908
rect 1976 2892 1992 2908
rect 2056 2892 2072 2908
rect 2136 2892 2152 2908
rect 2184 2892 2200 2908
rect 2344 2892 2360 2908
rect 2408 2892 2424 2908
rect 2472 2892 2488 2908
rect 2552 2912 2568 2928
rect 2584 2892 2600 2908
rect 2664 2912 2680 2928
rect 2760 2914 2776 2930
rect 2952 2912 2968 2928
rect 2984 2912 3000 2928
rect 3080 2912 3096 2928
rect 3144 2912 3160 2928
rect 3176 2912 3192 2928
rect 3208 2912 3224 2928
rect 3272 2912 3288 2928
rect 3384 2912 3400 2928
rect 3416 2912 3432 2928
rect 3448 2912 3464 2928
rect 3576 2912 3592 2928
rect 3784 2914 3800 2930
rect 3944 2912 3960 2928
rect 4008 2914 4024 2930
rect 4072 2912 4088 2928
rect 4264 2912 4280 2928
rect 4312 2914 4328 2930
rect 4424 2912 4440 2928
rect 4520 2912 4536 2928
rect 4552 2912 4568 2928
rect 4584 2912 4600 2928
rect 4648 2912 4664 2928
rect 4696 2912 4712 2928
rect 4744 2912 4776 2928
rect 4824 2912 4840 2928
rect 4872 2912 4888 2928
rect 4904 2912 4920 2928
rect 4984 2912 5000 2928
rect 5080 2912 5096 2928
rect 5112 2912 5128 2928
rect 5192 2912 5208 2928
rect 5352 2912 5368 2928
rect 5416 2914 5432 2930
rect 5496 2912 5512 2928
rect 2696 2892 2712 2908
rect 2968 2892 2984 2908
rect 3016 2892 3032 2908
rect 3208 2892 3224 2908
rect 3240 2892 3256 2908
rect 3272 2892 3288 2908
rect 4456 2892 4472 2908
rect 4520 2892 4536 2908
rect 4552 2892 4568 2908
rect 4664 2892 4680 2908
rect 4776 2892 4792 2908
rect 4808 2892 4824 2908
rect 4840 2892 4856 2908
rect 4920 2892 4936 2908
rect 5096 2892 5112 2908
rect 5224 2892 5240 2908
rect 5480 2892 5496 2908
rect 5512 2892 5528 2908
rect 5576 2892 5592 2908
rect 5640 2912 5656 2928
rect 5656 2892 5672 2908
rect 5768 2892 5784 2908
rect 5880 2892 5896 2908
rect 5928 2912 5944 2928
rect 6024 2912 6040 2928
rect 6136 2912 6152 2928
rect 6168 2932 6184 2948
rect 6248 2932 6264 2948
rect 6280 2932 6296 2948
rect 6360 2932 6392 2948
rect 6424 2932 6440 2948
rect 6536 2932 6568 2948
rect 6632 2932 6648 2948
rect 6664 2932 6680 2948
rect 6728 2932 6744 2948
rect 6808 2932 6824 2948
rect 6248 2912 6264 2928
rect 6104 2892 6120 2908
rect 6344 2912 6360 2928
rect 6440 2912 6456 2928
rect 6312 2892 6328 2908
rect 6408 2892 6424 2908
rect 6472 2892 6488 2908
rect 6520 2912 6536 2928
rect 6552 2912 6568 2928
rect 6616 2912 6632 2928
rect 6680 2912 6712 2928
rect 6744 2912 6760 2928
rect 6580 2892 6596 2908
rect 6600 2892 6616 2908
rect 184 2872 200 2888
rect 376 2872 392 2888
rect 1464 2872 1480 2888
rect 1496 2872 1512 2888
rect 1640 2872 1656 2888
rect 2024 2872 2040 2888
rect 2376 2872 2392 2888
rect 2680 2872 2696 2888
rect 5064 2872 5080 2888
rect 5272 2872 5288 2888
rect 360 2852 376 2868
rect 3368 2852 3384 2868
rect 5080 2852 5096 2868
rect 5496 2852 5512 2868
rect 200 2832 216 2848
rect 248 2832 264 2848
rect 936 2832 952 2848
rect 968 2832 984 2848
rect 1400 2832 1416 2848
rect 1448 2832 1464 2848
rect 1624 2832 1640 2848
rect 1688 2832 1704 2848
rect 1736 2832 1752 2848
rect 1784 2832 1800 2848
rect 1928 2832 1944 2848
rect 2040 2832 2056 2848
rect 2072 2832 2088 2848
rect 2328 2832 2344 2848
rect 2504 2832 2520 2848
rect 2904 2832 2920 2848
rect 3096 2832 3112 2848
rect 3304 2832 3320 2848
rect 3656 2832 3672 2848
rect 3880 2832 3896 2848
rect 4184 2832 4200 2848
rect 4504 2832 4520 2848
rect 4824 2832 4840 2848
rect 4872 2832 4888 2848
rect 5032 2832 5048 2848
rect 5256 2832 5272 2848
rect 5960 2832 5976 2848
rect 6216 2832 6232 2848
rect 6632 2832 6648 2848
rect 797 2802 833 2818
rect 2861 2802 2897 2818
rect 4909 2802 4945 2818
rect 1288 2772 1304 2788
rect 2296 2772 2312 2788
rect 2728 2772 2744 2788
rect 3320 2772 3336 2788
rect 3608 2772 3624 2788
rect 3784 2772 3800 2788
rect 4024 2772 4040 2788
rect 4440 2772 4456 2788
rect 4632 2772 4648 2788
rect 4856 2772 4872 2788
rect 5480 2772 5496 2788
rect 5672 2772 5688 2788
rect 5928 2772 5944 2788
rect 856 2752 872 2768
rect 1352 2752 1368 2768
rect 1528 2752 1544 2768
rect 1784 2752 1800 2768
rect 2920 2752 2936 2768
rect 5400 2752 5416 2768
rect 5768 2752 5784 2768
rect 8 2732 24 2748
rect 136 2732 152 2748
rect 680 2732 696 2748
rect 872 2732 888 2748
rect 1064 2732 1080 2748
rect 1176 2732 1192 2748
rect 1304 2732 1320 2748
rect 2104 2732 2120 2748
rect 3768 2732 3784 2748
rect 4008 2732 4024 2748
rect 4456 2732 4472 2748
rect 5400 2732 5416 2748
rect 6152 2732 6168 2748
rect 6296 2732 6312 2748
rect 104 2712 120 2728
rect 152 2712 168 2728
rect 440 2712 456 2728
rect 744 2712 760 2728
rect 40 2692 56 2708
rect 88 2692 104 2708
rect 120 2692 136 2708
rect 232 2692 248 2708
rect 280 2692 296 2708
rect 392 2692 408 2708
rect 472 2692 488 2708
rect 584 2692 600 2708
rect 616 2692 632 2708
rect 712 2692 728 2708
rect 984 2712 1000 2728
rect 856 2692 872 2708
rect 904 2692 920 2708
rect 936 2692 952 2708
rect 1032 2692 1048 2708
rect 1096 2712 1112 2728
rect 1128 2692 1144 2708
rect 1208 2712 1224 2728
rect 1272 2712 1288 2728
rect 1336 2712 1352 2728
rect 1384 2712 1400 2728
rect 1496 2712 1512 2728
rect 1704 2712 1720 2728
rect 1240 2692 1256 2708
rect 1288 2692 1304 2708
rect 1368 2692 1384 2708
rect 1416 2692 1432 2708
rect 56 2672 72 2688
rect 376 2672 392 2688
rect 408 2672 424 2688
rect 488 2672 504 2688
rect 696 2672 712 2688
rect 792 2672 808 2688
rect 920 2672 936 2688
rect 968 2672 984 2688
rect 1032 2672 1064 2688
rect 1144 2672 1176 2688
rect 1256 2672 1272 2688
rect 1368 2672 1384 2688
rect 1432 2672 1448 2688
rect 1464 2692 1480 2708
rect 1576 2692 1608 2708
rect 1656 2692 1672 2708
rect 1896 2712 1912 2728
rect 1816 2692 1848 2708
rect 1896 2692 1912 2708
rect 1932 2712 1948 2728
rect 2040 2712 2056 2728
rect 2136 2712 2152 2728
rect 2184 2712 2200 2728
rect 2232 2712 2264 2728
rect 2696 2712 2712 2728
rect 2856 2712 2872 2728
rect 2952 2712 2968 2728
rect 3032 2712 3048 2728
rect 3080 2712 3096 2728
rect 3416 2712 3432 2728
rect 3624 2712 3640 2728
rect 3644 2712 3660 2728
rect 3688 2712 3704 2728
rect 3800 2712 3816 2728
rect 4040 2712 4056 2728
rect 4104 2712 4120 2728
rect 4136 2712 4152 2728
rect 4200 2712 4216 2728
rect 4424 2712 4440 2728
rect 4488 2712 4504 2728
rect 4536 2712 4552 2728
rect 4900 2712 4916 2728
rect 4920 2712 4936 2728
rect 5016 2712 5032 2728
rect 1944 2692 1960 2708
rect 1976 2692 1992 2708
rect 2120 2692 2136 2708
rect 2360 2692 2376 2708
rect 2392 2692 2408 2708
rect 2504 2692 2520 2708
rect 2584 2692 2600 2708
rect 2696 2692 2712 2708
rect 2728 2692 2744 2708
rect 2760 2692 2776 2708
rect 1528 2672 1544 2688
rect 1560 2672 1576 2688
rect 1656 2672 1672 2688
rect 1752 2672 1768 2688
rect 1848 2672 1864 2688
rect 1960 2672 1976 2688
rect 2008 2672 2024 2688
rect 2072 2672 2088 2688
rect 2152 2672 2168 2688
rect 2200 2672 2216 2688
rect 2280 2672 2296 2688
rect 2328 2672 2344 2688
rect 2472 2672 2488 2688
rect 2568 2672 2584 2688
rect 2616 2672 2632 2688
rect 2680 2672 2696 2688
rect 2744 2672 2760 2688
rect 2808 2692 2824 2708
rect 2872 2692 2888 2708
rect 3096 2692 3128 2708
rect 3144 2692 3160 2708
rect 3208 2692 3224 2708
rect 3288 2692 3304 2708
rect 3352 2692 3368 2708
rect 3384 2692 3416 2708
rect 3480 2690 3496 2706
rect 3672 2692 3688 2708
rect 3736 2692 3752 2708
rect 3784 2692 3800 2708
rect 3816 2692 3832 2708
rect 3880 2692 3896 2708
rect 3928 2692 3944 2708
rect 4024 2692 4040 2708
rect 4072 2692 4088 2708
rect 4200 2692 4216 2708
rect 4232 2692 4264 2708
rect 4328 2692 4360 2708
rect 4408 2692 4424 2708
rect 4440 2692 4456 2708
rect 4520 2692 4536 2708
rect 4664 2692 4680 2708
rect 4760 2692 4776 2708
rect 4888 2692 4904 2708
rect 4968 2692 4984 2708
rect 5096 2692 5112 2708
rect 5160 2712 5176 2728
rect 5336 2712 5352 2728
rect 5416 2712 5432 2728
rect 5576 2712 5592 2728
rect 5596 2712 5612 2728
rect 5752 2712 5768 2728
rect 5832 2712 5848 2728
rect 6040 2712 6056 2728
rect 6104 2712 6136 2728
rect 6200 2712 6216 2728
rect 6504 2712 6520 2728
rect 6632 2712 6648 2728
rect 5208 2692 5224 2708
rect 5240 2692 5256 2708
rect 5288 2692 5304 2708
rect 5352 2692 5368 2708
rect 5384 2692 5400 2708
rect 5432 2692 5448 2708
rect 5528 2692 5544 2708
rect 5560 2692 5576 2708
rect 5608 2692 5624 2708
rect 5640 2692 5656 2708
rect 5720 2692 5736 2708
rect 5816 2692 5832 2708
rect 5848 2692 5880 2708
rect 5896 2692 5912 2708
rect 5992 2692 6008 2708
rect 6072 2692 6104 2708
rect 6152 2692 6168 2708
rect 6184 2692 6200 2708
rect 6248 2692 6264 2708
rect 2808 2672 2824 2688
rect 2904 2672 2920 2688
rect 2984 2672 3000 2688
rect 3064 2672 3080 2688
rect 3128 2672 3144 2688
rect 3160 2672 3176 2688
rect 3208 2672 3240 2688
rect 3272 2672 3288 2688
rect 3368 2672 3384 2688
rect 3736 2672 3752 2688
rect 3832 2672 3848 2688
rect 3864 2672 3880 2688
rect 3976 2672 3992 2688
rect 4056 2672 4072 2688
rect 4120 2672 4136 2688
rect 4168 2672 4184 2688
rect 4200 2672 4216 2688
rect 4248 2672 4264 2688
rect 4280 2672 4296 2688
rect 4312 2672 4328 2688
rect 4360 2672 4408 2688
rect 4536 2672 4552 2688
rect 4584 2676 4600 2692
rect 6392 2690 6408 2706
rect 6472 2692 6504 2708
rect 6536 2692 6552 2708
rect 4616 2672 4632 2688
rect 4744 2672 4760 2688
rect 4840 2672 4856 2688
rect 4872 2672 4888 2688
rect 4952 2672 4968 2688
rect 5048 2672 5064 2688
rect 5096 2672 5144 2688
rect 5192 2672 5208 2688
rect 5256 2672 5288 2688
rect 5432 2672 5448 2688
rect 5624 2672 5640 2688
rect 5704 2672 5720 2688
rect 5800 2672 5816 2688
rect 5880 2672 5896 2688
rect 5976 2672 5992 2688
rect 6056 2672 6072 2688
rect 6168 2672 6184 2688
rect 6200 2672 6216 2688
rect 6232 2672 6248 2688
rect 6376 2672 6392 2688
rect 6456 2672 6472 2688
rect 6520 2672 6536 2688
rect 6600 2692 6616 2708
rect 6696 2692 6712 2708
rect 6648 2672 6664 2688
rect 6712 2672 6728 2688
rect 2056 2652 2072 2668
rect 2360 2652 2376 2668
rect 2392 2652 2408 2668
rect 2456 2652 2488 2668
rect 2536 2652 2552 2668
rect 2600 2652 2616 2668
rect 2680 2652 2696 2668
rect 2760 2652 2776 2668
rect 2968 2652 2984 2668
rect 3480 2652 3496 2668
rect 5336 2652 5352 2668
rect 5480 2652 5528 2668
rect 6680 2652 6696 2668
rect 6728 2652 6760 2668
rect 344 2632 360 2648
rect 1624 2632 1640 2648
rect 1720 2632 1736 2648
rect 2104 2632 2120 2648
rect 2184 2632 2200 2648
rect 2232 2632 2264 2648
rect 2376 2632 2392 2648
rect 2888 2632 2904 2648
rect 3016 2632 3032 2648
rect 3048 2632 3064 2648
rect 3160 2632 3176 2648
rect 3256 2632 3272 2648
rect 3832 2632 3848 2648
rect 4312 2632 4328 2648
rect 5064 2632 5080 2648
rect 5320 2632 5336 2648
rect 5464 2632 5480 2648
rect 5928 2632 5944 2648
rect 6040 2632 6056 2648
rect 6264 2632 6280 2648
rect 1837 2602 1873 2618
rect 3885 2602 3921 2618
rect 5933 2602 5969 2618
rect 40 2572 56 2588
rect 88 2572 104 2588
rect 504 2572 520 2588
rect 712 2572 728 2588
rect 1880 2572 1896 2588
rect 2008 2572 2024 2588
rect 2168 2572 2184 2588
rect 2216 2572 2232 2588
rect 2280 2572 2296 2588
rect 2424 2572 2440 2588
rect 3544 2572 3560 2588
rect 3752 2572 3768 2588
rect 3800 2572 3816 2588
rect 3864 2572 3880 2588
rect 4056 2572 4072 2588
rect 4200 2572 4216 2588
rect 4376 2572 4392 2588
rect 4456 2572 4472 2588
rect 4728 2572 4744 2588
rect 4856 2572 4872 2588
rect 5192 2572 5208 2588
rect 5304 2572 5320 2588
rect 6232 2572 6248 2588
rect 6344 2572 6360 2588
rect 6424 2572 6440 2588
rect 6488 2572 6504 2588
rect 280 2552 296 2568
rect 2088 2552 2104 2568
rect 2264 2552 2280 2568
rect 2344 2552 2360 2568
rect 2376 2552 2392 2568
rect 2904 2552 2920 2568
rect 4648 2552 4680 2568
rect 5112 2552 5128 2568
rect 5208 2552 5224 2568
rect 5784 2552 5800 2568
rect 5864 2552 5880 2568
rect 5944 2552 5960 2568
rect 6760 2552 6776 2568
rect 8 2532 24 2548
rect 56 2532 72 2548
rect 152 2532 184 2548
rect 216 2532 232 2548
rect 440 2532 456 2548
rect 472 2532 504 2548
rect 536 2532 552 2548
rect 664 2532 680 2548
rect 728 2532 744 2548
rect 984 2532 1000 2548
rect 1128 2532 1144 2548
rect 1160 2532 1176 2548
rect 1192 2532 1208 2548
rect 1320 2532 1336 2548
rect 1496 2532 1512 2548
rect 1544 2532 1560 2548
rect 1592 2532 1608 2548
rect 1688 2532 1704 2548
rect 1720 2532 1736 2548
rect 1800 2532 1816 2548
rect 1864 2532 1880 2548
rect 1912 2532 1944 2548
rect 1976 2532 1992 2548
rect 2120 2532 2136 2548
rect 2200 2532 2216 2548
rect 2360 2532 2376 2548
rect 2392 2532 2408 2548
rect 2440 2532 2456 2548
rect 2552 2532 2568 2548
rect 2600 2532 2616 2548
rect 2632 2532 2648 2548
rect 2712 2532 2728 2548
rect 2776 2532 2792 2548
rect 2856 2532 2872 2548
rect 2904 2532 2920 2548
rect 2952 2532 2984 2548
rect 3048 2532 3064 2548
rect 3096 2532 3112 2548
rect 3160 2532 3176 2548
rect 3240 2532 3256 2548
rect 3336 2532 3352 2548
rect 3400 2532 3416 2548
rect 3448 2532 3464 2548
rect 3480 2532 3496 2548
rect 3512 2532 3544 2548
rect 3576 2532 3592 2548
rect 3608 2532 3624 2548
rect 3720 2532 3736 2548
rect 3768 2532 3784 2548
rect 3816 2532 3848 2548
rect 3912 2532 3928 2548
rect 4024 2532 4056 2548
rect 4136 2532 4152 2548
rect 40 2492 56 2508
rect 136 2512 152 2528
rect 200 2512 216 2528
rect 312 2512 344 2528
rect 456 2512 472 2528
rect 520 2512 536 2528
rect 104 2492 120 2508
rect 168 2492 184 2508
rect 424 2492 440 2508
rect 520 2492 536 2508
rect 568 2512 584 2528
rect 648 2512 664 2528
rect 680 2512 696 2528
rect 744 2512 760 2528
rect 712 2492 728 2508
rect 776 2492 792 2508
rect 840 2512 872 2528
rect 936 2512 952 2528
rect 1000 2512 1016 2528
rect 1112 2512 1128 2528
rect 1144 2512 1160 2528
rect 1272 2512 1288 2528
rect 1400 2512 1416 2528
rect 1512 2512 1528 2528
rect 952 2492 968 2508
rect 1176 2492 1192 2508
rect 1288 2492 1304 2508
rect 1560 2512 1576 2528
rect 1640 2512 1656 2528
rect 1672 2512 1688 2528
rect 1704 2512 1720 2528
rect 1784 2512 1800 2528
rect 1816 2512 1832 2528
rect 1560 2492 1576 2508
rect 1752 2492 1768 2508
rect 1960 2512 1976 2528
rect 2040 2512 2072 2528
rect 2136 2512 2152 2528
rect 2168 2512 2184 2528
rect 2200 2512 2216 2528
rect 2328 2512 2360 2528
rect 2504 2512 2520 2528
rect 2616 2512 2632 2528
rect 2680 2512 2696 2528
rect 2712 2512 2728 2528
rect 2760 2512 2776 2528
rect 2808 2512 2856 2528
rect 2952 2512 2968 2528
rect 2984 2512 3000 2528
rect 3016 2512 3032 2528
rect 3144 2512 3160 2528
rect 3208 2512 3224 2528
rect 2472 2492 2488 2508
rect 2584 2492 2600 2508
rect 2664 2492 2680 2508
rect 2728 2492 2744 2508
rect 2792 2492 2808 2508
rect 3016 2492 3032 2508
rect 3112 2492 3128 2508
rect 3224 2492 3240 2508
rect 3320 2512 3336 2528
rect 3368 2512 3400 2528
rect 3496 2512 3512 2528
rect 3528 2512 3544 2528
rect 3592 2512 3608 2528
rect 3624 2512 3656 2528
rect 3688 2512 3720 2528
rect 3896 2512 3912 2528
rect 3976 2512 3992 2528
rect 3288 2492 3304 2508
rect 3352 2492 3368 2508
rect 3416 2492 3432 2508
rect 3464 2492 3480 2508
rect 3656 2492 3672 2508
rect 3768 2492 3784 2508
rect 3960 2492 3976 2508
rect 4120 2512 4136 2528
rect 4216 2532 4232 2548
rect 4280 2532 4296 2548
rect 4344 2532 4360 2548
rect 4440 2532 4456 2548
rect 4488 2532 4520 2548
rect 4552 2532 4568 2548
rect 4168 2512 4184 2528
rect 4216 2512 4248 2528
rect 4296 2512 4312 2528
rect 4344 2512 4360 2528
rect 4408 2512 4424 2528
rect 4440 2512 4456 2528
rect 4520 2512 4536 2528
rect 4568 2512 4584 2528
rect 4680 2532 4696 2548
rect 4744 2532 4760 2548
rect 4808 2532 4824 2548
rect 4872 2532 4888 2548
rect 5016 2532 5032 2548
rect 5064 2532 5080 2548
rect 5224 2532 5256 2548
rect 5352 2532 5368 2548
rect 5448 2532 5464 2548
rect 5480 2532 5496 2548
rect 5544 2532 5560 2548
rect 5768 2532 5784 2548
rect 5800 2532 5816 2548
rect 5848 2532 5864 2548
rect 5976 2532 5992 2548
rect 6040 2532 6056 2548
rect 6200 2532 6232 2548
rect 6248 2532 6264 2548
rect 6280 2532 6296 2548
rect 6392 2532 6408 2548
rect 6456 2532 6472 2548
rect 6504 2532 6520 2548
rect 4696 2512 4712 2528
rect 4792 2512 4808 2528
rect 4824 2512 4840 2528
rect 4088 2492 4104 2508
rect 4200 2492 4216 2508
rect 4232 2492 4248 2508
rect 4264 2492 4280 2508
rect 4328 2492 4344 2508
rect 4376 2492 4408 2508
rect 4728 2492 4744 2508
rect 4872 2492 4888 2508
rect 4904 2492 4920 2508
rect 4968 2512 4984 2528
rect 5176 2512 5192 2528
rect 5336 2512 5352 2528
rect 5368 2512 5384 2528
rect 5416 2512 5432 2528
rect 5496 2512 5512 2528
rect 5528 2512 5544 2528
rect 5656 2512 5688 2528
rect 5752 2512 5768 2528
rect 5832 2512 5848 2528
rect 5912 2512 5928 2528
rect 5992 2512 6008 2528
rect 6056 2512 6072 2528
rect 6088 2512 6104 2528
rect 6168 2512 6184 2528
rect 6200 2512 6216 2528
rect 6264 2512 6280 2528
rect 6296 2512 6312 2528
rect 4984 2492 5000 2508
rect 5016 2492 5032 2508
rect 5272 2492 5288 2508
rect 5400 2492 5416 2508
rect 5800 2492 5816 2508
rect 6008 2492 6024 2508
rect 6072 2492 6088 2508
rect 6328 2492 6344 2508
rect 6392 2512 6408 2528
rect 6568 2512 6584 2528
rect 6664 2532 6680 2548
rect 6712 2532 6728 2548
rect 6632 2512 6648 2528
rect 6440 2492 6456 2508
rect 6488 2492 6504 2508
rect 6536 2492 6552 2508
rect 6712 2512 6728 2528
rect 6680 2492 6696 2508
rect 824 2472 840 2488
rect 1208 2472 1240 2488
rect 1256 2472 1272 2488
rect 1480 2472 1496 2488
rect 1624 2472 1640 2488
rect 1928 2472 1944 2488
rect 2520 2472 2536 2488
rect 2552 2472 2568 2488
rect 2760 2472 2776 2488
rect 2984 2472 3000 2488
rect 3736 2472 3752 2488
rect 3896 2472 3912 2488
rect 3928 2472 3944 2488
rect 4456 2472 4472 2488
rect 4552 2472 4568 2488
rect 4600 2472 4616 2488
rect 5912 2472 5928 2488
rect 6104 2472 6120 2488
rect 6136 2472 6152 2488
rect 6552 2472 6568 2488
rect 1624 2452 1640 2468
rect 3080 2452 3096 2468
rect 3432 2452 3448 2468
rect 408 2432 424 2448
rect 616 2432 632 2448
rect 904 2432 920 2448
rect 968 2432 984 2448
rect 1032 2432 1048 2448
rect 1080 2432 1096 2448
rect 1272 2432 1288 2448
rect 2424 2432 2440 2448
rect 2536 2432 2552 2448
rect 3176 2432 3192 2448
rect 4648 2432 4664 2448
rect 4968 2432 4984 2448
rect 5256 2432 5272 2448
rect 5368 2432 5384 2448
rect 5512 2432 5528 2448
rect 5736 2432 5752 2448
rect 5896 2432 5912 2448
rect 6088 2432 6104 2448
rect 6744 2432 6760 2448
rect 797 2402 833 2418
rect 2861 2402 2897 2418
rect 4909 2402 4945 2418
rect 520 2372 536 2388
rect 1496 2372 1512 2388
rect 1784 2372 1800 2388
rect 1992 2372 2008 2388
rect 2104 2372 2120 2388
rect 2184 2372 2216 2388
rect 2376 2372 2392 2388
rect 2488 2372 2504 2388
rect 2808 2372 2824 2388
rect 3400 2372 3416 2388
rect 4040 2372 4056 2388
rect 4232 2372 4248 2388
rect 4360 2372 4376 2388
rect 4424 2372 4440 2388
rect 4568 2372 4584 2388
rect 4760 2372 4776 2388
rect 5352 2372 5368 2388
rect 6120 2372 6136 2388
rect 6200 2372 6216 2388
rect 6792 2372 6808 2388
rect 3752 2352 3768 2368
rect 5064 2352 5080 2368
rect 24 2332 40 2348
rect 72 2332 88 2348
rect 152 2332 168 2348
rect 536 2332 552 2348
rect 1112 2332 1128 2348
rect 1432 2332 1448 2348
rect 1592 2332 1608 2348
rect 2168 2332 2184 2348
rect 2952 2332 2968 2348
rect 3176 2332 3192 2348
rect 3768 2332 3784 2348
rect 3800 2332 3816 2348
rect 40 2312 56 2328
rect 216 2312 232 2328
rect 312 2312 328 2328
rect 376 2312 392 2328
rect 408 2312 424 2328
rect 440 2312 456 2328
rect 504 2312 520 2328
rect 616 2312 632 2328
rect 648 2312 664 2328
rect 776 2312 792 2328
rect 984 2312 1000 2328
rect 1080 2312 1096 2328
rect 1144 2312 1160 2328
rect 1208 2312 1224 2328
rect 1576 2312 1592 2328
rect 88 2292 104 2308
rect 184 2292 232 2308
rect 344 2292 360 2308
rect 440 2292 456 2308
rect 488 2292 504 2308
rect 520 2292 536 2308
rect 584 2292 600 2308
rect 712 2292 728 2308
rect 760 2292 776 2308
rect 824 2292 840 2308
rect 920 2292 936 2308
rect 952 2292 968 2308
rect 1064 2292 1080 2308
rect 1096 2292 1112 2308
rect 1128 2292 1144 2308
rect 1176 2292 1192 2308
rect 1304 2290 1320 2306
rect 1368 2292 1384 2308
rect 1448 2292 1464 2308
rect 1512 2292 1528 2308
rect 1544 2292 1560 2308
rect 1656 2312 1672 2328
rect 1928 2312 1944 2328
rect 2072 2312 2088 2328
rect 2120 2312 2152 2328
rect 2216 2312 2232 2328
rect 2248 2312 2264 2328
rect 2424 2312 2440 2328
rect 2536 2312 2552 2328
rect 2728 2312 2744 2328
rect 3240 2312 3256 2328
rect 3304 2312 3320 2328
rect 1624 2292 1640 2308
rect 1672 2292 1704 2308
rect 1800 2292 1816 2308
rect 1976 2292 1992 2308
rect 2008 2292 2024 2308
rect 2152 2292 2168 2308
rect 2232 2292 2248 2308
rect 2312 2292 2328 2308
rect 2360 2292 2376 2308
rect 2408 2292 2424 2308
rect 2440 2292 2456 2308
rect 2488 2292 2504 2308
rect 2632 2290 2648 2306
rect 2696 2292 2712 2308
rect 2776 2292 2792 2308
rect 2856 2292 2872 2308
rect 2904 2292 2920 2308
rect 2936 2292 2952 2308
rect 3080 2290 3096 2306
rect 3208 2292 3240 2308
rect 3272 2292 3288 2308
rect 3368 2312 3384 2328
rect 3672 2312 3688 2328
rect 3400 2292 3416 2308
rect 3528 2292 3544 2308
rect 3640 2292 3656 2308
rect 3768 2292 3784 2308
rect 3848 2312 3864 2328
rect 4632 2312 4648 2328
rect 3880 2292 3896 2308
rect 3944 2292 3960 2308
rect 4008 2292 4024 2308
rect 4072 2292 4088 2308
rect 4184 2292 4216 2308
rect 4312 2292 4344 2308
rect 4392 2292 4408 2308
rect 4504 2292 4520 2308
rect 4600 2292 4616 2308
rect 5128 2312 5160 2328
rect 5288 2312 5304 2328
rect 5368 2312 5384 2328
rect 5416 2312 5432 2328
rect 5496 2312 5512 2328
rect 5560 2312 5576 2328
rect 5640 2312 5656 2328
rect 5752 2312 5768 2328
rect 5976 2312 5992 2328
rect 6056 2312 6072 2328
rect 6472 2312 6488 2328
rect 4680 2292 4696 2308
rect 4712 2292 4728 2308
rect 4776 2292 4792 2308
rect 4840 2292 4856 2308
rect 4968 2292 4984 2308
rect 5096 2292 5112 2308
rect 5144 2292 5192 2308
rect 5208 2292 5224 2308
rect 5288 2292 5304 2308
rect 5320 2292 5336 2308
rect 5416 2292 5448 2308
rect 5528 2292 5544 2308
rect 5560 2292 5592 2308
rect 5688 2292 5736 2308
rect 5768 2292 5784 2308
rect 5800 2292 5816 2308
rect 5928 2292 5944 2308
rect 5960 2292 5976 2308
rect 6040 2292 6056 2308
rect 6168 2292 6184 2308
rect 6344 2292 6360 2308
rect 6440 2292 6456 2308
rect 6600 2312 6616 2328
rect 6520 2292 6536 2308
rect 6568 2292 6600 2308
rect 8 2272 24 2288
rect 120 2272 136 2288
rect 168 2272 184 2288
rect 248 2272 280 2288
rect 296 2272 312 2288
rect 360 2272 376 2288
rect 424 2272 440 2288
rect 488 2272 504 2288
rect 568 2272 584 2288
rect 648 2272 664 2288
rect 680 2272 696 2288
rect 712 2272 728 2288
rect 840 2272 872 2288
rect 936 2272 952 2288
rect 1016 2272 1048 2288
rect 1064 2272 1080 2288
rect 1160 2272 1176 2288
rect 1192 2272 1208 2288
rect 1240 2272 1256 2288
rect 1464 2272 1480 2288
rect 1496 2272 1512 2288
rect 1528 2272 1544 2288
rect 1592 2272 1608 2288
rect 1640 2272 1656 2288
rect 1704 2272 1720 2288
rect 1752 2272 1768 2288
rect 2024 2272 2072 2288
rect 2088 2272 2104 2288
rect 2568 2272 2584 2288
rect 2664 2272 2680 2288
rect 2888 2272 2904 2288
rect 2936 2272 2952 2288
rect 3048 2272 3064 2288
rect 3112 2272 3128 2288
rect 3144 2272 3160 2288
rect 3192 2272 3208 2288
rect 3256 2272 3272 2288
rect 3352 2272 3368 2288
rect 3416 2272 3432 2288
rect 3496 2272 3512 2288
rect 3624 2272 3640 2288
rect 3720 2272 3736 2288
rect 3800 2272 3816 2288
rect 3896 2272 3912 2288
rect 4248 2272 4264 2288
rect 4536 2272 4552 2288
rect 4584 2272 4600 2288
rect 4664 2272 4680 2288
rect 4696 2272 4728 2288
rect 4792 2272 4824 2288
rect 4904 2272 4920 2288
rect 5080 2272 5096 2288
rect 5192 2272 5208 2288
rect 5224 2272 5240 2288
rect 5432 2272 5464 2288
rect 5480 2272 5496 2288
rect 5512 2272 5528 2288
rect 5608 2272 5624 2288
rect 5656 2272 5672 2288
rect 5688 2272 5704 2288
rect 5864 2288 5880 2292
rect 6664 2290 6680 2306
rect 5864 2276 5896 2288
rect 5880 2272 5896 2276
rect 5960 2272 5976 2288
rect 6040 2272 6056 2288
rect 6088 2272 6104 2288
rect 6392 2272 6408 2288
rect 6424 2272 6440 2288
rect 6536 2272 6568 2288
rect 6632 2272 6648 2288
rect 6776 2272 6792 2288
rect 440 2252 456 2268
rect 728 2252 744 2268
rect 1208 2252 1224 2268
rect 1304 2252 1320 2268
rect 1720 2252 1736 2268
rect 1880 2252 1912 2268
rect 1928 2252 1944 2268
rect 2328 2252 2344 2268
rect 2472 2252 2488 2268
rect 3976 2252 3992 2268
rect 4520 2252 4536 2268
rect 5368 2252 5384 2268
rect 5624 2252 5640 2268
rect 5816 2252 5832 2268
rect 6072 2252 6088 2268
rect 6488 2252 6504 2268
rect 72 2232 88 2248
rect 776 2232 792 2248
rect 2280 2232 2296 2248
rect 2344 2232 2360 2248
rect 2760 2232 2776 2248
rect 3176 2232 3192 2248
rect 3320 2232 3336 2248
rect 3608 2232 3624 2248
rect 4104 2232 4120 2248
rect 4152 2232 4168 2248
rect 4280 2232 4296 2248
rect 4360 2232 4376 2248
rect 4472 2232 4488 2248
rect 5064 2232 5080 2248
rect 5256 2232 5272 2248
rect 5832 2232 5848 2248
rect 5896 2232 5912 2248
rect 6232 2232 6248 2248
rect 1837 2202 1873 2218
rect 3885 2202 3921 2218
rect 5933 2202 5969 2218
rect 184 2172 200 2188
rect 472 2172 488 2188
rect 552 2172 568 2188
rect 1208 2172 1224 2188
rect 1432 2172 1448 2188
rect 1576 2172 1592 2188
rect 1704 2172 1720 2188
rect 1768 2172 1784 2188
rect 1960 2172 1976 2188
rect 2280 2172 2296 2188
rect 2408 2172 2424 2188
rect 3448 2172 3464 2188
rect 3656 2172 3672 2188
rect 3768 2172 3784 2188
rect 4008 2172 4024 2188
rect 4184 2172 4200 2188
rect 5720 2172 5736 2188
rect 5784 2172 5800 2188
rect 5880 2172 5896 2188
rect 6168 2172 6184 2188
rect 6504 2172 6520 2188
rect 6552 2172 6568 2188
rect 312 2152 344 2168
rect 1304 2152 1320 2168
rect 2328 2152 2344 2168
rect 2456 2152 2472 2168
rect 4072 2152 4104 2168
rect 4200 2152 4216 2168
rect 5144 2152 5160 2168
rect 6104 2152 6120 2168
rect 6232 2152 6248 2168
rect 6616 2152 6632 2168
rect 6664 2152 6680 2168
rect 200 2132 216 2148
rect 264 2132 280 2148
rect 392 2132 408 2148
rect 424 2132 456 2148
rect 536 2132 552 2148
rect 584 2132 600 2148
rect 648 2132 680 2148
rect 760 2132 776 2148
rect 872 2132 888 2148
rect 1464 2132 1528 2148
rect 1608 2132 1656 2148
rect 1752 2132 1768 2148
rect 1784 2132 1800 2148
rect 1928 2132 1944 2148
rect 1976 2132 2008 2148
rect 2120 2132 2136 2148
rect 2232 2132 2248 2148
rect 2264 2132 2280 2148
rect 2296 2132 2312 2148
rect 2360 2132 2376 2148
rect 2456 2132 2472 2148
rect 2648 2132 2664 2148
rect 2696 2132 2712 2148
rect 2728 2132 2744 2148
rect 2792 2132 2808 2148
rect 2888 2132 2904 2148
rect 2936 2132 2952 2148
rect 3032 2132 3048 2148
rect 3128 2132 3144 2148
rect 3208 2132 3224 2148
rect 3240 2132 3256 2148
rect 3336 2132 3352 2148
rect 3368 2132 3384 2148
rect 3400 2132 3416 2148
rect 3464 2132 3480 2148
rect 3512 2132 3544 2148
rect 3592 2132 3640 2148
rect 3656 2132 3672 2148
rect 3688 2132 3704 2148
rect 3768 2132 3784 2148
rect 3800 2132 3816 2148
rect 3848 2132 3864 2148
rect 3928 2132 3960 2148
rect 3992 2132 4008 2148
rect 4056 2132 4072 2148
rect 4168 2132 4184 2148
rect 4232 2132 4248 2148
rect 4312 2132 4328 2148
rect 4360 2132 4392 2148
rect 4424 2132 4456 2148
rect 4536 2132 4552 2148
rect 4648 2132 4664 2148
rect 4824 2132 4840 2148
rect 5080 2132 5096 2148
rect 5176 2132 5192 2148
rect 5368 2132 5384 2148
rect 5656 2132 5672 2148
rect 5832 2132 5864 2148
rect 5896 2132 5912 2148
rect 5928 2132 5944 2148
rect 6024 2132 6040 2148
rect 6056 2132 6072 2148
rect 6088 2132 6104 2148
rect 6136 2132 6152 2148
rect 6184 2132 6200 2148
rect 6296 2132 6312 2148
rect 6344 2132 6376 2148
rect 6424 2132 6440 2148
rect 6472 2132 6488 2148
rect 6600 2132 6616 2148
rect 6680 2132 6696 2148
rect 6744 2132 6760 2148
rect 72 2112 88 2128
rect 120 2112 136 2128
rect 216 2112 232 2128
rect 248 2112 264 2128
rect 280 2112 296 2128
rect 376 2112 392 2128
rect 408 2112 424 2128
rect 232 2092 248 2108
rect 520 2112 536 2128
rect 616 2112 648 2128
rect 680 2112 696 2128
rect 488 2092 504 2108
rect 552 2092 568 2108
rect 600 2092 616 2108
rect 712 2092 728 2108
rect 872 2112 888 2128
rect 920 2112 936 2128
rect 1048 2114 1064 2130
rect 1112 2112 1128 2128
rect 1240 2112 1256 2128
rect 1304 2114 1320 2130
rect 1448 2112 1464 2128
rect 1512 2112 1528 2128
rect 1544 2112 1560 2128
rect 1592 2112 1608 2128
rect 1656 2112 1688 2128
rect 1720 2112 1736 2128
rect 1800 2112 1816 2128
rect 1848 2112 1864 2128
rect 1896 2112 1912 2128
rect 1976 2112 1992 2128
rect 2008 2112 2024 2128
rect 2040 2092 2056 2108
rect 2072 2112 2104 2128
rect 2136 2112 2152 2128
rect 2216 2112 2232 2128
rect 2248 2112 2264 2128
rect 2328 2112 2344 2128
rect 2408 2112 2424 2128
rect 2520 2112 2536 2128
rect 2664 2114 2680 2130
rect 2744 2112 2760 2128
rect 2792 2112 2824 2128
rect 2952 2112 2968 2128
rect 3000 2112 3016 2128
rect 2148 2092 2164 2108
rect 2168 2092 2184 2108
rect 2204 2092 2220 2108
rect 2776 2092 2792 2108
rect 2840 2092 2856 2108
rect 2968 2092 2984 2108
rect 3016 2092 3032 2108
rect 3112 2112 3128 2128
rect 3144 2112 3160 2128
rect 3192 2112 3208 2128
rect 3288 2112 3304 2128
rect 3320 2112 3336 2128
rect 3352 2112 3368 2128
rect 3384 2112 3400 2128
rect 3416 2112 3432 2128
rect 3080 2092 3096 2108
rect 3144 2092 3160 2108
rect 3208 2092 3224 2108
rect 3304 2092 3320 2108
rect 3448 2092 3464 2108
rect 3512 2112 3544 2128
rect 3560 2112 3592 2128
rect 3608 2112 3624 2128
rect 3688 2112 3720 2128
rect 3816 2112 3832 2128
rect 3736 2092 3752 2108
rect 3864 2112 3880 2128
rect 3976 2112 3992 2128
rect 4008 2112 4024 2128
rect 4040 2112 4056 2128
rect 4168 2112 4184 2128
rect 4200 2112 4216 2128
rect 4328 2112 4344 2128
rect 4376 2112 4408 2128
rect 4456 2112 4472 2128
rect 4280 2092 4296 2108
rect 4424 2092 4440 2108
rect 4488 2092 4504 2108
rect 4568 2112 4584 2128
rect 4600 2112 4616 2128
rect 4744 2112 4760 2128
rect 4952 2112 4968 2128
rect 5000 2112 5016 2128
rect 5096 2112 5112 2128
rect 5144 2112 5160 2128
rect 5208 2112 5224 2128
rect 5256 2112 5272 2128
rect 5416 2112 5448 2128
rect 5592 2114 5608 2130
rect 4616 2092 4632 2108
rect 5224 2092 5240 2108
rect 5256 2092 5272 2108
rect 5304 2092 5320 2108
rect 5768 2092 5784 2108
rect 5816 2112 5832 2128
rect 5912 2112 5928 2128
rect 5880 2092 5896 2108
rect 6072 2112 6088 2128
rect 6120 2112 6152 2128
rect 6200 2112 6216 2128
rect 6264 2112 6296 2128
rect 6312 2112 6328 2128
rect 6344 2112 6360 2128
rect 6376 2112 6392 2128
rect 6424 2112 6440 2128
rect 6456 2112 6472 2128
rect 6536 2112 6552 2128
rect 6584 2112 6600 2128
rect 6696 2112 6728 2128
rect 5992 2092 6008 2108
rect 6040 2092 6056 2108
rect 6408 2092 6440 2108
rect 6552 2092 6568 2108
rect 2056 2072 2072 2088
rect 2536 2072 2552 2088
rect 2904 2072 2920 2088
rect 3272 2072 3288 2088
rect 4584 2072 4600 2088
rect 4664 2072 4680 2088
rect 5688 2072 5704 2088
rect 6104 2072 6120 2088
rect 3224 2052 3240 2068
rect 4632 2052 4648 2068
rect 5272 2052 5288 2068
rect 280 2032 296 2048
rect 744 2032 760 2048
rect 984 2032 1000 2048
rect 1176 2032 1192 2048
rect 1704 2032 1720 2048
rect 1880 2032 1896 2048
rect 3288 2032 3304 2048
rect 5064 2032 5080 2048
rect 6504 2032 6520 2048
rect 797 2002 833 2018
rect 2861 2002 2897 2018
rect 4909 2002 4945 2018
rect 408 1972 424 1988
rect 872 1972 888 1988
rect 1048 1972 1064 1988
rect 1128 1972 1144 1988
rect 2072 1972 2088 1988
rect 2328 1972 2344 1988
rect 2408 1972 2424 1988
rect 2504 1972 2520 1988
rect 3160 1972 3176 1988
rect 3544 1972 3560 1988
rect 3592 1972 3608 1988
rect 4008 1972 4024 1988
rect 4056 1972 4072 1988
rect 4392 1972 4408 1988
rect 4552 1972 4568 1988
rect 4888 1972 4904 1988
rect 4952 1972 4968 1988
rect 6648 1972 6664 1988
rect 264 1952 280 1968
rect 1336 1952 1352 1968
rect 200 1932 216 1948
rect 280 1932 296 1948
rect 760 1932 776 1948
rect 856 1932 872 1948
rect 1064 1932 1080 1948
rect 1304 1932 1320 1948
rect 1960 1932 1976 1948
rect 2184 1932 2200 1948
rect 2232 1932 2248 1948
rect 2264 1932 2280 1948
rect 2904 1932 2920 1948
rect 3240 1932 3256 1948
rect 3496 1932 3512 1948
rect 3528 1932 3544 1948
rect 4408 1932 4424 1948
rect 4872 1932 4888 1948
rect 5496 1932 5512 1948
rect 5528 1932 5544 1948
rect 6168 1932 6184 1948
rect 232 1912 248 1928
rect 452 1912 468 1928
rect 488 1912 504 1928
rect 552 1912 568 1928
rect 616 1912 632 1928
rect 636 1912 652 1928
rect 728 1912 744 1928
rect 776 1912 792 1928
rect 824 1912 840 1928
rect 936 1912 952 1928
rect 1032 1912 1048 1928
rect 1096 1912 1112 1928
rect 1400 1912 1432 1928
rect 1448 1912 1464 1928
rect 1528 1912 1544 1928
rect 2056 1912 2072 1928
rect 2088 1912 2104 1928
rect 2264 1912 2280 1928
rect 2600 1912 2616 1928
rect 2680 1912 2696 1928
rect 104 1892 136 1908
rect 264 1892 280 1908
rect 312 1892 328 1908
rect 392 1892 408 1908
rect 424 1892 440 1908
rect 536 1892 552 1908
rect 584 1892 600 1908
rect 648 1892 696 1908
rect 840 1892 856 1908
rect 904 1892 920 1908
rect 1016 1892 1032 1908
rect 1048 1892 1064 1908
rect 1128 1892 1144 1908
rect 1256 1892 1272 1908
rect 1368 1892 1400 1908
rect 1496 1892 1512 1908
rect 1560 1892 1576 1908
rect 1592 1892 1608 1908
rect 1656 1892 1672 1908
rect 1688 1892 1704 1908
rect 1768 1892 1784 1908
rect 1800 1892 1816 1908
rect 1832 1892 1848 1908
rect 1864 1892 1880 1908
rect 1960 1892 1976 1908
rect 2024 1892 2040 1908
rect 2072 1892 2088 1908
rect 2104 1892 2120 1908
rect 2168 1892 2184 1908
rect 2296 1892 2312 1908
rect 2424 1892 2440 1908
rect 2472 1892 2504 1908
rect 2552 1892 2568 1908
rect 2632 1892 2648 1908
rect 2664 1892 2680 1908
rect 2728 1912 2744 1928
rect 2840 1912 2856 1928
rect 2936 1912 2952 1928
rect 2760 1892 2776 1908
rect 200 1872 216 1888
rect 328 1872 376 1888
rect 424 1872 440 1888
rect 536 1872 568 1888
rect 600 1872 616 1888
rect 664 1872 696 1888
rect 728 1872 760 1888
rect 888 1872 904 1888
rect 952 1872 968 1888
rect 1000 1872 1016 1888
rect 1144 1872 1160 1888
rect 1352 1872 1368 1888
rect 1448 1872 1480 1888
rect 1512 1872 1528 1888
rect 1544 1872 1560 1888
rect 1576 1872 1608 1888
rect 1704 1872 1720 1888
rect 1784 1872 1800 1888
rect 1880 1872 1896 1888
rect 2120 1872 2136 1888
rect 2152 1872 2184 1888
rect 2216 1872 2232 1888
rect 2264 1872 2280 1888
rect 2376 1872 2392 1888
rect 2504 1872 2520 1888
rect 2536 1872 2552 1888
rect 2568 1872 2584 1888
rect 2616 1872 2632 1888
rect 2680 1872 2696 1888
rect 2776 1872 2792 1888
rect 2808 1892 2824 1908
rect 2856 1892 2872 1908
rect 3000 1912 3016 1928
rect 3064 1912 3080 1928
rect 3288 1912 3304 1928
rect 4104 1912 4120 1928
rect 4280 1912 4296 1928
rect 4324 1912 4340 1928
rect 4344 1912 4360 1928
rect 4520 1912 4536 1928
rect 4632 1912 4648 1928
rect 4776 1912 4792 1928
rect 3032 1892 3048 1908
rect 3096 1892 3112 1908
rect 3128 1892 3144 1908
rect 3176 1892 3192 1908
rect 3256 1892 3272 1908
rect 3336 1892 3352 1908
rect 3400 1890 3416 1906
rect 3464 1892 3480 1908
rect 3624 1892 3656 1908
rect 3688 1892 3704 1908
rect 3768 1892 3784 1908
rect 3832 1890 3848 1906
rect 3976 1892 3992 1908
rect 4040 1892 4056 1908
rect 4088 1892 4104 1908
rect 4168 1892 4184 1908
rect 4232 1892 4264 1908
rect 4280 1892 4296 1908
rect 4392 1892 4408 1908
rect 4456 1892 4472 1908
rect 4552 1892 4568 1908
rect 4600 1892 4616 1908
rect 4712 1892 4728 1908
rect 4744 1892 4760 1908
rect 4904 1912 4920 1928
rect 4968 1912 4984 1928
rect 5000 1912 5016 1928
rect 4808 1892 4840 1908
rect 4888 1892 4904 1908
rect 5048 1892 5064 1908
rect 5208 1912 5224 1928
rect 5272 1912 5288 1928
rect 5096 1892 5112 1908
rect 5160 1892 5176 1908
rect 5240 1892 5256 1908
rect 5352 1892 5368 1908
rect 5416 1912 5432 1928
rect 5560 1912 5576 1928
rect 5800 1912 5816 1928
rect 5928 1912 5944 1928
rect 5496 1892 5512 1908
rect 5544 1892 5560 1908
rect 5576 1892 5592 1908
rect 5656 1892 5672 1908
rect 5720 1892 5736 1908
rect 5752 1892 5768 1908
rect 5832 1892 5848 1908
rect 5880 1892 5896 1908
rect 6072 1912 6088 1928
rect 6152 1912 6168 1928
rect 6408 1912 6424 1928
rect 6456 1912 6472 1928
rect 6504 1912 6520 1928
rect 6632 1912 6648 1928
rect 6712 1912 6728 1928
rect 5976 1892 6008 1908
rect 6024 1892 6040 1908
rect 6104 1892 6136 1908
rect 6152 1892 6168 1908
rect 6232 1892 6264 1908
rect 6376 1892 6392 1908
rect 6536 1892 6552 1908
rect 6584 1892 6616 1908
rect 6696 1892 6712 1908
rect 2888 1872 2904 1888
rect 2952 1872 2968 1888
rect 3048 1872 3080 1888
rect 3112 1872 3128 1888
rect 3208 1872 3224 1888
rect 3256 1872 3272 1888
rect 3288 1872 3304 1888
rect 3320 1872 3336 1888
rect 3672 1872 3688 1888
rect 3768 1872 3784 1888
rect 3944 1872 3960 1888
rect 4104 1872 4120 1888
rect 4136 1872 4152 1888
rect 4232 1872 4248 1888
rect 4296 1872 4312 1888
rect 4440 1872 4456 1888
rect 4568 1872 4600 1888
rect 4648 1872 4664 1888
rect 4680 1872 4712 1888
rect 4728 1872 4744 1888
rect 4840 1872 4856 1888
rect 4984 1872 5000 1888
rect 5016 1872 5048 1888
rect 5112 1872 5128 1888
rect 5144 1872 5176 1888
rect 5224 1872 5240 1888
rect 5304 1872 5320 1888
rect 5336 1872 5352 1888
rect 5368 1872 5400 1888
rect 5448 1872 5464 1888
rect 5640 1872 5656 1888
rect 5704 1872 5720 1888
rect 5848 1872 5880 1888
rect 6008 1872 6024 1888
rect 6040 1872 6056 1888
rect 6088 1872 6120 1888
rect 6360 1872 6376 1888
rect 6424 1872 6440 1888
rect 6472 1872 6488 1888
rect 6584 1872 6600 1888
rect 6616 1872 6632 1888
rect 6808 1872 6824 1888
rect 392 1852 408 1868
rect 968 1852 984 1868
rect 1208 1852 1224 1868
rect 1640 1852 1656 1868
rect 1832 1852 1848 1868
rect 1896 1852 1912 1868
rect 1928 1852 1944 1868
rect 2344 1852 2360 1868
rect 2472 1852 2488 1868
rect 3560 1852 3576 1868
rect 4072 1852 4088 1868
rect 4360 1852 4376 1868
rect 4968 1852 4984 1868
rect 5464 1852 5480 1868
rect 5784 1852 5800 1868
rect 6408 1852 6424 1868
rect 6648 1852 6664 1868
rect 488 1832 504 1848
rect 1432 1832 1448 1848
rect 1736 1832 1752 1848
rect 1992 1832 2008 1848
rect 2152 1832 2168 1848
rect 2232 1832 2248 1848
rect 2600 1832 2616 1848
rect 2712 1832 2728 1848
rect 2840 1832 2856 1848
rect 2968 1832 2984 1848
rect 3592 1832 3608 1848
rect 3704 1832 3720 1848
rect 4184 1832 4200 1848
rect 4280 1832 4296 1848
rect 4376 1832 4392 1848
rect 4424 1832 4440 1848
rect 4488 1832 4504 1848
rect 4776 1832 4792 1848
rect 5080 1832 5096 1848
rect 5128 1832 5144 1848
rect 5208 1832 5224 1848
rect 5336 1832 5352 1848
rect 5512 1832 5528 1848
rect 5608 1832 5624 1848
rect 5688 1832 5704 1848
rect 5800 1832 5816 1848
rect 6456 1832 6472 1848
rect 6568 1832 6584 1848
rect 1837 1802 1873 1818
rect 3885 1802 3921 1818
rect 5933 1802 5969 1818
rect 184 1772 200 1788
rect 216 1772 232 1788
rect 456 1772 472 1788
rect 744 1772 760 1788
rect 872 1772 888 1788
rect 1096 1772 1112 1788
rect 1176 1772 1192 1788
rect 1304 1772 1320 1788
rect 1416 1772 1432 1788
rect 1736 1772 1752 1788
rect 2088 1772 2104 1788
rect 2248 1772 2264 1788
rect 2440 1772 2456 1788
rect 2488 1772 2504 1788
rect 3848 1772 3864 1788
rect 4056 1772 4072 1788
rect 4616 1772 4632 1788
rect 4872 1772 4888 1788
rect 5032 1772 5048 1788
rect 5096 1772 5112 1788
rect 5192 1772 5208 1788
rect 5464 1772 5480 1788
rect 5736 1772 5752 1788
rect 6696 1772 6712 1788
rect 200 1752 216 1768
rect 920 1752 936 1768
rect 1656 1752 1672 1768
rect 1880 1752 1896 1768
rect 2824 1752 2840 1768
rect 3000 1752 3016 1768
rect 3624 1752 3640 1768
rect 5112 1752 5128 1768
rect 5320 1752 5336 1768
rect 5480 1752 5512 1768
rect 5880 1752 5896 1768
rect 248 1732 264 1748
rect 280 1732 296 1748
rect 360 1732 376 1748
rect 424 1732 456 1748
rect 488 1732 504 1748
rect 584 1732 600 1748
rect 648 1732 680 1748
rect 760 1732 792 1748
rect 904 1732 920 1748
rect 936 1732 968 1748
rect 1064 1732 1080 1748
rect 1096 1732 1112 1748
rect 1128 1732 1144 1748
rect 1288 1732 1304 1748
rect 104 1712 136 1728
rect 232 1712 248 1728
rect 264 1712 280 1728
rect 344 1712 360 1728
rect 408 1712 424 1728
rect 488 1712 504 1728
rect 312 1692 328 1708
rect 376 1692 392 1708
rect 472 1692 488 1708
rect 536 1692 552 1708
rect 584 1712 600 1728
rect 632 1712 648 1728
rect 680 1712 696 1728
rect 600 1692 616 1708
rect 712 1692 728 1708
rect 792 1712 808 1728
rect 824 1692 840 1708
rect 968 1712 984 1728
rect 968 1692 984 1708
rect 1000 1692 1016 1708
rect 1064 1712 1096 1728
rect 1144 1712 1160 1728
rect 1224 1712 1240 1728
rect 1272 1712 1288 1728
rect 1304 1712 1320 1728
rect 1336 1712 1352 1728
rect 1368 1732 1384 1748
rect 1416 1732 1432 1748
rect 1448 1732 1480 1748
rect 1512 1732 1528 1748
rect 1576 1732 1592 1748
rect 1672 1732 1704 1748
rect 1864 1732 1880 1748
rect 1912 1732 1928 1748
rect 1976 1732 1992 1748
rect 2072 1732 2088 1748
rect 2104 1732 2120 1748
rect 2216 1732 2232 1748
rect 2248 1732 2264 1748
rect 2328 1732 2376 1748
rect 2392 1732 2408 1748
rect 2648 1732 2664 1748
rect 2760 1732 2808 1748
rect 2984 1732 3000 1748
rect 3016 1732 3032 1748
rect 3112 1732 3128 1748
rect 3192 1732 3208 1748
rect 3224 1732 3256 1748
rect 3368 1732 3384 1748
rect 3480 1732 3496 1748
rect 3656 1732 3672 1748
rect 3688 1732 3704 1748
rect 3768 1732 3784 1748
rect 3800 1732 3816 1748
rect 3976 1732 3992 1748
rect 4040 1732 4056 1748
rect 4088 1732 4120 1748
rect 4216 1732 4248 1748
rect 4296 1732 4312 1748
rect 4360 1732 4376 1748
rect 4408 1732 4424 1748
rect 4536 1732 4552 1748
rect 4600 1732 4616 1748
rect 4776 1732 4792 1748
rect 4856 1732 4872 1748
rect 4904 1732 4920 1748
rect 4968 1732 4984 1748
rect 1368 1712 1384 1728
rect 1496 1712 1512 1728
rect 1528 1712 1576 1728
rect 1592 1712 1608 1728
rect 1036 1692 1052 1708
rect 1400 1692 1432 1708
rect 1496 1692 1512 1708
rect 1560 1692 1576 1708
rect 1624 1692 1640 1708
rect 1704 1712 1720 1728
rect 1768 1712 1784 1728
rect 1848 1712 1864 1728
rect 1960 1712 1976 1728
rect 2040 1712 2072 1728
rect 2120 1712 2136 1728
rect 2152 1712 2168 1728
rect 2200 1712 2216 1728
rect 2264 1712 2280 1728
rect 2296 1712 2344 1728
rect 2408 1712 2424 1728
rect 2472 1712 2488 1728
rect 2616 1714 2632 1730
rect 2696 1712 2712 1728
rect 2744 1712 2760 1728
rect 2824 1712 2840 1728
rect 2856 1712 2872 1728
rect 2936 1712 2952 1728
rect 2968 1712 2984 1728
rect 3080 1712 3096 1728
rect 3128 1712 3144 1728
rect 3208 1712 3224 1728
rect 3256 1712 3288 1728
rect 1736 1692 1768 1708
rect 1928 1692 1944 1708
rect 2184 1692 2200 1708
rect 2280 1692 2296 1708
rect 2680 1692 2696 1708
rect 2840 1692 2856 1708
rect 2952 1692 2968 1708
rect 3048 1692 3064 1708
rect 3160 1692 3176 1708
rect 3304 1692 3320 1708
rect 3336 1712 3368 1728
rect 3416 1712 3432 1728
rect 3576 1712 3592 1728
rect 3704 1712 3720 1728
rect 3784 1712 3800 1728
rect 3816 1712 3832 1728
rect 3864 1712 3880 1728
rect 3960 1712 3976 1728
rect 4008 1712 4040 1728
rect 4120 1712 4152 1728
rect 3736 1692 3752 1708
rect 3880 1692 3896 1708
rect 3928 1692 3944 1708
rect 3960 1692 3976 1708
rect 3992 1692 4008 1708
rect 4056 1692 4072 1708
rect 4152 1692 4168 1708
rect 4216 1712 4232 1728
rect 4248 1712 4264 1728
rect 4296 1712 4328 1728
rect 4392 1712 4408 1728
rect 4424 1712 4440 1728
rect 4456 1712 4472 1728
rect 4488 1712 4504 1728
rect 4584 1712 4600 1728
rect 4712 1712 4728 1728
rect 4840 1712 4856 1728
rect 4984 1712 5000 1728
rect 5144 1732 5160 1748
rect 5512 1732 5528 1748
rect 5016 1712 5032 1728
rect 5064 1712 5096 1728
rect 5176 1712 5192 1728
rect 5256 1712 5272 1728
rect 5320 1714 5336 1730
rect 5400 1712 5416 1728
rect 5448 1712 5464 1728
rect 5560 1712 5576 1728
rect 5640 1732 5656 1748
rect 5736 1732 5752 1748
rect 5768 1732 5784 1748
rect 5800 1732 5816 1748
rect 5864 1732 5880 1748
rect 5896 1732 5912 1748
rect 6040 1732 6056 1748
rect 6088 1732 6120 1748
rect 6328 1732 6344 1748
rect 6408 1732 6424 1748
rect 6440 1732 6456 1748
rect 6616 1732 6632 1748
rect 6792 1732 6808 1748
rect 5624 1712 5640 1728
rect 5656 1712 5672 1728
rect 5720 1712 5736 1728
rect 5800 1712 5832 1728
rect 4188 1692 4204 1708
rect 4280 1692 4296 1708
rect 4344 1692 4360 1708
rect 4440 1692 4456 1708
rect 4504 1692 4520 1708
rect 4552 1692 4568 1708
rect 4808 1692 4824 1708
rect 4828 1692 4844 1708
rect 4952 1692 4968 1708
rect 5384 1692 5400 1708
rect 5528 1692 5544 1708
rect 5548 1692 5564 1708
rect 5828 1692 5844 1708
rect 5848 1692 5864 1708
rect 5928 1692 5944 1708
rect 5992 1712 6008 1728
rect 6072 1712 6088 1728
rect 6120 1712 6136 1728
rect 6232 1712 6264 1728
rect 6360 1712 6376 1728
rect 6472 1714 6488 1730
rect 6632 1712 6648 1728
rect 6728 1712 6744 1728
rect 6776 1712 6792 1728
rect 6040 1692 6056 1708
rect 6132 1692 6148 1708
rect 6152 1692 6168 1708
rect 6664 1692 6680 1708
rect 6744 1692 6760 1708
rect 1784 1672 1800 1688
rect 2168 1672 2184 1688
rect 2712 1672 2728 1688
rect 2952 1672 2968 1688
rect 3272 1672 3288 1688
rect 3400 1672 3432 1688
rect 3496 1672 3512 1688
rect 3528 1672 3544 1688
rect 3848 1672 3864 1688
rect 4472 1672 4488 1688
rect 4520 1672 4536 1688
rect 4872 1672 4888 1688
rect 5416 1672 5432 1688
rect 5944 1672 5960 1688
rect 6024 1672 6040 1688
rect 6168 1672 6184 1688
rect 1240 1652 1256 1668
rect 3416 1652 3432 1668
rect 5400 1652 5416 1668
rect 6600 1652 6616 1668
rect 408 1632 424 1648
rect 568 1632 584 1648
rect 1768 1632 1784 1648
rect 2008 1632 2024 1648
rect 2136 1632 2152 1648
rect 2360 1632 2376 1648
rect 2696 1632 2712 1648
rect 2872 1632 2888 1648
rect 2904 1632 2920 1648
rect 4584 1632 4600 1648
rect 5032 1632 5048 1648
rect 5688 1632 5704 1648
rect 797 1602 833 1618
rect 2861 1602 2897 1618
rect 4909 1602 4945 1618
rect 200 1572 216 1588
rect 1224 1572 1240 1588
rect 1368 1572 1384 1588
rect 1896 1572 1912 1588
rect 1976 1572 1992 1588
rect 2008 1572 2024 1588
rect 2456 1572 2472 1588
rect 2520 1572 2536 1588
rect 2968 1572 2984 1588
rect 3176 1572 3192 1588
rect 3288 1572 3304 1588
rect 3640 1572 3656 1588
rect 3864 1572 3880 1588
rect 4264 1572 4280 1588
rect 5224 1572 5240 1588
rect 5704 1572 5720 1588
rect 5992 1572 6008 1588
rect 6360 1572 6376 1588
rect 6424 1572 6440 1588
rect 6760 1572 6776 1588
rect 232 1532 248 1548
rect 376 1532 392 1548
rect 568 1532 584 1548
rect 904 1532 920 1548
rect 1416 1532 1432 1548
rect 2040 1532 2056 1548
rect 2952 1532 2968 1548
rect 3656 1532 3672 1548
rect 4168 1532 4184 1548
rect 4200 1532 4216 1548
rect 4344 1532 4360 1548
rect 4376 1532 4392 1548
rect 5608 1532 5624 1548
rect 6408 1532 6424 1548
rect 232 1492 248 1508
rect 312 1512 328 1528
rect 344 1492 360 1508
rect 424 1512 440 1528
rect 536 1512 552 1528
rect 600 1512 616 1528
rect 632 1512 648 1528
rect 696 1512 712 1528
rect 716 1512 732 1528
rect 760 1512 776 1528
rect 888 1512 904 1528
rect 456 1492 472 1508
rect 504 1492 520 1508
rect 584 1492 600 1508
rect 616 1492 632 1508
rect 680 1492 696 1508
rect 728 1492 760 1508
rect 808 1492 824 1508
rect 856 1492 872 1508
rect 936 1492 952 1508
rect 1016 1512 1032 1528
rect 1128 1512 1144 1528
rect 1048 1492 1064 1508
rect 8 1472 24 1488
rect 120 1472 136 1488
rect 264 1472 280 1488
rect 360 1472 392 1488
rect 472 1472 504 1488
rect 536 1472 552 1488
rect 632 1472 648 1488
rect 680 1472 696 1488
rect 744 1472 760 1488
rect 792 1472 808 1488
rect 824 1472 840 1488
rect 952 1472 984 1488
rect 1064 1472 1080 1488
rect 1096 1492 1112 1508
rect 1288 1512 1304 1528
rect 1352 1512 1368 1528
rect 1448 1512 1464 1528
rect 1512 1512 1528 1528
rect 1192 1492 1208 1508
rect 1320 1492 1352 1508
rect 1416 1492 1432 1508
rect 1480 1492 1496 1508
rect 1592 1492 1608 1508
rect 1656 1512 1672 1528
rect 2248 1512 2264 1528
rect 2312 1512 2328 1528
rect 1688 1492 1704 1508
rect 1768 1490 1784 1506
rect 1832 1492 1848 1508
rect 1976 1492 1992 1508
rect 2136 1490 2152 1506
rect 2216 1492 2232 1508
rect 2280 1492 2296 1508
rect 2376 1512 2392 1528
rect 2504 1512 2520 1528
rect 2536 1512 2552 1528
rect 2360 1492 2376 1508
rect 2408 1492 2424 1508
rect 2488 1492 2504 1508
rect 2520 1492 2536 1508
rect 2616 1492 2632 1508
rect 2680 1492 2712 1508
rect 2856 1492 2872 1508
rect 3032 1512 3048 1528
rect 3144 1512 3160 1528
rect 3112 1492 3128 1508
rect 3304 1512 3320 1528
rect 3432 1512 3448 1528
rect 3720 1512 3736 1528
rect 3848 1512 3864 1528
rect 3992 1512 4040 1528
rect 4136 1512 4152 1528
rect 4216 1512 4232 1528
rect 4456 1512 4472 1528
rect 4552 1512 4568 1528
rect 4616 1512 4632 1528
rect 4680 1512 4696 1528
rect 4776 1512 4792 1528
rect 5112 1512 5128 1528
rect 5176 1512 5192 1528
rect 5208 1512 5224 1528
rect 5288 1512 5304 1528
rect 5352 1512 5368 1528
rect 5384 1512 5400 1528
rect 5464 1512 5480 1528
rect 5496 1512 5512 1528
rect 5516 1512 5532 1528
rect 5800 1512 5816 1528
rect 5896 1512 5912 1528
rect 6024 1512 6040 1528
rect 6184 1512 6200 1528
rect 6456 1512 6472 1528
rect 6792 1512 6808 1528
rect 3208 1492 3224 1508
rect 3272 1492 3288 1508
rect 3336 1492 3352 1508
rect 3416 1492 3432 1508
rect 3464 1492 3480 1508
rect 3544 1492 3576 1508
rect 3688 1492 3720 1508
rect 3784 1492 3800 1508
rect 3816 1492 3848 1508
rect 3864 1492 3880 1508
rect 3960 1492 3976 1508
rect 4056 1492 4072 1508
rect 4120 1492 4136 1508
rect 4152 1492 4168 1508
rect 4296 1492 4312 1508
rect 4392 1492 4408 1508
rect 4472 1492 4488 1508
rect 4504 1492 4520 1508
rect 4584 1492 4600 1508
rect 4632 1492 4664 1508
rect 4680 1492 4696 1508
rect 4712 1492 4728 1508
rect 4744 1492 4760 1508
rect 4904 1492 4936 1508
rect 5000 1492 5016 1508
rect 5064 1492 5080 1508
rect 5096 1492 5112 1508
rect 5128 1492 5144 1508
rect 5160 1492 5176 1508
rect 5192 1492 5208 1508
rect 5256 1492 5272 1508
rect 5368 1492 5384 1508
rect 5448 1492 5464 1508
rect 5480 1492 5496 1508
rect 5752 1492 5768 1508
rect 5800 1492 5816 1508
rect 5864 1492 5880 1508
rect 6008 1492 6024 1508
rect 6040 1492 6056 1508
rect 6104 1492 6120 1508
rect 6184 1492 6232 1508
rect 6264 1492 6280 1508
rect 6296 1492 6312 1508
rect 6424 1492 6440 1508
rect 6568 1492 6584 1508
rect 6696 1492 6712 1508
rect 6760 1492 6776 1508
rect 1176 1472 1192 1488
rect 1256 1472 1272 1488
rect 1304 1472 1320 1488
rect 1384 1472 1400 1488
rect 1464 1472 1480 1488
rect 1544 1472 1560 1488
rect 1576 1472 1592 1488
rect 1608 1472 1624 1488
rect 1704 1472 1720 1488
rect 1736 1472 1752 1488
rect 1992 1472 2008 1488
rect 2168 1472 2184 1488
rect 2200 1472 2216 1488
rect 2264 1472 2280 1488
rect 2360 1472 2376 1488
rect 2424 1472 2440 1488
rect 2632 1472 2648 1488
rect 2776 1472 2792 1488
rect 2984 1472 3000 1488
rect 3080 1472 3112 1488
rect 3192 1472 3224 1488
rect 3352 1472 3384 1488
rect 3608 1472 3624 1488
rect 3672 1472 3688 1488
rect 3768 1472 3784 1488
rect 3800 1472 3816 1488
rect 3944 1472 3960 1488
rect 3992 1472 4008 1488
rect 4040 1472 4056 1488
rect 4072 1472 4120 1488
rect 4232 1472 4248 1488
rect 4312 1472 4328 1488
rect 4344 1472 4360 1488
rect 4424 1472 4440 1488
rect 4488 1472 4504 1488
rect 4520 1472 4536 1488
rect 4600 1472 4616 1488
rect 4664 1472 4680 1488
rect 4728 1472 4744 1488
rect 4792 1472 4808 1488
rect 5000 1472 5016 1488
rect 5080 1472 5096 1488
rect 5160 1472 5176 1488
rect 5240 1472 5256 1488
rect 5320 1472 5336 1488
rect 5368 1472 5384 1488
rect 5416 1472 5432 1488
rect 5544 1472 5560 1488
rect 5656 1472 5672 1488
rect 5736 1472 5752 1488
rect 5832 1472 5864 1488
rect 5960 1472 5976 1488
rect 5992 1472 6008 1488
rect 6072 1472 6088 1488
rect 6120 1472 6136 1488
rect 6232 1472 6248 1488
rect 6280 1472 6296 1488
rect 6312 1472 6328 1488
rect 6488 1472 6504 1488
rect 6520 1472 6536 1488
rect 6568 1472 6584 1488
rect 6744 1472 6760 1488
rect 88 1452 104 1468
rect 1384 1452 1400 1468
rect 3272 1452 3288 1468
rect 3592 1452 3608 1468
rect 3736 1452 3752 1468
rect 3896 1452 3912 1468
rect 5576 1452 5592 1468
rect 5816 1452 5832 1468
rect 6104 1452 6120 1468
rect 6168 1452 6184 1468
rect 6248 1452 6264 1468
rect 6616 1452 6632 1468
rect 24 1432 40 1448
rect 104 1432 120 1448
rect 168 1432 184 1448
rect 568 1432 584 1448
rect 760 1432 776 1448
rect 904 1432 920 1448
rect 984 1432 1000 1448
rect 1144 1432 1160 1448
rect 1288 1432 1304 1448
rect 1560 1432 1576 1448
rect 1640 1432 1656 1448
rect 2248 1432 2264 1448
rect 2344 1432 2360 1448
rect 2584 1432 2600 1448
rect 2728 1432 2744 1448
rect 3304 1432 3320 1448
rect 3432 1432 3448 1448
rect 3512 1432 3528 1448
rect 3752 1432 3768 1448
rect 4168 1432 4184 1448
rect 4392 1432 4408 1448
rect 5000 1432 5016 1448
rect 6328 1432 6344 1448
rect 6728 1432 6744 1448
rect 1837 1402 1873 1418
rect 3885 1402 3921 1418
rect 5933 1402 5969 1418
rect 600 1372 632 1388
rect 1688 1372 1704 1388
rect 1800 1372 1816 1388
rect 2056 1372 2072 1388
rect 2104 1372 2120 1388
rect 2184 1372 2200 1388
rect 2408 1372 2424 1388
rect 2520 1372 2536 1388
rect 3176 1372 3192 1388
rect 3512 1372 3528 1388
rect 4232 1372 4248 1388
rect 4600 1372 4616 1388
rect 5064 1372 5080 1388
rect 5416 1372 5432 1388
rect 5528 1372 5560 1388
rect 5640 1372 5656 1388
rect 5704 1372 5720 1388
rect 6104 1372 6120 1388
rect 6712 1372 6728 1388
rect 6792 1372 6808 1388
rect 104 1352 120 1368
rect 392 1352 408 1368
rect 1752 1352 1768 1368
rect 2344 1352 2360 1368
rect 3784 1352 3800 1368
rect 4072 1352 4088 1368
rect 4952 1352 4968 1368
rect 5000 1352 5016 1368
rect 5992 1352 6008 1368
rect 6152 1352 6168 1368
rect 6440 1352 6456 1368
rect 6696 1352 6712 1368
rect 8 1332 24 1348
rect 56 1332 72 1348
rect 136 1332 152 1348
rect 216 1332 232 1348
rect 312 1332 328 1348
rect 440 1332 456 1348
rect 776 1332 792 1348
rect 856 1332 872 1348
rect 888 1332 904 1348
rect 984 1332 1000 1348
rect 1080 1332 1096 1348
rect 1160 1332 1176 1348
rect 1304 1332 1320 1348
rect 1336 1332 1352 1348
rect 1432 1332 1448 1348
rect 1480 1332 1496 1348
rect 1544 1332 1560 1348
rect 1992 1332 2008 1348
rect 2040 1332 2056 1348
rect 2072 1332 2088 1348
rect 2136 1332 2152 1348
rect 2200 1332 2216 1348
rect 2296 1332 2312 1348
rect 2616 1332 2632 1348
rect 2712 1332 2728 1348
rect 2808 1332 2840 1348
rect 2936 1332 2952 1348
rect 2968 1332 2984 1348
rect 3064 1332 3080 1348
rect 3160 1332 3176 1348
rect 3288 1332 3304 1348
rect 3368 1332 3384 1348
rect 3480 1332 3528 1348
rect 3544 1332 3560 1348
rect 3576 1332 3592 1348
rect 3688 1332 3704 1348
rect 3720 1332 3736 1348
rect 3752 1332 3768 1348
rect 3944 1332 3960 1348
rect 4056 1332 4072 1348
rect 4104 1332 4120 1348
rect 4136 1332 4152 1348
rect 4216 1332 4232 1348
rect 4616 1332 4632 1348
rect 4680 1332 4696 1348
rect 4712 1332 4728 1348
rect 4776 1332 4792 1348
rect 5016 1332 5032 1348
rect 5128 1332 5160 1348
rect 5256 1332 5272 1348
rect 5384 1332 5400 1348
rect 5448 1332 5464 1348
rect 5480 1332 5496 1348
rect 5592 1332 5624 1348
rect 5688 1332 5704 1348
rect 5896 1332 5912 1348
rect 6008 1332 6040 1348
rect 6072 1332 6088 1348
rect 6200 1332 6232 1348
rect 40 1312 56 1328
rect 152 1312 168 1328
rect 248 1314 264 1330
rect 520 1312 536 1328
rect 744 1314 760 1330
rect 840 1312 856 1328
rect 904 1312 920 1328
rect 936 1312 952 1328
rect 184 1292 200 1308
rect 888 1292 904 1308
rect 920 1292 936 1308
rect 968 1292 984 1308
rect 1064 1312 1080 1328
rect 1192 1312 1224 1328
rect 1288 1312 1304 1328
rect 1352 1312 1368 1328
rect 1400 1312 1416 1328
rect 1496 1312 1528 1328
rect 1560 1312 1576 1328
rect 1624 1312 1640 1328
rect 1656 1312 1672 1328
rect 1736 1312 1752 1328
rect 1784 1312 1800 1328
rect 1912 1312 1928 1328
rect 2024 1312 2040 1328
rect 2104 1312 2120 1328
rect 2152 1312 2168 1328
rect 2264 1312 2280 1328
rect 2360 1312 2376 1328
rect 2440 1312 2456 1328
rect 2504 1312 2520 1328
rect 2584 1312 2616 1328
rect 2728 1312 2744 1328
rect 1032 1292 1048 1308
rect 1336 1292 1352 1308
rect 1432 1292 1448 1308
rect 1464 1292 1480 1308
rect 1528 1292 1544 1308
rect 1592 1292 1624 1308
rect 2104 1292 2120 1308
rect 2232 1292 2264 1308
rect 2376 1292 2392 1308
rect 2760 1292 2776 1308
rect 2808 1312 2824 1328
rect 2840 1312 2856 1328
rect 2984 1312 3000 1328
rect 3016 1312 3032 1328
rect 2872 1292 2888 1308
rect 3000 1292 3016 1308
rect 3144 1312 3160 1328
rect 3304 1314 3320 1330
rect 3384 1312 3416 1328
rect 3112 1292 3128 1308
rect 3432 1312 3496 1328
rect 3560 1312 3576 1328
rect 3592 1312 3608 1328
rect 3432 1292 3448 1308
rect 3624 1292 3640 1308
rect 3656 1312 3704 1328
rect 3912 1314 3928 1330
rect 3976 1312 3992 1328
rect 4040 1312 4056 1328
rect 4104 1312 4120 1328
rect 3720 1292 3736 1308
rect 4008 1292 4024 1308
rect 4088 1292 4104 1308
rect 4200 1312 4216 1328
rect 4312 1312 4328 1328
rect 4472 1314 4488 1330
rect 4536 1312 4552 1328
rect 4632 1312 4648 1328
rect 4664 1312 4680 1328
rect 4744 1312 4760 1328
rect 4840 1312 4856 1328
rect 5032 1312 5048 1328
rect 4168 1292 4184 1308
rect 5112 1312 5128 1328
rect 5144 1312 5160 1328
rect 5080 1292 5096 1308
rect 5160 1292 5176 1308
rect 5240 1312 5256 1328
rect 5272 1312 5288 1328
rect 5336 1312 5352 1328
rect 5400 1312 5416 1328
rect 5464 1312 5512 1328
rect 5576 1312 5592 1328
rect 5208 1292 5224 1308
rect 5528 1292 5544 1308
rect 5768 1312 5800 1328
rect 5656 1292 5672 1308
rect 5928 1292 5944 1308
rect 6040 1312 6056 1328
rect 6136 1312 6152 1328
rect 6184 1312 6200 1328
rect 6280 1312 6296 1328
rect 6392 1332 6408 1348
rect 6424 1332 6440 1348
rect 6472 1332 6488 1348
rect 6504 1332 6520 1348
rect 6584 1332 6600 1348
rect 6616 1332 6648 1348
rect 6728 1332 6744 1348
rect 6344 1312 6360 1328
rect 6072 1292 6088 1308
rect 6152 1292 6168 1308
rect 6248 1292 6264 1308
rect 6456 1312 6472 1328
rect 6488 1312 6504 1328
rect 6520 1312 6536 1328
rect 6392 1292 6408 1308
rect 6552 1292 6568 1308
rect 6600 1312 6616 1328
rect 6648 1312 6664 1328
rect 6744 1312 6760 1328
rect 6660 1292 6676 1308
rect 6680 1292 6696 1308
rect 6776 1292 6792 1308
rect 344 1272 360 1288
rect 952 1272 968 1288
rect 1272 1272 1288 1288
rect 1640 1272 1656 1288
rect 1864 1272 1880 1288
rect 2344 1272 2360 1288
rect 3032 1272 3048 1288
rect 3064 1272 3080 1288
rect 3816 1272 3832 1288
rect 5000 1272 5016 1288
rect 5304 1272 5320 1288
rect 168 1232 184 1248
rect 376 1232 392 1248
rect 408 1232 424 1248
rect 1000 1232 1016 1248
rect 1368 1232 1384 1248
rect 1560 1232 1576 1248
rect 2184 1232 2200 1248
rect 2472 1232 2488 1248
rect 2936 1232 2952 1248
rect 3016 1232 3032 1248
rect 4648 1232 4664 1248
rect 4968 1232 4984 1248
rect 5368 1232 5384 1248
rect 797 1202 833 1218
rect 2861 1202 2897 1218
rect 4909 1202 4945 1218
rect 40 1172 56 1188
rect 776 1172 792 1188
rect 1272 1172 1288 1188
rect 1368 1172 1384 1188
rect 1432 1172 1448 1188
rect 2040 1172 2056 1188
rect 2168 1172 2184 1188
rect 3048 1172 3064 1188
rect 3432 1172 3448 1188
rect 3624 1172 3640 1188
rect 3944 1172 3960 1188
rect 3992 1172 4008 1188
rect 4600 1172 4616 1188
rect 5064 1172 5080 1188
rect 5208 1172 5224 1188
rect 5752 1172 5768 1188
rect 5928 1172 5944 1188
rect 3176 1152 3192 1168
rect 40 1132 56 1148
rect 232 1132 248 1148
rect 1000 1132 1016 1148
rect 1448 1132 1464 1148
rect 1688 1132 1704 1148
rect 2328 1132 2344 1148
rect 3160 1132 3176 1148
rect 3832 1132 3848 1148
rect 4856 1132 4872 1148
rect 5080 1132 5096 1148
rect 5448 1132 5464 1148
rect 5768 1132 5784 1148
rect 5800 1132 5816 1148
rect 6232 1132 6248 1148
rect 56 1112 72 1128
rect 88 1112 104 1128
rect 152 1112 168 1128
rect 216 1112 232 1128
rect 264 1112 280 1128
rect 328 1112 344 1128
rect 40 1092 56 1108
rect 72 1092 88 1108
rect 136 1092 152 1108
rect 184 1092 200 1108
rect 280 1092 328 1108
rect 360 1092 376 1108
rect 424 1092 456 1108
rect 472 1092 488 1108
rect 568 1092 584 1108
rect 616 1092 632 1108
rect 680 1112 696 1128
rect 888 1112 904 1128
rect 1032 1112 1048 1128
rect 1304 1112 1320 1128
rect 1528 1112 1544 1128
rect 1656 1112 1672 1128
rect 2456 1112 2472 1128
rect 2664 1112 2680 1128
rect 728 1092 760 1108
rect 856 1092 872 1108
rect 968 1092 984 1108
rect 1016 1092 1032 1108
rect 1112 1092 1128 1108
rect 1160 1092 1176 1108
rect 1304 1092 1320 1108
rect 1336 1092 1352 1108
rect 1368 1092 1384 1108
rect 1464 1092 1480 1108
rect 1496 1092 1512 1108
rect 1544 1092 1576 1108
rect 88 1072 104 1088
rect 120 1072 152 1088
rect 200 1072 216 1088
rect 248 1072 264 1088
rect 312 1072 328 1088
rect 376 1072 392 1088
rect 424 1072 440 1088
rect 488 1072 504 1088
rect 568 1072 584 1088
rect 632 1072 648 1088
rect 728 1072 744 1088
rect 904 1072 920 1088
rect 968 1072 984 1088
rect 1288 1072 1304 1088
rect 1320 1072 1336 1088
rect 1352 1072 1368 1088
rect 1416 1072 1432 1088
rect 1464 1072 1480 1088
rect 1576 1072 1592 1088
rect 1640 1092 1656 1108
rect 1672 1092 1688 1108
rect 1704 1092 1720 1108
rect 1768 1090 1784 1106
rect 1832 1092 1848 1108
rect 1944 1092 1960 1108
rect 1976 1092 1992 1108
rect 2024 1092 2040 1108
rect 2072 1092 2104 1108
rect 2200 1092 2232 1108
rect 2360 1092 2376 1108
rect 2408 1092 2424 1108
rect 2488 1092 2504 1108
rect 2568 1092 2584 1108
rect 2632 1092 2648 1108
rect 2760 1112 2792 1128
rect 2872 1112 2888 1128
rect 3016 1112 3032 1128
rect 3192 1112 3208 1128
rect 3688 1112 3704 1128
rect 2712 1092 2728 1108
rect 2840 1092 2872 1108
rect 2904 1092 2920 1108
rect 2952 1092 2968 1108
rect 2984 1092 3000 1108
rect 3048 1092 3064 1108
rect 3080 1092 3096 1108
rect 3176 1092 3192 1108
rect 3288 1092 3304 1108
rect 3432 1092 3448 1108
rect 3512 1092 3528 1108
rect 3656 1092 3672 1108
rect 4040 1112 4056 1128
rect 4152 1112 4168 1128
rect 4248 1112 4264 1128
rect 4296 1112 4312 1128
rect 4328 1112 4344 1128
rect 4360 1112 4376 1128
rect 4952 1112 4968 1128
rect 4988 1112 5004 1128
rect 5128 1112 5144 1128
rect 5304 1112 5320 1128
rect 5400 1112 5416 1128
rect 5480 1112 5496 1128
rect 3752 1092 3768 1108
rect 3864 1092 3880 1108
rect 4024 1092 4040 1108
rect 4120 1092 4136 1108
rect 4232 1092 4248 1108
rect 4328 1092 4344 1108
rect 4424 1090 4440 1106
rect 4568 1092 4584 1108
rect 4632 1092 4648 1108
rect 4760 1092 4776 1108
rect 4808 1092 4824 1108
rect 4856 1092 4888 1108
rect 5080 1092 5096 1108
rect 5176 1092 5192 1108
rect 5240 1092 5256 1108
rect 5336 1092 5352 1108
rect 5416 1092 5432 1108
rect 5544 1092 5560 1108
rect 5592 1112 5608 1128
rect 5672 1112 5688 1128
rect 5736 1112 5752 1128
rect 5848 1112 5864 1128
rect 5976 1112 5992 1128
rect 6312 1112 6328 1128
rect 6360 1112 6376 1128
rect 6440 1112 6456 1128
rect 6600 1112 6616 1128
rect 5624 1092 5640 1108
rect 5656 1092 5672 1108
rect 5720 1092 5736 1108
rect 5752 1092 5768 1108
rect 5800 1092 5816 1108
rect 5880 1092 5896 1108
rect 6168 1092 6184 1108
rect 6200 1092 6216 1108
rect 6280 1092 6296 1108
rect 6328 1092 6344 1108
rect 6392 1092 6408 1108
rect 6472 1092 6488 1108
rect 6552 1092 6568 1108
rect 6632 1092 6648 1108
rect 6664 1092 6680 1108
rect 1960 1072 1976 1088
rect 1992 1072 2008 1088
rect 2280 1072 2296 1088
rect 2392 1072 2408 1088
rect 2504 1072 2520 1088
rect 2536 1072 2552 1088
rect 2632 1072 2648 1088
rect 2664 1072 2680 1088
rect 2824 1072 2840 1088
rect 2920 1072 2952 1088
rect 3000 1072 3016 1088
rect 3064 1072 3080 1088
rect 3640 1072 3656 1088
rect 3736 1072 3752 1088
rect 3800 1072 3816 1088
rect 4088 1072 4104 1088
rect 4200 1072 4216 1088
rect 4264 1072 4280 1088
rect 4392 1072 4408 1088
rect 4952 1072 4968 1088
rect 5016 1072 5032 1088
rect 5160 1072 5176 1088
rect 5288 1072 5304 1088
rect 5352 1072 5384 1088
rect 5528 1072 5544 1088
rect 5640 1072 5672 1088
rect 5704 1072 5720 1088
rect 5880 1072 5896 1088
rect 6024 1072 6056 1088
rect 6216 1072 6232 1088
rect 6264 1072 6280 1088
rect 6328 1072 6344 1088
rect 6456 1072 6472 1088
rect 6488 1072 6504 1088
rect 6536 1072 6552 1088
rect 392 1052 408 1068
rect 1400 1052 1416 1068
rect 2744 1052 2760 1068
rect 2776 1052 2792 1068
rect 2984 1052 3000 1068
rect 3336 1052 3352 1068
rect 3400 1052 3416 1068
rect 3496 1052 3512 1068
rect 4168 1052 4184 1068
rect 4488 1052 4504 1068
rect 4824 1052 4840 1068
rect 5048 1052 5064 1068
rect 5384 1052 5400 1068
rect 5832 1052 5848 1068
rect 6120 1052 6136 1068
rect 6200 1052 6216 1068
rect 6248 1052 6264 1068
rect 6504 1052 6520 1068
rect 6696 1052 6712 1068
rect 472 1032 488 1048
rect 648 1032 664 1048
rect 936 1032 952 1048
rect 1000 1032 1016 1048
rect 1224 1032 1240 1048
rect 1896 1032 1912 1048
rect 2120 1032 2136 1048
rect 2168 1032 2184 1048
rect 2248 1032 2264 1048
rect 2504 1032 2520 1048
rect 2584 1032 2600 1048
rect 3112 1032 3128 1048
rect 3208 1032 3224 1048
rect 3720 1032 3736 1048
rect 4040 1032 4056 1048
rect 4664 1032 4680 1048
rect 4712 1032 4728 1048
rect 4776 1032 4792 1048
rect 4904 1032 4920 1048
rect 5208 1032 5224 1048
rect 5272 1032 5288 1048
rect 5480 1032 5496 1048
rect 5576 1032 5592 1048
rect 5864 1032 5880 1048
rect 5928 1032 5944 1048
rect 5992 1032 6008 1048
rect 6056 1032 6072 1048
rect 6424 1032 6440 1048
rect 6520 1032 6536 1048
rect 1837 1002 1873 1018
rect 3885 1002 3921 1018
rect 5933 1002 5969 1018
rect 56 972 72 988
rect 584 972 600 988
rect 1160 972 1176 988
rect 1224 972 1240 988
rect 1272 972 1288 988
rect 1528 972 1544 988
rect 1608 972 1624 988
rect 1768 972 1784 988
rect 2136 972 2152 988
rect 2744 972 2760 988
rect 3000 972 3016 988
rect 3128 972 3144 988
rect 3192 972 3208 988
rect 3336 972 3352 988
rect 4184 972 4200 988
rect 4296 972 4312 988
rect 4488 972 4504 988
rect 4632 972 4648 988
rect 4760 972 4776 988
rect 4936 972 4952 988
rect 5080 972 5096 988
rect 5784 972 5800 988
rect 5944 972 5960 988
rect 8 952 24 968
rect 2312 952 2328 968
rect 2344 952 2360 968
rect 2440 952 2456 968
rect 2616 952 2632 968
rect 2680 952 2696 968
rect 3288 952 3304 968
rect 4072 952 4088 968
rect 4376 952 4392 968
rect 4440 952 4472 968
rect 4840 952 4856 968
rect 5000 952 5032 968
rect 5064 952 5080 968
rect 5304 952 5320 968
rect 5496 952 5512 968
rect 6600 952 6616 968
rect 72 932 104 948
rect 136 932 152 948
rect 184 932 216 948
rect 280 932 296 948
rect 312 932 328 948
rect 392 932 408 948
rect 664 932 680 948
rect 760 932 776 948
rect 792 932 824 948
rect 840 932 856 948
rect 872 932 888 948
rect 168 912 184 928
rect 216 912 232 928
rect 264 912 280 928
rect 376 912 392 928
rect 504 912 536 928
rect 600 912 616 928
rect 632 912 648 928
rect 40 892 56 908
rect 136 892 152 908
rect 228 892 244 908
rect 248 892 264 908
rect 344 892 360 908
rect 648 892 664 908
rect 744 912 760 928
rect 776 912 792 928
rect 920 912 936 928
rect 952 932 968 948
rect 1064 932 1080 948
rect 1128 932 1144 948
rect 1208 932 1224 948
rect 1384 932 1400 948
rect 1432 932 1464 948
rect 1544 932 1560 948
rect 1576 932 1592 948
rect 1608 932 1624 948
rect 1688 932 1704 948
rect 1752 932 1768 948
rect 1800 932 1816 948
rect 1880 932 1912 948
rect 2120 932 2136 948
rect 2152 932 2168 948
rect 2264 932 2280 948
rect 2408 932 2424 948
rect 2552 932 2568 948
rect 2824 932 2840 948
rect 2920 932 2936 948
rect 3016 932 3048 948
rect 3096 932 3112 948
rect 3144 932 3160 948
rect 3176 932 3192 948
rect 3272 932 3288 948
rect 3320 932 3336 948
rect 3384 932 3416 948
rect 3464 932 3480 948
rect 3560 932 3576 948
rect 3624 932 3640 948
rect 3816 932 3832 948
rect 3976 932 3992 948
rect 4008 932 4024 948
rect 4056 932 4072 948
rect 4088 932 4104 948
rect 4120 932 4136 948
rect 4232 932 4248 948
rect 4264 932 4280 948
rect 4312 932 4344 948
rect 4472 932 4488 948
rect 4536 932 4552 948
rect 4600 932 4616 948
rect 4680 932 4696 948
rect 4856 932 4872 948
rect 4920 932 4936 948
rect 4968 932 4984 948
rect 5032 932 5048 948
rect 5176 932 5192 948
rect 5320 932 5336 948
rect 5368 932 5400 948
rect 968 912 1000 928
rect 1064 912 1096 928
rect 1112 912 1128 928
rect 1192 912 1208 928
rect 1304 912 1320 928
rect 1368 912 1384 928
rect 1400 912 1416 928
rect 1464 912 1480 928
rect 712 892 728 908
rect 888 892 904 908
rect 1016 892 1032 908
rect 1036 892 1052 908
rect 1080 892 1096 908
rect 1240 892 1256 908
rect 1432 892 1448 908
rect 1496 892 1512 908
rect 1544 912 1576 928
rect 1672 912 1688 928
rect 1736 912 1752 928
rect 1848 912 1864 928
rect 1960 914 1976 930
rect 2024 912 2040 928
rect 2104 912 2120 928
rect 2168 912 2200 928
rect 2344 912 2360 928
rect 2376 912 2392 928
rect 2488 912 2504 928
rect 2616 914 2632 930
rect 2760 912 2776 928
rect 2824 912 2856 928
rect 2920 912 2952 928
rect 1640 892 1656 908
rect 1704 892 1720 908
rect 1724 892 1740 908
rect 1768 892 1784 908
rect 2056 892 2072 908
rect 2360 892 2376 908
rect 2472 892 2488 908
rect 2520 892 2536 908
rect 2872 892 2888 908
rect 2968 892 2984 908
rect 3048 912 3064 928
rect 3160 912 3176 928
rect 3080 892 3096 908
rect 3256 912 3272 928
rect 3304 912 3320 928
rect 3336 912 3352 928
rect 3368 912 3384 928
rect 3400 912 3416 928
rect 3432 912 3448 928
rect 3512 912 3528 928
rect 3640 912 3672 928
rect 3688 912 3704 928
rect 3720 912 3736 928
rect 3816 912 3832 928
rect 3976 912 3992 928
rect 4024 912 4040 928
rect 4104 912 4120 928
rect 4136 912 4168 928
rect 4216 912 4232 928
rect 4248 912 4264 928
rect 4312 912 4328 928
rect 3224 892 3240 908
rect 3496 892 3512 908
rect 3592 892 3624 908
rect 3672 892 3688 908
rect 3736 892 3752 908
rect 4024 892 4040 908
rect 4168 892 4184 908
rect 4360 892 4376 908
rect 4408 912 4424 928
rect 4488 912 4504 928
rect 4520 912 4536 928
rect 4568 912 4600 928
rect 4696 912 4712 928
rect 4792 912 4808 928
rect 4872 912 4888 928
rect 5048 912 5064 928
rect 5112 912 5128 928
rect 5160 912 5176 928
rect 5192 912 5224 928
rect 5256 912 5272 928
rect 5336 912 5352 928
rect 5400 912 5416 928
rect 5512 932 5528 948
rect 5576 932 5592 948
rect 5640 932 5656 948
rect 5704 932 5720 948
rect 5752 932 5768 948
rect 5816 932 5832 948
rect 5848 932 5864 948
rect 5928 932 5944 948
rect 5992 944 6024 948
rect 5976 932 6024 944
rect 6104 932 6120 948
rect 6248 932 6264 948
rect 6328 932 6344 948
rect 6376 932 6392 948
rect 6408 932 6424 948
rect 6472 932 6488 948
rect 6504 932 6520 948
rect 6536 932 6552 948
rect 6584 932 6600 948
rect 6696 932 6712 948
rect 5976 928 5992 932
rect 5464 912 5480 928
rect 5528 912 5544 928
rect 5592 912 5640 928
rect 4552 892 4568 908
rect 4760 892 4776 908
rect 4984 892 5000 908
rect 5128 892 5144 908
rect 5240 892 5256 908
rect 5368 892 5384 908
rect 5496 892 5512 908
rect 5560 892 5576 908
rect 5624 892 5640 908
rect 5688 892 5704 908
rect 5736 912 5752 928
rect 5848 912 5880 928
rect 6008 912 6024 928
rect 5896 892 5912 908
rect 6184 912 6200 928
rect 6232 912 6248 928
rect 6264 912 6280 928
rect 6072 892 6088 908
rect 6296 892 6312 908
rect 6360 912 6376 928
rect 6424 912 6440 928
rect 6472 912 6488 928
rect 6552 912 6568 928
rect 6680 912 6696 928
rect 6408 892 6424 908
rect 6456 892 6472 908
rect 6520 892 6536 908
rect 6584 892 6600 908
rect 120 872 136 888
rect 2088 872 2104 888
rect 2712 872 2728 888
rect 3704 872 3720 888
rect 3896 872 3912 888
rect 3928 872 3944 888
rect 6200 872 6216 888
rect 2488 852 2504 868
rect 2792 852 2808 868
rect 24 832 40 848
rect 104 832 120 848
rect 312 832 328 848
rect 1160 832 1176 848
rect 1272 832 1288 848
rect 1336 832 1352 848
rect 1880 832 1896 848
rect 2216 832 2232 848
rect 2344 832 2360 848
rect 3544 832 3560 848
rect 4632 832 4648 848
rect 4728 832 4744 848
rect 5304 832 5320 848
rect 5528 832 5544 848
rect 6024 832 6040 848
rect 6136 832 6152 848
rect 6440 832 6456 848
rect 797 802 833 818
rect 2861 802 2897 818
rect 4909 802 4945 818
rect 392 772 408 788
rect 1288 772 1304 788
rect 1352 772 1368 788
rect 1448 772 1464 788
rect 1576 772 1592 788
rect 1960 772 1976 788
rect 3016 772 3032 788
rect 3352 772 3368 788
rect 4616 772 4632 788
rect 5192 772 5208 788
rect 6056 772 6072 788
rect 6312 772 6328 788
rect 8 732 24 748
rect 184 732 200 748
rect 440 732 456 748
rect 872 732 888 748
rect 952 732 1000 748
rect 1032 732 1048 748
rect 1720 732 1736 748
rect 1944 732 1960 748
rect 2024 732 2040 748
rect 2328 732 2344 748
rect 3288 732 3304 748
rect 3768 732 3784 748
rect 4120 732 4136 748
rect 4712 732 4728 748
rect 4904 732 4920 748
rect 5576 732 5592 748
rect 6040 732 6056 748
rect 152 712 168 728
rect 40 692 56 708
rect 136 692 152 708
rect 168 692 184 708
rect 200 692 216 708
rect 264 690 280 706
rect 328 692 344 708
rect 440 692 456 708
rect 520 712 536 728
rect 568 692 584 708
rect 632 712 648 728
rect 936 712 952 728
rect 1192 712 1208 728
rect 1256 712 1272 728
rect 1496 712 1512 728
rect 1764 712 1780 728
rect 1784 712 1800 728
rect 1848 712 1864 728
rect 664 692 680 708
rect 792 692 808 708
rect 1000 692 1016 708
rect 1080 692 1096 708
rect 1112 692 1128 708
rect 1160 692 1176 708
rect 1208 692 1240 708
rect 1288 692 1304 708
rect 1336 692 1352 708
rect 1368 692 1384 708
rect 1400 692 1416 708
rect 1480 692 1496 708
rect 1528 692 1544 708
rect 1624 692 1640 708
rect 1752 692 1768 708
rect 1816 692 1832 708
rect 2056 712 2072 728
rect 1960 692 1976 708
rect 2008 692 2024 708
rect 2216 712 2232 728
rect 2088 692 2120 708
rect 2136 692 2152 708
rect 2200 692 2216 708
rect 2296 692 2312 708
rect 2376 692 2392 708
rect 2424 712 2440 728
rect 2648 712 2664 728
rect 2744 712 2760 728
rect 2776 712 2792 728
rect 2920 712 2936 728
rect 2472 692 2488 708
rect 2584 692 2600 708
rect 2616 692 2632 708
rect 2728 692 2744 708
rect 2824 692 2840 708
rect 3064 712 3080 728
rect 3208 712 3224 728
rect 3240 712 3256 728
rect 3272 712 3288 728
rect 3688 712 3704 728
rect 4104 712 4120 728
rect 4152 712 4168 728
rect 4216 712 4232 728
rect 4344 712 4360 728
rect 4408 712 4424 728
rect 4500 712 4516 728
rect 4520 712 4536 728
rect 4632 712 4648 728
rect 4744 712 4760 728
rect 4808 712 4824 728
rect 4920 712 4952 728
rect 5096 712 5112 728
rect 5256 712 5288 728
rect 5400 712 5416 728
rect 2968 692 2984 708
rect 3064 692 3096 708
rect 3144 692 3176 708
rect 3192 692 3208 708
rect 3224 692 3240 708
rect 3320 692 3336 708
rect 3384 692 3400 708
rect 3416 692 3432 708
rect 3528 692 3560 708
rect 3624 692 3640 708
rect 3720 692 3736 708
rect 3768 692 3784 708
rect 4008 692 4024 708
rect 4168 692 4200 708
rect 4248 692 4264 708
rect 4280 692 4296 708
rect 4376 692 4392 708
rect 4440 692 4456 708
rect 4488 692 4504 708
rect 4520 692 4536 708
rect 4568 692 4584 708
rect 4680 692 4696 708
rect 4776 692 4792 708
rect 4824 692 4840 708
rect 4920 692 4936 708
rect 5000 692 5016 708
rect 56 672 72 688
rect 456 672 504 688
rect 568 672 600 688
rect 680 672 696 688
rect 712 672 728 688
rect 920 672 936 688
rect 1064 672 1080 688
rect 1096 672 1112 688
rect 1144 672 1160 688
rect 1176 672 1192 688
rect 1240 672 1256 688
rect 1304 672 1336 688
rect 1384 672 1400 688
rect 1544 672 1560 688
rect 1672 672 1704 688
rect 1736 672 1752 688
rect 1800 672 1816 688
rect 1928 672 1944 688
rect 2008 672 2024 688
rect 2120 672 2152 688
rect 2184 672 2200 688
rect 2248 672 2264 688
rect 2312 672 2328 688
rect 2392 672 2408 688
rect 2456 672 2472 688
rect 2600 672 2616 688
rect 2680 672 2696 688
rect 2712 672 2728 688
rect 2776 672 2792 688
rect 2840 672 2856 688
rect 2888 672 2904 688
rect 2936 672 2952 688
rect 3032 672 3048 688
rect 3096 672 3112 688
rect 3128 672 3144 688
rect 3160 672 3176 688
rect 3224 672 3240 688
rect 3448 672 3464 688
rect 3672 672 3688 688
rect 3736 672 3768 688
rect 3880 672 3912 688
rect 4008 672 4024 688
rect 4104 672 4120 688
rect 4136 672 4152 688
rect 4264 672 4280 688
rect 4296 672 4312 688
rect 4392 672 4424 688
rect 4456 672 4488 688
rect 4584 672 4616 688
rect 4664 672 4712 688
rect 4760 672 4776 688
rect 4888 672 4904 688
rect 5064 692 5080 708
rect 5144 692 5176 708
rect 5304 692 5320 708
rect 5352 692 5368 708
rect 5416 692 5432 708
rect 5448 692 5480 708
rect 5528 712 5544 728
rect 5688 712 5704 728
rect 5752 712 5768 728
rect 5880 712 5896 728
rect 5944 712 5960 728
rect 6296 712 6312 728
rect 6504 712 6520 728
rect 6568 712 6584 728
rect 5624 692 5656 708
rect 5720 692 5752 708
rect 5784 692 5800 708
rect 5080 672 5096 688
rect 5144 672 5160 688
rect 5208 672 5224 688
rect 5320 672 5352 688
rect 5400 672 5416 688
rect 5464 672 5480 688
rect 5560 672 5576 688
rect 5608 672 5624 688
rect 5640 672 5656 688
rect 5704 672 5720 688
rect 5768 672 5784 688
rect 5848 692 5864 708
rect 5912 692 5928 708
rect 5992 692 6008 708
rect 6120 692 6152 708
rect 6264 692 6280 708
rect 6376 692 6408 708
rect 6536 692 6552 708
rect 6600 692 6616 708
rect 6648 692 6664 708
rect 6696 712 6712 728
rect 6728 692 6744 708
rect 5896 672 5912 688
rect 6248 672 6264 688
rect 6296 672 6312 688
rect 6472 672 6488 688
rect 6552 672 6568 688
rect 6616 672 6648 688
rect 6664 672 6680 688
rect 6744 672 6760 688
rect 104 652 120 668
rect 1160 652 1176 668
rect 1416 652 1432 668
rect 2152 652 2168 668
rect 2328 652 2344 668
rect 3000 652 3016 668
rect 3416 652 3432 668
rect 3864 652 3880 668
rect 4312 652 4344 668
rect 4872 652 4888 668
rect 5240 652 5256 668
rect 5512 652 5528 668
rect 5576 652 5592 668
rect 6040 652 6056 668
rect 600 632 616 648
rect 1496 632 1512 648
rect 1720 632 1736 648
rect 2216 632 2232 648
rect 2264 632 2280 648
rect 2504 632 2520 648
rect 2552 632 2568 648
rect 2696 632 2712 648
rect 2744 632 2760 648
rect 2792 632 2808 648
rect 3048 632 3064 648
rect 3112 632 3128 648
rect 3304 632 3320 648
rect 3608 632 3624 648
rect 3656 632 3672 648
rect 4344 632 4360 648
rect 4856 632 4872 648
rect 5096 632 5112 648
rect 5272 632 5288 648
rect 5384 632 5400 648
rect 5688 632 5704 648
rect 5880 632 5896 648
rect 6312 632 6328 648
rect 6504 632 6520 648
rect 6568 632 6584 648
rect 1837 602 1873 618
rect 3885 602 3921 618
rect 5933 602 5969 618
rect 744 572 760 588
rect 984 572 1000 588
rect 1080 572 1096 588
rect 1304 572 1320 588
rect 2360 572 2376 588
rect 2616 572 2632 588
rect 2904 572 2920 588
rect 3624 572 3640 588
rect 4072 572 4088 588
rect 4424 572 4440 588
rect 4664 572 4680 588
rect 4808 572 4824 588
rect 5080 572 5096 588
rect 5144 572 5160 588
rect 5224 572 5240 588
rect 5448 572 5464 588
rect 5912 572 5928 588
rect 6184 572 6200 588
rect 6408 572 6424 588
rect 6536 572 6552 588
rect 6728 572 6744 588
rect 56 552 88 568
rect 136 552 152 568
rect 1384 552 1400 568
rect 1928 552 1944 568
rect 2312 552 2328 568
rect 2632 552 2648 568
rect 2760 552 2776 568
rect 3000 552 3016 568
rect 3928 552 3944 568
rect 4264 552 4280 568
rect 4472 552 4488 568
rect 4712 552 4728 568
rect 5000 552 5016 568
rect 5672 552 5688 568
rect 5816 552 5832 568
rect 6424 552 6440 568
rect 6808 552 6824 568
rect 4744 548 4760 550
rect 8 532 24 548
rect 88 532 104 548
rect 184 532 200 548
rect 280 532 296 548
rect 376 532 424 548
rect 488 532 504 548
rect 552 532 568 548
rect 616 532 632 548
rect 776 532 792 548
rect 840 532 856 548
rect 936 532 952 548
rect 1016 532 1048 548
rect 1144 532 1160 548
rect 1176 532 1192 548
rect 1208 532 1224 548
rect 1288 532 1304 548
rect 1416 532 1432 548
rect 1512 532 1528 548
rect 1688 532 1704 548
rect 1800 532 1816 548
rect 2008 532 2024 548
rect 2056 532 2072 548
rect 2152 532 2168 548
rect 2184 532 2200 548
rect 2232 532 2248 548
rect 2296 532 2312 548
rect 2408 532 2424 548
rect 2456 532 2472 548
rect 2488 532 2504 548
rect 40 512 56 528
rect 168 512 216 528
rect 232 492 248 508
rect 312 512 328 528
rect 360 512 376 528
rect 472 512 504 528
rect 536 512 552 528
rect 664 512 680 528
rect 856 512 872 528
rect 904 512 920 528
rect 1016 512 1032 528
rect 1080 512 1096 528
rect 1128 512 1144 528
rect 1192 512 1208 528
rect 1256 512 1272 528
rect 1352 512 1368 528
rect 440 492 456 508
rect 504 492 520 508
rect 808 492 824 508
rect 920 492 936 508
rect 968 492 984 508
rect 1096 492 1112 508
rect 1160 492 1176 508
rect 1224 492 1240 508
rect 1496 512 1512 528
rect 1608 512 1624 528
rect 1816 512 1832 528
rect 1944 512 1960 528
rect 1976 512 1992 528
rect 2136 512 2152 528
rect 2168 512 2184 528
rect 2280 512 2296 528
rect 2344 512 2360 528
rect 2392 512 2408 528
rect 2424 512 2440 528
rect 2504 512 2520 528
rect 2600 532 2616 548
rect 3096 532 3112 548
rect 3192 532 3208 548
rect 2568 512 2584 528
rect 2648 512 2664 528
rect 2680 512 2696 528
rect 2760 514 2776 530
rect 3064 514 3080 530
rect 3144 512 3160 528
rect 3208 512 3224 528
rect 3336 532 3352 548
rect 3512 532 3528 548
rect 3576 532 3592 548
rect 3640 532 3656 548
rect 3672 532 3688 548
rect 3752 532 3768 548
rect 3784 532 3800 548
rect 3848 532 3880 548
rect 3944 532 3960 548
rect 3976 532 3992 548
rect 4040 532 4072 548
rect 4088 532 4104 548
rect 4120 532 4136 548
rect 4168 532 4200 548
rect 4232 532 4248 548
rect 4264 532 4280 548
rect 4296 532 4312 548
rect 4408 532 4424 548
rect 4440 532 4456 548
rect 4504 532 4520 548
rect 4552 532 4568 548
rect 4584 532 4600 548
rect 4728 534 4760 548
rect 4728 532 4744 534
rect 4792 532 4808 548
rect 4840 532 4856 548
rect 4904 532 4920 548
rect 4984 532 5000 548
rect 5016 532 5032 548
rect 5048 532 5064 548
rect 5112 532 5128 548
rect 5144 532 5160 548
rect 5192 532 5208 548
rect 5336 532 5352 548
rect 5528 532 5544 548
rect 5640 532 5672 548
rect 5688 532 5704 548
rect 5768 532 5784 548
rect 5816 532 5832 548
rect 5880 532 5896 548
rect 6024 532 6040 548
rect 6120 532 6136 548
rect 6232 532 6264 548
rect 6312 532 6328 548
rect 6424 532 6440 548
rect 6568 532 6584 548
rect 3272 512 3288 528
rect 3416 512 3448 528
rect 3528 512 3544 528
rect 3656 512 3672 528
rect 3688 512 3720 528
rect 3768 512 3800 528
rect 3832 512 3848 528
rect 3896 512 3912 528
rect 3960 512 3976 528
rect 3992 512 4008 528
rect 4040 512 4056 528
rect 4104 512 4120 528
rect 4152 512 4184 528
rect 4248 512 4264 528
rect 4312 512 4344 528
rect 4392 512 4408 528
rect 4456 512 4472 528
rect 4520 512 4552 528
rect 4568 512 4584 528
rect 4600 512 4616 528
rect 4632 512 4648 528
rect 4680 512 4696 528
rect 4744 512 4760 528
rect 4776 512 4792 528
rect 4872 512 4888 528
rect 4904 512 4920 528
rect 5032 512 5048 528
rect 5128 512 5144 528
rect 5192 512 5208 528
rect 5256 512 5272 528
rect 5352 512 5368 528
rect 5512 512 5528 528
rect 5544 512 5560 528
rect 1464 492 1480 508
rect 1960 492 1976 508
rect 1992 492 2024 508
rect 2104 492 2120 508
rect 2136 492 2152 508
rect 2184 492 2200 508
rect 2248 492 2264 508
rect 2600 492 2616 508
rect 2664 492 2680 508
rect 2696 492 2712 508
rect 3144 492 3176 508
rect 3284 492 3300 508
rect 3304 492 3320 508
rect 3560 492 3576 508
rect 3720 492 3752 508
rect 3800 492 3816 508
rect 4024 492 4040 508
rect 4120 492 4136 508
rect 4616 492 4632 508
rect 4808 492 4824 508
rect 4856 492 4872 508
rect 5064 492 5096 508
rect 5576 492 5592 508
rect 5656 512 5672 528
rect 5704 512 5736 528
rect 5768 512 5784 528
rect 5800 512 5816 528
rect 5864 512 5880 528
rect 6008 512 6024 528
rect 6136 512 6152 528
rect 5624 492 5640 508
rect 5688 492 5704 508
rect 5732 492 5748 508
rect 5752 492 5768 508
rect 5832 492 5848 508
rect 6168 492 6184 508
rect 6216 512 6248 528
rect 6280 512 6296 528
rect 6328 512 6344 528
rect 6376 512 6392 528
rect 6504 512 6520 528
rect 6616 512 6632 528
rect 6296 492 6312 508
rect 6360 492 6376 508
rect 6472 492 6488 508
rect 328 472 344 488
rect 712 472 728 488
rect 984 472 1000 488
rect 1992 472 2008 488
rect 3496 472 3512 488
rect 4200 472 4216 488
rect 4648 472 4664 488
rect 4680 472 4696 488
rect 5480 472 5496 488
rect 872 452 888 468
rect 1256 452 1272 468
rect 2344 452 2360 468
rect 3144 452 3160 468
rect 312 432 328 448
rect 1432 432 1448 448
rect 1528 432 1544 448
rect 4360 432 4376 448
rect 4472 432 4488 448
rect 4952 432 4968 448
rect 6744 432 6760 448
rect 797 402 833 418
rect 2861 402 2897 418
rect 4909 402 4945 418
rect 56 372 72 388
rect 88 372 104 388
rect 1496 372 1512 388
rect 2232 372 2248 388
rect 2664 372 2680 388
rect 4232 372 4248 388
rect 4520 372 4536 388
rect 4776 372 4792 388
rect 5592 372 5608 388
rect 5848 372 5864 388
rect 6696 372 6712 388
rect 6760 372 6776 388
rect 4248 352 4264 368
rect 5128 352 5144 368
rect 5768 352 5784 368
rect 488 332 504 348
rect 2488 332 2504 348
rect 4200 332 4216 348
rect 4744 332 4760 348
rect 4904 332 4920 348
rect 5736 332 5752 348
rect 6168 332 6184 348
rect 6440 332 6456 348
rect 6680 332 6696 348
rect 280 312 296 328
rect 424 312 440 328
rect 536 312 552 328
rect 600 312 616 328
rect 696 312 712 328
rect 200 292 216 308
rect 296 292 328 308
rect 344 292 360 308
rect 408 292 424 308
rect 440 292 456 308
rect 472 292 488 308
rect 568 292 600 308
rect 648 292 664 308
rect 712 292 728 308
rect 744 292 760 308
rect 776 312 792 328
rect 920 312 936 328
rect 808 292 824 308
rect 888 292 904 308
rect 1032 312 1048 328
rect 1000 292 1016 308
rect 1112 292 1128 308
rect 1240 312 1256 328
rect 1384 312 1400 328
rect 1160 292 1176 308
rect 1208 292 1224 308
rect 1288 292 1304 308
rect 1320 292 1352 308
rect 1432 312 1448 328
rect 1704 312 1720 328
rect 1992 312 2008 328
rect 2152 312 2168 328
rect 2276 312 2292 328
rect 2296 312 2312 328
rect 2344 312 2360 328
rect 2364 312 2380 328
rect 2436 312 2452 328
rect 2456 312 2472 328
rect 2520 312 2536 328
rect 2952 312 2968 328
rect 1464 292 1480 308
rect 1576 292 1592 308
rect 1624 292 1640 308
rect 1816 292 1832 308
rect 1976 292 1992 308
rect 2024 292 2040 308
rect 8 272 24 288
rect 248 272 264 288
rect 328 272 344 288
rect 360 272 376 288
rect 392 272 408 288
rect 472 272 488 288
rect 520 272 536 288
rect 584 272 600 288
rect 648 272 680 288
rect 712 272 728 288
rect 792 272 808 288
rect 856 272 888 288
rect 968 272 1000 288
rect 1064 272 1080 288
rect 1096 272 1112 288
rect 1176 272 1208 288
rect 1256 272 1272 288
rect 1304 272 1336 288
rect 1432 272 1448 288
rect 1528 272 1544 288
rect 1800 272 1816 288
rect 1928 272 1944 288
rect 2120 292 2136 308
rect 2184 292 2200 308
rect 2264 292 2280 308
rect 2424 292 2440 308
rect 2488 292 2504 308
rect 2568 292 2584 308
rect 2088 288 2104 292
rect 2648 292 2664 308
rect 2712 292 2744 308
rect 2792 292 2808 308
rect 2856 292 2872 308
rect 2920 292 2936 308
rect 2988 312 3004 328
rect 3256 312 3272 328
rect 3320 312 3336 328
rect 3416 312 3432 328
rect 3528 312 3544 328
rect 3672 312 3688 328
rect 3704 312 3720 328
rect 3736 312 3752 328
rect 3800 312 3816 328
rect 3832 312 3848 328
rect 3928 312 3944 328
rect 3992 312 4008 328
rect 4328 312 4344 328
rect 4584 312 4600 328
rect 3016 292 3048 308
rect 3096 292 3128 308
rect 3160 292 3176 308
rect 3192 292 3208 308
rect 3224 292 3240 308
rect 3288 292 3304 308
rect 3336 292 3352 308
rect 3368 292 3384 308
rect 3400 292 3416 308
rect 3432 292 3448 308
rect 3480 292 3512 308
rect 3544 292 3560 308
rect 3608 292 3624 308
rect 3640 292 3656 308
rect 3704 292 3720 308
rect 3752 292 3768 308
rect 3816 292 3832 308
rect 3864 292 3880 308
rect 3960 292 3976 308
rect 4120 292 4136 308
rect 4296 292 4312 308
rect 4440 292 4456 308
rect 4552 292 4568 308
rect 4808 312 4824 328
rect 4920 312 4936 328
rect 5032 312 5064 328
rect 5068 312 5084 328
rect 5240 312 5256 328
rect 4632 292 4648 308
rect 4680 292 4696 308
rect 4760 292 4776 308
rect 4840 292 4856 308
rect 4952 292 4968 308
rect 5000 292 5016 308
rect 5080 292 5112 308
rect 5176 292 5192 308
rect 5208 292 5224 308
rect 5512 312 5528 328
rect 5288 292 5304 308
rect 5320 292 5336 308
rect 5384 292 5400 308
rect 5448 292 5464 308
rect 5480 292 5496 308
rect 5560 312 5576 328
rect 5672 312 5688 328
rect 5576 292 5592 308
rect 5640 292 5656 308
rect 5704 292 5720 308
rect 5912 312 5928 328
rect 6744 312 6760 328
rect 2088 276 2120 288
rect 2104 272 2120 276
rect 2168 272 2184 288
rect 2216 272 2232 288
rect 2248 272 2264 288
rect 2392 272 2424 288
rect 2472 272 2488 288
rect 2584 272 2600 288
rect 2616 272 2648 288
rect 2696 272 2712 288
rect 2744 272 2760 288
rect 2776 272 2792 288
rect 2840 272 2856 288
rect 2904 272 2920 288
rect 3016 272 3032 288
rect 3048 272 3064 288
rect 3080 272 3112 288
rect 3128 272 3144 288
rect 3240 272 3256 288
rect 3272 272 3288 288
rect 3384 272 3400 288
rect 3464 272 3496 288
rect 3592 272 3608 288
rect 3624 272 3640 288
rect 3672 272 3704 288
rect 3752 272 3768 288
rect 3800 272 3816 288
rect 3848 272 3864 288
rect 3976 272 3992 288
rect 4024 272 4040 288
rect 4072 272 4088 288
rect 4280 272 4296 288
rect 4312 272 4328 288
rect 4392 272 4408 288
rect 4536 272 4552 288
rect 4616 272 4632 288
rect 4648 272 4680 288
rect 4760 272 4776 288
rect 4824 272 4840 288
rect 4936 272 4952 288
rect 4968 272 5000 288
rect 5096 272 5112 288
rect 5128 272 5144 288
rect 5160 272 5176 288
rect 5192 272 5208 288
rect 5304 272 5336 288
rect 5368 272 5384 288
rect 5432 272 5480 288
rect 5576 272 5592 288
rect 5624 272 5640 288
rect 5656 272 5672 288
rect 5688 272 5704 288
rect 5720 272 5736 288
rect 5896 292 5912 308
rect 6024 292 6040 308
rect 6088 292 6104 308
rect 6152 292 6168 308
rect 6264 292 6280 308
rect 6440 292 6472 308
rect 6504 292 6520 308
rect 6552 292 6568 308
rect 6648 292 6664 308
rect 6728 292 6744 308
rect 5816 272 5832 288
rect 5944 272 5960 288
rect 6104 272 6120 288
rect 6136 272 6152 288
rect 6344 272 6360 288
rect 2216 252 2232 268
rect 2328 252 2344 268
rect 2808 252 2824 268
rect 3192 252 3208 268
rect 4040 252 4056 268
rect 4264 252 4280 268
rect 4712 252 4728 268
rect 4744 252 4760 268
rect 5400 252 5416 268
rect 5608 252 5624 268
rect 5992 252 6008 268
rect 6136 252 6152 268
rect 6168 252 6184 268
rect 6488 272 6504 288
rect 6632 272 6648 288
rect 6776 272 6792 288
rect 6584 252 6600 268
rect 376 232 392 248
rect 488 232 504 248
rect 536 232 552 248
rect 696 232 712 248
rect 936 232 952 248
rect 1080 232 1096 248
rect 1128 232 1144 248
rect 1688 232 1704 248
rect 1944 232 1960 248
rect 1992 232 2008 248
rect 2552 232 2568 248
rect 2600 232 2616 248
rect 2760 232 2776 248
rect 2824 232 2840 248
rect 3064 232 3080 248
rect 3592 232 3608 248
rect 4872 232 4888 248
rect 5032 232 5048 248
rect 5256 232 5272 248
rect 5352 232 5368 248
rect 6056 232 6072 248
rect 6536 232 6552 248
rect 1837 202 1873 218
rect 3885 202 3921 218
rect 5933 202 5969 218
rect 408 172 424 188
rect 728 172 744 188
rect 776 172 792 188
rect 1640 172 1656 188
rect 1688 172 1704 188
rect 1752 172 1768 188
rect 1816 172 1832 188
rect 2424 172 2440 188
rect 2632 172 2648 188
rect 3048 172 3064 188
rect 3256 172 3272 188
rect 3656 172 3672 188
rect 3848 172 3864 188
rect 4360 172 4392 188
rect 4488 172 4504 188
rect 4520 172 4536 188
rect 4600 172 4616 188
rect 4632 172 4648 188
rect 5176 172 5208 188
rect 5512 172 5528 188
rect 5928 172 5960 188
rect 6024 172 6040 188
rect 6440 172 6456 188
rect 6632 172 6648 188
rect 6712 172 6728 188
rect 104 152 120 168
rect 136 152 152 168
rect 168 152 184 168
rect 248 152 264 168
rect 904 152 920 168
rect 1064 152 1080 168
rect 2152 152 2168 168
rect 2888 152 2904 168
rect 3176 152 3192 168
rect 3288 152 3304 168
rect 3992 152 4008 168
rect 5320 152 5336 168
rect 5448 152 5464 168
rect 5720 152 5736 168
rect 6248 152 6264 168
rect 6504 152 6520 168
rect 8 132 24 148
rect 56 132 72 148
rect 296 132 312 148
rect 424 132 440 148
rect 504 132 520 148
rect 616 132 632 148
rect 1048 132 1064 148
rect 1096 132 1112 148
rect 1160 132 1208 148
rect 1272 132 1288 148
rect 1336 132 1352 148
rect 1384 132 1400 148
rect 1528 132 1544 148
rect 1672 132 1688 148
rect 1704 132 1720 148
rect 1800 132 1816 148
rect 1960 132 1976 148
rect 2024 132 2040 148
rect 2120 132 2136 148
rect 2328 132 2344 148
rect 2360 132 2376 148
rect 2392 132 2408 148
rect 2424 132 2440 148
rect 2456 132 2472 148
rect 2504 132 2520 148
rect 2552 132 2568 148
rect 2616 132 2632 148
rect 2824 132 2840 148
rect 2952 132 2968 148
rect 2984 132 3000 148
rect 3240 132 3256 148
rect 3304 132 3320 148
rect 3400 132 3432 148
rect 3496 132 3512 148
rect 3688 132 3704 148
rect 40 112 56 128
rect 136 112 152 128
rect 184 112 216 128
rect 248 112 264 128
rect 312 112 328 128
rect 472 112 488 128
rect 600 114 616 130
rect 664 112 680 128
rect 904 114 920 130
rect 968 112 984 128
rect 1000 112 1016 128
rect 1032 112 1048 128
rect 1144 112 1160 128
rect 536 92 552 108
rect 1016 92 1032 108
rect 1112 92 1128 108
rect 1256 112 1288 128
rect 1304 112 1336 128
rect 1416 112 1432 128
rect 1448 112 1464 128
rect 1512 114 1528 130
rect 1656 112 1672 128
rect 1720 112 1736 128
rect 1848 112 1864 128
rect 1944 112 1960 128
rect 1992 112 2008 128
rect 2104 112 2120 128
rect 2264 112 2280 128
rect 2344 112 2360 128
rect 2376 112 2392 128
rect 2440 112 2456 128
rect 1224 92 1240 108
rect 1288 92 1304 108
rect 1352 92 1368 108
rect 2232 92 2248 108
rect 2280 92 2296 108
rect 2312 92 2328 108
rect 2488 92 2504 108
rect 2536 112 2568 128
rect 2696 112 2712 128
rect 2744 112 2760 128
rect 2856 112 2872 128
rect 2968 112 2984 128
rect 3000 112 3016 128
rect 3032 112 3048 128
rect 3128 112 3144 128
rect 3400 112 3416 128
rect 3432 112 3448 128
rect 3528 114 3544 130
rect 3720 114 3736 130
rect 3864 112 3880 128
rect 4008 132 4024 148
rect 4072 132 4088 148
rect 4104 132 4136 148
rect 4168 132 4184 148
rect 4200 132 4216 148
rect 4472 132 4488 148
rect 4504 132 4520 148
rect 4616 132 4632 148
rect 4872 132 4904 148
rect 4968 132 4984 148
rect 5432 132 5448 148
rect 5464 132 5480 148
rect 5560 132 5592 148
rect 5624 132 5640 148
rect 5656 132 5672 148
rect 5688 132 5704 148
rect 5768 132 5784 148
rect 5864 132 5880 148
rect 6008 132 6024 148
rect 6072 132 6088 148
rect 6136 132 6152 148
rect 6344 132 6360 148
rect 6680 132 6712 148
rect 4088 112 4104 128
rect 4136 112 4152 128
rect 4248 112 4264 128
rect 4456 112 4472 128
rect 4552 112 4584 128
rect 2824 92 2840 108
rect 3032 92 3048 108
rect 3272 92 3288 108
rect 3384 92 3400 108
rect 3444 92 3460 108
rect 3464 92 3480 108
rect 4168 92 4184 108
rect 4408 92 4424 108
rect 4472 92 4488 108
rect 4696 112 4712 128
rect 4760 114 4776 130
rect 4856 112 4872 128
rect 4920 112 4936 128
rect 4952 112 4968 128
rect 4984 112 5000 128
rect 5064 112 5080 128
rect 5112 112 5128 128
rect 5320 114 5336 130
rect 5400 112 5432 128
rect 5544 112 5560 128
rect 5592 112 5608 128
rect 5624 112 5640 128
rect 5672 112 5688 128
rect 5704 112 5720 128
rect 5800 114 5816 130
rect 6056 112 6072 128
rect 6120 112 6136 128
rect 6168 112 6216 128
rect 6328 112 6344 128
rect 6520 112 6536 128
rect 6648 112 6664 128
rect 4824 92 4840 108
rect 4844 92 4860 108
rect 5384 92 5400 108
rect 5624 92 5640 108
rect 5976 92 5992 108
rect 488 72 504 88
rect 984 72 1000 88
rect 1432 72 1448 88
rect 6072 72 6088 88
rect 472 52 488 68
rect 2264 52 2280 68
rect 344 32 360 48
rect 1880 32 1896 48
rect 3976 32 3992 48
rect 797 2 833 18
rect 2861 2 2897 18
rect 4909 2 4945 18
<< metal2 >>
rect 13 4728 19 4732
rect 56 4697 67 4703
rect 61 4688 67 4697
rect 173 4668 179 4863
rect 221 4828 227 4863
rect 189 4668 195 4812
rect 349 4788 355 4863
rect 397 4828 403 4863
rect 493 4857 515 4863
rect 264 4737 275 4743
rect 269 4708 275 4737
rect 301 4697 312 4703
rect 301 4688 307 4697
rect 365 4668 371 4812
rect 440 4737 451 4743
rect 445 4708 451 4737
rect 477 4697 488 4703
rect 477 4688 483 4697
rect 509 4683 515 4857
rect 525 4857 547 4863
rect 525 4788 531 4857
rect 573 4788 579 4863
rect 621 4737 632 4743
rect 621 4708 627 4737
rect 541 4688 547 4692
rect 493 4677 515 4683
rect 493 4588 499 4677
rect 701 4668 707 4863
rect 781 4688 787 4863
rect 829 4857 851 4863
rect 845 4788 851 4857
rect 893 4688 899 4863
rect 909 4737 920 4743
rect 909 4708 915 4737
rect 957 4688 963 4863
rect 1085 4788 1091 4863
rect 973 4697 984 4703
rect 13 4528 19 4532
rect 61 4523 67 4532
rect 56 4517 67 4523
rect 269 4528 275 4532
rect 237 4488 243 4514
rect 541 4523 547 4532
rect 573 4528 579 4572
rect 536 4517 547 4523
rect 45 4328 51 4332
rect 173 4308 179 4312
rect 88 4297 99 4303
rect 93 4288 99 4297
rect 253 4168 259 4272
rect 13 4028 19 4032
rect 141 3988 147 4114
rect 13 3928 19 3932
rect 56 3897 67 3903
rect 61 3888 67 3897
rect 173 3868 179 3892
rect 61 3748 67 3852
rect 189 3788 195 3892
rect 237 3788 243 3912
rect 269 3888 275 4512
rect 589 4488 595 4532
rect 701 4528 707 4532
rect 605 4368 611 4432
rect 621 4368 627 4472
rect 509 4348 515 4352
rect 429 4268 435 4272
rect 445 4268 451 4292
rect 301 4068 307 4112
rect 317 4048 323 4112
rect 397 4108 403 4232
rect 429 4228 435 4252
rect 445 4123 451 4252
rect 477 4188 483 4312
rect 605 4288 611 4292
rect 653 4288 659 4312
rect 669 4308 675 4372
rect 685 4308 691 4332
rect 717 4328 723 4352
rect 445 4117 456 4123
rect 413 4108 419 4112
rect 381 4028 387 4032
rect 333 3788 339 3932
rect 365 3928 371 4012
rect 365 3908 371 3912
rect 381 3868 387 3872
rect 61 3468 67 3732
rect 109 3508 115 3512
rect 205 3508 211 3732
rect 237 3708 243 3712
rect 269 3668 275 3712
rect 317 3648 323 3732
rect 365 3568 371 3612
rect 45 3328 51 3352
rect 61 3328 67 3452
rect 125 3328 131 3332
rect 141 3328 147 3372
rect 77 3308 83 3312
rect 61 3283 67 3292
rect 61 3277 83 3283
rect 77 3248 83 3277
rect 56 3237 67 3243
rect 61 3106 67 3237
rect 93 3088 99 3312
rect 157 3308 163 3352
rect 189 3188 195 3292
rect 13 2728 19 2732
rect 29 2543 35 2892
rect 93 2708 99 3052
rect 125 3048 131 3092
rect 205 3088 211 3472
rect 237 3468 243 3512
rect 285 3508 291 3512
rect 237 3348 243 3412
rect 221 3188 227 3272
rect 109 2868 115 2912
rect 125 2848 131 2912
rect 189 2888 195 2912
rect 205 2908 211 3072
rect 237 3068 243 3312
rect 253 3128 259 3292
rect 269 2988 275 3392
rect 301 3348 307 3532
rect 349 3488 355 3512
rect 365 3508 371 3552
rect 381 3488 387 3852
rect 413 3828 419 3872
rect 429 3788 435 3892
rect 397 3728 403 3732
rect 413 3728 419 3732
rect 397 3688 403 3712
rect 429 3708 435 3732
rect 445 3568 451 3872
rect 461 3748 467 3872
rect 477 3808 483 3892
rect 493 3888 499 4192
rect 509 4108 515 4172
rect 509 3908 515 4092
rect 525 4088 531 4132
rect 525 3908 531 3972
rect 541 3828 547 4272
rect 605 4248 611 4272
rect 621 4168 627 4272
rect 685 4228 691 4272
rect 589 3988 595 4092
rect 557 3908 563 3912
rect 621 3888 627 4152
rect 733 4128 739 4632
rect 749 4528 755 4572
rect 925 4548 931 4672
rect 973 4528 979 4697
rect 1037 4697 1048 4703
rect 1037 4688 1043 4697
rect 989 4668 995 4672
rect 1005 4528 1011 4532
rect 1069 4508 1075 4514
rect 1101 4488 1107 4672
rect 1133 4588 1139 4712
rect 1181 4608 1187 4692
rect 1197 4588 1203 4712
rect 1133 4548 1139 4552
rect 749 4328 755 4352
rect 765 4148 771 4472
rect 829 4308 835 4332
rect 845 4328 851 4352
rect 861 4308 867 4372
rect 877 4368 883 4432
rect 973 4348 979 4352
rect 669 4088 675 4112
rect 685 4048 691 4112
rect 797 4108 803 4272
rect 877 4228 883 4292
rect 893 4288 899 4332
rect 909 4308 915 4312
rect 973 4308 979 4332
rect 1005 4328 1011 4332
rect 1053 4328 1059 4432
rect 1101 4428 1107 4472
rect 1085 4328 1091 4392
rect 1133 4388 1139 4532
rect 1149 4508 1155 4512
rect 1181 4488 1187 4492
rect 1229 4388 1235 4532
rect 1245 4488 1251 4492
rect 1245 4428 1251 4472
rect 1101 4308 1107 4312
rect 941 4288 947 4292
rect 1053 4288 1059 4292
rect 957 4208 963 4272
rect 973 4248 979 4272
rect 1037 4208 1043 4272
rect 653 3948 659 4012
rect 685 3968 691 4032
rect 749 3908 755 3912
rect 637 3888 643 3892
rect 461 3688 467 3712
rect 397 3508 403 3512
rect 429 3508 435 3512
rect 413 3488 419 3492
rect 445 3488 451 3552
rect 477 3548 483 3732
rect 525 3728 531 3752
rect 557 3748 563 3792
rect 573 3788 579 3872
rect 557 3728 563 3732
rect 493 3628 499 3692
rect 509 3548 515 3692
rect 509 3528 515 3532
rect 477 3508 483 3512
rect 365 3348 371 3352
rect 381 3348 387 3472
rect 285 3288 291 3312
rect 285 3168 291 3272
rect 285 3108 291 3152
rect 301 3148 307 3332
rect 317 3268 323 3312
rect 397 3283 403 3312
rect 397 3277 408 3283
rect 317 3088 323 3192
rect 333 3188 339 3232
rect 429 3208 435 3472
rect 445 3428 451 3472
rect 461 3408 467 3492
rect 445 3308 451 3352
rect 477 3288 483 3432
rect 493 3308 499 3312
rect 509 3308 515 3392
rect 525 3368 531 3412
rect 541 3323 547 3712
rect 573 3528 579 3532
rect 557 3508 563 3512
rect 589 3508 595 3872
rect 621 3868 627 3872
rect 653 3788 659 3832
rect 685 3788 691 3892
rect 765 3888 771 4092
rect 861 4088 867 4132
rect 877 4128 883 4132
rect 909 4128 915 4172
rect 1053 4163 1059 4272
rect 1101 4248 1107 4272
rect 1101 4168 1107 4232
rect 1053 4157 1075 4163
rect 925 4148 931 4152
rect 957 4068 963 4132
rect 973 4108 979 4112
rect 989 3988 995 4132
rect 1005 4128 1011 4132
rect 1037 4108 1043 4112
rect 1021 4088 1027 4092
rect 1069 4088 1075 4157
rect 1117 4148 1123 4292
rect 1133 4228 1139 4312
rect 1213 4308 1219 4312
rect 1149 4288 1155 4292
rect 1165 4288 1171 4292
rect 1261 4288 1267 4652
rect 1389 4648 1395 4652
rect 1389 4588 1395 4592
rect 1293 4548 1299 4552
rect 1277 4508 1283 4512
rect 1357 4428 1363 4492
rect 1293 4306 1299 4312
rect 1389 4308 1395 4532
rect 1421 4428 1427 4532
rect 1437 4528 1443 4652
rect 1464 4537 1475 4543
rect 1197 4268 1203 4272
rect 1229 4243 1235 4252
rect 1229 4237 1251 4243
rect 1245 4188 1251 4237
rect 1293 4188 1299 4252
rect 1213 4148 1219 4152
rect 1229 4148 1235 4152
rect 1085 4128 1091 4132
rect 1101 4008 1107 4132
rect 701 3728 707 3872
rect 717 3868 723 3872
rect 781 3848 787 3892
rect 845 3848 851 3892
rect 1085 3888 1091 3972
rect 1101 3948 1107 3972
rect 1101 3888 1107 3892
rect 621 3548 627 3712
rect 653 3528 659 3632
rect 653 3503 659 3512
rect 648 3497 659 3503
rect 573 3348 579 3372
rect 589 3348 595 3352
rect 621 3348 627 3472
rect 637 3408 643 3472
rect 541 3317 552 3323
rect 525 3268 531 3292
rect 589 3288 595 3332
rect 605 3328 611 3332
rect 669 3328 675 3532
rect 685 3428 691 3512
rect 701 3388 707 3712
rect 749 3708 755 3832
rect 893 3788 899 3872
rect 957 3868 963 3872
rect 973 3848 979 3872
rect 781 3668 787 3712
rect 797 3688 803 3712
rect 797 3643 803 3672
rect 781 3637 803 3643
rect 717 3508 723 3512
rect 733 3488 739 3632
rect 749 3488 755 3492
rect 717 3477 728 3483
rect 637 3308 643 3312
rect 413 3088 419 3152
rect 221 2968 227 2972
rect 301 2968 307 3072
rect 269 2888 275 2892
rect 285 2888 291 2912
rect 301 2848 307 2932
rect 205 2788 211 2832
rect 56 2697 67 2703
rect 61 2688 67 2697
rect 109 2683 115 2712
rect 93 2677 115 2683
rect 45 2588 51 2652
rect 93 2588 99 2677
rect 24 2537 35 2543
rect 13 2288 19 2532
rect 45 2508 51 2532
rect 61 2328 67 2532
rect 109 2508 115 2512
rect 45 2268 51 2312
rect 93 2288 99 2292
rect 125 2288 131 2672
rect 141 2668 147 2732
rect 237 2708 243 2712
rect 141 2528 147 2572
rect 157 2508 163 2532
rect 173 2508 179 2512
rect 205 2508 211 2512
rect 157 2483 163 2492
rect 157 2477 179 2483
rect 173 2308 179 2477
rect 221 2408 227 2532
rect 253 2428 259 2832
rect 285 2708 291 2832
rect 285 2568 291 2692
rect 317 2623 323 3072
rect 445 3048 451 3072
rect 333 2928 339 2932
rect 349 2928 355 2932
rect 381 2888 387 2972
rect 429 2948 435 2992
rect 397 2908 403 2912
rect 424 2897 435 2903
rect 381 2688 387 2832
rect 392 2677 403 2683
rect 301 2617 323 2623
rect 205 2308 211 2332
rect 221 2328 227 2332
rect 173 2288 179 2292
rect 189 2248 195 2292
rect 77 2128 83 2232
rect 221 2188 227 2292
rect 253 2228 259 2272
rect 285 2168 291 2552
rect 301 2328 307 2617
rect 333 2528 339 2592
rect 317 2388 323 2512
rect 349 2508 355 2632
rect 317 2328 323 2332
rect 301 2288 307 2312
rect 333 2168 339 2492
rect 349 2308 355 2452
rect 125 2128 131 2152
rect 317 2148 323 2152
rect 109 1908 115 1952
rect 125 1908 131 2112
rect 253 2088 259 2112
rect 285 2108 291 2112
rect 205 1928 211 1932
rect 125 1728 131 1892
rect 205 1868 211 1872
rect 221 1788 227 2072
rect 237 1908 243 1912
rect 269 1888 275 1892
rect 285 1848 291 1932
rect 317 1908 323 1912
rect 349 1908 355 2292
rect 365 2288 371 2292
rect 381 2188 387 2312
rect 397 2228 403 2677
rect 429 2648 435 2897
rect 445 2548 451 2712
rect 477 2708 483 3132
rect 493 3108 499 3232
rect 525 3148 531 3252
rect 621 3188 627 3232
rect 541 3068 547 3092
rect 525 2928 531 3052
rect 541 2948 547 2952
rect 605 2948 611 3112
rect 701 3108 707 3152
rect 717 3128 723 3477
rect 749 3468 755 3472
rect 733 3088 739 3332
rect 781 3108 787 3637
rect 829 3428 835 3512
rect 829 3348 835 3372
rect 797 3328 803 3332
rect 845 3328 851 3752
rect 941 3688 947 3832
rect 1021 3668 1027 3712
rect 861 3508 867 3512
rect 877 3488 883 3552
rect 909 3468 915 3552
rect 909 3428 915 3452
rect 877 3308 883 3412
rect 925 3383 931 3492
rect 941 3488 947 3492
rect 973 3488 979 3592
rect 989 3508 995 3552
rect 1037 3548 1043 3712
rect 1021 3448 1027 3532
rect 1037 3488 1043 3492
rect 1053 3468 1059 3872
rect 1069 3788 1075 3812
rect 1085 3608 1091 3872
rect 1117 3788 1123 4132
rect 1197 4028 1203 4112
rect 1229 4028 1235 4132
rect 1261 4108 1267 4152
rect 1277 4068 1283 4132
rect 1341 4108 1347 4112
rect 1181 3908 1187 3912
rect 1197 3908 1203 4012
rect 1245 3908 1251 4032
rect 1277 3988 1283 4032
rect 1357 3968 1363 4292
rect 1421 4268 1427 4412
rect 1453 4388 1459 4472
rect 1469 4388 1475 4537
rect 1485 4388 1491 4472
rect 1421 4228 1427 4232
rect 1421 4168 1427 4212
rect 1437 4208 1443 4272
rect 1453 4188 1459 4192
rect 1437 4108 1443 4132
rect 1389 4088 1395 4092
rect 1453 4088 1459 4092
rect 1469 4068 1475 4372
rect 1501 4288 1507 4863
rect 1677 4788 1683 4863
rect 1709 4857 1731 4863
rect 1629 4697 1640 4703
rect 1517 4603 1523 4692
rect 1517 4597 1539 4603
rect 1533 4588 1539 4597
rect 1517 4528 1523 4572
rect 1565 4528 1571 4632
rect 1597 4628 1603 4692
rect 1629 4688 1635 4697
rect 1709 4688 1715 4857
rect 1917 4788 1923 4863
rect 2429 4788 2435 4863
rect 3085 4788 3091 4863
rect 3501 4828 3507 4863
rect 5229 4788 5235 4863
rect 5437 4788 5443 4863
rect 5613 4788 5619 4863
rect 6301 4788 6307 4863
rect 6477 4788 6483 4863
rect 6573 4788 6579 4863
rect 6621 4828 6627 4863
rect 6589 4788 6595 4812
rect 3352 4737 3363 4743
rect 2237 4728 2243 4732
rect 2173 4706 2179 4712
rect 1992 4697 2003 4703
rect 1725 4648 1731 4652
rect 1837 4648 1843 4692
rect 1997 4688 2003 4697
rect 2472 4697 2483 4703
rect 2477 4688 2483 4697
rect 2637 4688 2643 4692
rect 1693 4588 1699 4632
rect 1997 4588 2003 4632
rect 1565 4508 1571 4512
rect 1533 4488 1539 4492
rect 1581 4428 1587 4532
rect 1517 4208 1523 4232
rect 1533 4228 1539 4232
rect 1485 4028 1491 4112
rect 1501 4108 1507 4132
rect 1517 4108 1523 4172
rect 1549 4128 1555 4292
rect 1565 4148 1571 4272
rect 1613 4188 1619 4532
rect 1645 4448 1651 4492
rect 1661 4306 1667 4372
rect 1581 4168 1587 4172
rect 1613 4108 1619 4152
rect 1661 4148 1667 4232
rect 1693 4148 1699 4512
rect 1709 4428 1715 4532
rect 1789 4528 1795 4532
rect 1757 4448 1763 4492
rect 1805 4388 1811 4512
rect 1821 4468 1827 4532
rect 1981 4528 1987 4572
rect 1901 4488 1907 4492
rect 1805 4368 1811 4372
rect 1805 4348 1811 4352
rect 1757 4323 1763 4332
rect 1757 4317 1779 4323
rect 1624 4097 1635 4103
rect 1421 3988 1427 4012
rect 1421 3968 1427 3972
rect 1309 3928 1315 3932
rect 1149 3808 1155 3892
rect 1165 3828 1171 3872
rect 1149 3768 1155 3792
rect 1213 3748 1219 3832
rect 1261 3828 1267 3872
rect 1277 3848 1283 3892
rect 1117 3628 1123 3632
rect 973 3388 979 3432
rect 925 3377 936 3383
rect 893 3348 899 3352
rect 989 3348 995 3392
rect 1005 3388 1011 3392
rect 1037 3328 1043 3412
rect 845 3288 851 3292
rect 909 3268 915 3312
rect 941 3288 947 3292
rect 1005 3288 1011 3292
rect 813 3128 819 3132
rect 904 3117 931 3123
rect 813 3108 819 3112
rect 925 3103 931 3117
rect 925 3097 936 3103
rect 637 3068 643 3072
rect 733 3068 739 3072
rect 493 2888 499 2892
rect 477 2588 483 2692
rect 493 2668 499 2672
rect 509 2588 515 2632
rect 477 2548 483 2552
rect 445 2528 451 2532
rect 461 2528 467 2532
rect 461 2303 467 2512
rect 456 2297 467 2303
rect 477 2288 483 2532
rect 493 2508 499 2532
rect 525 2528 531 2892
rect 541 2883 547 2912
rect 589 2908 595 2912
rect 541 2877 563 2883
rect 557 2568 563 2877
rect 589 2708 595 2752
rect 541 2503 547 2532
rect 536 2497 547 2503
rect 605 2428 611 2932
rect 621 2908 627 2932
rect 653 2848 659 2912
rect 621 2608 627 2692
rect 621 2588 627 2592
rect 653 2528 659 2832
rect 669 2548 675 2952
rect 781 2948 787 3092
rect 861 3048 867 3072
rect 893 3028 899 3072
rect 925 2968 931 3032
rect 973 3028 979 3112
rect 685 2728 691 2732
rect 701 2688 707 2852
rect 717 2748 723 2892
rect 861 2788 867 2912
rect 717 2708 723 2732
rect 653 2468 659 2512
rect 552 2337 563 2343
rect 477 2188 483 2252
rect 493 2248 499 2272
rect 509 2268 515 2312
rect 525 2308 531 2312
rect 317 1868 323 1892
rect 365 1888 371 2092
rect 381 1988 387 2112
rect 413 1988 419 2112
rect 397 1908 403 1932
rect 429 1928 435 2132
rect 445 2108 451 2132
rect 493 2108 499 2172
rect 525 2148 531 2252
rect 557 2188 563 2337
rect 589 2308 595 2412
rect 621 2343 627 2432
rect 669 2368 675 2532
rect 685 2528 691 2552
rect 621 2337 643 2343
rect 573 2268 579 2272
rect 621 2248 627 2312
rect 605 2188 611 2232
rect 541 2148 547 2152
rect 525 2128 531 2132
rect 557 2108 563 2112
rect 605 2108 611 2172
rect 637 2128 643 2337
rect 653 2288 659 2292
rect 685 2228 691 2272
rect 701 2228 707 2672
rect 749 2668 755 2712
rect 845 2688 851 2732
rect 909 2708 915 2712
rect 925 2688 931 2952
rect 989 2948 995 3072
rect 941 2763 947 2832
rect 941 2757 963 2763
rect 797 2668 803 2672
rect 717 2588 723 2652
rect 749 2648 755 2652
rect 733 2548 739 2552
rect 749 2528 755 2532
rect 845 2508 851 2512
rect 717 2328 723 2432
rect 717 2308 723 2312
rect 765 2308 771 2452
rect 781 2348 787 2492
rect 829 2468 835 2472
rect 717 2228 723 2272
rect 669 2148 675 2192
rect 765 2188 771 2292
rect 653 2088 659 2132
rect 461 1928 467 1932
rect 493 1928 499 1932
rect 557 1928 563 1932
rect 429 1908 435 1912
rect 541 1908 547 1912
rect 589 1908 595 1972
rect 525 1883 531 1892
rect 605 1888 611 1892
rect 525 1877 536 1883
rect 189 1768 195 1772
rect 237 1728 243 1752
rect 253 1748 259 1752
rect 285 1748 291 1812
rect 109 1588 115 1712
rect 125 1568 131 1712
rect 237 1708 243 1712
rect 13 1488 19 1492
rect 125 1488 131 1532
rect 13 1328 19 1332
rect 29 1168 35 1432
rect 109 1368 115 1432
rect 173 1428 179 1432
rect 61 1323 67 1332
rect 56 1317 67 1323
rect 45 1188 51 1272
rect 61 988 67 1112
rect 93 1108 99 1112
rect 77 1088 83 1092
rect 109 1083 115 1332
rect 125 1088 131 1392
rect 141 1348 147 1352
rect 221 1348 227 1552
rect 269 1508 275 1712
rect 285 1588 291 1732
rect 269 1468 275 1472
rect 285 1348 291 1572
rect 317 1528 323 1692
rect 333 1688 339 1872
rect 365 1828 371 1872
rect 365 1748 371 1752
rect 413 1728 419 1792
rect 429 1768 435 1872
rect 477 1837 488 1843
rect 461 1788 467 1832
rect 333 1408 339 1672
rect 349 1668 355 1712
rect 349 1508 355 1592
rect 365 1488 371 1652
rect 413 1528 419 1632
rect 429 1568 435 1732
rect 445 1728 451 1732
rect 445 1508 451 1712
rect 477 1708 483 1837
rect 493 1708 499 1712
rect 461 1508 467 1652
rect 381 1488 387 1492
rect 477 1488 483 1632
rect 493 1488 499 1692
rect 525 1648 531 1877
rect 621 1868 627 1912
rect 669 1908 675 1912
rect 685 1908 691 2112
rect 717 1988 723 2092
rect 829 2043 835 2292
rect 845 2288 851 2352
rect 877 2148 883 2572
rect 909 2428 915 2432
rect 925 2403 931 2672
rect 957 2608 963 2757
rect 973 2728 979 2832
rect 989 2828 995 2932
rect 1005 2928 1011 3252
rect 1021 3048 1027 3112
rect 1053 3083 1059 3452
rect 1069 3408 1075 3512
rect 1085 3388 1091 3492
rect 1101 3468 1107 3472
rect 1133 3348 1139 3592
rect 1069 3328 1075 3332
rect 1117 3268 1123 3312
rect 1149 3268 1155 3712
rect 1181 3688 1187 3732
rect 1261 3688 1267 3812
rect 1277 3808 1283 3832
rect 1181 3508 1187 3672
rect 1197 3508 1203 3512
rect 1213 3388 1219 3672
rect 1357 3588 1363 3952
rect 1517 3908 1523 3912
rect 1389 3868 1395 3892
rect 1501 3868 1507 3892
rect 1533 3888 1539 3972
rect 1549 3908 1555 3912
rect 1581 3908 1587 4032
rect 1565 3868 1571 3872
rect 1469 3748 1475 3832
rect 1453 3688 1459 3732
rect 1245 3328 1251 3372
rect 1341 3328 1347 3432
rect 1181 3308 1187 3312
rect 1048 3077 1059 3083
rect 1037 2988 1043 3072
rect 1053 3028 1059 3032
rect 1069 2948 1075 3232
rect 1096 3117 1139 3123
rect 1133 3108 1139 3117
rect 1149 3108 1155 3112
rect 1133 3008 1139 3072
rect 1149 2948 1155 2952
rect 1165 2948 1171 3132
rect 1181 3108 1187 3152
rect 1245 3148 1251 3152
rect 1213 3108 1219 3112
rect 1229 3108 1235 3132
rect 1245 3108 1251 3132
rect 1181 3008 1187 3092
rect 1197 3068 1203 3072
rect 1037 2928 1043 2932
rect 1117 2928 1123 2932
rect 1229 2928 1235 3032
rect 973 2688 979 2712
rect 973 2543 979 2672
rect 989 2648 995 2712
rect 973 2537 984 2543
rect 1005 2528 1011 2912
rect 1005 2508 1011 2512
rect 909 2397 931 2403
rect 909 2228 915 2397
rect 941 2328 947 2412
rect 941 2288 947 2312
rect 973 2308 979 2432
rect 989 2328 995 2452
rect 1021 2448 1027 2912
rect 1085 2908 1091 2912
rect 1101 2888 1107 2912
rect 1165 2908 1171 2912
rect 1053 2688 1059 2752
rect 1101 2648 1107 2712
rect 1133 2708 1139 2732
rect 1165 2668 1171 2672
rect 1133 2548 1139 2552
rect 1085 2368 1091 2432
rect 1117 2428 1123 2512
rect 1181 2508 1187 2592
rect 1197 2588 1203 2812
rect 1213 2648 1219 2712
rect 1229 2708 1235 2912
rect 1261 2708 1267 3072
rect 1309 2908 1315 3092
rect 1325 3048 1331 3072
rect 1341 3068 1347 3112
rect 1341 2968 1347 2972
rect 1325 2948 1331 2952
rect 1357 2828 1363 3492
rect 1389 3403 1395 3472
rect 1373 3397 1395 3403
rect 1373 3328 1379 3397
rect 1453 3348 1459 3632
rect 1469 3528 1475 3732
rect 1501 3708 1507 3832
rect 1517 3748 1523 3792
rect 1581 3728 1587 3792
rect 1512 3697 1523 3703
rect 1485 3508 1491 3572
rect 1469 3488 1475 3492
rect 1405 3108 1411 3132
rect 1437 3128 1443 3232
rect 1437 3088 1443 3112
rect 1421 2988 1427 3052
rect 1453 2988 1459 3332
rect 1517 3303 1523 3697
rect 1581 3648 1587 3672
rect 1533 3528 1539 3632
rect 1581 3528 1587 3632
rect 1597 3608 1603 4032
rect 1613 3988 1619 4032
rect 1629 4008 1635 4097
rect 1661 4088 1667 4112
rect 1677 4068 1683 4132
rect 1709 4128 1715 4212
rect 1725 4148 1731 4312
rect 1741 4148 1747 4312
rect 1757 4188 1763 4292
rect 1773 4288 1779 4317
rect 1789 4148 1795 4172
rect 1821 4168 1827 4452
rect 1901 4448 1907 4472
rect 1805 4148 1811 4152
rect 1821 4128 1827 4132
rect 1709 4068 1715 4072
rect 1613 3708 1619 3732
rect 1629 3708 1635 3712
rect 1645 3628 1651 3892
rect 1661 3868 1667 3912
rect 1661 3728 1667 3832
rect 1677 3788 1683 4052
rect 1725 3988 1731 4112
rect 1805 4088 1811 4112
rect 1837 4088 1843 4092
rect 1853 4088 1859 4092
rect 1741 3948 1747 4072
rect 1709 3928 1715 3932
rect 1709 3763 1715 3912
rect 1853 3908 1859 4032
rect 1869 3968 1875 4132
rect 1885 4048 1891 4292
rect 1901 4148 1907 4412
rect 1917 4388 1923 4492
rect 1965 4388 1971 4452
rect 2029 4428 2035 4532
rect 2093 4528 2099 4532
rect 2029 4408 2035 4412
rect 1997 4328 2003 4372
rect 2093 4368 2099 4512
rect 2109 4488 2115 4512
rect 2125 4448 2131 4492
rect 2141 4388 2147 4412
rect 1917 4188 1923 4272
rect 1949 4268 1955 4272
rect 1949 4248 1955 4252
rect 1997 4148 2003 4152
rect 2013 4128 2019 4272
rect 2029 4208 2035 4292
rect 2061 4228 2067 4312
rect 2141 4308 2147 4352
rect 2173 4348 2179 4472
rect 2189 4448 2195 4492
rect 2221 4363 2227 4532
rect 2237 4388 2243 4592
rect 2221 4357 2243 4363
rect 2205 4288 2211 4312
rect 2237 4288 2243 4357
rect 2253 4328 2259 4532
rect 2269 4528 2275 4652
rect 2445 4548 2451 4652
rect 2717 4648 2723 4672
rect 2573 4548 2579 4632
rect 2701 4628 2707 4632
rect 2749 4628 2755 4712
rect 2797 4608 2803 4692
rect 2813 4648 2819 4712
rect 2973 4688 2979 4692
rect 2941 4588 2947 4612
rect 3021 4588 3027 4632
rect 2557 4528 2563 4532
rect 2493 4508 2499 4512
rect 2269 4428 2275 4432
rect 2269 4328 2275 4412
rect 2285 4388 2291 4432
rect 2317 4348 2323 4472
rect 2525 4468 2531 4492
rect 2573 4408 2579 4532
rect 2621 4528 2627 4532
rect 2653 4528 2659 4572
rect 2621 4428 2627 4492
rect 2637 4488 2643 4512
rect 2397 4308 2403 4332
rect 2109 4248 2115 4272
rect 2125 4268 2131 4272
rect 2077 4148 2083 4192
rect 1949 4088 1955 4092
rect 1901 3908 1907 4052
rect 1933 3928 1939 3972
rect 1949 3908 1955 4072
rect 1725 3843 1731 3872
rect 1741 3868 1747 3892
rect 1821 3888 1827 3892
rect 1805 3868 1811 3872
rect 1773 3843 1779 3852
rect 1725 3837 1779 3843
rect 1789 3808 1795 3832
rect 1709 3757 1720 3763
rect 1693 3648 1699 3752
rect 1709 3748 1715 3757
rect 1741 3748 1747 3752
rect 1773 3708 1779 3712
rect 1597 3468 1603 3492
rect 1629 3488 1635 3512
rect 1677 3508 1683 3512
rect 1533 3437 1544 3443
rect 1533 3348 1539 3437
rect 1549 3368 1555 3392
rect 1501 3297 1523 3303
rect 1485 3128 1491 3292
rect 1501 3188 1507 3297
rect 1501 2988 1507 3012
rect 1437 2908 1443 2972
rect 1453 2928 1459 2952
rect 1533 2928 1539 3332
rect 1549 2948 1555 3352
rect 1565 3048 1571 3092
rect 1581 2988 1587 3352
rect 1629 3328 1635 3432
rect 1661 3343 1667 3472
rect 1693 3448 1699 3632
rect 1757 3508 1763 3512
rect 1773 3488 1779 3492
rect 1709 3388 1715 3452
rect 1741 3388 1747 3452
rect 1805 3448 1811 3712
rect 1837 3708 1843 3752
rect 1885 3748 1891 3872
rect 1805 3428 1811 3432
rect 1821 3408 1827 3432
rect 1805 3368 1811 3372
rect 1885 3368 1891 3452
rect 1901 3408 1907 3712
rect 1933 3708 1939 3752
rect 1949 3748 1955 3772
rect 1965 3728 1971 3892
rect 1981 3888 1987 4112
rect 1997 3888 2003 3932
rect 2029 3888 2035 3952
rect 2061 3903 2067 4112
rect 2077 4108 2083 4112
rect 2077 4028 2083 4092
rect 2093 4088 2099 4232
rect 2125 4108 2131 4212
rect 2141 4148 2147 4172
rect 2157 3988 2163 4252
rect 2205 4148 2211 4272
rect 2237 4188 2243 4272
rect 2285 4188 2291 4212
rect 2221 4117 2232 4123
rect 2173 4103 2179 4112
rect 2221 4103 2227 4117
rect 2285 4108 2291 4112
rect 2301 4108 2307 4292
rect 2317 4268 2323 4272
rect 2381 4268 2387 4292
rect 2413 4288 2419 4312
rect 2488 4297 2499 4303
rect 2413 4268 2419 4272
rect 2461 4248 2467 4272
rect 2349 4208 2355 4232
rect 2317 4128 2323 4152
rect 2173 4097 2227 4103
rect 2285 4028 2291 4092
rect 2333 4088 2339 4132
rect 2349 4128 2355 4192
rect 2397 4128 2403 4132
rect 2429 4108 2435 4112
rect 2088 3917 2099 3923
rect 2061 3897 2083 3903
rect 1997 3848 2003 3852
rect 2013 3788 2019 3832
rect 2013 3708 2019 3712
rect 2029 3708 2035 3732
rect 2045 3688 2051 3712
rect 2061 3688 2067 3832
rect 2077 3828 2083 3897
rect 2093 3788 2099 3917
rect 2109 3888 2115 3892
rect 2109 3848 2115 3872
rect 2125 3868 2131 3872
rect 2093 3768 2099 3772
rect 2141 3748 2147 3932
rect 2205 3908 2211 3972
rect 2333 3948 2339 4072
rect 2445 4048 2451 4132
rect 2461 4128 2467 4132
rect 2477 4128 2483 4192
rect 2493 4183 2499 4297
rect 2525 4188 2531 4332
rect 2541 4308 2547 4312
rect 2557 4188 2563 4332
rect 2493 4177 2504 4183
rect 2573 4148 2579 4192
rect 2605 4168 2611 4312
rect 2557 4108 2563 4112
rect 2525 4068 2531 4092
rect 2301 3908 2307 3912
rect 2397 3906 2403 4032
rect 2189 3888 2195 3892
rect 2077 3728 2083 3732
rect 1917 3488 1923 3492
rect 1949 3488 1955 3492
rect 1981 3488 1987 3572
rect 2157 3548 2163 3652
rect 2013 3508 2019 3512
rect 1949 3388 1955 3472
rect 2013 3388 2019 3472
rect 2093 3428 2099 3532
rect 2109 3468 2115 3492
rect 2061 3388 2067 3392
rect 2093 3388 2099 3412
rect 1656 3337 1667 3343
rect 1597 3148 1603 3312
rect 1661 3308 1667 3312
rect 1693 3268 1699 3312
rect 1613 3108 1619 3172
rect 1645 3068 1651 3072
rect 1597 2928 1603 2932
rect 1533 2908 1539 2912
rect 1629 2908 1635 2912
rect 1645 2888 1651 2992
rect 1405 2808 1411 2832
rect 1309 2748 1315 2752
rect 1277 2728 1283 2732
rect 1293 2708 1299 2732
rect 1352 2717 1379 2723
rect 1373 2708 1379 2717
rect 1197 2548 1203 2572
rect 1213 2548 1219 2632
rect 1245 2528 1251 2692
rect 1261 2668 1267 2672
rect 1261 2503 1267 2652
rect 1389 2648 1395 2712
rect 1405 2588 1411 2792
rect 1421 2668 1427 2692
rect 1245 2497 1267 2503
rect 1069 2308 1075 2332
rect 1085 2308 1091 2312
rect 957 2248 963 2292
rect 1101 2288 1107 2292
rect 925 2128 931 2152
rect 1021 2148 1027 2272
rect 1069 2228 1075 2272
rect 1117 2268 1123 2332
rect 1149 2328 1155 2452
rect 1229 2448 1235 2472
rect 1229 2388 1235 2412
rect 1165 2303 1171 2352
rect 1181 2308 1187 2312
rect 1149 2297 1171 2303
rect 829 2037 851 2043
rect 733 1928 739 1972
rect 749 1968 755 2032
rect 589 1748 595 1772
rect 589 1708 595 1712
rect 605 1708 611 1812
rect 637 1728 643 1792
rect 653 1748 659 1892
rect 749 1888 755 1932
rect 829 1928 835 1952
rect 845 1928 851 2037
rect 877 1988 883 2112
rect 781 1888 787 1912
rect 845 1888 851 1892
rect 669 1868 675 1872
rect 669 1748 675 1832
rect 877 1788 883 1932
rect 941 1928 947 1972
rect 893 1888 899 1892
rect 1005 1888 1011 1952
rect 1021 1908 1027 2032
rect 1053 1988 1059 2114
rect 1069 1968 1075 2212
rect 1117 2128 1123 2152
rect 1037 1928 1043 1932
rect 1053 1888 1059 1892
rect 957 1868 963 1872
rect 973 1868 979 1872
rect 541 1528 547 1692
rect 605 1648 611 1692
rect 573 1548 579 1632
rect 669 1523 675 1732
rect 765 1728 771 1732
rect 685 1668 691 1712
rect 653 1517 675 1523
rect 589 1508 595 1512
rect 189 1308 195 1312
rect 253 1288 259 1314
rect 141 1108 147 1172
rect 104 1077 115 1083
rect 93 948 99 1072
rect 125 968 131 1072
rect 45 908 51 912
rect 13 728 19 732
rect 29 668 35 832
rect 56 697 67 703
rect 61 688 67 697
rect 93 588 99 932
rect 141 928 147 932
rect 157 903 163 1112
rect 173 928 179 1232
rect 189 1108 195 1152
rect 221 1108 227 1112
rect 189 1088 195 1092
rect 253 1088 259 1252
rect 333 1128 339 1172
rect 317 1108 323 1112
rect 205 1008 211 1072
rect 189 948 195 992
rect 205 948 211 972
rect 269 928 275 1032
rect 301 1008 307 1092
rect 317 1068 323 1072
rect 285 948 291 952
rect 317 948 323 952
rect 349 923 355 1272
rect 381 1268 387 1472
rect 493 1468 499 1472
rect 365 1108 371 1232
rect 381 1188 387 1232
rect 333 917 355 923
rect 173 908 179 912
rect 152 897 163 903
rect 237 888 243 892
rect 253 848 259 892
rect 109 728 115 832
rect 269 788 275 912
rect 173 708 179 712
rect 189 688 195 732
rect 317 728 323 832
rect 333 708 339 917
rect 349 848 355 892
rect 365 708 371 1092
rect 381 1088 387 1152
rect 413 1083 419 1232
rect 445 1108 451 1112
rect 413 1077 424 1083
rect 397 1048 403 1052
rect 397 948 403 972
rect 381 928 387 932
rect 445 748 451 832
rect 189 548 195 552
rect 285 548 291 572
rect 13 528 19 532
rect 45 528 51 532
rect 173 528 179 532
rect 317 528 323 532
rect 61 388 67 512
rect 93 388 99 472
rect 13 288 19 312
rect 13 128 19 132
rect 61 123 67 132
rect 56 117 67 123
rect 173 -43 179 152
rect 189 128 195 512
rect 333 488 339 592
rect 381 548 387 712
rect 461 688 467 1152
rect 493 1128 499 1452
rect 509 1128 515 1492
rect 541 1488 547 1492
rect 605 1448 611 1512
rect 525 1328 531 1432
rect 637 1408 643 1472
rect 605 1388 611 1392
rect 573 1108 579 1132
rect 621 1108 627 1132
rect 477 1028 483 1032
rect 493 948 499 1072
rect 573 1008 579 1072
rect 637 1008 643 1072
rect 653 1068 659 1517
rect 685 1508 691 1632
rect 701 1528 707 1692
rect 765 1648 771 1712
rect 781 1668 787 1732
rect 749 1508 755 1532
rect 685 1348 691 1472
rect 525 848 531 912
rect 573 748 579 992
rect 637 928 643 932
rect 653 908 659 1032
rect 669 888 675 932
rect 685 928 691 1112
rect 733 1108 739 1492
rect 797 1488 803 1572
rect 749 1468 755 1472
rect 781 1348 787 1352
rect 749 1308 755 1314
rect 781 1188 787 1272
rect 813 1248 819 1492
rect 829 1488 835 1512
rect 861 1508 867 1752
rect 909 1748 915 1852
rect 925 1768 931 1832
rect 1005 1808 1011 1872
rect 1069 1788 1075 1932
rect 1101 1928 1107 2032
rect 1133 1908 1139 1912
rect 1149 1888 1155 2297
rect 1213 2288 1219 2312
rect 1197 2228 1203 2272
rect 1181 2008 1187 2032
rect 1101 1788 1107 1872
rect 1181 1788 1187 1872
rect 1181 1768 1187 1772
rect 909 1608 915 1732
rect 893 1528 899 1552
rect 893 1508 899 1512
rect 941 1508 947 1592
rect 957 1528 963 1732
rect 973 1728 979 1732
rect 1069 1668 1075 1712
rect 1085 1708 1091 1712
rect 973 1528 979 1632
rect 1101 1628 1107 1732
rect 1133 1728 1139 1732
rect 1101 1588 1107 1612
rect 1021 1528 1027 1532
rect 1133 1528 1139 1532
rect 829 1303 835 1472
rect 845 1388 851 1492
rect 973 1488 979 1512
rect 1053 1488 1059 1492
rect 845 1328 851 1372
rect 893 1348 899 1392
rect 909 1328 915 1432
rect 893 1308 899 1312
rect 829 1297 851 1303
rect 845 1168 851 1297
rect 957 1288 963 1432
rect 973 1423 979 1472
rect 973 1417 995 1423
rect 973 1308 979 1372
rect 989 1348 995 1417
rect 989 1328 995 1332
rect 749 1108 755 1132
rect 893 1128 899 1212
rect 861 1108 867 1112
rect 717 908 723 912
rect 525 728 531 732
rect 573 708 579 732
rect 589 708 595 872
rect 733 868 739 1072
rect 765 948 771 1032
rect 781 928 787 972
rect 797 948 803 952
rect 909 948 915 1072
rect 749 868 755 912
rect 797 843 803 932
rect 781 837 803 843
rect 477 688 483 692
rect 589 688 595 692
rect 461 668 467 672
rect 573 668 579 672
rect 413 548 419 572
rect 493 548 499 552
rect 557 548 563 652
rect 605 608 611 632
rect 365 488 371 512
rect 205 308 211 432
rect 285 328 291 332
rect 301 308 307 332
rect 333 288 339 312
rect 349 308 355 332
rect 365 288 371 352
rect 381 283 387 532
rect 413 368 419 532
rect 477 528 483 532
rect 493 508 499 512
rect 509 488 515 492
rect 541 428 547 512
rect 413 308 419 332
rect 429 328 435 352
rect 461 337 488 343
rect 461 303 467 337
rect 477 308 483 312
rect 456 297 467 303
rect 525 288 531 372
rect 541 328 547 352
rect 573 328 579 472
rect 573 308 579 312
rect 589 308 595 352
rect 605 328 611 332
rect 381 277 392 283
rect 253 248 259 272
rect 253 143 259 152
rect 253 137 275 143
rect 269 -37 275 137
rect 301 123 307 132
rect 381 128 387 232
rect 413 188 419 272
rect 477 268 483 272
rect 621 248 627 532
rect 637 508 643 712
rect 669 708 675 732
rect 685 688 691 692
rect 717 688 723 832
rect 781 728 787 837
rect 669 468 675 512
rect 717 488 723 672
rect 749 588 755 612
rect 781 548 787 712
rect 797 708 803 732
rect 845 688 851 932
rect 925 928 931 1112
rect 957 1068 963 1192
rect 1005 1148 1011 1232
rect 1037 1228 1043 1292
rect 1053 1288 1059 1472
rect 1101 1428 1107 1492
rect 1181 1488 1187 1572
rect 1149 1388 1155 1432
rect 1197 1368 1203 1492
rect 1213 1388 1219 1852
rect 1229 1728 1235 2372
rect 1245 2328 1251 2497
rect 1277 2468 1283 2512
rect 1293 2508 1299 2532
rect 1245 2128 1251 2132
rect 1277 2128 1283 2432
rect 1309 2168 1315 2252
rect 1325 2103 1331 2532
rect 1405 2468 1411 2512
rect 1453 2508 1459 2832
rect 1469 2708 1475 2732
rect 1469 2428 1475 2692
rect 1501 2648 1507 2712
rect 1501 2548 1507 2552
rect 1517 2528 1523 2772
rect 1597 2728 1603 2812
rect 1533 2688 1539 2712
rect 1597 2708 1603 2712
rect 1581 2608 1587 2692
rect 1373 2308 1379 2312
rect 1309 2097 1331 2103
rect 1309 1948 1315 2097
rect 1261 1908 1267 1932
rect 1373 1908 1379 2252
rect 1453 2248 1459 2292
rect 1469 2288 1475 2392
rect 1501 2388 1507 2432
rect 1517 2328 1523 2512
rect 1549 2503 1555 2532
rect 1565 2528 1571 2572
rect 1597 2508 1603 2532
rect 1549 2497 1560 2503
rect 1517 2288 1523 2292
rect 1533 2288 1539 2352
rect 1597 2348 1603 2352
rect 1453 2183 1459 2232
rect 1448 2177 1459 2183
rect 1469 2168 1475 2272
rect 1501 2188 1507 2272
rect 1549 2268 1555 2292
rect 1405 1968 1411 2112
rect 1453 2048 1459 2112
rect 1469 1968 1475 2132
rect 1485 2048 1491 2092
rect 1501 2028 1507 2132
rect 1549 2128 1555 2132
rect 1517 2028 1523 2112
rect 1565 2088 1571 2312
rect 1581 2248 1587 2312
rect 1613 2228 1619 2772
rect 1661 2768 1667 3132
rect 1677 3108 1683 3132
rect 1693 2968 1699 3252
rect 1725 3128 1731 3332
rect 1741 3308 1747 3312
rect 1805 3308 1811 3332
rect 1869 3328 1875 3352
rect 1885 3328 1891 3352
rect 1869 3188 1875 3312
rect 1917 3308 1923 3312
rect 2013 3288 2019 3332
rect 1837 3128 1843 3152
rect 1757 3108 1763 3112
rect 1837 3108 1843 3112
rect 1917 3108 1923 3152
rect 1997 3128 2003 3232
rect 1709 3088 1715 3092
rect 1741 3068 1747 3072
rect 1805 3068 1811 3092
rect 1997 3063 2003 3112
rect 2013 3108 2019 3272
rect 2045 3168 2051 3312
rect 2093 3308 2099 3352
rect 2173 3348 2179 3492
rect 2205 3368 2211 3472
rect 2221 3468 2227 3872
rect 2269 3588 2275 3892
rect 2285 3868 2291 3872
rect 2285 3528 2291 3532
rect 2237 3508 2243 3512
rect 2125 3308 2131 3332
rect 2061 3288 2067 3292
rect 2093 3248 2099 3292
rect 2029 3088 2035 3152
rect 1997 3057 2008 3063
rect 1709 2988 1715 3052
rect 1789 3008 1795 3032
rect 1693 2903 1699 2952
rect 1709 2948 1715 2972
rect 1725 2968 1731 2972
rect 1885 2968 1891 3052
rect 1789 2928 1795 2952
rect 1688 2897 1699 2903
rect 1805 2888 1811 2892
rect 1661 2708 1667 2752
rect 1709 2648 1715 2712
rect 1629 2628 1635 2632
rect 1645 2543 1651 2612
rect 1629 2537 1651 2543
rect 1629 2488 1635 2537
rect 1661 2368 1667 2632
rect 1725 2608 1731 2632
rect 1677 2488 1683 2512
rect 1693 2448 1699 2532
rect 1661 2328 1667 2352
rect 1629 2288 1635 2292
rect 1693 2288 1699 2292
rect 1709 2288 1715 2312
rect 1693 2263 1699 2272
rect 1693 2257 1715 2263
rect 1645 2148 1651 2152
rect 1613 2128 1619 2132
rect 1661 2128 1667 2192
rect 1709 2188 1715 2257
rect 1725 2128 1731 2252
rect 1597 2088 1603 2112
rect 1405 1928 1411 1952
rect 1389 1908 1395 1912
rect 1373 1748 1379 1832
rect 1325 1717 1336 1723
rect 1229 1648 1235 1712
rect 1277 1708 1283 1712
rect 1229 1588 1235 1612
rect 1293 1508 1299 1512
rect 1309 1488 1315 1532
rect 1325 1508 1331 1717
rect 1373 1588 1379 1712
rect 1389 1628 1395 1872
rect 1405 1848 1411 1912
rect 1421 1888 1427 1912
rect 1565 1908 1571 1912
rect 1517 1888 1523 1892
rect 1453 1868 1459 1872
rect 1549 1868 1555 1872
rect 1597 1868 1603 1872
rect 1405 1708 1411 1792
rect 1421 1788 1427 1832
rect 1437 1703 1443 1832
rect 1432 1697 1443 1703
rect 1357 1528 1363 1532
rect 1165 1348 1171 1352
rect 1069 1288 1075 1312
rect 973 1108 979 1112
rect 957 948 963 1052
rect 973 968 979 1072
rect 1021 1068 1027 1092
rect 1037 1028 1043 1112
rect 1117 1048 1123 1092
rect 973 928 979 932
rect 893 908 899 912
rect 925 828 931 872
rect 877 708 883 732
rect 925 688 931 812
rect 957 748 963 872
rect 973 868 979 912
rect 989 888 995 912
rect 1069 908 1075 912
rect 1021 788 1027 892
rect 989 728 995 732
rect 1005 708 1011 712
rect 845 588 851 672
rect 845 548 851 572
rect 861 528 867 552
rect 909 508 915 512
rect 925 508 931 572
rect 941 508 947 532
rect 973 508 979 592
rect 1021 548 1027 752
rect 1037 748 1043 892
rect 1085 888 1091 892
rect 1069 688 1075 832
rect 1085 708 1091 732
rect 1101 688 1107 952
rect 1117 868 1123 912
rect 1133 808 1139 932
rect 1117 708 1123 712
rect 1149 688 1155 1332
rect 1165 1108 1171 1332
rect 1213 1328 1219 1372
rect 1261 1348 1267 1472
rect 1293 1368 1299 1432
rect 1309 1428 1315 1472
rect 1325 1408 1331 1492
rect 1389 1488 1395 1612
rect 1469 1528 1475 1732
rect 1517 1728 1523 1732
rect 1533 1728 1539 1732
rect 1565 1728 1571 1752
rect 1581 1748 1587 1752
rect 1613 1748 1619 2112
rect 1677 2108 1683 2112
rect 1661 1908 1667 1932
rect 1693 1908 1699 1952
rect 1709 1928 1715 2032
rect 1645 1848 1651 1852
rect 1677 1848 1683 1892
rect 1677 1748 1683 1832
rect 1709 1803 1715 1872
rect 1725 1828 1731 2112
rect 1741 1888 1747 2832
rect 1789 2808 1795 2832
rect 1821 2748 1827 2912
rect 1933 2908 1939 2912
rect 1949 2908 1955 3012
rect 2029 3008 2035 3032
rect 1757 2528 1763 2572
rect 1757 2508 1763 2512
rect 1773 2383 1779 2732
rect 1789 2528 1795 2692
rect 1821 2628 1827 2692
rect 1837 2648 1843 2692
rect 1853 2688 1859 2812
rect 1821 2588 1827 2612
rect 1885 2588 1891 2872
rect 1933 2828 1939 2832
rect 1965 2748 1971 2912
rect 2061 2908 2067 3132
rect 2093 3103 2099 3232
rect 2141 3228 2147 3332
rect 2205 3328 2211 3352
rect 2253 3348 2259 3452
rect 2237 3328 2243 3332
rect 2173 3317 2184 3323
rect 2157 3268 2163 3312
rect 2173 3308 2179 3317
rect 2269 3323 2275 3412
rect 2285 3388 2291 3492
rect 2301 3348 2307 3672
rect 2317 3588 2323 3832
rect 2429 3768 2435 3992
rect 2525 3988 2531 4012
rect 2461 3908 2467 3912
rect 2557 3908 2563 4092
rect 2589 4088 2595 4132
rect 2605 4128 2611 4152
rect 2637 4108 2643 4332
rect 2637 4068 2643 4092
rect 2653 3948 2659 4292
rect 2669 4268 2675 4532
rect 2701 4288 2707 4532
rect 2797 4528 2803 4532
rect 2733 4468 2739 4492
rect 2733 4428 2739 4452
rect 2717 4288 2723 4372
rect 2749 4328 2755 4332
rect 2765 4328 2771 4332
rect 2669 4168 2675 4252
rect 2685 4128 2691 4192
rect 2669 4088 2675 4092
rect 2701 4068 2707 4132
rect 2605 3908 2611 3912
rect 2509 3837 2520 3843
rect 2461 3768 2467 3772
rect 2509 3768 2515 3837
rect 2557 3768 2563 3872
rect 2397 3728 2403 3752
rect 2509 3748 2515 3752
rect 2653 3748 2659 3772
rect 2669 3768 2675 4052
rect 2701 3888 2707 4052
rect 2733 3908 2739 4292
rect 2781 4288 2787 4352
rect 2797 4348 2803 4452
rect 2797 4308 2803 4312
rect 2781 4208 2787 4272
rect 2797 4188 2803 4232
rect 2829 4228 2835 4512
rect 2845 4328 2851 4572
rect 2877 4508 2883 4532
rect 2909 4508 2915 4512
rect 2877 4288 2883 4372
rect 2925 4368 2931 4532
rect 3005 4528 3011 4532
rect 2973 4508 2979 4512
rect 2941 4448 2947 4492
rect 2941 4308 2947 4392
rect 3005 4368 3011 4512
rect 3037 4488 3043 4632
rect 3101 4628 3107 4632
rect 3101 4588 3107 4612
rect 3245 4568 3251 4612
rect 3309 4588 3315 4692
rect 3357 4588 3363 4737
rect 3421 4608 3427 4632
rect 3085 4508 3091 4512
rect 3053 4448 3059 4492
rect 3117 4488 3123 4552
rect 3149 4508 3155 4532
rect 3213 4528 3219 4532
rect 3245 4528 3251 4552
rect 2957 4328 2963 4332
rect 3000 4317 3011 4323
rect 2893 4248 2899 4292
rect 2989 4288 2995 4292
rect 3005 4288 3011 4317
rect 3021 4288 3027 4412
rect 3037 4308 3043 4312
rect 3101 4308 3107 4372
rect 3053 4288 3059 4292
rect 3069 4288 3075 4292
rect 2749 4048 2755 4132
rect 2749 3908 2755 3912
rect 2744 3877 2755 3883
rect 2749 3868 2755 3877
rect 2669 3748 2675 3752
rect 2621 3728 2627 3732
rect 2413 3708 2419 3712
rect 2333 3688 2339 3692
rect 2365 3528 2371 3532
rect 2349 3468 2355 3492
rect 2264 3317 2275 3323
rect 2237 3288 2243 3292
rect 2109 3128 2115 3212
rect 2205 3188 2211 3212
rect 2301 3168 2307 3332
rect 2333 3288 2339 3292
rect 2349 3268 2355 3312
rect 2365 3308 2371 3412
rect 2381 3308 2387 3332
rect 2365 3288 2371 3292
rect 2093 3097 2115 3103
rect 2077 3088 2083 3092
rect 2077 2963 2083 3072
rect 2077 2957 2099 2963
rect 1981 2888 1987 2892
rect 2045 2763 2051 2832
rect 2077 2788 2083 2832
rect 2029 2757 2051 2763
rect 1912 2717 1932 2723
rect 1805 2548 1811 2552
rect 1901 2528 1907 2692
rect 1917 2548 1923 2632
rect 1949 2568 1955 2692
rect 1965 2688 1971 2692
rect 1981 2668 1987 2692
rect 1933 2528 1939 2532
rect 1789 2408 1795 2512
rect 1773 2377 1784 2383
rect 1773 2188 1779 2272
rect 1757 2148 1763 2152
rect 1789 2148 1795 2232
rect 1805 2108 1811 2112
rect 1805 2088 1811 2092
rect 1805 1908 1811 2032
rect 1821 2028 1827 2512
rect 1997 2388 2003 2732
rect 2013 2588 2019 2652
rect 2029 2528 2035 2757
rect 2045 2728 2051 2732
rect 2077 2688 2083 2732
rect 2061 2528 2067 2652
rect 2093 2568 2099 2957
rect 2109 2888 2115 3097
rect 2125 2968 2131 3032
rect 2157 2988 2163 3112
rect 2173 3088 2179 3092
rect 2189 3048 2195 3072
rect 2205 2988 2211 3052
rect 2221 2948 2227 2952
rect 2200 2937 2211 2943
rect 2109 2748 2115 2872
rect 2125 2828 2131 2932
rect 2125 2708 2131 2752
rect 2141 2728 2147 2732
rect 2157 2688 2163 2832
rect 2189 2728 2195 2852
rect 2205 2848 2211 2937
rect 2237 2928 2243 3112
rect 2301 3068 2307 3092
rect 2253 2948 2259 3032
rect 2205 2688 2211 2752
rect 2109 2588 2115 2632
rect 2045 2488 2051 2512
rect 2061 2488 2067 2512
rect 2109 2388 2115 2452
rect 2125 2428 2131 2532
rect 2141 2528 2147 2592
rect 2173 2588 2179 2612
rect 2221 2588 2227 2912
rect 2237 2728 2243 2732
rect 2253 2728 2259 2852
rect 2269 2828 2275 2952
rect 2301 2908 2307 2972
rect 2317 2948 2323 3032
rect 2349 2988 2355 3092
rect 2381 3088 2387 3272
rect 2397 3028 2403 3632
rect 2413 3488 2419 3692
rect 2493 3688 2499 3712
rect 2589 3668 2595 3712
rect 2653 3708 2659 3712
rect 2429 3468 2435 3472
rect 2413 3308 2419 3352
rect 2413 3208 2419 3292
rect 2429 3188 2435 3292
rect 2429 3108 2435 3112
rect 2445 3088 2451 3612
rect 2509 3508 2515 3532
rect 2541 3508 2547 3632
rect 2605 3628 2611 3632
rect 2461 3388 2467 3472
rect 2461 3368 2467 3372
rect 2477 3328 2483 3492
rect 2493 3308 2499 3472
rect 2509 3348 2515 3472
rect 2557 3408 2563 3472
rect 2525 3328 2531 3352
rect 2573 3268 2579 3492
rect 2605 3428 2611 3452
rect 2621 3248 2627 3472
rect 2557 3228 2563 3232
rect 2285 2688 2291 2872
rect 2301 2788 2307 2892
rect 2317 2888 2323 2912
rect 2349 2888 2355 2892
rect 2381 2888 2387 2952
rect 2397 2928 2403 2952
rect 2429 2948 2435 3052
rect 2216 2537 2227 2543
rect 2189 2517 2200 2523
rect 2189 2503 2195 2517
rect 2221 2503 2227 2537
rect 2173 2497 2195 2503
rect 2205 2497 2227 2503
rect 2173 2468 2179 2497
rect 2189 2388 2195 2452
rect 2205 2388 2211 2497
rect 2237 2408 2243 2632
rect 2253 2448 2259 2632
rect 2285 2588 2291 2652
rect 2269 2568 2275 2572
rect 1901 2268 1907 2332
rect 1944 2317 2003 2323
rect 1997 2303 2003 2317
rect 1997 2297 2008 2303
rect 2029 2268 2035 2272
rect 1885 2248 1891 2252
rect 1901 2128 1907 2252
rect 1933 2248 1939 2252
rect 1965 2188 1971 2212
rect 1933 2148 1939 2152
rect 1981 2148 1987 2232
rect 1997 2148 2003 2232
rect 1944 2137 1955 2143
rect 1741 1808 1747 1832
rect 1709 1797 1731 1803
rect 1725 1783 1731 1797
rect 1725 1777 1736 1783
rect 1597 1728 1603 1732
rect 1549 1703 1555 1712
rect 1512 1697 1555 1703
rect 1565 1648 1571 1692
rect 1389 1428 1395 1452
rect 1309 1348 1315 1392
rect 1421 1348 1427 1492
rect 1437 1348 1443 1452
rect 1453 1428 1459 1512
rect 1485 1508 1491 1592
rect 1517 1528 1523 1532
rect 1469 1408 1475 1472
rect 1485 1348 1491 1432
rect 1197 1248 1203 1312
rect 1293 1308 1299 1312
rect 1341 1308 1347 1312
rect 1277 1288 1283 1292
rect 1229 1048 1235 1052
rect 1165 988 1171 1032
rect 1213 948 1219 992
rect 1229 988 1235 1012
rect 1213 888 1219 932
rect 1245 908 1251 1012
rect 1165 728 1171 832
rect 1197 728 1203 772
rect 1213 768 1219 872
rect 1261 748 1267 1252
rect 1277 1188 1283 1212
rect 1293 1088 1299 1152
rect 1309 1128 1315 1212
rect 1325 1103 1331 1272
rect 1357 1108 1363 1312
rect 1469 1308 1475 1312
rect 1373 1188 1379 1212
rect 1437 1188 1443 1292
rect 1485 1208 1491 1332
rect 1501 1328 1507 1392
rect 1533 1363 1539 1612
rect 1549 1488 1555 1492
rect 1581 1488 1587 1672
rect 1597 1668 1603 1712
rect 1629 1648 1635 1692
rect 1677 1588 1683 1732
rect 1709 1728 1715 1732
rect 1661 1528 1667 1532
rect 1693 1523 1699 1712
rect 1757 1708 1763 1752
rect 1773 1728 1779 1752
rect 1741 1588 1747 1692
rect 1789 1688 1795 1712
rect 1693 1517 1715 1523
rect 1565 1368 1571 1432
rect 1597 1428 1603 1492
rect 1613 1488 1619 1512
rect 1533 1357 1555 1363
rect 1549 1348 1555 1357
rect 1533 1248 1539 1292
rect 1549 1288 1555 1332
rect 1565 1328 1571 1332
rect 1613 1308 1619 1432
rect 1629 1328 1635 1352
rect 1645 1288 1651 1432
rect 1693 1408 1699 1492
rect 1709 1488 1715 1517
rect 1773 1506 1779 1632
rect 1821 1488 1827 2012
rect 1853 1888 1859 2112
rect 1885 1948 1891 2032
rect 1885 1888 1891 1932
rect 1901 1748 1907 1852
rect 1917 1748 1923 1872
rect 1853 1728 1859 1732
rect 1869 1688 1875 1732
rect 1901 1588 1907 1732
rect 1949 1708 1955 2137
rect 1981 2108 1987 2112
rect 1997 1988 2003 2132
rect 2013 2128 2019 2252
rect 2077 2248 2083 2312
rect 2125 2308 2131 2312
rect 2141 2288 2147 2312
rect 2157 2308 2163 2352
rect 2093 2228 2099 2272
rect 2205 2248 2211 2272
rect 2221 2248 2227 2312
rect 2253 2308 2259 2312
rect 2125 2148 2131 2192
rect 2141 2128 2147 2172
rect 2221 2128 2227 2192
rect 2269 2183 2275 2512
rect 2317 2388 2323 2872
rect 2333 2703 2339 2832
rect 2381 2808 2387 2872
rect 2365 2708 2371 2792
rect 2397 2708 2403 2912
rect 2413 2768 2419 2892
rect 2333 2697 2355 2703
rect 2333 2668 2339 2672
rect 2349 2588 2355 2697
rect 2365 2668 2371 2692
rect 2429 2588 2435 2932
rect 2445 2868 2451 2912
rect 2381 2568 2387 2572
rect 2349 2548 2355 2552
rect 2365 2548 2371 2552
rect 2397 2548 2403 2572
rect 2445 2548 2451 2672
rect 2461 2668 2467 3032
rect 2477 2888 2483 2892
rect 2493 2868 2499 3072
rect 2525 3068 2531 3072
rect 2541 3068 2547 3092
rect 2557 3088 2563 3112
rect 2589 3068 2595 3172
rect 2621 3168 2627 3212
rect 2621 3088 2627 3152
rect 2637 3108 2643 3692
rect 2653 3448 2659 3452
rect 2653 3428 2659 3432
rect 2669 3148 2675 3632
rect 2685 3588 2691 3812
rect 2701 3728 2707 3732
rect 2717 3728 2723 3792
rect 2749 3688 2755 3852
rect 2765 3788 2771 4132
rect 2781 3928 2787 3952
rect 2797 3908 2803 4172
rect 2829 4148 2835 4212
rect 2877 4168 2883 4212
rect 2941 4208 2947 4272
rect 3053 4228 3059 4272
rect 3069 4248 3075 4272
rect 2877 4148 2883 4152
rect 2813 4088 2819 4092
rect 2893 4068 2899 4132
rect 2909 3988 2915 4112
rect 2925 4048 2931 4152
rect 3037 4148 3043 4152
rect 2957 4128 2963 4132
rect 2957 4088 2963 4112
rect 2989 4108 2995 4112
rect 2845 3928 2851 3972
rect 2909 3883 2915 3972
rect 2925 3888 2931 4032
rect 3053 4028 3059 4212
rect 3101 4148 3107 4272
rect 3117 4148 3123 4412
rect 3213 4388 3219 4512
rect 3245 4368 3251 4432
rect 3133 4328 3139 4332
rect 3165 4328 3171 4332
rect 3181 4268 3187 4292
rect 3213 4288 3219 4312
rect 3245 4288 3251 4352
rect 3261 4308 3267 4532
rect 3309 4428 3315 4532
rect 3325 4508 3331 4512
rect 3341 4428 3347 4532
rect 3389 4468 3395 4492
rect 3405 4383 3411 4592
rect 3517 4588 3523 4712
rect 3549 4706 3555 4712
rect 3629 4588 3635 4732
rect 3645 4588 3651 4692
rect 3693 4588 3699 4712
rect 3869 4706 3875 4752
rect 3901 4668 3907 4672
rect 3437 4548 3443 4552
rect 3565 4548 3571 4552
rect 3709 4548 3715 4552
rect 3501 4528 3507 4532
rect 3453 4468 3459 4492
rect 3549 4448 3555 4532
rect 3389 4377 3411 4383
rect 3293 4348 3299 4352
rect 3277 4308 3283 4312
rect 3181 4188 3187 4252
rect 3197 4228 3203 4272
rect 3341 4208 3347 4332
rect 3357 4208 3363 4272
rect 3080 4137 3091 4143
rect 3085 4128 3091 4137
rect 3069 4068 3075 4072
rect 2941 3908 2947 3912
rect 2893 3877 2915 3883
rect 2765 3768 2771 3772
rect 2765 3668 2771 3712
rect 2749 3588 2755 3612
rect 2701 3488 2707 3492
rect 2749 3488 2755 3492
rect 2701 3468 2707 3472
rect 2765 3428 2771 3512
rect 2765 3368 2771 3412
rect 2685 3288 2691 3314
rect 2701 3108 2707 3132
rect 2717 3108 2723 3332
rect 2733 3108 2739 3112
rect 2621 3028 2627 3052
rect 2637 2948 2643 2992
rect 2685 2948 2691 3072
rect 2733 3068 2739 3092
rect 2765 2968 2771 3092
rect 2477 2668 2483 2672
rect 2477 2608 2483 2652
rect 2333 2528 2339 2532
rect 2317 2308 2323 2352
rect 2333 2268 2339 2472
rect 2349 2348 2355 2512
rect 2429 2428 2435 2432
rect 2445 2428 2451 2532
rect 2381 2388 2387 2412
rect 2285 2208 2291 2232
rect 2365 2228 2371 2292
rect 2413 2288 2419 2292
rect 2269 2177 2280 2183
rect 2269 2148 2275 2152
rect 2013 2108 2019 2112
rect 2077 2108 2083 2112
rect 2189 2097 2204 2103
rect 2045 2068 2051 2092
rect 2157 2063 2163 2092
rect 2173 2088 2179 2092
rect 2157 2057 2179 2063
rect 1965 1928 1971 1932
rect 2013 1903 2019 2052
rect 2077 1988 2083 2012
rect 2077 1908 2083 1912
rect 2013 1897 2024 1903
rect 1965 1808 1971 1892
rect 1997 1848 2003 1852
rect 1965 1728 1971 1732
rect 1933 1648 1939 1692
rect 1965 1608 1971 1712
rect 1981 1668 1987 1732
rect 1997 1688 2003 1832
rect 2029 1728 2035 1892
rect 2045 1728 2051 1892
rect 2093 1788 2099 1912
rect 2109 1908 2115 2052
rect 2173 1908 2179 2057
rect 2189 1948 2195 2097
rect 2077 1748 2083 1752
rect 2109 1748 2115 1892
rect 2125 1868 2131 1872
rect 2157 1868 2163 1872
rect 1981 1588 1987 1632
rect 2013 1628 2019 1632
rect 2045 1628 2051 1712
rect 2061 1603 2067 1712
rect 2045 1597 2067 1603
rect 2013 1588 2019 1592
rect 2045 1568 2051 1597
rect 2045 1508 2051 1532
rect 1693 1388 1699 1392
rect 1741 1388 1747 1472
rect 1981 1428 1987 1492
rect 1997 1468 2003 1472
rect 1805 1388 1811 1412
rect 2045 1348 2051 1472
rect 2061 1388 2067 1392
rect 2077 1368 2083 1732
rect 1661 1328 1667 1332
rect 1741 1328 1747 1332
rect 1917 1328 1923 1332
rect 1464 1137 1491 1143
rect 1469 1108 1475 1112
rect 1320 1097 1331 1103
rect 1485 1103 1491 1137
rect 1533 1128 1539 1232
rect 1485 1097 1496 1103
rect 1277 988 1283 992
rect 1309 948 1315 1092
rect 1325 1028 1331 1072
rect 1357 1048 1363 1072
rect 1373 1068 1379 1092
rect 1405 988 1411 1052
rect 1421 1008 1427 1072
rect 1469 1068 1475 1072
rect 1565 1068 1571 1092
rect 1533 988 1539 1012
rect 1549 988 1555 992
rect 1341 828 1347 832
rect 1261 728 1267 732
rect 1309 688 1315 792
rect 1357 788 1363 972
rect 1373 928 1379 932
rect 1373 908 1379 912
rect 1389 808 1395 932
rect 1405 868 1411 912
rect 1437 908 1443 912
rect 1453 883 1459 932
rect 1469 928 1475 972
rect 1549 948 1555 972
rect 1501 908 1507 932
rect 1565 928 1571 992
rect 1613 988 1619 1092
rect 1645 1088 1651 1092
rect 1661 1028 1667 1112
rect 1581 948 1587 952
rect 1613 888 1619 932
rect 1645 908 1651 932
rect 1677 928 1683 1052
rect 1693 1028 1699 1132
rect 1741 1088 1747 1312
rect 1789 1268 1795 1312
rect 2029 1288 2035 1312
rect 1869 1108 1875 1272
rect 1981 1108 1987 1232
rect 2045 1188 2051 1332
rect 2077 1188 2083 1332
rect 2029 1108 2035 1112
rect 2045 1108 2051 1172
rect 2093 1108 2099 1712
rect 2109 1608 2115 1732
rect 2125 1728 2131 1792
rect 2157 1728 2163 1832
rect 2173 1688 2179 1872
rect 2205 1808 2211 2072
rect 2237 1948 2243 2092
rect 2253 2068 2259 2112
rect 2269 2008 2275 2132
rect 2333 2088 2339 2112
rect 2333 1988 2339 1992
rect 2269 1948 2275 1952
rect 2365 1948 2371 2132
rect 2397 2128 2403 2232
rect 2413 2188 2419 2212
rect 2413 1988 2419 1992
rect 2429 1948 2435 2112
rect 2445 2008 2451 2292
rect 2461 2263 2467 2532
rect 2477 2508 2483 2532
rect 2493 2503 2499 2832
rect 2509 2828 2515 2832
rect 2509 2668 2515 2692
rect 2525 2608 2531 2932
rect 2541 2928 2547 2932
rect 2557 2868 2563 2912
rect 2589 2888 2595 2892
rect 2573 2688 2579 2732
rect 2589 2628 2595 2692
rect 2637 2688 2643 2932
rect 2621 2668 2627 2672
rect 2669 2668 2675 2912
rect 2685 2828 2691 2872
rect 2733 2788 2739 2912
rect 2765 2908 2771 2914
rect 2712 2717 2723 2723
rect 2717 2708 2723 2717
rect 2733 2708 2739 2752
rect 2749 2688 2755 2792
rect 2781 2788 2787 3872
rect 2893 3808 2899 3877
rect 2957 3868 2963 3932
rect 2973 3908 2979 3932
rect 2989 3868 2995 3912
rect 3005 3908 3011 3952
rect 3021 3888 3027 4012
rect 3117 3968 3123 4132
rect 2893 3768 2899 3792
rect 3021 3788 3027 3872
rect 3037 3788 3043 3952
rect 3085 3928 3091 3932
rect 3133 3928 3139 4172
rect 3165 4108 3171 4112
rect 3197 4108 3203 4112
rect 3165 4068 3171 4092
rect 3213 4088 3219 4132
rect 3261 4108 3267 4112
rect 3213 3963 3219 4072
rect 3229 3988 3235 4092
rect 3277 3988 3283 4132
rect 3325 4128 3331 4172
rect 3389 4168 3395 4377
rect 3421 4168 3427 4192
rect 3453 4188 3459 4392
rect 3485 4308 3491 4312
rect 3581 4268 3587 4512
rect 3661 4428 3667 4532
rect 3677 4448 3683 4532
rect 3709 4468 3715 4472
rect 3565 4183 3571 4232
rect 3565 4177 3587 4183
rect 3373 4103 3379 4112
rect 3324 4097 3379 4103
rect 3213 3957 3235 3963
rect 3149 3928 3155 3932
rect 3165 3928 3171 3932
rect 3133 3908 3139 3912
rect 3053 3888 3059 3892
rect 3197 3888 3203 3912
rect 3053 3808 3059 3872
rect 2829 3748 2835 3752
rect 2797 3608 2803 3632
rect 2925 3608 2931 3632
rect 2957 3548 2963 3692
rect 2925 3508 2931 3512
rect 2941 3488 2947 3512
rect 2797 3308 2803 3432
rect 2893 3408 2899 3432
rect 2973 3428 2979 3472
rect 2989 3448 2995 3712
rect 3005 3668 3011 3732
rect 3037 3588 3043 3732
rect 3069 3708 3075 3712
rect 3085 3703 3091 3712
rect 3085 3697 3096 3703
rect 3133 3628 3139 3872
rect 3229 3788 3235 3957
rect 3245 3888 3251 3952
rect 3213 3728 3219 3752
rect 3293 3748 3299 4092
rect 3341 3908 3347 4032
rect 3389 3823 3395 4032
rect 3469 3908 3475 4092
rect 3485 4068 3491 4112
rect 3501 4088 3507 4112
rect 3565 4088 3571 4112
rect 3581 4088 3587 4177
rect 3629 4143 3635 4212
rect 3645 4168 3651 4312
rect 3661 4268 3667 4412
rect 3677 4308 3683 4372
rect 3725 4308 3731 4652
rect 3757 4468 3763 4512
rect 3773 4388 3779 4452
rect 3789 4348 3795 4532
rect 3837 4528 3843 4592
rect 3869 4548 3875 4552
rect 3805 4408 3811 4512
rect 3821 4508 3827 4512
rect 3725 4288 3731 4292
rect 3624 4137 3640 4143
rect 3661 4048 3667 4252
rect 3725 4148 3731 4152
rect 3469 3888 3475 3892
rect 3389 3817 3411 3823
rect 3309 3788 3315 3792
rect 3149 3648 3155 3712
rect 3277 3688 3283 3712
rect 3101 3588 3107 3612
rect 3021 3528 3027 3532
rect 3149 3528 3155 3592
rect 3181 3568 3187 3632
rect 3245 3568 3251 3672
rect 3357 3568 3363 3632
rect 3192 3537 3208 3543
rect 3165 3508 3171 3512
rect 3021 3488 3027 3492
rect 3069 3468 3075 3492
rect 2813 3328 2819 3352
rect 2861 3348 2867 3372
rect 2845 3108 2851 3132
rect 2797 3008 2803 3072
rect 2797 2708 2803 2932
rect 2813 2708 2819 2952
rect 2829 2748 2835 3072
rect 2861 2968 2867 3012
rect 2909 2968 2915 3332
rect 2925 3188 2931 3312
rect 2941 3048 2947 3132
rect 2989 3108 2995 3432
rect 3085 3388 3091 3412
rect 3101 3363 3107 3472
rect 3133 3468 3139 3492
rect 3085 3357 3107 3363
rect 3021 3248 3027 3292
rect 3021 3148 3027 3232
rect 3053 3108 3059 3312
rect 3085 3308 3091 3357
rect 3085 3168 3091 3292
rect 3069 3108 3075 3132
rect 3037 3088 3043 3092
rect 2957 3028 2963 3072
rect 3053 3068 3059 3072
rect 2909 2828 2915 2832
rect 2925 2768 2931 2872
rect 2941 2868 2947 2932
rect 2957 2928 2963 2992
rect 3005 2948 3011 3052
rect 3053 2988 3059 2992
rect 3101 2988 3107 3232
rect 3117 3128 3123 3312
rect 3133 3103 3139 3192
rect 3117 3097 3139 3103
rect 3037 2968 3043 2972
rect 2989 2908 2995 2912
rect 3069 2888 3075 2952
rect 3101 2948 3107 2972
rect 3085 2928 3091 2932
rect 3085 2908 3091 2912
rect 2957 2728 2963 2812
rect 3101 2808 3107 2832
rect 2605 2648 2611 2652
rect 2685 2648 2691 2652
rect 2557 2548 2563 2592
rect 2701 2537 2712 2543
rect 2589 2508 2595 2512
rect 2493 2497 2515 2503
rect 2493 2288 2499 2292
rect 2461 2257 2472 2263
rect 2472 2157 2483 2163
rect 2461 2128 2467 2132
rect 2477 2088 2483 2157
rect 2509 1988 2515 2497
rect 2541 2428 2547 2432
rect 2605 2248 2611 2532
rect 2701 2528 2707 2537
rect 2765 2528 2771 2552
rect 2797 2548 2803 2652
rect 2829 2548 2835 2572
rect 2877 2568 2883 2692
rect 2909 2668 2915 2672
rect 2925 2657 2968 2663
rect 2925 2643 2931 2657
rect 2904 2637 2931 2643
rect 2957 2548 2963 2572
rect 2973 2548 2979 2552
rect 2829 2528 2835 2532
rect 2621 2488 2627 2512
rect 2669 2488 2675 2492
rect 2637 2306 2643 2412
rect 2701 2408 2707 2512
rect 2717 2468 2723 2512
rect 2813 2503 2819 2512
rect 2845 2503 2851 2512
rect 2813 2497 2851 2503
rect 2733 2388 2739 2492
rect 2797 2488 2803 2492
rect 2861 2488 2867 2532
rect 2909 2508 2915 2532
rect 2989 2528 2995 2652
rect 3005 2637 3016 2643
rect 3005 2528 3011 2637
rect 2813 2468 2819 2472
rect 2733 2328 2739 2372
rect 2781 2308 2787 2432
rect 2813 2388 2819 2452
rect 2813 2368 2819 2372
rect 2701 2288 2707 2292
rect 2701 2148 2707 2272
rect 2253 1917 2264 1923
rect 2205 1728 2211 1792
rect 2237 1728 2243 1832
rect 2253 1788 2259 1917
rect 2269 1848 2275 1872
rect 2317 1768 2323 1772
rect 2253 1748 2259 1752
rect 2317 1728 2323 1752
rect 2333 1748 2339 1932
rect 2381 1888 2387 1932
rect 2429 1908 2435 1932
rect 2557 1908 2563 2052
rect 2621 1928 2627 2132
rect 2605 1908 2611 1912
rect 2477 1868 2483 1892
rect 2349 1848 2355 1852
rect 2365 1788 2371 1852
rect 2365 1748 2371 1772
rect 2189 1708 2195 1712
rect 2285 1648 2291 1692
rect 2349 1668 2355 1732
rect 2109 1388 2115 1572
rect 2141 1506 2147 1632
rect 2205 1488 2211 1492
rect 2221 1488 2227 1492
rect 2269 1488 2275 1552
rect 2285 1508 2291 1572
rect 2317 1528 2323 1632
rect 2349 1588 2355 1652
rect 2365 1548 2371 1632
rect 2381 1528 2387 1832
rect 2397 1728 2403 1732
rect 2413 1728 2419 1832
rect 2493 1808 2499 1892
rect 2541 1848 2547 1872
rect 2445 1788 2451 1792
rect 2493 1788 2499 1792
rect 2461 1588 2467 1772
rect 2365 1508 2371 1512
rect 2173 1443 2179 1472
rect 2173 1437 2195 1443
rect 2109 1328 2115 1352
rect 2125 1337 2136 1343
rect 2109 1188 2115 1292
rect 2125 1268 2131 1337
rect 1965 1088 1971 1092
rect 1997 1048 2003 1072
rect 1773 988 1779 1012
rect 1693 928 1699 932
rect 1437 877 1459 883
rect 1405 828 1411 852
rect 1341 708 1347 732
rect 1384 697 1400 703
rect 1037 648 1043 652
rect 1037 548 1043 632
rect 637 283 643 412
rect 653 308 659 432
rect 669 368 675 372
rect 941 368 947 492
rect 989 468 995 472
rect 669 288 675 352
rect 717 308 723 312
rect 637 277 648 283
rect 717 268 723 272
rect 301 117 312 123
rect 253 -43 275 -37
rect 349 -43 355 32
rect 429 -43 435 132
rect 493 88 499 232
rect 541 108 547 232
rect 621 148 627 232
rect 669 128 675 152
rect 605 68 611 114
rect 701 88 707 232
rect 733 188 739 332
rect 941 328 947 352
rect 749 308 755 312
rect 781 188 787 312
rect 813 308 819 312
rect 861 288 867 312
rect 781 148 787 172
rect 797 108 803 272
rect 877 268 883 272
rect 893 228 899 292
rect 925 248 931 312
rect 973 288 979 312
rect 909 168 915 172
rect 941 68 947 232
rect 989 228 995 272
rect 989 188 995 212
rect 1021 188 1027 512
rect 1053 408 1059 572
rect 1053 328 1059 392
rect 1069 388 1075 672
rect 1085 588 1091 592
rect 1101 588 1107 672
rect 1117 588 1123 612
rect 1133 528 1139 612
rect 1149 548 1155 552
rect 1165 523 1171 652
rect 1245 608 1251 672
rect 1309 623 1315 672
rect 1293 617 1315 623
rect 1405 657 1416 663
rect 1213 548 1219 552
rect 1181 528 1187 532
rect 1197 528 1203 532
rect 1149 517 1171 523
rect 1085 468 1091 512
rect 1101 468 1107 492
rect 1037 248 1043 312
rect 1005 128 1011 152
rect 1037 148 1043 212
rect 1053 148 1059 312
rect 1069 288 1075 372
rect 1149 348 1155 517
rect 1229 508 1235 572
rect 1293 548 1299 617
rect 1309 588 1315 592
rect 1261 528 1267 532
rect 1165 468 1171 492
rect 1101 288 1107 312
rect 1165 308 1171 312
rect 1069 208 1075 272
rect 1085 168 1091 232
rect 1117 208 1123 292
rect 1101 148 1107 192
rect 1037 128 1043 132
rect 1149 128 1155 292
rect 1181 288 1187 332
rect 1245 328 1251 352
rect 1197 288 1203 312
rect 1261 288 1267 372
rect 1277 288 1283 532
rect 1293 348 1299 532
rect 1309 288 1315 392
rect 1325 308 1331 432
rect 1341 328 1347 512
rect 1341 308 1347 312
rect 1277 203 1283 272
rect 1325 268 1331 272
rect 1357 248 1363 512
rect 1405 448 1411 657
rect 1421 548 1427 572
rect 1437 568 1443 877
rect 1453 868 1459 877
rect 1453 788 1459 812
rect 1501 683 1507 712
rect 1549 688 1555 812
rect 1581 788 1587 832
rect 1613 768 1619 872
rect 1485 677 1507 683
rect 1389 328 1395 352
rect 1261 197 1283 203
rect 1181 148 1187 152
rect 1261 148 1267 197
rect 1277 148 1283 197
rect 1165 128 1171 132
rect 1277 128 1283 132
rect 1021 108 1027 112
rect 1277 108 1283 112
rect 1293 108 1299 232
rect 1341 148 1347 172
rect 1389 148 1395 152
rect 1421 148 1427 532
rect 1469 508 1475 552
rect 1437 328 1443 432
rect 1453 283 1459 492
rect 1469 328 1475 492
rect 1485 448 1491 677
rect 1501 568 1507 632
rect 1613 588 1619 752
rect 1629 708 1635 872
rect 1693 868 1699 912
rect 1709 908 1715 932
rect 1740 897 1768 903
rect 1805 828 1811 932
rect 1853 908 1859 912
rect 1885 848 1891 852
rect 1693 688 1699 812
rect 1773 728 1779 732
rect 1789 728 1795 732
rect 1853 728 1859 732
rect 1757 688 1763 692
rect 1821 688 1827 692
rect 1741 668 1747 672
rect 1805 628 1811 672
rect 1805 548 1811 552
rect 1613 388 1619 512
rect 1581 308 1587 312
rect 1805 308 1811 532
rect 1885 508 1891 832
rect 1901 548 1907 932
rect 1965 788 1971 914
rect 1933 688 1939 752
rect 1949 648 1955 732
rect 2013 708 2019 992
rect 2029 928 2035 952
rect 2061 728 2067 892
rect 1965 688 1971 692
rect 1965 508 1971 532
rect 1997 508 2003 592
rect 1821 308 1827 432
rect 1981 308 1987 352
rect 1997 328 2003 472
rect 2077 368 2083 1092
rect 2125 1028 2131 1032
rect 2141 988 2147 1312
rect 2173 1188 2179 1412
rect 2189 1408 2195 1437
rect 2189 1388 2195 1392
rect 2205 1348 2211 1352
rect 2253 1308 2259 1432
rect 2173 1008 2179 1032
rect 2189 968 2195 1232
rect 2205 1108 2211 1152
rect 2285 1108 2291 1112
rect 2221 1088 2227 1092
rect 2285 1088 2291 1092
rect 2109 928 2115 932
rect 2125 928 2131 932
rect 2093 888 2099 892
rect 2109 708 2115 712
rect 2125 688 2131 832
rect 2157 828 2163 932
rect 2173 908 2179 912
rect 2189 688 2195 812
rect 2205 708 2211 892
rect 2221 888 2227 912
rect 2221 748 2227 832
rect 2237 768 2243 1072
rect 2253 1048 2259 1052
rect 2221 708 2227 712
rect 2141 648 2147 672
rect 2157 668 2163 672
rect 2109 508 2115 552
rect 2141 528 2147 572
rect 2157 468 2163 532
rect 2173 528 2179 632
rect 2189 548 2195 632
rect 2221 608 2227 632
rect 2237 548 2243 752
rect 2253 708 2259 1032
rect 2317 968 2323 1452
rect 2349 1383 2355 1432
rect 2381 1388 2387 1512
rect 2413 1488 2419 1492
rect 2429 1468 2435 1472
rect 2477 1468 2483 1712
rect 2557 1568 2563 1892
rect 2573 1888 2579 1892
rect 2621 1888 2627 1912
rect 2637 1908 2643 1932
rect 2605 1748 2611 1832
rect 2653 1748 2659 2132
rect 2696 1917 2707 1923
rect 2685 1888 2691 1892
rect 2701 1888 2707 1917
rect 2733 1888 2739 1912
rect 2749 1868 2755 2112
rect 2765 1968 2771 2232
rect 2781 2088 2787 2092
rect 2813 1948 2819 2112
rect 2765 1908 2771 1932
rect 2781 1848 2787 1872
rect 2621 1648 2627 1714
rect 2653 1568 2659 1732
rect 2685 1708 2691 1732
rect 2701 1728 2707 1732
rect 2717 1688 2723 1832
rect 2813 1823 2819 1892
rect 2797 1817 2819 1823
rect 2749 1808 2755 1812
rect 2749 1728 2755 1792
rect 2797 1768 2803 1817
rect 2813 1808 2819 1817
rect 2829 1768 2835 2412
rect 2845 2308 2851 2452
rect 2957 2388 2963 2512
rect 3021 2508 3027 2512
rect 2909 2308 2915 2312
rect 2957 2308 2963 2332
rect 3021 2308 3027 2492
rect 3037 2468 3043 2712
rect 3069 2688 3075 2792
rect 3085 2728 3091 2752
rect 3101 2708 3107 2732
rect 3117 2708 3123 3097
rect 3149 2948 3155 3112
rect 3165 3088 3171 3432
rect 3181 3308 3187 3432
rect 3181 3148 3187 3232
rect 3181 3108 3187 3132
rect 3197 3108 3203 3112
rect 3133 2888 3139 2932
rect 3165 2928 3171 3072
rect 3213 3068 3219 3472
rect 3229 3348 3235 3352
rect 3245 3328 3251 3552
rect 3261 3528 3267 3532
rect 3261 3428 3267 3512
rect 3357 3508 3363 3512
rect 3336 3497 3347 3503
rect 3341 3488 3347 3497
rect 3373 3488 3379 3792
rect 3389 3648 3395 3712
rect 3405 3708 3411 3817
rect 3485 3748 3491 3752
rect 3405 3528 3411 3532
rect 3309 3448 3315 3472
rect 3229 3288 3235 3312
rect 3277 3308 3283 3332
rect 3293 3328 3299 3412
rect 3309 3328 3315 3332
rect 3325 3328 3331 3472
rect 3245 3108 3251 3292
rect 3293 3188 3299 3312
rect 3293 3128 3299 3132
rect 3245 3088 3251 3092
rect 3245 3003 3251 3072
rect 3261 3008 3267 3092
rect 3229 2997 3251 3003
rect 3197 2923 3203 2992
rect 3229 2948 3235 2997
rect 3293 2948 3299 3092
rect 3309 3088 3315 3092
rect 3325 3008 3331 3092
rect 3341 3028 3347 3332
rect 3373 3308 3379 3432
rect 3421 3408 3427 3632
rect 3437 3508 3443 3652
rect 3421 3348 3427 3352
rect 3405 3208 3411 3312
rect 3437 3288 3443 3312
rect 3453 3268 3459 3472
rect 3469 3428 3475 3432
rect 3485 3408 3491 3712
rect 3501 3348 3507 4032
rect 3533 4028 3539 4032
rect 3517 3868 3523 3892
rect 3533 3868 3539 3972
rect 3629 3888 3635 4032
rect 3661 3988 3667 4032
rect 3677 4008 3683 4112
rect 3709 4008 3715 4092
rect 3677 3888 3683 3992
rect 3725 3968 3731 4132
rect 3741 3948 3747 4032
rect 3757 3988 3763 4272
rect 3549 3768 3555 3832
rect 3581 3748 3587 3772
rect 3597 3728 3603 3792
rect 3629 3708 3635 3832
rect 3677 3748 3683 3752
rect 3693 3688 3699 3892
rect 3709 3868 3715 3872
rect 3757 3848 3763 3912
rect 3773 3908 3779 4292
rect 3805 4228 3811 4352
rect 3821 4328 3827 4332
rect 3821 4268 3827 4272
rect 3789 4148 3795 4192
rect 3805 4148 3811 4212
rect 3821 4128 3827 4132
rect 3805 4103 3811 4112
rect 3805 4097 3827 4103
rect 3789 3908 3795 3912
rect 3805 3888 3811 4012
rect 3821 3928 3827 4097
rect 3709 3728 3715 3772
rect 3725 3688 3731 3832
rect 3821 3768 3827 3912
rect 3837 3823 3843 4292
rect 3869 4208 3875 4532
rect 3901 4528 3907 4532
rect 3949 4448 3955 4672
rect 3997 4588 4003 4712
rect 4109 4568 4115 4612
rect 4125 4588 4131 4692
rect 4109 4548 4115 4552
rect 4141 4548 4147 4672
rect 4189 4668 4195 4692
rect 4285 4628 4291 4672
rect 4301 4588 4307 4732
rect 4333 4588 4339 4692
rect 4365 4588 4371 4732
rect 4381 4708 4387 4712
rect 4413 4568 4419 4712
rect 4253 4548 4259 4552
rect 4013 4488 4019 4532
rect 4029 4468 4035 4492
rect 4061 4448 4067 4512
rect 4077 4508 4083 4532
rect 3917 4328 3923 4332
rect 3885 4308 3891 4312
rect 3869 4148 3875 4192
rect 3933 4188 3939 4292
rect 3949 4248 3955 4312
rect 3965 4283 3971 4312
rect 3965 4277 3987 4283
rect 3949 4148 3955 4152
rect 3853 4028 3859 4092
rect 3853 4008 3859 4012
rect 3869 4008 3875 4112
rect 3901 4108 3907 4112
rect 3901 4088 3907 4092
rect 3853 3988 3859 3992
rect 3869 3888 3875 3972
rect 3901 3868 3907 3892
rect 3917 3888 3923 4132
rect 3965 3888 3971 4132
rect 3981 4108 3987 4277
rect 3997 4148 4003 4292
rect 4029 4288 4035 4432
rect 4077 4368 4083 4492
rect 4093 4348 4099 4512
rect 4221 4508 4227 4532
rect 4269 4508 4275 4512
rect 4173 4468 4179 4492
rect 4013 4268 4019 4272
rect 4029 4228 4035 4272
rect 4093 4148 4099 4272
rect 4125 4208 4131 4272
rect 4189 4248 4195 4292
rect 4125 4188 4131 4192
rect 4141 4148 4147 4172
rect 4077 4128 4083 4132
rect 3981 4088 3987 4092
rect 3837 3817 3859 3823
rect 3853 3748 3859 3817
rect 3933 3788 3939 3872
rect 3965 3828 3971 3872
rect 3869 3728 3875 3732
rect 3981 3728 3987 3852
rect 3997 3848 4003 3912
rect 4013 3883 4019 4092
rect 4029 3908 4035 4112
rect 4045 3888 4051 3912
rect 4013 3877 4035 3883
rect 4029 3748 4035 3877
rect 4061 3868 4067 3912
rect 4093 3908 4099 4132
rect 4109 4068 4115 4112
rect 4173 4108 4179 4112
rect 4093 3868 4099 3892
rect 4109 3888 4115 3972
rect 4157 3948 4163 3992
rect 3597 3348 3603 3472
rect 3629 3348 3635 3612
rect 3741 3568 3747 3632
rect 3757 3628 3763 3632
rect 3981 3608 3987 3712
rect 3997 3688 4003 3732
rect 4077 3728 4083 3752
rect 4125 3748 4131 3892
rect 4141 3868 4147 3932
rect 4189 3728 4195 4232
rect 4205 4188 4211 4472
rect 4237 4468 4243 4492
rect 4221 4228 4227 4352
rect 4237 4308 4243 4432
rect 4285 4323 4291 4532
rect 4301 4508 4307 4552
rect 4269 4317 4291 4323
rect 4237 4288 4243 4292
rect 4269 4288 4275 4317
rect 4285 4248 4291 4292
rect 4221 3968 4227 4212
rect 4237 4128 4243 4232
rect 4285 4083 4291 4232
rect 4269 4077 4291 4083
rect 4221 3888 4227 3952
rect 4237 3888 4243 4032
rect 4221 3808 4227 3872
rect 4125 3708 4131 3712
rect 4061 3688 4067 3692
rect 3773 3557 3784 3563
rect 3693 3528 3699 3532
rect 3661 3468 3667 3472
rect 3677 3368 3683 3492
rect 3709 3448 3715 3512
rect 3773 3508 3779 3557
rect 3565 3328 3571 3332
rect 3517 3228 3523 3232
rect 3533 3208 3539 3292
rect 3549 3288 3555 3312
rect 3549 3248 3555 3272
rect 3565 3188 3571 3312
rect 3597 3308 3603 3312
rect 3613 3308 3619 3312
rect 3373 3088 3379 3152
rect 3357 2968 3363 2972
rect 3405 2948 3411 3012
rect 3437 2948 3443 3032
rect 3453 3028 3459 3072
rect 3485 3063 3491 3072
rect 3469 3057 3491 3063
rect 3469 2988 3475 3057
rect 3389 2928 3395 2932
rect 3197 2917 3208 2923
rect 3149 2908 3155 2912
rect 3181 2908 3187 2912
rect 3053 2628 3059 2632
rect 3053 2548 3059 2572
rect 3101 2548 3107 2672
rect 3117 2568 3123 2692
rect 3133 2688 3139 2852
rect 3149 2808 3155 2892
rect 3149 2708 3155 2732
rect 3165 2688 3171 2752
rect 3101 2508 3107 2532
rect 3149 2528 3155 2552
rect 3117 2488 3123 2492
rect 3037 2428 3043 2452
rect 2925 2297 2936 2303
rect 2861 2268 2867 2292
rect 2893 2288 2899 2292
rect 2845 2108 2851 2112
rect 2893 2068 2899 2132
rect 2925 1948 2931 2297
rect 2941 2168 2947 2272
rect 3037 2148 3043 2312
rect 3085 2306 3091 2372
rect 3149 2348 3155 2512
rect 3165 2508 3171 2532
rect 3181 2388 3187 2432
rect 3197 2328 3203 2917
rect 3261 2917 3272 2923
rect 3213 2708 3219 2812
rect 3229 2688 3235 2872
rect 3213 2628 3219 2672
rect 3261 2668 3267 2917
rect 3277 2688 3283 2812
rect 3309 2788 3315 2832
rect 3325 2788 3331 2852
rect 3405 2768 3411 2932
rect 3421 2728 3427 2912
rect 3437 2908 3443 2932
rect 3437 2788 3443 2892
rect 3485 2748 3491 3032
rect 3501 3028 3507 3092
rect 3533 3048 3539 3052
rect 3501 2928 3507 3012
rect 3565 3008 3571 3172
rect 3597 3108 3603 3112
rect 3629 3088 3635 3332
rect 3645 3328 3651 3352
rect 3693 3348 3699 3352
rect 3709 3328 3715 3332
rect 3661 3308 3667 3312
rect 3693 3188 3699 3252
rect 3725 3108 3731 3452
rect 3789 3388 3795 3492
rect 3837 3388 3843 3392
rect 3853 3283 3859 3452
rect 3917 3448 3923 3512
rect 3949 3368 3955 3492
rect 3965 3488 3971 3512
rect 3997 3488 4003 3512
rect 4045 3508 4051 3552
rect 3965 3348 3971 3352
rect 3949 3328 3955 3332
rect 3869 3308 3875 3312
rect 3901 3288 3907 3292
rect 3848 3277 3859 3283
rect 3933 3263 3939 3312
rect 3933 3257 3955 3263
rect 3805 3108 3811 3192
rect 3933 3188 3939 3232
rect 3901 3108 3907 3112
rect 3752 3097 3763 3103
rect 3677 3088 3683 3092
rect 3629 3028 3635 3032
rect 3389 2688 3395 2692
rect 3213 2588 3219 2612
rect 3245 2548 3251 2592
rect 3213 2468 3219 2512
rect 3229 2468 3235 2492
rect 3261 2408 3267 2632
rect 3533 2628 3539 2992
rect 3565 2948 3571 2952
rect 3661 2948 3667 3072
rect 3581 2728 3587 2912
rect 3661 2828 3667 2832
rect 3597 2808 3603 2812
rect 3549 2588 3555 2692
rect 3453 2548 3459 2572
rect 3485 2548 3491 2552
rect 3533 2548 3539 2572
rect 3149 2288 3155 2312
rect 2941 2028 2947 2132
rect 3117 2128 3123 2172
rect 3133 2148 3139 2212
rect 2957 2108 2963 2112
rect 3005 2088 3011 2112
rect 3085 2108 3091 2112
rect 3165 2108 3171 2312
rect 3213 2308 3219 2352
rect 3229 2308 3235 2332
rect 3197 2288 3203 2292
rect 3261 2288 3267 2352
rect 3277 2308 3283 2532
rect 3325 2528 3331 2532
rect 3325 2508 3331 2512
rect 3293 2488 3299 2492
rect 3325 2408 3331 2492
rect 3021 2068 3027 2092
rect 3085 2088 3091 2092
rect 3149 2088 3155 2092
rect 2845 1928 2851 1932
rect 2845 1888 2851 1912
rect 2861 1868 2867 1892
rect 2845 1743 2851 1832
rect 2829 1737 2851 1743
rect 2765 1728 2771 1732
rect 2829 1728 2835 1737
rect 2861 1728 2867 1852
rect 2893 1788 2899 1872
rect 2493 1508 2499 1512
rect 2509 1483 2515 1512
rect 2525 1508 2531 1532
rect 2701 1528 2707 1612
rect 2765 1548 2771 1712
rect 2861 1708 2867 1712
rect 2861 1688 2867 1692
rect 2909 1568 2915 1632
rect 2493 1477 2515 1483
rect 2429 1448 2435 1452
rect 2413 1388 2419 1432
rect 2349 1377 2371 1383
rect 2365 1343 2371 1377
rect 2365 1337 2387 1343
rect 2381 1308 2387 1337
rect 2349 1288 2355 1292
rect 2477 1248 2483 1252
rect 2365 1108 2371 1112
rect 2461 1108 2467 1112
rect 2317 788 2323 952
rect 2333 748 2339 972
rect 2413 968 2419 1092
rect 2445 968 2451 1052
rect 2477 968 2483 1232
rect 2493 1228 2499 1477
rect 2509 1188 2515 1312
rect 2541 1208 2547 1512
rect 2621 1508 2627 1512
rect 2701 1508 2707 1512
rect 2685 1488 2691 1492
rect 2781 1488 2787 1552
rect 2861 1508 2867 1552
rect 2589 1428 2595 1432
rect 2589 1328 2595 1392
rect 2605 1328 2611 1352
rect 2925 1348 2931 1852
rect 2941 1828 2947 1912
rect 2957 1888 2963 2052
rect 2957 1868 2963 1872
rect 2941 1728 2947 1752
rect 2973 1743 2979 1832
rect 2989 1748 2995 2012
rect 3165 1988 3171 2092
rect 3181 2088 3187 2232
rect 3197 2128 3203 2232
rect 3309 2228 3315 2312
rect 3341 2268 3347 2532
rect 3549 2523 3555 2552
rect 3581 2548 3587 2612
rect 3597 2528 3603 2792
rect 3629 2728 3635 2732
rect 3693 2728 3699 2752
rect 3677 2688 3683 2692
rect 3544 2517 3555 2523
rect 3373 2508 3379 2512
rect 3501 2508 3507 2512
rect 3357 2488 3363 2492
rect 3469 2488 3475 2492
rect 3405 2388 3411 2472
rect 3469 2468 3475 2472
rect 3357 2288 3363 2312
rect 3533 2308 3539 2352
rect 3597 2328 3603 2512
rect 3613 2388 3619 2532
rect 3629 2508 3635 2512
rect 3645 2488 3651 2512
rect 3661 2468 3667 2492
rect 3677 2468 3683 2672
rect 3709 2528 3715 2672
rect 3725 2628 3731 3092
rect 3757 3068 3763 3097
rect 3805 3048 3811 3092
rect 3837 2983 3843 3032
rect 3949 3028 3955 3257
rect 3965 3088 3971 3152
rect 3997 3108 4003 3272
rect 4013 3128 4019 3252
rect 3981 3088 3987 3092
rect 4029 3088 4035 3092
rect 3821 2977 3843 2983
rect 3821 2948 3827 2977
rect 3821 2928 3827 2932
rect 3741 2708 3747 2832
rect 3789 2788 3795 2914
rect 3757 2737 3768 2743
rect 3741 2668 3747 2672
rect 3757 2588 3763 2737
rect 3805 2588 3811 2712
rect 3837 2688 3843 2812
rect 3869 2688 3875 2872
rect 3885 2748 3891 2832
rect 3885 2708 3891 2732
rect 3933 2688 3939 2692
rect 3869 2588 3875 2632
rect 3773 2548 3779 2552
rect 3837 2548 3843 2552
rect 3725 2528 3731 2532
rect 3693 2508 3699 2512
rect 3629 2328 3635 2392
rect 3629 2288 3635 2312
rect 3405 2277 3416 2283
rect 3213 2148 3219 2172
rect 3245 2148 3251 2172
rect 3213 2108 3219 2112
rect 3261 2068 3267 2152
rect 3325 2143 3331 2232
rect 3341 2148 3347 2152
rect 3405 2148 3411 2277
rect 3309 2137 3331 2143
rect 3309 2108 3315 2137
rect 3336 2117 3347 2123
rect 3341 2108 3347 2117
rect 3069 1928 3075 1932
rect 3005 1888 3011 1912
rect 3037 1908 3043 1912
rect 3101 1908 3107 1972
rect 3181 1908 3187 1952
rect 3053 1768 3059 1872
rect 2957 1737 2979 1743
rect 2957 1708 2963 1737
rect 2957 1548 2963 1672
rect 2973 1588 2979 1712
rect 2941 1348 2947 1392
rect 2973 1348 2979 1532
rect 2989 1388 2995 1472
rect 3021 1408 3027 1732
rect 3069 1703 3075 1872
rect 3101 1808 3107 1892
rect 3213 1888 3219 1952
rect 3261 1908 3267 2052
rect 3325 1968 3331 1972
rect 3325 1888 3331 1952
rect 3341 1948 3347 2092
rect 3373 1968 3379 2132
rect 3405 2088 3411 2132
rect 3421 2128 3427 2252
rect 3453 2188 3459 2212
rect 3469 2128 3475 2132
rect 3341 1908 3347 1932
rect 3197 1848 3203 1852
rect 3085 1728 3091 1792
rect 3117 1748 3123 1752
rect 3064 1697 3075 1703
rect 3053 1523 3059 1692
rect 3117 1648 3123 1732
rect 3133 1728 3139 1812
rect 3197 1748 3203 1832
rect 3245 1748 3251 1872
rect 3261 1788 3267 1872
rect 3048 1517 3059 1523
rect 3117 1508 3123 1632
rect 3085 1488 3091 1492
rect 3069 1348 3075 1372
rect 2493 1028 2499 1092
rect 2509 1088 2515 1092
rect 2573 1088 2579 1092
rect 2349 888 2355 912
rect 2381 908 2387 912
rect 2365 868 2371 892
rect 2413 848 2419 932
rect 2253 668 2259 672
rect 2253 568 2259 652
rect 2269 548 2275 632
rect 2173 488 2179 512
rect 2189 508 2195 512
rect 1805 288 1811 292
rect 2109 288 2115 332
rect 1448 277 1459 283
rect 1533 168 1539 272
rect 1645 188 1651 192
rect 1533 148 1539 152
rect 1325 128 1331 132
rect 1661 128 1667 212
rect 1677 148 1683 272
rect 1933 268 1939 272
rect 2157 268 2163 312
rect 2189 308 2195 412
rect 2237 408 2243 532
rect 2285 528 2291 692
rect 2349 608 2355 832
rect 2365 588 2371 832
rect 2429 728 2435 952
rect 2509 923 2515 1032
rect 2621 968 2627 1332
rect 2717 1308 2723 1332
rect 2829 1308 2835 1332
rect 2765 1268 2771 1292
rect 2877 1268 2883 1292
rect 2973 1168 2979 1332
rect 3069 1328 3075 1332
rect 2989 1208 2995 1312
rect 3005 1308 3011 1312
rect 3021 1283 3027 1312
rect 3005 1277 3027 1283
rect 3005 1248 3011 1277
rect 3048 1277 3064 1283
rect 3032 1237 3043 1243
rect 3021 1208 3027 1212
rect 2637 1108 2643 1132
rect 2717 1108 2723 1112
rect 2781 1108 2787 1112
rect 2669 1088 2675 1092
rect 2557 948 2563 952
rect 2504 917 2515 923
rect 2525 828 2531 892
rect 2621 868 2627 914
rect 2525 748 2531 812
rect 2429 708 2435 712
rect 2461 688 2467 692
rect 2397 648 2403 672
rect 2317 568 2323 572
rect 2301 548 2307 552
rect 2413 548 2419 672
rect 2477 608 2483 692
rect 2509 608 2515 632
rect 2349 528 2355 532
rect 2253 428 2259 452
rect 2253 328 2259 412
rect 2349 368 2355 452
rect 2413 348 2419 532
rect 2429 528 2435 592
rect 2461 528 2467 532
rect 2461 368 2467 512
rect 2477 468 2483 572
rect 2509 528 2515 552
rect 2461 328 2467 332
rect 2221 288 2227 312
rect 2253 288 2259 312
rect 1693 248 1699 252
rect 1693 188 1699 212
rect 1709 148 1715 192
rect 1821 188 1827 232
rect 1949 208 1955 232
rect 1949 168 1955 192
rect 1725 128 1731 152
rect 1805 148 1811 152
rect 2029 148 2035 252
rect 2157 168 2163 252
rect 2125 148 2131 152
rect 2173 148 2179 272
rect 1965 123 1971 132
rect 1997 128 2003 132
rect 2269 128 2275 192
rect 1960 117 1971 123
rect 1309 108 1315 112
rect 1437 68 1443 72
rect 2109 68 2115 112
rect 2285 108 2291 232
rect 2301 228 2307 312
rect 2397 288 2403 292
rect 2477 288 2483 452
rect 2509 408 2515 412
rect 2509 303 2515 392
rect 2541 388 2547 752
rect 2637 728 2643 1072
rect 2749 1068 2755 1092
rect 2829 1088 2835 1152
rect 3021 1128 3027 1192
rect 3037 1128 3043 1237
rect 3053 1208 3059 1252
rect 3053 1188 3059 1192
rect 2845 1088 2851 1092
rect 2749 988 2755 1052
rect 2717 888 2723 952
rect 2717 808 2723 872
rect 2813 848 2819 992
rect 2829 948 2835 1072
rect 2845 928 2851 1072
rect 2877 1068 2883 1112
rect 2989 1108 2995 1112
rect 3085 1108 3091 1132
rect 2877 928 2883 932
rect 2829 888 2835 912
rect 2877 908 2883 912
rect 2749 728 2755 732
rect 2589 708 2595 712
rect 2605 688 2611 712
rect 2653 703 2659 712
rect 2637 697 2659 703
rect 2621 688 2627 692
rect 2637 648 2643 697
rect 2717 688 2723 712
rect 2685 668 2691 672
rect 2557 448 2563 632
rect 2573 528 2579 572
rect 2637 568 2643 632
rect 2616 537 2627 543
rect 2605 508 2611 512
rect 2621 508 2627 537
rect 2701 523 2707 632
rect 2733 588 2739 692
rect 2749 628 2755 632
rect 2696 517 2707 523
rect 2557 408 2563 432
rect 2589 388 2595 472
rect 2504 297 2515 303
rect 2365 148 2371 252
rect 2413 188 2419 272
rect 2429 188 2435 192
rect 2397 148 2403 152
rect 2461 148 2467 152
rect 2317 108 2323 132
rect 2381 128 2387 132
rect 2493 128 2499 272
rect 2525 248 2531 312
rect 2541 143 2547 372
rect 2573 308 2579 312
rect 2589 288 2595 372
rect 2621 288 2627 472
rect 2669 388 2675 412
rect 2733 388 2739 572
rect 2765 568 2771 792
rect 2781 688 2787 712
rect 2813 703 2819 832
rect 2829 788 2835 872
rect 2813 697 2824 703
rect 2845 688 2851 792
rect 2893 688 2899 692
rect 2909 688 2915 1092
rect 3053 1088 3059 1092
rect 3069 1088 3075 1092
rect 2925 1048 2931 1072
rect 2925 983 2931 1032
rect 2941 1008 2947 1072
rect 3005 1048 3011 1072
rect 3005 988 3011 992
rect 2925 977 2947 983
rect 2925 948 2931 952
rect 2941 928 2947 977
rect 3021 948 3027 952
rect 3037 948 3043 1032
rect 3053 948 3059 1052
rect 3101 948 3107 1332
rect 3117 1208 3123 1292
rect 3133 1123 3139 1712
rect 3165 1688 3171 1692
rect 3149 1528 3155 1672
rect 3165 1588 3171 1592
rect 3181 1588 3187 1592
rect 3165 1348 3171 1572
rect 3213 1508 3219 1692
rect 3229 1548 3235 1732
rect 3277 1728 3283 1792
rect 3261 1708 3267 1712
rect 3293 1708 3299 1872
rect 3373 1848 3379 1952
rect 3405 1906 3411 2032
rect 3421 1768 3427 2112
rect 3501 1948 3507 2272
rect 3645 2248 3651 2292
rect 3517 2148 3523 2172
rect 3544 2137 3555 2143
rect 3549 2128 3555 2137
rect 3581 2128 3587 2172
rect 3597 2148 3603 2192
rect 3613 2148 3619 2232
rect 3661 2188 3667 2412
rect 3821 2408 3827 2532
rect 3517 2108 3523 2112
rect 3533 2008 3539 2112
rect 3565 2108 3571 2112
rect 3629 2108 3635 2132
rect 3661 2068 3667 2132
rect 3677 2128 3683 2312
rect 3725 2288 3731 2392
rect 3693 2148 3699 2192
rect 3709 2128 3715 2212
rect 3773 2188 3779 2292
rect 3837 2288 3843 2532
rect 3901 2528 3907 2552
rect 3933 2528 3939 2672
rect 3965 2548 3971 3072
rect 4077 2988 4083 3632
rect 4125 3408 4131 3692
rect 4189 3688 4195 3712
rect 4221 3648 4227 3652
rect 4157 3588 4163 3592
rect 4221 3548 4227 3632
rect 4253 3608 4259 3712
rect 4269 3628 4275 4077
rect 4285 3928 4291 4012
rect 4301 3988 4307 4132
rect 4317 4088 4323 4112
rect 4333 4048 4339 4532
rect 4397 4448 4403 4512
rect 4349 4388 4355 4412
rect 4397 4328 4403 4412
rect 4445 4368 4451 4672
rect 4621 4668 4627 4672
rect 4653 4648 4659 4652
rect 4461 4608 4467 4632
rect 4493 4448 4499 4512
rect 4525 4408 4531 4512
rect 4429 4328 4435 4332
rect 4365 4228 4371 4272
rect 4381 4148 4387 4272
rect 4349 4068 4355 4092
rect 4381 4088 4387 4112
rect 4397 4088 4403 4292
rect 4445 4288 4451 4332
rect 4429 4148 4435 4192
rect 4413 4108 4419 4132
rect 4445 4128 4451 4272
rect 4461 4128 4467 4292
rect 4429 4108 4435 4112
rect 4445 4048 4451 4112
rect 4493 4108 4499 4312
rect 4541 4308 4547 4312
rect 4557 4288 4563 4612
rect 4573 4508 4579 4632
rect 4621 4528 4627 4532
rect 4637 4448 4643 4532
rect 4669 4528 4675 4632
rect 4685 4568 4691 4632
rect 4701 4608 4707 4652
rect 4717 4548 4723 4552
rect 4621 4348 4627 4352
rect 4573 4288 4579 4292
rect 4509 4188 4515 4212
rect 4525 4208 4531 4272
rect 4541 4168 4547 4172
rect 4557 4148 4563 4272
rect 4589 4228 4595 4312
rect 4605 4308 4611 4312
rect 4669 4288 4675 4352
rect 4701 4348 4707 4512
rect 4733 4508 4739 4632
rect 4749 4588 4755 4712
rect 4845 4708 4851 4732
rect 4776 4697 4787 4703
rect 4749 4528 4755 4552
rect 4701 4306 4707 4312
rect 4749 4248 4755 4512
rect 4685 4188 4691 4212
rect 4589 4148 4595 4152
rect 4525 4128 4531 4132
rect 4317 4008 4323 4032
rect 4301 3748 4307 3952
rect 4397 3928 4403 3992
rect 4525 3968 4531 4112
rect 4573 4088 4579 4112
rect 4605 4068 4611 4112
rect 4637 4068 4643 4092
rect 4653 4048 4659 4112
rect 4749 4108 4755 4132
rect 4317 3908 4323 3912
rect 4381 3908 4387 3912
rect 4525 3908 4531 3952
rect 4317 3788 4323 3812
rect 4333 3708 4339 3872
rect 4349 3808 4355 3872
rect 4429 3868 4435 3872
rect 4445 3808 4451 3892
rect 4461 3888 4467 3892
rect 4509 3848 4515 3872
rect 4541 3868 4547 3872
rect 4573 3868 4579 4032
rect 4637 3908 4643 3932
rect 4509 3788 4515 3832
rect 4525 3788 4531 3852
rect 4621 3848 4627 3872
rect 4653 3868 4659 3872
rect 4557 3743 4563 3832
rect 4685 3828 4691 3872
rect 4637 3748 4643 3812
rect 4701 3748 4707 3892
rect 4717 3828 4723 4092
rect 4749 3928 4755 4092
rect 4557 3737 4579 3743
rect 4173 3368 4179 3472
rect 4189 3348 4195 3372
rect 4093 3108 4099 3172
rect 4125 3088 4131 3312
rect 4221 3308 4227 3512
rect 4269 3508 4275 3612
rect 4285 3488 4291 3532
rect 4301 3508 4307 3652
rect 4397 3528 4403 3712
rect 4269 3448 4275 3472
rect 4317 3468 4323 3472
rect 4253 3308 4259 3352
rect 4285 3348 4291 3392
rect 4333 3368 4339 3512
rect 4365 3488 4371 3512
rect 4541 3488 4547 3612
rect 4557 3508 4563 3712
rect 4573 3708 4579 3737
rect 4749 3743 4755 3912
rect 4765 3888 4771 4672
rect 4781 4628 4787 4697
rect 4813 4648 4819 4672
rect 4813 4528 4819 4572
rect 4861 4528 4867 4592
rect 4877 4548 4883 4632
rect 4893 4608 4899 4712
rect 4909 4563 4915 4732
rect 4957 4728 4963 4732
rect 5181 4708 5187 4772
rect 5309 4688 5315 4692
rect 5053 4668 5059 4672
rect 5245 4628 5251 4632
rect 4893 4557 4915 4563
rect 4781 4448 4787 4492
rect 4781 4428 4787 4432
rect 4829 4428 4835 4472
rect 4845 4308 4851 4392
rect 4861 4388 4867 4452
rect 4893 4328 4899 4557
rect 4973 4548 4979 4552
rect 5069 4548 5075 4612
rect 4909 4528 4915 4532
rect 4989 4528 4995 4532
rect 5021 4448 5027 4492
rect 5037 4488 5043 4532
rect 4829 4248 4835 4272
rect 4781 3968 4787 4192
rect 4845 4188 4851 4212
rect 4797 4108 4803 4132
rect 4845 4128 4851 4172
rect 4877 4148 4883 4272
rect 4877 4088 4883 4132
rect 4765 3788 4771 3872
rect 4781 3788 4787 3952
rect 4797 3908 4803 3912
rect 4813 3903 4819 3912
rect 4813 3897 4835 3903
rect 4813 3788 4819 3872
rect 4829 3863 4835 3897
rect 4861 3888 4867 3992
rect 4893 3948 4899 4312
rect 4925 4108 4931 4172
rect 4941 4168 4947 4272
rect 4877 3888 4883 3892
rect 4893 3863 4899 3872
rect 4829 3857 4899 3863
rect 4877 3748 4883 3752
rect 4749 3737 4771 3743
rect 4701 3728 4707 3732
rect 4653 3508 4659 3612
rect 4765 3528 4771 3737
rect 4813 3688 4819 3692
rect 4845 3688 4851 3732
rect 4813 3508 4819 3532
rect 4845 3508 4851 3672
rect 4589 3428 4595 3492
rect 4637 3488 4643 3492
rect 4861 3488 4867 3712
rect 4893 3708 4899 3752
rect 4909 3748 4915 3852
rect 4925 3728 4931 3932
rect 4941 3908 4947 3912
rect 4957 3888 4963 3892
rect 4973 3768 4979 4312
rect 5053 4308 5059 4512
rect 5085 4468 5091 4492
rect 5085 4308 5091 4392
rect 5101 4368 5107 4492
rect 5133 4348 5139 4512
rect 5149 4508 5155 4512
rect 5165 4508 5171 4512
rect 5016 4297 5027 4303
rect 4989 4288 4995 4292
rect 5005 4128 5011 4272
rect 5021 4168 5027 4297
rect 5165 4306 5171 4392
rect 5069 4208 5075 4292
rect 5021 4128 5027 4132
rect 5037 4128 5043 4172
rect 5101 4148 5107 4292
rect 5149 4188 5155 4192
rect 5133 4128 5139 4132
rect 5101 4108 5107 4112
rect 4989 3923 4995 3932
rect 4989 3917 5000 3923
rect 4989 3748 4995 3917
rect 5021 3908 5027 4032
rect 5085 3928 5091 4052
rect 5117 3968 5123 4112
rect 5117 3928 5123 3952
rect 4877 3508 4883 3532
rect 4269 3328 4275 3332
rect 4237 3288 4243 3292
rect 4285 3248 4291 3332
rect 4333 3208 4339 3332
rect 4397 3328 4403 3332
rect 4413 3308 4419 3332
rect 4429 3328 4435 3332
rect 4509 3328 4515 3332
rect 4525 3308 4531 3352
rect 4349 3268 4355 3292
rect 4125 2988 4131 3032
rect 4173 2988 4179 2992
rect 4109 2968 4115 2972
rect 4109 2948 4115 2952
rect 4013 2783 4019 2914
rect 4077 2908 4083 2912
rect 4125 2908 4131 2952
rect 4173 2828 4179 2892
rect 4013 2777 4024 2783
rect 3981 2568 3987 2672
rect 4013 2648 4019 2732
rect 4029 2708 4035 2712
rect 4045 2663 4051 2712
rect 4077 2708 4083 2772
rect 4109 2688 4115 2712
rect 4125 2688 4131 2752
rect 4045 2657 4067 2663
rect 4045 2588 4051 2592
rect 4061 2588 4067 2657
rect 4045 2548 4051 2572
rect 3805 2148 3811 2152
rect 3853 2148 3859 2312
rect 3901 2288 3907 2372
rect 3949 2308 3955 2512
rect 4093 2508 4099 2672
rect 4141 2548 4147 2692
rect 4173 2688 4179 2812
rect 4189 2588 4195 2832
rect 4205 2728 4211 2732
rect 4205 2708 4211 2712
rect 4221 2688 4227 3112
rect 4253 3088 4259 3092
rect 4269 2928 4275 3092
rect 4333 3048 4339 3072
rect 4349 3068 4355 3092
rect 4397 2988 4403 3292
rect 4461 3268 4467 3292
rect 4573 3288 4579 3332
rect 4589 3288 4595 3292
rect 4605 3288 4611 3432
rect 4621 3328 4627 3412
rect 4701 3408 4707 3432
rect 4749 3368 4755 3472
rect 4445 3108 4451 3232
rect 4461 3088 4467 3112
rect 4493 3108 4499 3112
rect 4509 3088 4515 3272
rect 4525 3128 4531 3152
rect 4541 3108 4547 3152
rect 4445 2968 4451 3072
rect 4477 2968 4483 3012
rect 4509 3008 4515 3072
rect 4253 2708 4259 2852
rect 4285 2748 4291 2932
rect 4317 2808 4323 2914
rect 4381 2768 4387 2932
rect 4525 2928 4531 3092
rect 4573 3088 4579 3172
rect 4621 3108 4627 3252
rect 4637 3208 4643 3232
rect 4637 3123 4643 3192
rect 4653 3148 4659 3332
rect 4669 3228 4675 3312
rect 4701 3308 4707 3312
rect 4717 3188 4723 3332
rect 4733 3288 4739 3332
rect 4792 3317 4803 3323
rect 4797 3308 4803 3317
rect 4829 3288 4835 3332
rect 4877 3308 4883 3352
rect 4637 3117 4659 3123
rect 4653 3108 4659 3117
rect 4669 3088 4675 3152
rect 4717 3108 4723 3152
rect 4765 3108 4771 3112
rect 4573 2948 4579 2992
rect 4589 2948 4595 3032
rect 4637 2983 4643 3072
rect 4781 3048 4787 3072
rect 4797 3068 4803 3072
rect 4632 2977 4643 2983
rect 4653 2948 4659 2992
rect 4669 2988 4675 3032
rect 4733 2948 4739 2972
rect 4429 2908 4435 2912
rect 4205 2588 4211 2632
rect 4221 2548 4227 2672
rect 4125 2528 4131 2532
rect 4237 2528 4243 2692
rect 4285 2688 4291 2732
rect 4333 2708 4339 2712
rect 4349 2648 4355 2692
rect 4397 2688 4403 2812
rect 4509 2808 4515 2832
rect 4589 2828 4595 2912
rect 4605 2888 4611 2932
rect 4749 2928 4755 2952
rect 4445 2788 4451 2792
rect 4509 2748 4515 2792
rect 4637 2788 4643 2872
rect 4317 2628 4323 2632
rect 4125 2488 4131 2512
rect 4221 2483 4227 2512
rect 4269 2508 4275 2572
rect 4349 2548 4355 2592
rect 4381 2588 4387 2632
rect 4413 2588 4419 2692
rect 4429 2648 4435 2712
rect 4445 2688 4451 2692
rect 4221 2477 4243 2483
rect 4045 2388 4051 2392
rect 4077 2388 4083 2432
rect 4237 2388 4243 2477
rect 4013 2308 4019 2312
rect 4077 2308 4083 2372
rect 4237 2348 4243 2372
rect 4189 2248 4195 2292
rect 3933 2148 3939 2192
rect 3549 1988 3555 2012
rect 3597 1988 3603 1992
rect 3597 1968 3603 1972
rect 3645 1908 3651 2032
rect 3693 1908 3699 2112
rect 3709 1908 3715 2112
rect 3741 2108 3747 2112
rect 3773 2008 3779 2132
rect 3469 1788 3475 1892
rect 3629 1868 3635 1892
rect 3773 1888 3779 1892
rect 3565 1848 3571 1852
rect 3357 1728 3363 1732
rect 3341 1688 3347 1712
rect 3293 1588 3299 1612
rect 3197 1328 3203 1472
rect 3149 1308 3155 1312
rect 3197 1248 3203 1312
rect 3213 1208 3219 1452
rect 3277 1388 3283 1452
rect 3293 1348 3299 1552
rect 3309 1508 3315 1512
rect 3341 1508 3347 1652
rect 3373 1648 3379 1732
rect 3469 1688 3475 1772
rect 3565 1768 3571 1792
rect 3373 1488 3379 1632
rect 3405 1608 3411 1672
rect 3453 1643 3459 1672
rect 3469 1643 3475 1672
rect 3453 1637 3475 1643
rect 3469 1568 3475 1637
rect 3485 1603 3491 1732
rect 3501 1688 3507 1692
rect 3485 1597 3507 1603
rect 3421 1508 3427 1532
rect 3437 1468 3443 1512
rect 3309 1368 3315 1432
rect 3437 1403 3443 1432
rect 3421 1397 3443 1403
rect 3373 1348 3379 1352
rect 3389 1288 3395 1312
rect 3421 1303 3427 1397
rect 3437 1328 3443 1372
rect 3469 1368 3475 1492
rect 3501 1408 3507 1597
rect 3533 1568 3539 1672
rect 3581 1668 3587 1712
rect 3597 1668 3603 1832
rect 3709 1828 3715 1832
rect 3773 1788 3779 1872
rect 3629 1768 3635 1772
rect 3661 1748 3667 1772
rect 3805 1748 3811 2132
rect 3853 2128 3859 2132
rect 3821 2108 3827 2112
rect 3869 2108 3875 2112
rect 3869 2088 3875 2092
rect 3645 1588 3651 1612
rect 3661 1548 3667 1552
rect 3565 1508 3571 1532
rect 3693 1508 3699 1732
rect 3709 1728 3715 1732
rect 3741 1688 3747 1692
rect 3709 1508 3715 1552
rect 3725 1528 3731 1672
rect 3773 1668 3779 1732
rect 3821 1728 3827 1812
rect 3933 1808 3939 1872
rect 3965 1828 3971 2192
rect 4013 2128 4019 2152
rect 4013 1988 4019 2092
rect 3981 1908 3987 1912
rect 3821 1708 3827 1712
rect 3885 1708 3891 1772
rect 3965 1768 3971 1812
rect 3981 1768 3987 1792
rect 3965 1728 3971 1752
rect 3981 1748 3987 1752
rect 4029 1728 4035 2232
rect 4109 2208 4115 2232
rect 4045 1948 4051 2112
rect 4061 1988 4067 2132
rect 4093 2088 4099 2152
rect 4157 2068 4163 2232
rect 4189 2188 4195 2212
rect 4205 2208 4211 2292
rect 4205 2168 4211 2172
rect 4173 2148 4179 2152
rect 4093 1908 4099 2052
rect 4141 1988 4147 1992
rect 4141 1888 4147 1972
rect 4173 1908 4179 2092
rect 4205 1908 4211 2112
rect 4077 1808 4083 1852
rect 4109 1788 4115 1872
rect 4109 1748 4115 1752
rect 3965 1688 3971 1692
rect 3773 1568 3779 1652
rect 3853 1628 3859 1672
rect 4045 1668 4051 1732
rect 4125 1728 4131 1812
rect 4221 1748 4227 2152
rect 4237 1908 4243 1912
rect 4253 1908 4259 2272
rect 4269 2108 4275 2492
rect 4301 2488 4307 2512
rect 4381 2508 4387 2512
rect 4413 2488 4419 2512
rect 4301 2448 4307 2472
rect 4365 2388 4371 2452
rect 4397 2308 4403 2472
rect 4429 2388 4435 2572
rect 4445 2548 4451 2632
rect 4461 2588 4467 2732
rect 4541 2703 4547 2712
rect 4536 2697 4547 2703
rect 4653 2697 4664 2703
rect 4509 2628 4515 2652
rect 4493 2548 4499 2552
rect 4509 2548 4515 2612
rect 4445 2448 4451 2512
rect 4525 2448 4531 2512
rect 4557 2383 4563 2472
rect 4573 2428 4579 2512
rect 4589 2408 4595 2676
rect 4653 2568 4659 2697
rect 4701 2688 4707 2912
rect 4765 2908 4771 2912
rect 4797 2903 4803 3052
rect 4813 2988 4819 3012
rect 4861 2988 4867 3092
rect 4877 3048 4883 3052
rect 4893 3028 4899 3692
rect 4973 3688 4979 3692
rect 4973 3608 4979 3672
rect 5021 3568 5027 3732
rect 5037 3728 5043 3912
rect 5117 3888 5123 3892
rect 5133 3888 5139 3932
rect 5149 3908 5155 3912
rect 5069 3848 5075 3852
rect 5053 3628 5059 3832
rect 5085 3748 5091 3852
rect 5165 3848 5171 4252
rect 5181 4188 5187 4612
rect 5245 4548 5251 4592
rect 5341 4588 5347 4712
rect 5629 4708 5635 4772
rect 6669 4737 6680 4743
rect 6397 4708 6403 4732
rect 6669 4708 6675 4737
rect 5480 4697 5491 4703
rect 5357 4588 5363 4692
rect 5485 4688 5491 4697
rect 5565 4697 5576 4703
rect 5533 4648 5539 4692
rect 5565 4688 5571 4697
rect 6344 4697 6355 4703
rect 5645 4668 5651 4672
rect 5933 4668 5939 4672
rect 5437 4548 5443 4552
rect 5485 4548 5491 4552
rect 5549 4548 5555 4612
rect 5197 4528 5203 4532
rect 5197 4448 5203 4512
rect 5213 4508 5219 4532
rect 5229 4488 5235 4512
rect 5261 4468 5267 4492
rect 5277 4268 5283 4532
rect 5373 4528 5379 4532
rect 5293 4488 5299 4512
rect 5325 4468 5331 4492
rect 5357 4308 5363 4312
rect 5293 4248 5299 4252
rect 5181 4148 5187 4172
rect 5181 4048 5187 4112
rect 5213 4108 5219 4132
rect 5213 3928 5219 4092
rect 5229 3988 5235 4172
rect 5181 3908 5187 3912
rect 5181 3888 5187 3892
rect 5149 3828 5155 3832
rect 5085 3728 5091 3732
rect 5165 3648 5171 3712
rect 5101 3528 5107 3612
rect 5133 3508 5139 3612
rect 5165 3488 5171 3592
rect 5197 3548 5203 3892
rect 5229 3528 5235 3752
rect 5181 3488 5187 3492
rect 4925 3388 4931 3432
rect 5069 3408 5075 3472
rect 5149 3468 5155 3472
rect 5197 3468 5203 3472
rect 5048 3377 5075 3383
rect 5053 3348 5059 3352
rect 5069 3343 5075 3377
rect 5133 3348 5139 3432
rect 5181 3388 5187 3432
rect 5229 3388 5235 3412
rect 5069 3337 5096 3343
rect 4957 3328 4963 3332
rect 4973 3228 4979 3332
rect 5149 3328 5155 3332
rect 5053 3188 5059 3312
rect 5085 3308 5091 3312
rect 5117 3248 5123 3312
rect 4973 3168 4979 3172
rect 5149 3128 5155 3312
rect 4861 2948 4867 2972
rect 4909 2928 4915 3052
rect 4792 2897 4803 2903
rect 4829 2868 4835 2912
rect 4925 2908 4931 2912
rect 4941 2843 4947 3052
rect 4957 2948 4963 3092
rect 4989 3068 4995 3092
rect 5005 3088 5011 3092
rect 5037 3088 5043 3092
rect 5021 2968 5027 3072
rect 4941 2837 4963 2843
rect 4749 2768 4755 2772
rect 4749 2688 4755 2752
rect 4701 2588 4707 2672
rect 4765 2628 4771 2692
rect 4733 2588 4739 2612
rect 4557 2377 4568 2383
rect 4509 2308 4515 2312
rect 4605 2308 4611 2332
rect 4637 2328 4643 2392
rect 4653 2328 4659 2432
rect 4669 2348 4675 2552
rect 4749 2548 4755 2572
rect 4829 2568 4835 2832
rect 4861 2788 4867 2812
rect 4877 2703 4883 2832
rect 4957 2728 4963 2837
rect 4925 2708 4931 2712
rect 4973 2708 4979 2952
rect 5037 2848 5043 2912
rect 5053 2908 5059 3112
rect 5165 3108 5171 3232
rect 5197 3208 5203 3312
rect 5213 3208 5219 3332
rect 5245 3228 5251 4152
rect 5277 4108 5283 4112
rect 5261 3868 5267 3892
rect 5261 3748 5267 3792
rect 5261 3728 5267 3732
rect 5261 3348 5267 3412
rect 5277 3328 5283 4092
rect 5293 3888 5299 4232
rect 5309 4188 5315 4272
rect 5325 4248 5331 4292
rect 5357 4248 5363 4272
rect 5325 4188 5331 4232
rect 5309 4068 5315 4092
rect 5309 3788 5315 3912
rect 5325 3908 5331 4112
rect 5341 3948 5347 4032
rect 5357 3908 5363 4232
rect 5373 4208 5379 4492
rect 5421 4468 5427 4512
rect 5453 4508 5459 4532
rect 5645 4528 5651 4652
rect 6013 4588 6019 4692
rect 6349 4688 6355 4697
rect 6429 4697 6440 4703
rect 6077 4637 6088 4643
rect 5917 4548 5923 4552
rect 5997 4548 6003 4552
rect 6077 4548 6083 4637
rect 6221 4548 6227 4672
rect 5773 4528 5779 4532
rect 5853 4517 5864 4523
rect 5469 4488 5475 4512
rect 5405 4308 5411 4412
rect 5485 4388 5491 4492
rect 5421 4308 5427 4332
rect 5501 4308 5507 4392
rect 5533 4388 5539 4432
rect 5389 4268 5395 4272
rect 5405 4248 5411 4292
rect 5421 4288 5427 4292
rect 5373 4088 5379 4132
rect 5389 4128 5395 4192
rect 5421 4188 5427 4232
rect 5437 4208 5443 4292
rect 5453 4288 5459 4292
rect 5485 4268 5491 4272
rect 5501 4243 5507 4292
rect 5517 4268 5523 4272
rect 5517 4248 5523 4252
rect 5485 4237 5507 4243
rect 5405 4128 5411 4132
rect 5421 4128 5427 4172
rect 5437 4068 5443 4092
rect 5453 4088 5459 4092
rect 5485 3908 5491 4237
rect 5533 4228 5539 4292
rect 5517 4168 5523 4192
rect 5549 4128 5555 4312
rect 5581 4308 5587 4432
rect 5661 4388 5667 4472
rect 5821 4468 5827 4512
rect 5597 4268 5603 4372
rect 5773 4308 5779 4312
rect 5613 4288 5619 4292
rect 5565 4068 5571 4112
rect 5517 3908 5523 3972
rect 5293 3708 5299 3712
rect 5309 3668 5315 3752
rect 5325 3748 5331 3772
rect 5389 3728 5395 3872
rect 5437 3848 5443 3892
rect 5437 3748 5443 3752
rect 5261 3308 5267 3312
rect 5261 3228 5267 3292
rect 5325 3248 5331 3492
rect 5101 3068 5107 3072
rect 5117 2928 5123 3012
rect 5037 2828 5043 2832
rect 5053 2728 5059 2892
rect 5085 2868 5091 2872
rect 5133 2768 5139 3032
rect 5149 2988 5155 3032
rect 5181 2888 5187 2932
rect 5197 2928 5203 3072
rect 4861 2697 4883 2703
rect 4749 2528 4755 2532
rect 4733 2428 4739 2492
rect 4797 2448 4803 2512
rect 4765 2388 4771 2412
rect 4637 2308 4643 2312
rect 4717 2308 4723 2352
rect 4317 2288 4323 2292
rect 4541 2288 4547 2292
rect 4477 2248 4483 2252
rect 4285 2188 4291 2232
rect 4365 2148 4371 2232
rect 4381 2148 4387 2152
rect 4317 2108 4323 2132
rect 4333 2108 4339 2112
rect 4285 2068 4291 2092
rect 4269 1917 4280 1923
rect 4253 1888 4259 1892
rect 4237 1868 4243 1872
rect 4269 1808 4275 1917
rect 4285 1868 4291 1892
rect 4301 1888 4307 1932
rect 4333 1928 4339 1932
rect 4365 1928 4371 2132
rect 4397 2128 4403 2132
rect 4429 2128 4435 2132
rect 4381 2088 4387 2112
rect 4429 2068 4435 2092
rect 4445 2028 4451 2132
rect 4461 2128 4467 2132
rect 4061 1708 4067 1712
rect 3853 1528 3859 1592
rect 3869 1588 3875 1652
rect 3677 1488 3683 1492
rect 3517 1408 3523 1432
rect 3501 1348 3507 1392
rect 3549 1348 3555 1372
rect 3421 1297 3432 1303
rect 3149 1148 3155 1152
rect 3117 1117 3139 1123
rect 3117 1068 3123 1117
rect 3117 1028 3123 1032
rect 3133 988 3139 1092
rect 3149 948 3155 1132
rect 3165 1088 3171 1132
rect 3053 928 3059 932
rect 2925 908 2931 912
rect 3085 888 3091 892
rect 3021 788 3027 792
rect 3069 748 3075 752
rect 3101 748 3107 932
rect 3149 768 3155 932
rect 3165 928 3171 1032
rect 3197 988 3203 1112
rect 3293 1108 3299 1152
rect 3341 1048 3347 1052
rect 3277 948 3283 1012
rect 3341 988 3347 992
rect 3069 728 3075 732
rect 2925 708 2931 712
rect 2781 648 2787 672
rect 2797 628 2803 632
rect 2909 588 2915 632
rect 2925 568 2931 692
rect 2941 688 2947 712
rect 3085 708 3091 712
rect 3037 688 3043 692
rect 3005 648 3011 652
rect 3037 628 3043 672
rect 3005 568 3011 612
rect 2557 168 2563 232
rect 2541 137 2552 143
rect 2493 108 2499 112
rect 2557 108 2563 112
rect 2605 108 2611 232
rect 2621 148 2627 252
rect 2637 248 2643 272
rect 2637 188 2643 232
rect 2653 128 2659 292
rect 2701 288 2707 312
rect 2733 308 2739 372
rect 2717 248 2723 292
rect 2749 288 2755 332
rect 2797 308 2803 332
rect 2861 308 2867 312
rect 2909 288 2915 452
rect 2925 308 2931 432
rect 2957 328 2963 372
rect 3037 363 3043 572
rect 3053 508 3059 632
rect 3069 588 3075 692
rect 3133 688 3139 732
rect 3149 708 3155 732
rect 3165 708 3171 852
rect 3181 728 3187 932
rect 3229 888 3235 892
rect 3197 708 3203 732
rect 3229 708 3235 832
rect 3293 748 3299 952
rect 3325 948 3331 952
rect 3341 928 3347 952
rect 3373 928 3379 1252
rect 3405 1008 3411 1052
rect 3405 948 3411 952
rect 3373 908 3379 912
rect 3389 808 3395 932
rect 3405 908 3411 912
rect 3277 708 3283 712
rect 3325 708 3331 712
rect 3101 648 3107 672
rect 3133 668 3139 672
rect 3165 668 3171 672
rect 3117 588 3123 632
rect 3101 548 3107 552
rect 3149 528 3155 572
rect 3197 548 3203 572
rect 3213 528 3219 632
rect 3309 548 3315 632
rect 3341 548 3347 552
rect 3277 528 3283 532
rect 3069 468 3075 514
rect 3037 357 3059 363
rect 2989 328 2995 332
rect 3021 308 3027 312
rect 3037 308 3043 332
rect 3053 288 3059 357
rect 3085 288 3091 412
rect 3101 308 3107 372
rect 3117 308 3123 352
rect 3133 288 3139 512
rect 3261 328 3267 332
rect 3293 308 3299 452
rect 3389 448 3395 692
rect 3405 648 3411 892
rect 3421 708 3427 1172
rect 3437 1068 3443 1092
rect 3437 768 3443 912
rect 3453 688 3459 1032
rect 3469 968 3475 1312
rect 3517 1168 3523 1332
rect 3565 1328 3571 1452
rect 3581 1348 3587 1392
rect 3581 1288 3587 1332
rect 3597 1328 3603 1352
rect 3517 1108 3523 1112
rect 3501 988 3507 1052
rect 3469 928 3475 932
rect 3533 923 3539 1192
rect 3565 948 3571 1032
rect 3597 1023 3603 1312
rect 3613 1248 3619 1472
rect 3693 1468 3699 1492
rect 3789 1488 3795 1492
rect 3693 1448 3699 1452
rect 3629 1308 3635 1352
rect 3677 1328 3683 1412
rect 3757 1388 3763 1432
rect 3757 1348 3763 1372
rect 3736 1337 3747 1343
rect 3661 1308 3667 1312
rect 3693 1308 3699 1312
rect 3613 1048 3619 1232
rect 3629 1188 3635 1212
rect 3741 1168 3747 1337
rect 3581 1017 3603 1023
rect 3528 917 3539 923
rect 3581 848 3587 1017
rect 3629 948 3635 952
rect 3645 928 3651 1072
rect 3693 1068 3699 1112
rect 3741 1088 3747 1152
rect 3773 1128 3779 1472
rect 3805 1448 3811 1472
rect 3869 1468 3875 1492
rect 3901 1488 3907 1492
rect 3949 1488 3955 1652
rect 3965 1528 3971 1572
rect 3997 1528 4003 1612
rect 3965 1508 3971 1512
rect 4045 1488 4051 1552
rect 4061 1488 4067 1492
rect 4077 1488 4083 1532
rect 4109 1488 4115 1712
rect 4125 1648 4131 1692
rect 4125 1508 4131 1632
rect 4141 1628 4147 1712
rect 4204 1697 4211 1703
rect 4205 1548 4211 1697
rect 4221 1668 4227 1712
rect 4237 1608 4243 1732
rect 4253 1728 4259 1732
rect 4173 1528 4179 1532
rect 4157 1488 4163 1492
rect 4237 1488 4243 1512
rect 3901 1468 3907 1472
rect 3757 1088 3763 1092
rect 3613 908 3619 912
rect 3645 888 3651 912
rect 3677 908 3683 1052
rect 3725 983 3731 1032
rect 3741 1008 3747 1072
rect 3725 977 3747 983
rect 3725 928 3731 952
rect 3741 908 3747 977
rect 3709 888 3715 892
rect 3549 808 3555 832
rect 3805 768 3811 1072
rect 3821 948 3827 1272
rect 3549 708 3555 712
rect 3693 708 3699 712
rect 3533 688 3539 692
rect 3741 688 3747 732
rect 3757 688 3763 692
rect 3421 648 3427 652
rect 3453 603 3459 672
rect 3613 648 3619 652
rect 3437 597 3459 603
rect 3421 528 3427 532
rect 3437 528 3443 597
rect 3176 297 3192 303
rect 2781 248 2787 272
rect 2813 268 2819 272
rect 2717 228 2723 232
rect 2701 128 2707 132
rect 2749 128 2755 132
rect 2765 88 2771 232
rect 2781 208 2787 232
rect 2829 228 2835 232
rect 2861 128 2867 232
rect 2957 148 2963 272
rect 3021 268 3027 272
rect 3053 268 3059 272
rect 3197 268 3203 272
rect 3229 248 3235 292
rect 2989 148 2995 212
rect 2973 128 2979 132
rect 3005 128 3011 232
rect 3053 188 3059 192
rect 3037 88 3043 92
rect 3069 88 3075 232
rect 3181 168 3187 172
rect 3245 163 3251 272
rect 3261 188 3267 272
rect 3293 228 3299 272
rect 3309 208 3315 372
rect 3325 308 3331 312
rect 3373 308 3379 332
rect 3421 308 3427 312
rect 3341 268 3347 292
rect 3389 288 3395 292
rect 3405 288 3411 292
rect 3245 157 3267 163
rect 1885 -43 1891 32
rect 3245 -43 3251 132
rect 3261 128 3267 157
rect 3293 148 3299 152
rect 3309 148 3315 192
rect 3421 188 3427 292
rect 3469 288 3475 612
rect 3485 308 3491 552
rect 3501 488 3507 492
rect 3517 448 3523 532
rect 3533 528 3539 632
rect 3549 608 3555 632
rect 3661 608 3667 632
rect 3645 528 3651 532
rect 3661 528 3667 592
rect 3677 548 3683 572
rect 3533 448 3539 512
rect 3533 328 3539 372
rect 3501 308 3507 312
rect 3549 308 3555 472
rect 3693 388 3699 512
rect 3725 508 3731 572
rect 3789 548 3795 692
rect 3805 568 3811 752
rect 3741 508 3747 532
rect 3757 528 3763 532
rect 3773 528 3779 532
rect 3837 528 3843 772
rect 3853 628 3859 1272
rect 3869 1228 3875 1452
rect 3949 1448 3955 1472
rect 3949 1348 3955 1352
rect 3997 1268 4003 1452
rect 4045 1448 4051 1472
rect 4109 1428 4115 1472
rect 4253 1468 4259 1712
rect 4285 1708 4291 1832
rect 4301 1748 4307 1872
rect 4317 1728 4323 1892
rect 4269 1588 4275 1612
rect 4269 1548 4275 1572
rect 4301 1508 4307 1592
rect 4317 1588 4323 1712
rect 4349 1708 4355 1912
rect 4365 1848 4371 1852
rect 4365 1648 4371 1732
rect 4365 1628 4371 1632
rect 4381 1608 4387 1832
rect 4413 1748 4419 1912
rect 4445 1888 4451 1972
rect 4461 1908 4467 2032
rect 4477 2008 4483 2232
rect 4701 2228 4707 2272
rect 4541 2148 4547 2192
rect 4653 2148 4659 2172
rect 4493 2068 4499 2092
rect 4525 1928 4531 2072
rect 4541 1988 4547 2132
rect 4573 2108 4579 2112
rect 4589 2068 4595 2072
rect 4653 2068 4659 2132
rect 4557 1988 4563 2052
rect 4557 1888 4563 1892
rect 4605 1888 4611 1892
rect 4573 1868 4579 1872
rect 4429 1823 4435 1832
rect 4429 1817 4451 1823
rect 4429 1728 4435 1792
rect 4445 1708 4451 1817
rect 4493 1768 4499 1832
rect 4589 1828 4595 1872
rect 4637 1808 4643 1912
rect 4717 1908 4723 1912
rect 4733 1888 4739 1972
rect 4765 1948 4771 2272
rect 4781 2088 4787 2292
rect 4797 2288 4803 2392
rect 4813 2328 4819 2532
rect 4829 2528 4835 2532
rect 4845 2408 4851 2672
rect 4861 2648 4867 2697
rect 4893 2688 4899 2692
rect 4861 2588 4867 2612
rect 4845 2308 4851 2372
rect 4829 2128 4835 2132
rect 4765 1903 4771 1932
rect 4781 1928 4787 2032
rect 4829 1908 4835 1992
rect 4760 1897 4771 1903
rect 4621 1788 4627 1792
rect 4173 1428 4179 1432
rect 4045 1328 4051 1372
rect 4077 1368 4083 1392
rect 4125 1343 4131 1392
rect 4120 1337 4131 1343
rect 3997 1188 4003 1252
rect 3869 1108 3875 1112
rect 4029 1108 4035 1252
rect 4125 1248 4131 1337
rect 4173 1308 4179 1332
rect 4205 1168 4211 1312
rect 4221 1288 4227 1332
rect 4045 1128 4051 1152
rect 4045 1083 4051 1112
rect 4029 1077 4051 1083
rect 4029 928 4035 1077
rect 4045 1048 4051 1052
rect 3933 888 3939 912
rect 3981 888 3987 912
rect 4045 903 4051 1032
rect 4061 948 4067 1132
rect 4125 1108 4131 1152
rect 4125 1088 4131 1092
rect 4157 1008 4163 1112
rect 4189 1077 4200 1083
rect 4093 948 4099 952
rect 4125 948 4131 972
rect 4040 897 4051 903
rect 3901 728 3907 872
rect 4061 748 4067 932
rect 4109 928 4115 932
rect 4141 888 4147 912
rect 4173 908 4179 1052
rect 4189 988 4195 1077
rect 4221 1068 4227 1272
rect 4269 1243 4275 1432
rect 4269 1237 4291 1243
rect 4237 1108 4243 1112
rect 4253 1048 4259 1112
rect 4269 1008 4275 1072
rect 4269 948 4275 952
rect 4189 808 4195 932
rect 4221 908 4227 912
rect 4237 868 4243 932
rect 4269 848 4275 932
rect 4109 728 4115 732
rect 3901 688 3907 712
rect 4013 708 4019 712
rect 4141 688 4147 772
rect 3885 668 3891 672
rect 3853 548 3859 612
rect 3869 608 3875 652
rect 3869 588 3875 592
rect 3581 317 3619 323
rect 3581 308 3587 317
rect 3613 308 3619 317
rect 3645 308 3651 312
rect 3549 288 3555 292
rect 3597 288 3603 292
rect 3405 68 3411 112
rect 3421 108 3427 132
rect 3437 128 3443 232
rect 3485 228 3491 272
rect 3501 148 3507 152
rect 3597 108 3603 232
rect 3661 188 3667 332
rect 3741 328 3747 372
rect 3688 317 3704 323
rect 3741 308 3747 312
rect 3757 308 3763 472
rect 3789 468 3795 512
rect 3805 408 3811 492
rect 3901 488 3907 512
rect 3949 508 3955 532
rect 3965 528 3971 552
rect 3981 528 3987 532
rect 3997 448 4003 512
rect 4013 448 4019 672
rect 4077 588 4083 652
rect 4093 608 4099 672
rect 4157 668 4163 712
rect 4173 708 4179 712
rect 4189 708 4195 792
rect 4269 788 4275 792
rect 4093 548 4099 592
rect 4093 528 4099 532
rect 4109 528 4115 552
rect 4173 548 4179 672
rect 4253 648 4259 692
rect 4269 688 4275 772
rect 4285 708 4291 1237
rect 4301 1208 4307 1492
rect 4317 1488 4323 1512
rect 4381 1488 4387 1532
rect 4461 1488 4467 1512
rect 4477 1508 4483 1612
rect 4429 1468 4435 1472
rect 4317 1328 4323 1412
rect 4397 1308 4403 1432
rect 4477 1388 4483 1492
rect 4525 1488 4531 1632
rect 4541 1528 4547 1732
rect 4557 1708 4563 1772
rect 4589 1728 4595 1772
rect 4605 1748 4611 1752
rect 4557 1628 4563 1692
rect 4653 1648 4659 1872
rect 4589 1608 4595 1632
rect 4557 1528 4563 1592
rect 4589 1508 4595 1572
rect 4621 1528 4627 1592
rect 4685 1528 4691 1592
rect 4653 1508 4659 1512
rect 4493 1468 4499 1472
rect 4477 1308 4483 1314
rect 4493 1188 4499 1452
rect 4541 1328 4547 1412
rect 4301 1168 4307 1172
rect 4301 1128 4307 1152
rect 4333 1028 4339 1092
rect 4397 1088 4403 1132
rect 4589 1128 4595 1492
rect 4669 1488 4675 1512
rect 4685 1488 4691 1492
rect 4701 1468 4707 1872
rect 4733 1768 4739 1872
rect 4749 1788 4755 1892
rect 4781 1808 4787 1832
rect 4845 1828 4851 1872
rect 4781 1748 4787 1772
rect 4749 1548 4755 1552
rect 4717 1508 4723 1512
rect 4749 1508 4755 1532
rect 4781 1528 4787 1712
rect 4813 1708 4819 1792
rect 4845 1728 4851 1812
rect 4861 1748 4867 2552
rect 4877 2508 4883 2532
rect 4877 2368 4883 2492
rect 4893 2408 4899 2672
rect 4909 2468 4915 2492
rect 4957 2428 4963 2672
rect 5021 2648 5027 2712
rect 5101 2708 5107 2732
rect 5165 2728 5171 2752
rect 5021 2628 5027 2632
rect 4973 2528 4979 2552
rect 4989 2508 4995 2532
rect 5032 2497 5043 2503
rect 4973 2308 4979 2432
rect 4909 2148 4915 2272
rect 4957 2108 4963 2112
rect 4909 2043 4915 2092
rect 4893 2037 4915 2043
rect 4893 1988 4899 2037
rect 4957 1988 4963 2072
rect 5005 2008 5011 2112
rect 5037 2068 5043 2497
rect 5053 2268 5059 2672
rect 5117 2648 5123 2672
rect 5069 2568 5075 2632
rect 5117 2568 5123 2632
rect 5181 2528 5187 2872
rect 5197 2868 5203 2912
rect 5197 2688 5203 2832
rect 5213 2808 5219 3192
rect 5341 3188 5347 3312
rect 5357 3168 5363 3232
rect 5357 3148 5363 3152
rect 5229 3068 5235 3132
rect 5245 3108 5251 3132
rect 5261 3108 5267 3112
rect 5341 3108 5347 3112
rect 5357 3068 5363 3072
rect 5229 2908 5235 2912
rect 5245 2908 5251 3032
rect 5277 2928 5283 3052
rect 5293 2988 5299 3052
rect 5309 3048 5315 3052
rect 5373 2948 5379 3392
rect 5389 3328 5395 3632
rect 5405 3428 5411 3432
rect 5421 3388 5427 3732
rect 5453 3708 5459 3712
rect 5485 3708 5491 3832
rect 5517 3788 5523 3872
rect 5533 3868 5539 4052
rect 5581 4028 5587 4232
rect 5597 3888 5603 4012
rect 5613 3928 5619 4252
rect 5645 4188 5651 4192
rect 5661 4028 5667 4132
rect 5677 4128 5683 4172
rect 5693 4063 5699 4292
rect 5725 4277 5736 4283
rect 5709 4188 5715 4272
rect 5725 4268 5731 4277
rect 5725 4148 5731 4252
rect 5757 4248 5763 4292
rect 5789 4283 5795 4312
rect 5805 4308 5811 4312
rect 5821 4308 5827 4452
rect 5837 4328 5843 4452
rect 5853 4348 5859 4517
rect 5901 4448 5907 4492
rect 5789 4277 5800 4283
rect 5757 4228 5763 4232
rect 5709 4088 5715 4092
rect 5693 4057 5715 4063
rect 5677 3928 5683 3932
rect 5693 3928 5699 3932
rect 5613 3908 5619 3912
rect 5709 3908 5715 4057
rect 5725 4028 5731 4132
rect 5741 4128 5747 4212
rect 5805 4208 5811 4272
rect 5821 4268 5827 4272
rect 5805 4168 5811 4192
rect 5837 4188 5843 4312
rect 5869 4308 5875 4392
rect 5933 4368 5939 4512
rect 5997 4388 6003 4472
rect 6061 4468 6067 4512
rect 5885 4328 5891 4332
rect 5853 4148 5859 4272
rect 5853 4068 5859 4132
rect 5885 4128 5891 4132
rect 5533 3788 5539 3832
rect 5453 3628 5459 3692
rect 5501 3608 5507 3712
rect 5693 3708 5699 3892
rect 5725 3748 5731 3932
rect 5757 3908 5763 4052
rect 5869 4008 5875 4112
rect 5901 4088 5907 4112
rect 5917 4108 5923 4292
rect 5933 4288 5939 4352
rect 6029 4328 6035 4372
rect 6077 4328 6083 4532
rect 6093 4508 6099 4512
rect 6125 4408 6131 4512
rect 6141 4488 6147 4492
rect 6173 4468 6179 4512
rect 5949 4068 5955 4132
rect 5917 3988 5923 4012
rect 5773 3888 5779 3892
rect 5885 3888 5891 3892
rect 5853 3748 5859 3872
rect 5965 3868 5971 4152
rect 5981 4128 5987 4272
rect 5997 4248 6003 4292
rect 6109 4288 6115 4352
rect 6125 4268 6131 4392
rect 6189 4368 6195 4532
rect 6253 4530 6259 4632
rect 6381 4583 6387 4692
rect 6429 4688 6435 4697
rect 6525 4697 6536 4703
rect 6493 4588 6499 4692
rect 6525 4688 6531 4697
rect 6632 4697 6643 4703
rect 6637 4688 6643 4697
rect 6749 4668 6755 4863
rect 6381 4577 6392 4583
rect 6461 4508 6467 4512
rect 6653 4508 6659 4512
rect 6349 4488 6355 4492
rect 6621 4308 6627 4472
rect 6685 4388 6691 4512
rect 6813 4328 6819 4332
rect 6125 4168 6131 4232
rect 6125 4148 6131 4152
rect 6109 4137 6120 4143
rect 5997 4128 6003 4132
rect 6045 4128 6051 4132
rect 5981 3988 5987 4012
rect 5997 3988 6003 4112
rect 6013 4108 6019 4112
rect 6061 4088 6067 4132
rect 6109 4108 6115 4137
rect 6173 4128 6179 4132
rect 6189 4128 6195 4252
rect 6237 4188 6243 4292
rect 6413 4168 6419 4292
rect 6733 4297 6744 4303
rect 6285 4148 6291 4152
rect 6333 4148 6339 4152
rect 5997 3848 6003 3972
rect 6029 3908 6035 3992
rect 6045 3868 6051 4032
rect 6125 4028 6131 4112
rect 6157 4108 6163 4112
rect 6093 3908 6099 3932
rect 5613 3588 5619 3592
rect 5693 3588 5699 3692
rect 5741 3637 5752 3643
rect 5741 3523 5747 3637
rect 5885 3588 5891 3714
rect 5981 3648 5987 3712
rect 6013 3568 6019 3632
rect 5741 3517 5763 3523
rect 5453 3328 5459 3412
rect 5469 3408 5475 3492
rect 5485 3468 5491 3492
rect 5757 3488 5763 3517
rect 5805 3517 5816 3523
rect 5693 3448 5699 3472
rect 5469 3388 5475 3392
rect 5565 3328 5571 3332
rect 5581 3328 5587 3392
rect 5613 3348 5619 3432
rect 5629 3328 5635 3332
rect 5421 3248 5427 3272
rect 5421 3128 5427 3232
rect 5453 3128 5459 3312
rect 5469 3268 5475 3312
rect 5501 3308 5507 3312
rect 5549 3308 5555 3312
rect 5565 3148 5571 3312
rect 5645 3308 5651 3312
rect 5613 3288 5619 3292
rect 5389 3108 5395 3112
rect 5597 3108 5603 3232
rect 5213 2688 5219 2692
rect 5197 2648 5203 2672
rect 5197 2588 5203 2612
rect 5229 2548 5235 2892
rect 5277 2888 5283 2892
rect 5245 2708 5251 2752
rect 5261 2708 5267 2832
rect 5277 2688 5283 2872
rect 5293 2668 5299 2692
rect 5245 2548 5251 2632
rect 5101 2368 5107 2472
rect 5101 2308 5107 2352
rect 5133 2308 5139 2312
rect 5149 2308 5155 2312
rect 5165 2308 5171 2312
rect 5181 2308 5187 2412
rect 5053 2208 5059 2252
rect 5069 2108 5075 2232
rect 5101 2128 5107 2272
rect 5149 2168 5155 2292
rect 5181 2263 5187 2292
rect 5197 2288 5203 2492
rect 5213 2308 5219 2312
rect 5229 2268 5235 2272
rect 5181 2257 5203 2263
rect 4877 1788 4883 1932
rect 4973 1908 4979 1912
rect 5053 1908 5059 1952
rect 4893 1888 4899 1892
rect 5101 1888 5107 1892
rect 5117 1888 5123 1992
rect 5149 1888 5155 2092
rect 5165 1908 5171 2192
rect 5181 2128 5187 2132
rect 5197 2028 5203 2257
rect 5245 2228 5251 2532
rect 5277 2508 5283 2652
rect 5309 2588 5315 2792
rect 5357 2788 5363 2912
rect 5389 2908 5395 3032
rect 5421 3008 5427 3092
rect 5549 3083 5555 3092
rect 5613 3088 5619 3192
rect 5661 3188 5667 3332
rect 5677 3288 5683 3312
rect 5629 3108 5635 3132
rect 5533 3077 5555 3083
rect 5533 3068 5539 3077
rect 5421 2868 5427 2914
rect 5517 2908 5523 3032
rect 5485 2788 5491 2872
rect 5533 2808 5539 3052
rect 5549 3048 5555 3052
rect 5549 2948 5555 3012
rect 5565 3008 5571 3072
rect 5549 2848 5555 2932
rect 5581 2908 5587 3072
rect 5597 2988 5603 3032
rect 5613 2968 5619 2972
rect 5629 2948 5635 3032
rect 5661 3008 5667 3092
rect 5645 2948 5651 2972
rect 5693 2948 5699 3432
rect 5757 3328 5763 3472
rect 5773 3388 5779 3472
rect 5789 3388 5795 3452
rect 5709 3308 5715 3312
rect 5709 3208 5715 3292
rect 5725 3188 5731 3272
rect 5741 3148 5747 3312
rect 5789 3288 5795 3292
rect 5773 3188 5779 3192
rect 5741 3128 5747 3132
rect 5805 3128 5811 3517
rect 5853 3483 5859 3532
rect 5869 3528 5875 3532
rect 5832 3477 5859 3483
rect 5837 3348 5843 3352
rect 5853 3343 5859 3452
rect 5933 3448 5939 3492
rect 5981 3488 5987 3552
rect 5869 3388 5875 3432
rect 5848 3337 5859 3343
rect 5821 3108 5827 3112
rect 5709 3028 5715 3072
rect 5789 2988 5795 3072
rect 5837 2983 5843 3272
rect 5869 3208 5875 3292
rect 5885 3228 5891 3312
rect 5933 3308 5939 3332
rect 5949 3328 5955 3352
rect 5981 3328 5987 3472
rect 5997 3368 6003 3392
rect 6013 3363 6019 3552
rect 6029 3508 6035 3792
rect 6061 3768 6067 3832
rect 6125 3768 6131 3832
rect 6157 3768 6163 3872
rect 6189 3808 6195 4112
rect 6269 3928 6275 4112
rect 6317 3988 6323 4112
rect 6349 4088 6355 4092
rect 6237 3823 6243 3892
rect 6221 3817 6243 3823
rect 6221 3788 6227 3817
rect 6061 3708 6067 3712
rect 6157 3648 6163 3752
rect 6184 3737 6195 3743
rect 6189 3728 6195 3737
rect 6237 3728 6243 3792
rect 6285 3748 6291 3852
rect 6317 3828 6323 3972
rect 6429 3908 6435 4272
rect 6557 4208 6563 4290
rect 6557 4188 6563 4192
rect 6621 4148 6627 4292
rect 6701 4188 6707 4292
rect 6733 4288 6739 4297
rect 6477 4128 6483 4132
rect 6749 4128 6755 4192
rect 6445 3968 6451 4112
rect 6605 4108 6611 4114
rect 6621 3928 6627 4052
rect 6637 3928 6643 4072
rect 6349 3848 6355 3852
rect 6157 3548 6163 3612
rect 6173 3608 6179 3712
rect 6221 3708 6227 3712
rect 6109 3517 6120 3523
rect 6029 3468 6035 3472
rect 6013 3357 6024 3363
rect 6029 3348 6035 3352
rect 5901 3148 5907 3172
rect 5901 3088 5907 3132
rect 5917 3108 5923 3152
rect 5933 3048 5939 3292
rect 5949 3128 5955 3172
rect 5832 2977 5843 2983
rect 5805 2948 5811 2972
rect 5341 2668 5347 2712
rect 5341 2608 5347 2652
rect 5357 2548 5363 2672
rect 5405 2628 5411 2732
rect 5421 2708 5427 2712
rect 5437 2708 5443 2752
rect 5533 2708 5539 2752
rect 5437 2648 5443 2672
rect 5485 2648 5491 2652
rect 5469 2608 5475 2632
rect 5501 2608 5507 2652
rect 5421 2528 5427 2552
rect 5384 2517 5395 2523
rect 5277 2488 5283 2492
rect 5261 2328 5267 2432
rect 5277 2288 5283 2472
rect 5261 2128 5267 2232
rect 5293 2168 5299 2292
rect 5213 2108 5219 2112
rect 5309 2108 5315 2452
rect 5325 2288 5331 2292
rect 5341 2248 5347 2512
rect 5389 2468 5395 2517
rect 5405 2508 5411 2512
rect 5357 2388 5363 2412
rect 5373 2328 5379 2432
rect 5405 2308 5411 2492
rect 5437 2308 5443 2572
rect 5549 2548 5555 2772
rect 5581 2728 5587 2792
rect 5597 2728 5603 2932
rect 5645 2888 5651 2912
rect 5661 2908 5667 2912
rect 5677 2788 5683 2892
rect 5613 2648 5619 2692
rect 5485 2508 5491 2532
rect 5533 2528 5539 2532
rect 5501 2428 5507 2512
rect 5517 2428 5523 2432
rect 5373 2268 5379 2292
rect 5421 2288 5427 2292
rect 5453 2288 5459 2312
rect 5501 2288 5507 2312
rect 5533 2308 5539 2392
rect 5581 2308 5587 2592
rect 5613 2348 5619 2632
rect 5629 2368 5635 2672
rect 5645 2568 5651 2692
rect 5693 2608 5699 2932
rect 5837 2763 5843 2952
rect 5853 2948 5859 3012
rect 5885 2928 5891 2992
rect 5885 2908 5891 2912
rect 5933 2788 5939 2832
rect 5965 2788 5971 2832
rect 5837 2757 5859 2763
rect 5837 2728 5843 2732
rect 5853 2708 5859 2757
rect 5805 2688 5811 2692
rect 5821 2688 5827 2692
rect 5869 2688 5875 2692
rect 5885 2688 5891 2712
rect 5981 2708 5987 3312
rect 6045 3288 6051 3492
rect 6061 3368 6067 3472
rect 6077 3428 6083 3432
rect 6109 3368 6115 3517
rect 6157 3508 6163 3532
rect 6013 3228 6019 3232
rect 6029 3188 6035 3232
rect 6061 3208 6067 3312
rect 6093 3308 6099 3352
rect 6040 3097 6051 3103
rect 6045 2988 6051 3097
rect 6061 3028 6067 3112
rect 6077 2948 6083 3152
rect 6093 3088 6099 3172
rect 6109 3108 6115 3212
rect 6093 2968 6099 3072
rect 6029 2888 6035 2912
rect 6077 2908 6083 2932
rect 6109 2908 6115 3052
rect 6125 2888 6131 3492
rect 6173 3488 6179 3572
rect 6189 3488 6195 3692
rect 6253 3548 6259 3732
rect 6221 3528 6227 3532
rect 6285 3528 6291 3732
rect 6301 3728 6307 3752
rect 6301 3508 6307 3552
rect 6317 3543 6323 3732
rect 6333 3568 6339 3712
rect 6365 3708 6371 3832
rect 6397 3748 6403 3852
rect 6429 3748 6435 3752
rect 6445 3728 6451 3792
rect 6461 3708 6467 3732
rect 6349 3588 6355 3632
rect 6477 3628 6483 3712
rect 6317 3537 6339 3543
rect 6157 3388 6163 3452
rect 6189 3448 6195 3472
rect 6317 3408 6323 3492
rect 6333 3488 6339 3537
rect 6173 3348 6179 3352
rect 6333 3348 6339 3472
rect 6349 3428 6355 3552
rect 6381 3508 6387 3592
rect 6381 3468 6387 3472
rect 6429 3448 6435 3512
rect 6493 3488 6499 3852
rect 6525 3748 6531 3752
rect 6525 3708 6531 3732
rect 6173 3283 6179 3332
rect 6205 3328 6211 3332
rect 6269 3328 6275 3332
rect 6349 3328 6355 3412
rect 6365 3368 6371 3392
rect 6397 3388 6403 3392
rect 6461 3388 6467 3472
rect 6493 3328 6499 3352
rect 6509 3348 6515 3432
rect 6525 3328 6531 3332
rect 6541 3328 6547 3812
rect 6557 3788 6563 3912
rect 6589 3908 6595 3912
rect 6669 3908 6675 4112
rect 6717 3897 6728 3903
rect 6573 3788 6579 3872
rect 6589 3688 6595 3732
rect 6605 3648 6611 3712
rect 6637 3528 6643 3632
rect 6653 3463 6659 3892
rect 6717 3888 6723 3897
rect 6669 3748 6675 3872
rect 6685 3768 6691 3792
rect 6733 3723 6739 3732
rect 6733 3717 6744 3723
rect 6653 3457 6675 3463
rect 6189 3308 6195 3312
rect 6221 3308 6227 3312
rect 6173 3277 6195 3283
rect 6141 2928 6147 3192
rect 6173 3108 6179 3252
rect 6141 2868 6147 2912
rect 6157 2908 6163 3072
rect 6173 2988 6179 2992
rect 6173 2948 6179 2972
rect 6189 2768 6195 3277
rect 6269 3168 6275 3312
rect 6429 3308 6435 3312
rect 6317 3128 6323 3232
rect 6365 3088 6371 3092
rect 6237 3068 6243 3072
rect 6205 2988 6211 3032
rect 6269 2948 6275 2952
rect 6285 2948 6291 3052
rect 6317 3043 6323 3072
rect 6301 3037 6323 3043
rect 6253 2908 6259 2912
rect 5709 2628 5715 2672
rect 5517 2288 5523 2292
rect 5229 2068 5235 2092
rect 5277 2068 5283 2072
rect 5309 2048 5315 2092
rect 5213 1928 5219 2032
rect 5229 1888 5235 2012
rect 5000 1877 5011 1883
rect 4957 1708 4963 1832
rect 4973 1748 4979 1852
rect 4989 1728 4995 1752
rect 4829 1688 4835 1692
rect 4957 1588 4963 1692
rect 4925 1508 4931 1552
rect 4733 1488 4739 1492
rect 4797 1428 4803 1472
rect 4989 1428 4995 1712
rect 5005 1508 5011 1877
rect 5021 1748 5027 1872
rect 5037 1788 5043 1852
rect 5101 1788 5107 1792
rect 5005 1448 5011 1472
rect 5005 1368 5011 1432
rect 5021 1388 5027 1712
rect 5085 1668 5091 1712
rect 5037 1388 5043 1632
rect 5069 1508 5075 1512
rect 5101 1508 5107 1632
rect 5133 1528 5139 1832
rect 5197 1788 5203 1872
rect 5149 1748 5155 1772
rect 5213 1768 5219 1832
rect 5149 1728 5155 1732
rect 5181 1708 5187 1712
rect 5229 1643 5235 1872
rect 5277 1848 5283 1912
rect 5229 1637 5251 1643
rect 5229 1588 5235 1612
rect 5176 1497 5187 1503
rect 5085 1383 5091 1472
rect 5080 1377 5091 1383
rect 4685 1348 4691 1352
rect 4621 1328 4627 1332
rect 4637 1328 4643 1332
rect 4429 1106 4435 1112
rect 4493 1028 4499 1052
rect 4301 988 4307 1012
rect 4461 1008 4467 1012
rect 4461 968 4467 992
rect 4493 988 4499 992
rect 4317 948 4323 952
rect 4333 928 4339 932
rect 4413 908 4419 912
rect 4477 828 4483 932
rect 4525 928 4531 952
rect 4541 948 4547 992
rect 4605 968 4611 1052
rect 4621 1028 4627 1312
rect 4637 1108 4643 1252
rect 4637 988 4643 1072
rect 4605 948 4611 952
rect 4493 868 4499 912
rect 4541 888 4547 932
rect 4557 808 4563 892
rect 4301 688 4307 712
rect 4349 708 4355 712
rect 4445 708 4451 772
rect 4573 748 4579 912
rect 4589 768 4595 912
rect 4509 728 4515 732
rect 4525 728 4531 732
rect 4525 688 4531 692
rect 4333 668 4339 672
rect 4397 668 4403 672
rect 4253 628 4259 632
rect 4029 508 4035 512
rect 4045 488 4051 512
rect 4125 508 4131 512
rect 3816 317 3832 323
rect 3944 317 3992 323
rect 3693 288 3699 292
rect 3805 288 3811 292
rect 3869 248 3875 292
rect 3965 288 3971 292
rect 3981 288 3987 292
rect 3853 188 3859 192
rect 3693 148 3699 152
rect 3981 148 3987 272
rect 4013 208 4019 392
rect 4029 288 4035 372
rect 4077 288 4083 432
rect 4157 328 4163 512
rect 4173 348 4179 512
rect 4189 468 4195 532
rect 4237 508 4243 532
rect 4253 528 4259 572
rect 4301 548 4307 572
rect 4333 528 4339 532
rect 4397 528 4403 572
rect 4413 548 4419 592
rect 4445 548 4451 632
rect 4477 608 4483 672
rect 4477 568 4483 572
rect 4461 448 4467 512
rect 4125 288 4131 292
rect 4205 288 4211 332
rect 4285 288 4291 332
rect 4333 328 4339 332
rect 4045 228 4051 252
rect 4013 148 4019 192
rect 4077 148 4083 152
rect 4125 148 4131 152
rect 4141 128 4147 232
rect 4205 148 4211 272
rect 4253 128 4259 132
rect 3469 88 3475 92
rect 3869 -43 3875 112
rect 4301 48 4307 292
rect 4317 268 4323 272
rect 4365 248 4371 432
rect 4477 428 4483 432
rect 4365 188 4371 192
rect 4381 188 4387 192
rect 4397 148 4403 272
rect 4413 108 4419 332
rect 4445 308 4451 352
rect 4493 188 4499 592
rect 4509 548 4515 632
rect 4541 628 4547 712
rect 4573 708 4579 732
rect 4605 688 4611 792
rect 4621 788 4627 892
rect 4637 743 4643 832
rect 4621 737 4643 743
rect 4541 528 4547 612
rect 4589 548 4595 552
rect 4621 548 4627 737
rect 4653 668 4659 1232
rect 4669 728 4675 1032
rect 4685 948 4691 1032
rect 4701 928 4707 1192
rect 4765 1108 4771 1132
rect 4813 1128 4819 1212
rect 4845 1188 4851 1312
rect 5005 1308 5011 1352
rect 5021 1348 5027 1372
rect 5133 1348 5139 1432
rect 5149 1348 5155 1392
rect 4861 1148 4867 1272
rect 5117 1248 5123 1312
rect 5165 1308 5171 1472
rect 4872 1137 4883 1143
rect 4813 1108 4819 1112
rect 4877 1108 4883 1137
rect 4957 1088 4963 1112
rect 4973 1088 4979 1232
rect 4989 1128 4995 1132
rect 5133 1128 5139 1152
rect 5021 1068 5027 1072
rect 4781 1048 4787 1052
rect 4717 1008 4723 1032
rect 4685 708 4691 792
rect 4717 763 4723 992
rect 4765 988 4771 992
rect 4733 828 4739 832
rect 4781 808 4787 1032
rect 4797 928 4803 1012
rect 4941 988 4947 1052
rect 4717 757 4739 763
rect 4701 688 4707 732
rect 4669 588 4675 612
rect 4557 468 4563 532
rect 4685 528 4691 652
rect 4717 548 4723 552
rect 4733 548 4739 757
rect 4749 668 4755 712
rect 4797 703 4803 912
rect 4829 848 4835 872
rect 4813 728 4819 732
rect 4829 708 4835 832
rect 4792 697 4803 703
rect 4765 688 4771 692
rect 4845 668 4851 952
rect 4925 928 4931 932
rect 4877 908 4883 912
rect 4920 737 4947 743
rect 4941 728 4947 737
rect 4877 697 4920 703
rect 4877 668 4883 697
rect 4893 668 4899 672
rect 4989 648 4995 892
rect 5005 808 5011 952
rect 5053 928 5059 1052
rect 5085 988 5091 1092
rect 5053 908 5059 912
rect 5117 888 5123 912
rect 5005 788 5011 792
rect 5005 708 5011 772
rect 4813 588 4819 592
rect 4845 548 4851 592
rect 4781 528 4787 532
rect 4589 517 4600 523
rect 4573 508 4579 512
rect 4525 388 4531 432
rect 4557 308 4563 392
rect 4589 328 4595 517
rect 4637 508 4643 512
rect 4621 488 4627 492
rect 4525 188 4531 252
rect 4589 168 4595 312
rect 4637 308 4643 312
rect 4653 288 4659 412
rect 4685 308 4691 392
rect 4605 188 4611 272
rect 4669 208 4675 272
rect 4733 228 4739 452
rect 4749 348 4755 512
rect 4781 428 4787 512
rect 4861 508 4867 632
rect 4845 428 4851 432
rect 4765 308 4771 392
rect 4781 388 4787 392
rect 4749 228 4755 252
rect 4765 208 4771 272
rect 4813 228 4819 312
rect 4845 308 4851 412
rect 4877 368 4883 512
rect 4909 488 4915 512
rect 4957 368 4963 432
rect 4909 348 4915 352
rect 4925 308 4931 312
rect 4829 288 4835 292
rect 4957 288 4963 292
rect 4973 288 4979 612
rect 5021 548 5027 652
rect 4989 368 4995 532
rect 5037 528 5043 712
rect 5069 708 5075 732
rect 5149 728 5155 1292
rect 5181 1188 5187 1497
rect 5197 1408 5203 1492
rect 5213 1488 5219 1512
rect 5245 1508 5251 1637
rect 5261 1508 5267 1512
rect 5245 1488 5251 1492
rect 5245 1368 5251 1472
rect 5181 1108 5187 1112
rect 5165 928 5171 972
rect 5181 948 5187 952
rect 5197 928 5203 1352
rect 5277 1328 5283 1792
rect 5309 1748 5315 1872
rect 5325 1768 5331 2112
rect 5357 1928 5363 2152
rect 5373 2148 5379 2252
rect 5437 2188 5443 2272
rect 5437 2088 5443 2112
rect 5421 1928 5427 1992
rect 5357 1908 5363 1912
rect 5341 1808 5347 1832
rect 5293 1448 5299 1512
rect 5213 1288 5219 1292
rect 5245 1248 5251 1312
rect 5309 1288 5315 1732
rect 5325 1668 5331 1714
rect 5357 1648 5363 1892
rect 5373 1848 5379 1872
rect 5389 1708 5395 1752
rect 5405 1728 5411 1792
rect 5421 1748 5427 1912
rect 5453 1888 5459 2212
rect 5485 2128 5491 2272
rect 5517 2208 5523 2272
rect 5565 2268 5571 2292
rect 5512 1937 5528 1943
rect 5549 1908 5555 1992
rect 5565 1943 5571 2232
rect 5629 2208 5635 2252
rect 5645 2188 5651 2312
rect 5661 2288 5667 2312
rect 5661 2268 5667 2272
rect 5677 2243 5683 2512
rect 5757 2508 5763 2512
rect 5693 2308 5699 2352
rect 5709 2308 5715 2492
rect 5789 2448 5795 2552
rect 5837 2548 5843 2572
rect 5853 2548 5859 2572
rect 5869 2568 5875 2612
rect 5805 2528 5811 2532
rect 5837 2528 5843 2532
rect 5901 2503 5907 2692
rect 5917 2637 5928 2643
rect 5917 2528 5923 2637
rect 5917 2508 5923 2512
rect 5885 2497 5907 2503
rect 5741 2428 5747 2432
rect 5805 2308 5811 2492
rect 5885 2388 5891 2497
rect 5901 2408 5907 2432
rect 5949 2368 5955 2552
rect 5981 2548 5987 2672
rect 5981 2428 5987 2532
rect 5997 2528 6003 2692
rect 6013 2508 6019 2512
rect 5981 2328 5987 2412
rect 5933 2308 5939 2312
rect 5773 2288 5779 2292
rect 5869 2268 5875 2276
rect 5661 2237 5683 2243
rect 5661 2148 5667 2237
rect 5789 2188 5795 2192
rect 5821 2148 5827 2252
rect 5837 2148 5843 2232
rect 5853 2148 5859 2232
rect 5885 2188 5891 2272
rect 5965 2268 5971 2272
rect 5901 2148 5907 2232
rect 5981 2148 5987 2312
rect 6029 2163 6035 2732
rect 6045 2728 6051 2732
rect 6093 2708 6099 2712
rect 6045 2588 6051 2632
rect 6061 2628 6067 2672
rect 6077 2648 6083 2692
rect 6109 2628 6115 2712
rect 6125 2708 6131 2712
rect 6205 2708 6211 2712
rect 6109 2608 6115 2612
rect 6045 2548 6051 2552
rect 6061 2528 6067 2592
rect 6077 2508 6083 2512
rect 6157 2488 6163 2692
rect 6173 2668 6179 2672
rect 6205 2608 6211 2672
rect 6221 2648 6227 2832
rect 6253 2708 6259 2892
rect 6301 2748 6307 3037
rect 6381 2968 6387 3292
rect 6397 2988 6403 3292
rect 6541 3208 6547 3312
rect 6557 3188 6563 3452
rect 6573 3308 6579 3372
rect 6653 3348 6659 3432
rect 6669 3428 6675 3457
rect 6589 3328 6595 3332
rect 6637 3128 6643 3232
rect 6653 3148 6659 3332
rect 6669 3328 6675 3412
rect 6717 3408 6723 3512
rect 6749 3388 6755 3476
rect 6781 3468 6787 4032
rect 6813 3928 6819 3932
rect 6813 3728 6819 3732
rect 6749 3348 6755 3352
rect 6781 3348 6787 3432
rect 6717 3308 6723 3312
rect 6701 3128 6707 3292
rect 6413 3028 6419 3032
rect 6381 2948 6387 2952
rect 6349 2708 6355 2912
rect 6237 2623 6243 2632
rect 6269 2628 6275 2632
rect 6221 2617 6243 2623
rect 6205 2548 6211 2572
rect 6221 2548 6227 2617
rect 6253 2548 6259 2592
rect 6285 2548 6291 2652
rect 6045 2308 6051 2352
rect 6061 2328 6067 2472
rect 6125 2388 6131 2452
rect 6173 2323 6179 2512
rect 6205 2388 6211 2472
rect 6173 2317 6195 2323
rect 6061 2228 6067 2272
rect 6093 2268 6099 2272
rect 6093 2248 6099 2252
rect 6173 2208 6179 2292
rect 6189 2183 6195 2317
rect 6269 2308 6275 2512
rect 6285 2448 6291 2532
rect 6301 2528 6307 2692
rect 6349 2588 6355 2672
rect 6365 2668 6371 2932
rect 6413 2908 6419 3012
rect 6477 2968 6483 3032
rect 6493 2988 6499 3072
rect 6413 2808 6419 2892
rect 6509 2888 6515 3092
rect 6541 2948 6547 3012
rect 6637 2968 6643 3012
rect 6557 2948 6563 2952
rect 6637 2948 6643 2952
rect 6669 2948 6675 2972
rect 6525 2908 6531 2912
rect 6333 2528 6339 2552
rect 6301 2488 6307 2512
rect 6333 2508 6339 2512
rect 6381 2428 6387 2672
rect 6397 2548 6403 2612
rect 6429 2588 6435 2732
rect 6477 2708 6483 2872
rect 6557 2848 6563 2912
rect 6589 2883 6595 2892
rect 6573 2877 6595 2883
rect 6477 2568 6483 2692
rect 6509 2688 6515 2712
rect 6541 2708 6547 2712
rect 6525 2588 6531 2672
rect 6184 2177 6195 2183
rect 6029 2157 6051 2163
rect 5565 1937 5587 1943
rect 5565 1908 5571 1912
rect 5581 1908 5587 1937
rect 5645 1888 5651 2132
rect 5661 1908 5667 2012
rect 5693 2008 5699 2072
rect 5773 2048 5779 2092
rect 5821 2088 5827 2112
rect 5917 2088 5923 2112
rect 6045 2108 6051 2157
rect 6109 2148 6115 2152
rect 6141 2148 6147 2172
rect 5997 2088 6003 2092
rect 5453 1808 5459 1872
rect 5501 1768 5507 1832
rect 5517 1768 5523 1832
rect 5613 1768 5619 1832
rect 5645 1748 5651 1872
rect 5661 1788 5667 1892
rect 5709 1888 5715 1972
rect 5725 1908 5731 1932
rect 5805 1908 5811 1912
rect 5693 1748 5699 1832
rect 5528 1737 5555 1743
rect 5549 1723 5555 1737
rect 5629 1728 5635 1732
rect 5549 1717 5560 1723
rect 5373 1508 5379 1632
rect 5453 1628 5459 1712
rect 5501 1528 5507 1712
rect 5533 1708 5539 1712
rect 5549 1688 5555 1692
rect 5629 1588 5635 1712
rect 5325 1248 5331 1472
rect 5373 1428 5379 1472
rect 5389 1468 5395 1512
rect 5453 1508 5459 1512
rect 5421 1388 5427 1392
rect 5213 1188 5219 1232
rect 5245 1108 5251 1192
rect 5213 948 5219 1032
rect 5261 928 5267 1232
rect 5309 1088 5315 1112
rect 5224 917 5235 923
rect 5197 788 5203 812
rect 5149 708 5155 712
rect 5165 708 5171 712
rect 5229 708 5235 917
rect 5245 908 5251 912
rect 5261 888 5267 912
rect 5261 728 5267 812
rect 5277 788 5283 1032
rect 5293 908 5299 1072
rect 5341 1008 5347 1092
rect 5357 1088 5363 1372
rect 5389 1128 5395 1332
rect 5453 1328 5459 1332
rect 5469 1328 5475 1472
rect 5485 1408 5491 1492
rect 5645 1488 5651 1732
rect 5661 1708 5667 1712
rect 5693 1568 5699 1632
rect 5709 1588 5715 1812
rect 5741 1788 5747 1892
rect 5837 1828 5843 1892
rect 5869 1888 5875 1972
rect 5885 1908 5891 1932
rect 5837 1788 5843 1812
rect 5725 1728 5731 1772
rect 5869 1768 5875 1872
rect 5773 1748 5779 1752
rect 5661 1488 5667 1512
rect 5533 1388 5539 1432
rect 5549 1388 5555 1472
rect 5581 1388 5587 1452
rect 5485 1348 5491 1352
rect 5501 1328 5507 1332
rect 5405 1148 5411 1312
rect 5485 1308 5491 1312
rect 5405 1128 5411 1132
rect 5485 1128 5491 1152
rect 5357 1028 5363 1072
rect 5373 1068 5379 1072
rect 5325 948 5331 972
rect 5341 928 5347 992
rect 5357 988 5363 1012
rect 5389 948 5395 1052
rect 5373 928 5379 932
rect 5309 748 5315 832
rect 5277 728 5283 732
rect 5229 688 5235 692
rect 5085 588 5091 672
rect 5101 548 5107 632
rect 5149 628 5155 672
rect 5149 588 5155 592
rect 5197 548 5203 552
rect 5213 548 5219 672
rect 5229 588 5235 632
rect 5069 508 5075 532
rect 5085 508 5091 512
rect 5005 308 5011 472
rect 5133 408 5139 512
rect 5149 468 5155 532
rect 5037 328 5043 352
rect 5084 317 5107 323
rect 5053 308 5059 312
rect 5101 308 5107 317
rect 4637 168 4643 172
rect 4829 148 4835 272
rect 4477 128 4483 132
rect 3981 28 3987 32
rect 3949 -43 3955 12
rect 4413 -37 4419 92
rect 4461 48 4467 112
rect 4413 -43 4435 -37
rect 4461 -43 4467 32
rect 4509 -43 4515 132
rect 4557 -43 4563 112
rect 4573 108 4579 112
rect 4621 -43 4627 132
rect 4701 128 4707 132
rect 4861 128 4867 172
rect 4877 148 4883 232
rect 4893 148 4899 272
rect 4941 263 4947 272
rect 4989 263 4995 272
rect 4941 257 4995 263
rect 4925 128 4931 252
rect 5005 188 5011 292
rect 5101 248 5107 272
rect 5133 268 5139 272
rect 5165 248 5171 272
rect 5048 237 5075 243
rect 4973 148 4979 152
rect 5069 128 5075 237
rect 5101 128 5107 232
rect 5181 223 5187 292
rect 5197 288 5203 392
rect 5245 368 5251 552
rect 5261 528 5267 692
rect 5325 688 5331 852
rect 5341 768 5347 912
rect 5405 728 5411 752
rect 5421 728 5427 1092
rect 5405 703 5411 712
rect 5405 697 5416 703
rect 5405 668 5411 672
rect 5437 663 5443 892
rect 5469 808 5475 912
rect 5485 903 5491 1032
rect 5501 988 5507 1312
rect 5533 1308 5539 1352
rect 5597 1348 5603 1472
rect 5645 1388 5651 1412
rect 5693 1408 5699 1552
rect 5613 1348 5619 1372
rect 5709 1368 5715 1372
rect 5725 1368 5731 1712
rect 5741 1708 5747 1732
rect 5773 1528 5779 1732
rect 5821 1728 5827 1732
rect 5805 1668 5811 1712
rect 5853 1708 5859 1712
rect 5837 1688 5843 1692
rect 5853 1568 5859 1692
rect 5885 1648 5891 1752
rect 5901 1708 5907 1732
rect 5757 1508 5763 1512
rect 5853 1508 5859 1532
rect 5885 1523 5891 1632
rect 5917 1608 5923 2072
rect 5933 1928 5939 1952
rect 5933 1868 5939 1912
rect 5997 1888 6003 1892
rect 6013 1888 6019 1972
rect 6029 1928 6035 2072
rect 6093 2068 6099 2132
rect 6141 2108 6147 2112
rect 6093 1988 6099 2052
rect 6093 1948 6099 1952
rect 6029 1908 6035 1912
rect 6013 1788 6019 1872
rect 5933 1708 5939 1712
rect 5885 1517 5896 1523
rect 5869 1508 5875 1512
rect 5805 1488 5811 1492
rect 5853 1488 5859 1492
rect 5821 1448 5827 1452
rect 5581 1308 5587 1312
rect 5597 1268 5603 1332
rect 5693 1308 5699 1332
rect 5773 1328 5779 1392
rect 5789 1328 5795 1372
rect 5837 1308 5843 1472
rect 5549 1108 5555 1132
rect 5597 1128 5603 1132
rect 5629 1108 5635 1232
rect 5661 1108 5667 1132
rect 5517 968 5523 992
rect 5581 988 5587 1032
rect 5517 948 5523 952
rect 5533 928 5539 972
rect 5581 948 5587 952
rect 5629 928 5635 1092
rect 5645 948 5651 1072
rect 5693 948 5699 1292
rect 5757 1188 5763 1232
rect 5853 1128 5859 1152
rect 5869 1128 5875 1492
rect 5901 1388 5907 1512
rect 5901 1308 5907 1332
rect 5917 1308 5923 1572
rect 5933 1468 5939 1692
rect 5997 1588 6003 1712
rect 6029 1703 6035 1892
rect 6045 1888 6051 1892
rect 6093 1888 6099 1932
rect 6109 1908 6115 2072
rect 6125 1888 6131 1892
rect 6109 1848 6115 1872
rect 6189 1868 6195 2132
rect 6269 2128 6275 2192
rect 6301 2148 6307 2232
rect 6349 2188 6355 2292
rect 6429 2288 6435 2432
rect 6445 2308 6451 2472
rect 6477 2348 6483 2552
rect 6493 2508 6499 2512
rect 6541 2508 6547 2552
rect 6573 2528 6579 2877
rect 6637 2788 6643 2832
rect 6637 2728 6643 2732
rect 6637 2528 6643 2692
rect 6669 2568 6675 2932
rect 6685 2908 6691 2912
rect 6701 2768 6707 2912
rect 6701 2708 6707 2712
rect 6717 2708 6723 3292
rect 6765 3188 6771 3292
rect 6749 3048 6755 3112
rect 6733 2968 6739 3032
rect 6781 2968 6787 3072
rect 6733 2923 6739 2932
rect 6813 2928 6819 2932
rect 6733 2917 6744 2923
rect 6717 2568 6723 2672
rect 6669 2528 6675 2532
rect 6477 2308 6483 2312
rect 6093 1748 6099 1812
rect 6109 1748 6115 1752
rect 6045 1728 6051 1732
rect 6013 1697 6035 1703
rect 6013 1588 6019 1697
rect 6013 1508 6019 1572
rect 6029 1528 6035 1552
rect 6045 1508 6051 1552
rect 5997 1368 6003 1472
rect 5933 1308 5939 1352
rect 6013 1348 6019 1372
rect 6061 1323 6067 1732
rect 6077 1728 6083 1732
rect 6125 1728 6131 1792
rect 6141 1528 6147 1692
rect 6157 1668 6163 1692
rect 6173 1688 6179 1692
rect 6205 1608 6211 2112
rect 6301 2108 6307 2132
rect 6349 2088 6355 2112
rect 6237 1908 6243 1992
rect 6237 1728 6243 1892
rect 6365 1888 6371 2132
rect 6381 2128 6387 2212
rect 6429 2168 6435 2272
rect 6381 1908 6387 2112
rect 6429 2108 6435 2112
rect 6365 1768 6371 1872
rect 6381 1828 6387 1892
rect 6429 1888 6435 1912
rect 6445 1768 6451 2292
rect 6509 2188 6515 2372
rect 6557 2308 6563 2472
rect 6573 2368 6579 2512
rect 6749 2463 6755 2652
rect 6733 2457 6755 2463
rect 6573 2308 6579 2332
rect 6605 2328 6611 2372
rect 6461 2128 6467 2132
rect 6477 2068 6483 2132
rect 6509 1968 6515 2032
rect 6509 1928 6515 1932
rect 6525 1928 6531 2292
rect 6637 2288 6643 2412
rect 6557 2268 6563 2272
rect 6541 2128 6547 2192
rect 6605 2148 6611 2152
rect 6621 2128 6627 2152
rect 6461 1908 6467 1912
rect 6589 1908 6595 2112
rect 6637 2008 6643 2272
rect 6653 1988 6659 2212
rect 6701 2128 6707 2132
rect 6717 2128 6723 2392
rect 6701 1948 6707 2112
rect 6477 1848 6483 1872
rect 6541 1868 6547 1892
rect 6605 1888 6611 1892
rect 6461 1808 6467 1832
rect 6573 1748 6579 1832
rect 6589 1828 6595 1872
rect 6621 1848 6627 1872
rect 6637 1848 6643 1912
rect 6733 1888 6739 2457
rect 6749 2388 6755 2432
rect 6765 2228 6771 2552
rect 6797 2388 6803 2532
rect 6653 1868 6659 1872
rect 6413 1728 6419 1732
rect 6253 1688 6259 1712
rect 6109 1508 6115 1512
rect 6077 1488 6083 1492
rect 6109 1468 6115 1492
rect 6125 1448 6131 1472
rect 6173 1468 6179 1592
rect 6365 1588 6371 1712
rect 6477 1588 6483 1714
rect 6669 1708 6675 1792
rect 6701 1788 6707 1832
rect 6205 1508 6211 1512
rect 6173 1408 6179 1452
rect 6189 1448 6195 1492
rect 6237 1488 6243 1532
rect 6269 1508 6275 1512
rect 6285 1488 6291 1492
rect 6301 1488 6307 1492
rect 6317 1488 6323 1572
rect 6413 1548 6419 1552
rect 6429 1508 6435 1512
rect 6253 1448 6259 1452
rect 6173 1388 6179 1392
rect 6221 1348 6227 1412
rect 6077 1328 6083 1332
rect 6141 1328 6147 1332
rect 6056 1317 6067 1323
rect 5933 1228 5939 1292
rect 5709 1008 5715 1072
rect 5725 1068 5731 1092
rect 5757 1088 5763 1092
rect 5645 928 5651 932
rect 5485 897 5496 903
rect 5469 708 5475 792
rect 5533 768 5539 832
rect 5533 728 5539 732
rect 5453 683 5459 692
rect 5453 677 5464 683
rect 5437 657 5459 663
rect 5341 548 5347 592
rect 5357 528 5363 632
rect 5389 628 5395 632
rect 5453 588 5459 657
rect 5261 508 5267 512
rect 5213 308 5219 352
rect 5245 328 5251 352
rect 5197 228 5203 272
rect 5176 217 5187 223
rect 5181 188 5187 217
rect 5245 208 5251 312
rect 5293 308 5299 312
rect 5261 228 5267 232
rect 5197 188 5203 192
rect 5293 188 5299 292
rect 5309 288 5315 392
rect 5389 383 5395 572
rect 5389 377 5411 383
rect 5405 368 5411 377
rect 5389 308 5395 352
rect 5336 297 5347 303
rect 5117 128 5123 152
rect 5309 128 5315 272
rect 5325 268 5331 272
rect 5341 228 5347 297
rect 5373 248 5379 272
rect 5357 208 5363 232
rect 5389 228 5395 292
rect 5405 268 5411 352
rect 4765 108 4771 114
rect 4829 108 4835 112
rect 4989 108 4995 112
rect 5325 108 5331 114
rect 5389 108 5395 192
rect 5421 128 5427 472
rect 5437 288 5443 512
rect 5453 308 5459 372
rect 5469 288 5475 632
rect 5517 528 5523 572
rect 5533 548 5539 552
rect 5549 528 5555 912
rect 5565 868 5571 892
rect 5565 688 5571 852
rect 5597 648 5603 912
rect 5613 728 5619 912
rect 5693 908 5699 912
rect 5629 708 5635 872
rect 5645 708 5651 832
rect 5613 628 5619 672
rect 5629 588 5635 692
rect 5661 608 5667 892
rect 5693 828 5699 892
rect 5709 688 5715 932
rect 5725 908 5731 1052
rect 5789 988 5795 1072
rect 5805 1048 5811 1092
rect 5837 1068 5843 1072
rect 5885 1068 5891 1072
rect 5981 1048 5987 1112
rect 6061 1108 6067 1317
rect 6077 1268 6083 1292
rect 5917 1037 5928 1043
rect 5821 948 5827 1032
rect 5853 948 5859 1012
rect 5869 943 5875 1032
rect 5869 937 5891 943
rect 5757 868 5763 932
rect 5821 768 5827 932
rect 5853 908 5859 912
rect 5757 728 5763 732
rect 5789 708 5795 712
rect 5853 708 5859 872
rect 5661 563 5667 592
rect 5677 568 5683 652
rect 5645 557 5667 563
rect 5645 548 5651 557
rect 5693 528 5699 532
rect 5725 528 5731 692
rect 5773 668 5779 672
rect 5773 548 5779 632
rect 5821 568 5827 632
rect 5629 517 5640 523
rect 5533 468 5539 492
rect 5485 308 5491 412
rect 5549 408 5555 512
rect 5629 508 5635 517
rect 5661 508 5667 512
rect 5709 488 5715 512
rect 5805 508 5811 512
rect 5741 488 5747 492
rect 5437 148 5443 192
rect 5453 168 5459 272
rect 5469 268 5475 272
rect 5469 148 5475 212
rect 5517 188 5523 192
rect 5533 123 5539 392
rect 5581 328 5587 432
rect 5597 388 5603 452
rect 5821 428 5827 532
rect 5869 528 5875 912
rect 5885 728 5891 937
rect 5901 908 5907 912
rect 5917 828 5923 1037
rect 5949 968 5955 972
rect 5997 948 6003 1032
rect 6013 948 6019 952
rect 5917 708 5923 772
rect 5949 728 5955 932
rect 6013 888 6019 912
rect 6029 863 6035 1072
rect 6045 1008 6051 1072
rect 6125 1068 6131 1252
rect 6061 1028 6067 1032
rect 6109 928 6115 932
rect 6141 928 6147 1312
rect 6157 1308 6163 1312
rect 6189 1208 6195 1312
rect 6205 1288 6211 1332
rect 6173 1108 6179 1192
rect 6221 1168 6227 1332
rect 6301 1328 6307 1472
rect 6461 1468 6467 1512
rect 6493 1488 6499 1652
rect 6701 1488 6707 1492
rect 6333 1348 6339 1432
rect 6349 1328 6355 1392
rect 6381 1303 6387 1452
rect 6445 1348 6451 1352
rect 6477 1348 6483 1352
rect 6509 1348 6515 1392
rect 6381 1297 6392 1303
rect 6253 1288 6259 1292
rect 6205 1108 6211 1132
rect 6221 1088 6227 1112
rect 6269 1088 6275 1152
rect 6365 1128 6371 1212
rect 6253 948 6259 1012
rect 6269 928 6275 992
rect 6013 857 6035 863
rect 5901 668 5907 672
rect 5917 588 5923 592
rect 5997 588 6003 692
rect 5677 328 5683 412
rect 5565 163 5571 312
rect 5581 308 5587 312
rect 5629 288 5635 312
rect 5693 288 5699 312
rect 5709 288 5715 292
rect 5565 157 5587 163
rect 5581 148 5587 157
rect 5661 148 5667 272
rect 5693 148 5699 252
rect 5725 168 5731 272
rect 5837 268 5843 492
rect 5869 448 5875 512
rect 5885 488 5891 532
rect 5997 528 6003 572
rect 6013 548 6019 857
rect 6029 723 6035 832
rect 6061 788 6067 852
rect 6109 788 6115 912
rect 6141 808 6147 832
rect 6269 828 6275 832
rect 6029 717 6051 723
rect 6029 548 6035 692
rect 6045 668 6051 717
rect 6141 708 6147 712
rect 6173 548 6179 752
rect 6269 708 6275 812
rect 6189 588 6195 672
rect 6237 548 6243 552
rect 6285 548 6291 1092
rect 6317 1068 6323 1112
rect 6333 1108 6339 1112
rect 6317 968 6323 1052
rect 6301 908 6307 912
rect 6301 728 6307 732
rect 6333 668 6339 852
rect 6013 508 6019 512
rect 6029 368 6035 532
rect 6141 408 6147 512
rect 6173 508 6179 532
rect 6221 528 6227 532
rect 6237 448 6243 512
rect 6253 488 6259 532
rect 6285 508 6291 512
rect 6301 508 6307 572
rect 6317 568 6323 632
rect 5837 168 5843 252
rect 5773 148 5779 152
rect 5869 148 5875 352
rect 5533 117 5544 123
rect 5405 108 5411 112
rect 5421 108 5427 112
rect 5597 108 5603 112
rect 5677 108 5683 112
rect 5917 108 5923 312
rect 6029 308 6035 332
rect 6093 308 6099 372
rect 6317 328 6323 532
rect 6333 528 6339 652
rect 6333 428 6339 512
rect 6109 288 6115 292
rect 5949 248 5955 272
rect 5997 268 6003 272
rect 6029 188 6035 232
rect 5933 168 5939 172
rect 6061 148 6067 232
rect 6173 143 6179 252
rect 6189 148 6195 292
rect 6269 288 6275 292
rect 6349 288 6355 1092
rect 6365 928 6371 1112
rect 6381 1048 6387 1297
rect 6429 1268 6435 1332
rect 6525 1328 6531 1332
rect 6461 1308 6467 1312
rect 6493 1188 6499 1312
rect 6557 1308 6563 1312
rect 6557 1288 6563 1292
rect 6397 1108 6403 1112
rect 6477 1108 6483 1132
rect 6493 1088 6499 1152
rect 6557 1108 6563 1172
rect 6573 1108 6579 1472
rect 6621 1388 6627 1452
rect 6701 1368 6707 1452
rect 6717 1388 6723 1872
rect 6733 1468 6739 1712
rect 6749 1708 6755 1852
rect 6765 1588 6771 1812
rect 6797 1748 6803 2052
rect 6749 1488 6755 1532
rect 6733 1368 6739 1432
rect 6781 1423 6787 1712
rect 6765 1417 6787 1423
rect 6621 1303 6627 1332
rect 6605 1297 6627 1303
rect 6605 1268 6611 1297
rect 6605 1128 6611 1252
rect 6669 1108 6675 1292
rect 6701 1188 6707 1352
rect 6381 948 6387 952
rect 6413 948 6419 972
rect 6429 948 6435 1032
rect 6461 908 6467 1032
rect 6477 888 6483 912
rect 6493 868 6499 1072
rect 6509 948 6515 1052
rect 6525 928 6531 1032
rect 6445 748 6451 832
rect 6509 728 6515 732
rect 6397 688 6403 692
rect 6413 588 6419 712
rect 6429 568 6435 632
rect 6477 568 6483 672
rect 6365 508 6371 532
rect 6157 137 6179 143
rect 5949 -43 5955 12
rect 6013 -37 6019 132
rect 6061 28 6067 112
rect 6077 108 6083 132
rect 6141 123 6147 132
rect 6136 117 6147 123
rect 5997 -43 6019 -37
rect 6029 -43 6035 12
rect 6077 -43 6083 72
rect 6157 -37 6163 137
rect 6189 128 6195 132
rect 6157 -43 6179 -37
rect 6253 -43 6259 152
rect 6349 148 6355 272
rect 6429 248 6435 532
rect 6509 528 6515 532
rect 6456 337 6467 343
rect 6461 308 6467 337
rect 6493 297 6504 303
rect 6493 288 6499 297
rect 6509 148 6515 152
rect 6525 128 6531 852
rect 6541 708 6547 872
rect 6557 848 6563 912
rect 6589 908 6595 912
rect 6605 708 6611 832
rect 6637 688 6643 972
rect 6701 948 6707 1052
rect 6685 928 6691 932
rect 6733 723 6739 1332
rect 6765 1168 6771 1417
rect 6797 1388 6803 1512
rect 6813 888 6819 1872
rect 6733 717 6755 723
rect 6653 708 6659 712
rect 6541 677 6552 683
rect 6541 588 6547 677
rect 6573 548 6579 552
rect 6621 528 6627 632
rect 6637 588 6643 672
rect 6653 508 6659 692
rect 6749 688 6755 717
rect 6701 388 6707 672
rect 6589 268 6595 352
rect 6637 297 6648 303
rect 6637 288 6643 297
rect 6541 -43 6547 232
rect 6701 148 6707 272
rect 6717 188 6723 412
rect 6749 368 6755 432
rect 6765 388 6771 392
rect 6781 288 6787 872
rect 6685 128 6691 132
<< m3contact >>
rect 8 4712 24 4728
rect 136 4692 152 4708
rect 184 4812 200 4828
rect 216 4812 232 4828
rect 360 4812 376 4828
rect 392 4812 408 4828
rect 248 4692 264 4708
rect 424 4692 440 4708
rect 632 4692 648 4708
rect 104 4652 120 4668
rect 136 4652 152 4668
rect 536 4672 552 4688
rect 584 4672 600 4688
rect 797 4802 833 4818
rect 792 4772 808 4788
rect 840 4772 856 4788
rect 936 4692 952 4708
rect 1112 4732 1128 4748
rect 1160 4732 1176 4748
rect 888 4672 904 4688
rect 920 4672 936 4688
rect 952 4672 968 4688
rect 568 4572 584 4588
rect 632 4572 648 4588
rect 456 4532 472 4548
rect 8 4512 24 4528
rect 264 4512 280 4528
rect 360 4512 376 4528
rect 424 4514 440 4528
rect 424 4512 440 4514
rect 696 4532 712 4548
rect 232 4472 248 4488
rect 40 4312 56 4328
rect 168 4312 184 4328
rect 8 4252 40 4268
rect 136 4252 152 4268
rect 8 4012 24 4028
rect 136 3972 152 3988
rect 8 3912 24 3928
rect 232 3912 248 3928
rect 56 3852 72 3868
rect 168 3852 184 3868
rect 296 4472 312 4488
rect 584 4472 600 4488
rect 664 4372 680 4388
rect 504 4352 520 4368
rect 600 4352 632 4368
rect 584 4332 600 4348
rect 408 4312 424 4328
rect 456 4312 468 4328
rect 468 4312 472 4328
rect 648 4312 664 4328
rect 280 4292 296 4308
rect 376 4272 392 4288
rect 424 4252 456 4268
rect 360 4232 376 4248
rect 296 4052 312 4068
rect 424 4212 440 4228
rect 488 4292 504 4308
rect 520 4292 536 4308
rect 632 4292 648 4308
rect 712 4352 728 4368
rect 680 4332 696 4348
rect 536 4272 552 4288
rect 600 4272 616 4288
rect 488 4192 504 4208
rect 472 4172 488 4188
rect 472 4132 488 4148
rect 408 4092 424 4108
rect 424 4072 440 4088
rect 408 4052 424 4068
rect 312 4032 328 4048
rect 360 4012 392 4028
rect 312 3972 328 3988
rect 296 3912 312 3928
rect 312 3892 328 3908
rect 360 3912 376 3928
rect 440 3912 456 3928
rect 392 3892 408 3908
rect 376 3852 392 3868
rect 248 3732 264 3748
rect 88 3712 104 3728
rect 184 3552 200 3568
rect 104 3512 120 3528
rect 232 3712 248 3728
rect 280 3712 296 3728
rect 296 3692 312 3708
rect 264 3652 280 3668
rect 360 3692 376 3708
rect 312 3632 328 3648
rect 360 3612 376 3628
rect 360 3552 376 3568
rect 216 3532 232 3548
rect 264 3532 280 3548
rect 296 3532 312 3548
rect 248 3512 264 3528
rect 280 3512 296 3528
rect 200 3492 216 3508
rect 184 3472 200 3488
rect 40 3352 56 3368
rect 136 3372 152 3388
rect 104 3352 120 3368
rect 88 3332 104 3348
rect 168 3352 184 3368
rect 56 3312 72 3328
rect 88 3312 104 3328
rect 120 3312 136 3328
rect 72 3292 88 3308
rect 24 3272 40 3288
rect 72 3232 88 3248
rect 152 3292 168 3308
rect 184 3292 200 3308
rect 88 3052 104 3068
rect 24 2892 40 2908
rect 8 2712 24 2728
rect 232 3452 248 3468
rect 232 3412 248 3428
rect 264 3392 280 3408
rect 248 3372 264 3388
rect 216 3292 232 3308
rect 216 3272 232 3288
rect 120 3032 136 3048
rect 184 2912 200 2928
rect 104 2852 120 2868
rect 248 3292 264 3308
rect 248 3112 264 3128
rect 232 3052 248 3068
rect 408 3812 424 3828
rect 440 3872 456 3888
rect 392 3732 408 3748
rect 424 3732 440 3748
rect 408 3712 424 3728
rect 424 3692 440 3708
rect 392 3672 408 3688
rect 504 4172 520 4188
rect 520 4072 536 4088
rect 520 3972 536 3988
rect 504 3892 520 3908
rect 504 3872 520 3888
rect 600 4232 616 4248
rect 680 4212 696 4228
rect 616 4152 632 4168
rect 552 4132 568 4148
rect 584 4092 600 4108
rect 552 3892 568 3908
rect 744 4572 760 4588
rect 936 4572 952 4588
rect 984 4672 1000 4688
rect 1000 4532 1016 4548
rect 968 4512 984 4528
rect 1064 4492 1080 4508
rect 1144 4692 1160 4708
rect 1176 4592 1192 4608
rect 1256 4706 1272 4708
rect 1256 4692 1272 4706
rect 1320 4692 1336 4708
rect 1464 4692 1480 4708
rect 1384 4652 1400 4668
rect 1432 4652 1448 4668
rect 1128 4572 1144 4588
rect 1240 4572 1256 4588
rect 1128 4552 1144 4568
rect 760 4472 776 4488
rect 1096 4472 1112 4488
rect 744 4352 760 4368
rect 744 4292 760 4308
rect 744 4172 760 4188
rect 1048 4432 1064 4448
rect 797 4402 833 4418
rect 856 4372 872 4388
rect 840 4352 856 4368
rect 824 4332 840 4348
rect 872 4352 888 4368
rect 936 4352 952 4368
rect 968 4352 984 4368
rect 888 4332 904 4348
rect 968 4332 984 4348
rect 1000 4332 1016 4348
rect 792 4272 808 4288
rect 760 4132 776 4148
rect 728 4112 744 4128
rect 664 4072 680 4088
rect 1096 4412 1112 4428
rect 1080 4392 1096 4408
rect 1144 4492 1160 4508
rect 1176 4472 1192 4488
rect 1240 4472 1256 4488
rect 1240 4412 1256 4428
rect 1128 4372 1144 4388
rect 1224 4372 1240 4388
rect 1176 4332 1192 4348
rect 1016 4312 1032 4328
rect 1048 4312 1064 4328
rect 1096 4312 1112 4328
rect 1128 4312 1144 4328
rect 1144 4312 1160 4328
rect 1208 4312 1224 4328
rect 1224 4312 1240 4328
rect 904 4292 920 4308
rect 1112 4292 1128 4308
rect 936 4272 952 4288
rect 1048 4272 1064 4288
rect 872 4212 888 4228
rect 968 4232 984 4248
rect 952 4192 968 4208
rect 1032 4192 1048 4208
rect 904 4172 920 4188
rect 824 4132 840 4148
rect 856 4132 888 4148
rect 760 4092 776 4108
rect 792 4092 808 4108
rect 824 4092 840 4108
rect 680 4032 696 4048
rect 648 4012 664 4028
rect 680 3952 696 3968
rect 648 3932 664 3948
rect 632 3892 648 3908
rect 744 3892 760 3908
rect 568 3872 584 3888
rect 536 3812 552 3828
rect 472 3792 488 3808
rect 552 3792 568 3808
rect 520 3752 536 3768
rect 456 3732 472 3748
rect 472 3732 488 3748
rect 456 3672 472 3688
rect 440 3552 456 3568
rect 392 3512 408 3528
rect 424 3512 440 3528
rect 408 3492 424 3508
rect 552 3712 568 3728
rect 488 3612 504 3628
rect 472 3532 488 3548
rect 504 3532 520 3548
rect 472 3512 488 3528
rect 312 3472 328 3488
rect 344 3472 360 3488
rect 360 3352 376 3368
rect 328 3332 344 3348
rect 376 3332 392 3348
rect 408 3332 424 3348
rect 280 3272 296 3288
rect 280 3152 296 3168
rect 408 3312 424 3328
rect 360 3292 376 3308
rect 312 3252 328 3268
rect 328 3232 344 3248
rect 312 3192 328 3208
rect 296 3132 312 3148
rect 440 3412 456 3428
rect 504 3472 520 3488
rect 472 3432 488 3448
rect 456 3392 472 3408
rect 440 3352 456 3368
rect 520 3412 536 3428
rect 504 3392 520 3408
rect 520 3352 536 3368
rect 568 3532 584 3548
rect 552 3512 568 3528
rect 616 3852 632 3868
rect 648 3832 664 3848
rect 920 4152 936 4168
rect 1096 4232 1112 4248
rect 936 4132 952 4148
rect 1000 4132 1016 4148
rect 888 4092 904 4108
rect 840 4072 856 4088
rect 968 4092 984 4108
rect 952 4052 968 4068
rect 797 4002 833 4018
rect 1032 4092 1048 4108
rect 1048 4092 1064 4108
rect 1096 4152 1112 4168
rect 1144 4292 1160 4308
rect 1400 4632 1416 4648
rect 1384 4592 1400 4608
rect 1288 4552 1304 4568
rect 1288 4532 1304 4548
rect 1384 4532 1400 4548
rect 1320 4512 1336 4528
rect 1272 4492 1288 4508
rect 1352 4412 1368 4428
rect 1288 4312 1304 4328
rect 1448 4472 1464 4488
rect 1416 4412 1432 4428
rect 1384 4292 1400 4308
rect 1160 4272 1176 4288
rect 1192 4272 1208 4288
rect 1224 4252 1240 4268
rect 1288 4252 1304 4268
rect 1128 4212 1144 4228
rect 1208 4152 1240 4168
rect 1256 4152 1272 4168
rect 1080 4132 1096 4148
rect 1128 4132 1144 4148
rect 1016 4072 1032 4088
rect 1064 4072 1080 4088
rect 1096 3992 1112 4008
rect 984 3972 1000 3988
rect 1080 3972 1112 3988
rect 808 3912 824 3928
rect 904 3912 920 3928
rect 1016 3912 1032 3928
rect 792 3892 808 3908
rect 984 3892 1000 3908
rect 760 3872 776 3888
rect 680 3772 696 3788
rect 712 3852 728 3868
rect 1096 3932 1112 3948
rect 872 3872 904 3888
rect 1096 3872 1112 3888
rect 776 3832 792 3848
rect 840 3832 856 3848
rect 696 3712 712 3728
rect 616 3532 632 3548
rect 664 3532 680 3548
rect 648 3512 664 3528
rect 584 3492 600 3508
rect 552 3472 568 3488
rect 568 3452 584 3468
rect 568 3372 584 3388
rect 584 3352 600 3368
rect 648 3432 664 3448
rect 632 3392 648 3408
rect 600 3332 632 3348
rect 648 3332 664 3348
rect 488 3292 504 3308
rect 680 3412 696 3428
rect 952 3852 968 3868
rect 968 3832 984 3848
rect 840 3752 856 3768
rect 744 3692 760 3708
rect 792 3672 808 3688
rect 776 3652 792 3668
rect 728 3632 744 3648
rect 712 3512 728 3528
rect 744 3492 760 3508
rect 696 3372 712 3388
rect 632 3292 648 3308
rect 584 3272 600 3288
rect 520 3252 536 3268
rect 696 3252 712 3268
rect 424 3192 440 3208
rect 408 3152 424 3168
rect 360 3112 376 3128
rect 392 3092 408 3108
rect 472 3132 488 3148
rect 296 3072 312 3088
rect 216 2972 232 2988
rect 296 2952 312 2968
rect 216 2932 232 2948
rect 280 2912 296 2928
rect 200 2892 216 2908
rect 264 2872 296 2888
rect 120 2832 136 2848
rect 280 2832 312 2848
rect 200 2772 216 2788
rect 120 2692 136 2708
rect 40 2652 56 2668
rect 120 2672 136 2688
rect 40 2532 56 2548
rect 24 2332 40 2348
rect 104 2512 120 2528
rect 72 2332 88 2348
rect 56 2312 72 2328
rect 152 2712 168 2728
rect 232 2712 248 2728
rect 136 2652 152 2668
rect 136 2572 152 2588
rect 168 2532 184 2548
rect 168 2512 184 2528
rect 152 2492 168 2508
rect 200 2492 216 2508
rect 152 2332 168 2348
rect 440 3032 456 3048
rect 424 2992 440 3008
rect 376 2972 392 2988
rect 344 2932 360 2948
rect 328 2912 344 2928
rect 328 2892 344 2908
rect 456 2932 472 2948
rect 440 2912 456 2928
rect 392 2892 408 2908
rect 360 2852 376 2868
rect 376 2832 392 2848
rect 392 2692 408 2708
rect 248 2412 264 2428
rect 216 2392 232 2408
rect 200 2332 232 2348
rect 168 2292 184 2308
rect 88 2272 104 2288
rect 40 2252 56 2268
rect 184 2232 200 2248
rect 264 2272 280 2288
rect 248 2212 264 2228
rect 184 2172 200 2188
rect 216 2172 232 2188
rect 328 2592 344 2608
rect 328 2492 360 2508
rect 312 2372 328 2388
rect 312 2332 328 2348
rect 296 2312 312 2328
rect 312 2312 328 2328
rect 344 2452 360 2468
rect 360 2292 376 2308
rect 120 2152 136 2168
rect 280 2152 296 2168
rect 184 2132 200 2148
rect 264 2132 280 2148
rect 312 2132 328 2148
rect 216 2112 232 2128
rect 104 1952 120 1968
rect 232 2092 248 2108
rect 280 2092 296 2108
rect 216 2072 232 2088
rect 248 2072 264 2088
rect 200 1912 216 1928
rect 200 1852 216 1868
rect 296 2032 312 2048
rect 264 1952 280 1968
rect 232 1892 248 1908
rect 264 1872 280 1888
rect 312 1912 328 1928
rect 408 2672 424 2688
rect 424 2632 440 2648
rect 616 3172 632 3188
rect 696 3152 712 3168
rect 520 3132 536 3148
rect 600 3132 616 3148
rect 600 3112 616 3128
rect 520 3052 552 3068
rect 536 2952 552 2968
rect 760 3472 776 3488
rect 744 3452 760 3468
rect 712 3112 728 3128
rect 712 3092 728 3108
rect 797 3602 833 3618
rect 824 3412 840 3428
rect 824 3372 840 3388
rect 920 3712 936 3728
rect 904 3692 920 3708
rect 984 3772 1000 3788
rect 920 3652 936 3668
rect 1016 3652 1032 3668
rect 968 3592 984 3608
rect 872 3552 888 3568
rect 904 3552 920 3568
rect 856 3512 872 3528
rect 936 3492 952 3508
rect 888 3432 904 3448
rect 872 3412 888 3428
rect 904 3412 920 3428
rect 792 3312 808 3328
rect 984 3552 1000 3568
rect 1032 3532 1048 3548
rect 1000 3512 1016 3528
rect 952 3472 968 3488
rect 1032 3472 1048 3488
rect 1064 3832 1080 3848
rect 1064 3812 1080 3828
rect 1160 4092 1176 4108
rect 1336 4132 1352 4148
rect 1304 4092 1320 4108
rect 1336 4092 1352 4108
rect 1272 4052 1288 4068
rect 1240 4032 1256 4048
rect 1272 4032 1288 4048
rect 1192 4012 1208 4028
rect 1224 4012 1240 4028
rect 1128 3912 1132 3928
rect 1132 3912 1144 3928
rect 1176 3912 1192 3928
rect 1464 4372 1496 4388
rect 1448 4292 1464 4308
rect 1432 4272 1448 4288
rect 1416 4252 1432 4268
rect 1416 4212 1432 4228
rect 1432 4192 1464 4208
rect 1368 4152 1384 4168
rect 1416 4152 1432 4168
rect 1384 4132 1400 4148
rect 1416 4112 1432 4128
rect 1432 4092 1448 4108
rect 1384 4072 1400 4088
rect 1448 4072 1464 4088
rect 1480 4312 1496 4328
rect 1560 4632 1576 4648
rect 1512 4572 1528 4588
rect 2861 4802 2897 4818
rect 3496 4812 3512 4828
rect 4909 4802 4945 4818
rect 6584 4812 6600 4828
rect 6616 4812 6632 4828
rect 5176 4772 5192 4788
rect 5224 4772 5240 4788
rect 5624 4772 5640 4788
rect 3864 4752 3880 4768
rect 4024 4752 4040 4768
rect 2728 4732 2744 4748
rect 2776 4732 2792 4748
rect 2168 4712 2184 4728
rect 2232 4712 2248 4728
rect 3336 4712 3352 4728
rect 2360 4706 2376 4708
rect 1720 4652 1736 4668
rect 2360 4692 2376 4706
rect 2504 4692 2520 4708
rect 2584 4692 2600 4708
rect 1880 4672 1896 4688
rect 2200 4672 2216 4688
rect 2392 4672 2408 4688
rect 2632 4672 2648 4688
rect 2264 4652 2280 4668
rect 2440 4652 2456 4668
rect 1832 4632 1848 4648
rect 1992 4632 2008 4648
rect 1592 4612 1608 4628
rect 1837 4602 1873 4618
rect 2232 4592 2248 4608
rect 1592 4572 1608 4588
rect 1688 4572 1704 4588
rect 1976 4572 1992 4588
rect 2216 4572 2232 4588
rect 1608 4532 1624 4548
rect 1688 4532 1704 4548
rect 1784 4532 1800 4548
rect 1832 4532 1848 4548
rect 1928 4532 1944 4548
rect 1528 4492 1544 4508
rect 1560 4492 1576 4508
rect 1576 4412 1592 4428
rect 1544 4292 1560 4308
rect 1528 4212 1544 4228
rect 1512 4192 1528 4208
rect 1512 4172 1528 4188
rect 1464 4052 1480 4068
rect 1528 4132 1544 4148
rect 1560 4272 1576 4288
rect 1640 4432 1656 4448
rect 1656 4372 1672 4388
rect 1640 4252 1656 4268
rect 1656 4232 1672 4248
rect 1576 4172 1592 4188
rect 1608 4172 1624 4188
rect 1608 4152 1624 4168
rect 1560 4132 1576 4148
rect 1720 4492 1736 4508
rect 1752 4432 1768 4448
rect 1704 4412 1720 4428
rect 2072 4532 2088 4548
rect 2088 4532 2104 4548
rect 2136 4532 2152 4548
rect 1912 4492 1928 4508
rect 1896 4472 1912 4488
rect 1816 4452 1832 4468
rect 1736 4372 1752 4388
rect 1800 4352 1816 4368
rect 1800 4332 1816 4348
rect 1736 4312 1752 4328
rect 1704 4212 1720 4228
rect 1656 4132 1672 4148
rect 1688 4132 1704 4148
rect 1496 4092 1512 4108
rect 1576 4032 1592 4048
rect 1608 4032 1624 4048
rect 1416 4012 1432 4028
rect 1480 4012 1496 4028
rect 1528 3972 1544 3988
rect 1352 3952 1368 3968
rect 1416 3952 1432 3968
rect 1304 3932 1320 3948
rect 1176 3892 1192 3908
rect 1192 3892 1208 3908
rect 1192 3872 1208 3888
rect 1224 3872 1240 3888
rect 1160 3812 1176 3828
rect 1144 3792 1160 3808
rect 1112 3772 1128 3788
rect 1144 3752 1160 3768
rect 1336 3852 1352 3868
rect 1272 3832 1288 3848
rect 1256 3812 1272 3828
rect 1208 3732 1224 3748
rect 1112 3612 1128 3628
rect 1080 3592 1096 3608
rect 1128 3592 1144 3608
rect 1112 3552 1128 3568
rect 1048 3452 1064 3468
rect 968 3432 984 3448
rect 1016 3432 1032 3448
rect 1032 3412 1048 3428
rect 984 3392 1016 3408
rect 888 3352 904 3368
rect 984 3332 1000 3348
rect 904 3312 920 3328
rect 792 3292 808 3308
rect 840 3292 856 3308
rect 840 3272 856 3288
rect 952 3292 968 3308
rect 936 3272 952 3288
rect 1000 3272 1016 3288
rect 904 3252 920 3268
rect 1000 3252 1016 3268
rect 797 3202 833 3218
rect 920 3152 936 3168
rect 808 3112 824 3128
rect 776 3092 792 3108
rect 904 3092 920 3108
rect 728 3072 744 3088
rect 632 3052 648 3068
rect 728 3052 744 3068
rect 616 2972 632 2988
rect 664 2952 680 2968
rect 568 2932 584 2948
rect 616 2932 632 2948
rect 648 2932 664 2948
rect 584 2912 600 2928
rect 520 2892 536 2908
rect 488 2872 504 2888
rect 488 2652 504 2668
rect 504 2632 520 2648
rect 472 2572 488 2588
rect 472 2552 488 2568
rect 456 2532 472 2548
rect 440 2512 456 2528
rect 424 2492 440 2508
rect 408 2432 424 2448
rect 408 2312 424 2328
rect 440 2312 456 2328
rect 552 2892 568 2908
rect 584 2892 600 2908
rect 584 2752 600 2768
rect 552 2552 568 2568
rect 488 2492 504 2508
rect 568 2512 584 2528
rect 648 2912 664 2928
rect 648 2832 664 2848
rect 616 2592 632 2608
rect 616 2572 632 2588
rect 856 3032 872 3048
rect 920 3032 936 3048
rect 888 3012 904 3028
rect 968 3012 984 3028
rect 968 2972 984 2988
rect 920 2952 936 2968
rect 712 2912 728 2928
rect 680 2892 696 2908
rect 712 2892 728 2908
rect 696 2852 712 2868
rect 680 2712 696 2728
rect 797 2802 833 2818
rect 856 2772 872 2788
rect 856 2752 872 2768
rect 712 2732 728 2748
rect 840 2732 856 2748
rect 872 2732 888 2748
rect 680 2552 696 2568
rect 648 2452 664 2468
rect 584 2412 616 2428
rect 520 2372 536 2388
rect 520 2312 536 2328
rect 488 2292 504 2308
rect 424 2272 440 2288
rect 472 2272 488 2288
rect 440 2252 456 2268
rect 472 2252 488 2268
rect 392 2212 408 2228
rect 504 2252 536 2268
rect 488 2232 504 2248
rect 376 2172 392 2188
rect 488 2172 504 2188
rect 392 2132 408 2148
rect 424 2132 440 2148
rect 360 2092 376 2108
rect 344 1892 360 1908
rect 376 1972 392 1988
rect 392 1932 408 1948
rect 664 2352 680 2368
rect 568 2252 584 2268
rect 600 2232 632 2248
rect 600 2172 616 2188
rect 536 2152 552 2168
rect 520 2132 536 2148
rect 584 2132 600 2148
rect 552 2112 568 2128
rect 648 2312 664 2328
rect 648 2292 664 2308
rect 904 2712 920 2728
rect 856 2692 872 2708
rect 984 2932 1000 2948
rect 936 2692 952 2708
rect 792 2672 808 2688
rect 840 2672 856 2688
rect 712 2652 728 2668
rect 744 2652 760 2668
rect 792 2652 808 2668
rect 744 2632 760 2648
rect 872 2572 888 2588
rect 728 2552 744 2568
rect 744 2532 760 2548
rect 856 2512 872 2528
rect 712 2492 728 2508
rect 840 2492 856 2508
rect 760 2452 776 2468
rect 712 2432 728 2448
rect 712 2312 728 2328
rect 824 2452 840 2468
rect 797 2402 833 2418
rect 840 2352 856 2368
rect 776 2332 792 2348
rect 776 2312 792 2328
rect 728 2252 744 2268
rect 680 2212 728 2228
rect 664 2192 680 2208
rect 776 2232 792 2248
rect 760 2172 776 2188
rect 760 2132 776 2148
rect 616 2112 632 2128
rect 440 2092 456 2108
rect 648 2072 664 2088
rect 584 1972 600 1988
rect 456 1932 472 1948
rect 488 1932 504 1948
rect 552 1932 568 1948
rect 424 1912 440 1928
rect 536 1912 552 1928
rect 552 1912 568 1928
rect 632 1912 636 1928
rect 636 1912 648 1928
rect 664 1912 680 1928
rect 520 1892 536 1908
rect 536 1892 552 1908
rect 600 1892 616 1908
rect 344 1872 360 1888
rect 424 1872 440 1888
rect 312 1852 328 1868
rect 280 1832 296 1848
rect 280 1812 296 1828
rect 184 1752 200 1768
rect 200 1752 216 1768
rect 232 1752 264 1768
rect 104 1572 120 1588
rect 232 1692 248 1708
rect 200 1572 216 1588
rect 120 1552 136 1568
rect 216 1552 232 1568
rect 120 1532 136 1548
rect 8 1492 24 1508
rect 88 1452 104 1468
rect 8 1312 24 1328
rect 168 1412 184 1428
rect 120 1392 136 1408
rect 104 1332 120 1348
rect 40 1272 56 1288
rect 24 1152 40 1168
rect 40 1132 56 1148
rect 40 1092 56 1108
rect 88 1092 104 1108
rect 72 1072 88 1088
rect 136 1352 152 1368
rect 232 1532 248 1548
rect 280 1572 296 1588
rect 232 1492 248 1508
rect 264 1492 280 1508
rect 264 1452 280 1468
rect 392 1852 408 1868
rect 360 1812 376 1828
rect 408 1792 424 1808
rect 360 1752 376 1768
rect 456 1832 472 1848
rect 424 1752 440 1768
rect 328 1672 344 1688
rect 312 1512 328 1528
rect 376 1692 392 1708
rect 344 1652 376 1668
rect 344 1592 360 1608
rect 376 1532 392 1548
rect 440 1712 456 1728
rect 424 1552 440 1568
rect 408 1512 424 1528
rect 488 1732 504 1748
rect 488 1692 504 1708
rect 456 1652 472 1668
rect 472 1632 488 1648
rect 376 1492 392 1508
rect 440 1492 456 1508
rect 552 1872 568 1888
rect 856 2272 872 2288
rect 904 2412 920 2428
rect 1080 3492 1096 3508
rect 1064 3392 1080 3408
rect 1096 3452 1112 3468
rect 1064 3312 1080 3328
rect 1240 3712 1256 3728
rect 1272 3792 1288 3808
rect 1176 3672 1192 3688
rect 1208 3672 1224 3688
rect 1256 3672 1272 3688
rect 1192 3512 1208 3528
rect 1336 3632 1352 3648
rect 1512 3912 1528 3928
rect 1544 3912 1560 3928
rect 1384 3852 1400 3868
rect 1496 3852 1512 3868
rect 1560 3852 1576 3868
rect 1496 3832 1512 3848
rect 1384 3712 1400 3728
rect 1448 3672 1464 3688
rect 1448 3632 1464 3648
rect 1352 3572 1368 3588
rect 1336 3432 1352 3448
rect 1208 3372 1224 3388
rect 1240 3372 1256 3388
rect 1176 3292 1192 3308
rect 1112 3252 1128 3268
rect 1144 3252 1160 3268
rect 1064 3232 1080 3248
rect 1016 3032 1032 3048
rect 1048 3012 1064 3028
rect 1032 2972 1048 2988
rect 1176 3152 1192 3168
rect 1240 3152 1256 3168
rect 1160 3132 1176 3148
rect 1096 3092 1112 3108
rect 1128 3092 1160 3108
rect 1144 3032 1160 3048
rect 1128 2992 1144 3008
rect 1224 3132 1256 3148
rect 1272 3112 1288 3128
rect 1336 3112 1352 3128
rect 1208 3092 1224 3108
rect 1256 3092 1272 3108
rect 1256 3072 1272 3088
rect 1192 3052 1208 3068
rect 1224 3032 1240 3048
rect 1176 2992 1192 3008
rect 1192 2952 1208 2968
rect 1144 2932 1160 2948
rect 1032 2912 1048 2928
rect 1112 2912 1128 2928
rect 984 2812 1000 2828
rect 968 2712 984 2728
rect 952 2592 968 2608
rect 984 2632 1000 2648
rect 952 2512 968 2528
rect 952 2492 968 2508
rect 1000 2492 1016 2508
rect 984 2452 1000 2468
rect 936 2412 952 2428
rect 936 2312 952 2328
rect 920 2292 936 2308
rect 1048 2892 1064 2908
rect 1080 2892 1096 2908
rect 1160 2892 1176 2908
rect 1096 2872 1112 2888
rect 1192 2812 1208 2828
rect 1048 2752 1064 2768
rect 1032 2692 1048 2708
rect 1064 2732 1080 2748
rect 1128 2732 1144 2748
rect 1176 2732 1192 2748
rect 1032 2672 1048 2688
rect 1144 2672 1160 2688
rect 1160 2652 1176 2668
rect 1096 2632 1112 2648
rect 1176 2592 1192 2608
rect 1128 2552 1144 2568
rect 1160 2532 1176 2548
rect 1160 2512 1176 2528
rect 1016 2432 1032 2448
rect 1032 2432 1048 2448
rect 1288 2932 1304 2948
rect 1320 3032 1336 3048
rect 1336 2972 1352 2988
rect 1320 2952 1336 2968
rect 1336 2912 1352 2928
rect 1304 2892 1320 2908
rect 1512 3792 1528 3808
rect 1576 3792 1592 3808
rect 1528 3712 1544 3728
rect 1480 3572 1496 3588
rect 1464 3512 1480 3528
rect 1464 3472 1480 3488
rect 1496 3372 1512 3388
rect 1400 3132 1416 3148
rect 1432 3112 1448 3128
rect 1400 3052 1416 3068
rect 1560 3692 1576 3708
rect 1576 3672 1592 3688
rect 1640 4072 1656 4088
rect 1656 4072 1672 4088
rect 1768 4272 1784 4288
rect 1784 4172 1800 4188
rect 1896 4432 1912 4448
rect 1896 4412 1912 4428
rect 1837 4202 1873 4218
rect 1800 4152 1832 4168
rect 1816 4132 1832 4148
rect 1672 4052 1688 4068
rect 1704 4052 1720 4068
rect 1624 3992 1640 4008
rect 1608 3752 1624 3768
rect 1624 3712 1640 3728
rect 1608 3692 1624 3708
rect 1656 3852 1672 3868
rect 1736 4072 1752 4088
rect 1800 4072 1816 4088
rect 1832 4072 1864 4088
rect 1720 3972 1736 3988
rect 1848 4032 1864 4048
rect 1704 3932 1720 3948
rect 1736 3932 1752 3948
rect 1688 3872 1704 3888
rect 1672 3772 1688 3788
rect 1688 3752 1704 3768
rect 1992 4472 2008 4488
rect 1960 4452 1976 4468
rect 2152 4512 2168 4528
rect 2040 4472 2072 4488
rect 2024 4412 2040 4428
rect 2024 4392 2040 4408
rect 1992 4372 2008 4388
rect 2104 4472 2120 4488
rect 2168 4472 2184 4488
rect 2120 4432 2136 4448
rect 2136 4412 2152 4428
rect 2088 4352 2104 4368
rect 2136 4352 2152 4368
rect 1976 4292 1992 4308
rect 1912 4272 1928 4288
rect 1944 4252 1960 4268
rect 1944 4232 1960 4248
rect 1992 4152 2008 4168
rect 2184 4432 2200 4448
rect 2200 4312 2216 4328
rect 2280 4572 2296 4588
rect 2568 4632 2584 4648
rect 2712 4632 2728 4648
rect 2760 4692 2776 4708
rect 2696 4612 2712 4628
rect 2744 4612 2760 4628
rect 2904 4706 2920 4708
rect 2904 4692 2920 4706
rect 3048 4692 3064 4708
rect 3224 4706 3240 4708
rect 3224 4692 3240 4706
rect 3288 4692 3304 4708
rect 2968 4672 2984 4688
rect 3256 4672 3272 4688
rect 2808 4632 2824 4648
rect 3016 4632 3032 4648
rect 2936 4612 2952 4628
rect 2792 4592 2808 4608
rect 2648 4572 2664 4588
rect 2840 4572 2856 4588
rect 2472 4532 2488 4548
rect 2552 4532 2568 4548
rect 2616 4532 2632 4548
rect 2392 4512 2408 4528
rect 2488 4492 2504 4508
rect 2264 4432 2280 4448
rect 2264 4412 2280 4428
rect 2280 4372 2296 4388
rect 2520 4452 2536 4468
rect 2680 4532 2696 4548
rect 2760 4532 2776 4548
rect 2808 4532 2824 4548
rect 2600 4512 2616 4528
rect 2632 4512 2648 4528
rect 2616 4412 2632 4428
rect 2568 4392 2584 4408
rect 2584 4372 2600 4388
rect 2600 4372 2616 4388
rect 2312 4332 2328 4348
rect 2392 4332 2408 4348
rect 2632 4332 2648 4348
rect 2248 4312 2264 4328
rect 2408 4312 2424 4328
rect 2440 4312 2456 4328
rect 2296 4292 2312 4308
rect 2232 4272 2248 4288
rect 2120 4252 2136 4268
rect 2152 4252 2168 4268
rect 2104 4232 2120 4248
rect 2056 4212 2072 4228
rect 2024 4192 2040 4208
rect 2072 4192 2088 4208
rect 2008 4112 2024 4128
rect 1944 4072 1960 4088
rect 1896 4052 1912 4068
rect 1880 4032 1896 4048
rect 1864 3952 1880 3968
rect 1928 3972 1944 3988
rect 1752 3872 1768 3888
rect 1816 3872 1832 3888
rect 1864 3872 1880 3888
rect 1880 3872 1896 3888
rect 1736 3852 1752 3868
rect 1800 3852 1816 3868
rect 1784 3792 1800 3808
rect 1837 3802 1873 3818
rect 1672 3732 1688 3748
rect 1736 3752 1752 3768
rect 1768 3752 1784 3768
rect 1832 3752 1848 3768
rect 1704 3732 1720 3748
rect 1784 3732 1800 3748
rect 1768 3712 1784 3728
rect 1816 3712 1832 3728
rect 1640 3612 1656 3628
rect 1592 3592 1608 3608
rect 1528 3512 1544 3528
rect 1560 3512 1576 3528
rect 1576 3512 1592 3528
rect 1624 3512 1640 3528
rect 1672 3512 1688 3528
rect 1640 3492 1656 3508
rect 1592 3452 1608 3468
rect 1560 3432 1576 3448
rect 1624 3432 1640 3448
rect 1544 3392 1560 3408
rect 1576 3352 1592 3368
rect 1528 3332 1544 3348
rect 1464 3232 1480 3248
rect 1480 3112 1496 3128
rect 1464 3032 1480 3048
rect 1496 3012 1512 3028
rect 1416 2972 1464 2988
rect 1368 2912 1384 2928
rect 1448 2952 1464 2968
rect 1560 3292 1576 3308
rect 1560 3032 1576 3048
rect 1752 3512 1768 3528
rect 1752 3492 1768 3508
rect 1768 3492 1784 3508
rect 1720 3472 1736 3488
rect 1704 3452 1720 3468
rect 1736 3452 1752 3468
rect 1688 3432 1704 3448
rect 1944 3772 1960 3788
rect 1928 3752 1944 3768
rect 1880 3732 1896 3748
rect 1800 3432 1816 3448
rect 1800 3412 1816 3428
rect 1816 3392 1832 3408
rect 1837 3402 1873 3418
rect 1800 3372 1816 3388
rect 2024 4092 2040 4108
rect 2024 3952 2040 3968
rect 1992 3932 2008 3948
rect 2072 4092 2088 4108
rect 2120 4212 2136 4228
rect 2136 4172 2152 4188
rect 2088 4072 2104 4088
rect 2072 4012 2088 4028
rect 2280 4212 2296 4228
rect 2232 4172 2248 4188
rect 2200 4112 2216 4128
rect 2280 4112 2296 4128
rect 2472 4272 2488 4288
rect 2312 4252 2328 4268
rect 2376 4252 2392 4268
rect 2408 4252 2424 4268
rect 2456 4232 2472 4248
rect 2344 4192 2360 4208
rect 2472 4192 2488 4208
rect 2312 4152 2328 4168
rect 2296 4092 2312 4108
rect 2312 4092 2328 4108
rect 2216 4072 2232 4088
rect 2248 4072 2264 4088
rect 2264 4032 2280 4048
rect 2344 4112 2360 4128
rect 2376 4112 2392 4128
rect 2392 4112 2408 4128
rect 2424 4112 2440 4128
rect 2344 4092 2360 4108
rect 2360 4092 2364 4108
rect 2364 4092 2376 4108
rect 2408 4092 2424 4108
rect 2328 4072 2344 4088
rect 2280 4012 2296 4028
rect 2200 3972 2216 3988
rect 2136 3932 2152 3948
rect 1976 3872 1992 3888
rect 1992 3832 2008 3848
rect 2008 3772 2024 3788
rect 1976 3732 1992 3748
rect 2024 3732 2040 3748
rect 1960 3712 1976 3728
rect 2008 3692 2024 3708
rect 2072 3812 2088 3828
rect 2104 3872 2120 3888
rect 2120 3852 2136 3868
rect 2104 3832 2120 3848
rect 2088 3752 2104 3768
rect 2536 4312 2552 4328
rect 2600 4312 2616 4328
rect 2568 4192 2584 4208
rect 2552 4172 2568 4188
rect 2600 4152 2616 4168
rect 2456 4112 2472 4128
rect 2552 4092 2568 4108
rect 2520 4052 2536 4068
rect 2392 4032 2408 4048
rect 2440 4032 2456 4048
rect 2328 3932 2344 3948
rect 2296 3912 2312 3928
rect 2520 4012 2536 4028
rect 2424 3992 2440 4008
rect 2184 3872 2200 3888
rect 2232 3872 2248 3888
rect 2072 3732 2088 3748
rect 2120 3712 2136 3728
rect 2200 3714 2216 3728
rect 2200 3712 2216 3714
rect 2088 3692 2104 3708
rect 1960 3672 1976 3688
rect 2040 3672 2056 3688
rect 2152 3652 2168 3668
rect 1976 3572 1992 3588
rect 1944 3492 1960 3508
rect 2088 3532 2104 3548
rect 2152 3532 2168 3548
rect 2008 3512 2024 3528
rect 2040 3492 2056 3508
rect 1912 3472 1928 3488
rect 1944 3472 1960 3488
rect 1896 3392 1912 3408
rect 2104 3452 2120 3468
rect 2088 3412 2104 3428
rect 2056 3392 2072 3408
rect 2008 3372 2024 3388
rect 1800 3352 1816 3368
rect 1864 3352 1880 3368
rect 2088 3352 2104 3368
rect 1672 3332 1688 3348
rect 1624 3312 1640 3328
rect 1624 3292 1640 3308
rect 1656 3292 1672 3308
rect 1688 3252 1704 3268
rect 1608 3172 1624 3188
rect 1592 3132 1608 3148
rect 1656 3132 1688 3148
rect 1624 3052 1640 3068
rect 1640 3052 1656 3068
rect 1624 3032 1640 3048
rect 1640 2992 1656 3008
rect 1560 2912 1576 2928
rect 1592 2912 1608 2928
rect 1528 2892 1544 2908
rect 1624 2892 1640 2908
rect 1464 2872 1480 2888
rect 1496 2872 1512 2888
rect 1624 2832 1640 2848
rect 1352 2812 1368 2828
rect 1400 2792 1416 2808
rect 1288 2772 1304 2788
rect 1304 2752 1320 2768
rect 1352 2752 1368 2768
rect 1272 2732 1304 2748
rect 1224 2692 1240 2708
rect 1256 2692 1272 2708
rect 1208 2632 1224 2648
rect 1192 2572 1208 2588
rect 1208 2532 1224 2548
rect 1368 2672 1384 2688
rect 1256 2652 1272 2668
rect 1240 2512 1256 2528
rect 1384 2632 1400 2648
rect 1432 2672 1448 2688
rect 1416 2652 1432 2668
rect 1400 2572 1416 2588
rect 1288 2532 1304 2548
rect 1208 2472 1224 2488
rect 1144 2452 1160 2468
rect 1112 2412 1128 2428
rect 1080 2352 1096 2368
rect 1064 2332 1080 2348
rect 968 2292 984 2308
rect 1080 2292 1096 2308
rect 1032 2272 1048 2288
rect 1096 2272 1112 2288
rect 952 2232 968 2248
rect 904 2212 920 2228
rect 920 2152 936 2168
rect 1224 2432 1240 2448
rect 1224 2412 1240 2428
rect 1224 2372 1240 2388
rect 1160 2352 1176 2368
rect 1128 2292 1144 2308
rect 1176 2312 1192 2328
rect 1112 2252 1128 2268
rect 1064 2212 1080 2228
rect 1016 2132 1032 2148
rect 712 1972 744 1988
rect 797 2002 833 2018
rect 744 1952 760 1968
rect 824 1952 840 1968
rect 744 1932 760 1948
rect 760 1932 776 1948
rect 680 1892 696 1908
rect 616 1852 632 1868
rect 600 1812 616 1828
rect 584 1772 600 1788
rect 632 1792 648 1808
rect 984 2032 1000 2048
rect 1016 2032 1032 2048
rect 936 1972 952 1988
rect 856 1932 872 1948
rect 872 1932 888 1948
rect 840 1912 856 1928
rect 696 1872 712 1888
rect 728 1872 744 1888
rect 776 1872 792 1888
rect 840 1872 856 1888
rect 664 1852 680 1868
rect 664 1832 680 1848
rect 1000 1952 1016 1968
rect 888 1892 904 1908
rect 904 1892 920 1908
rect 1112 2152 1128 2168
rect 1096 2032 1112 2048
rect 1064 1952 1080 1968
rect 1032 1932 1048 1948
rect 968 1872 984 1888
rect 1048 1872 1064 1888
rect 904 1852 920 1868
rect 952 1852 968 1868
rect 744 1772 760 1788
rect 856 1752 872 1768
rect 536 1692 552 1708
rect 584 1692 600 1708
rect 520 1632 536 1648
rect 600 1632 616 1648
rect 584 1512 600 1528
rect 632 1512 648 1528
rect 760 1712 776 1728
rect 696 1692 712 1708
rect 712 1692 728 1708
rect 680 1652 696 1668
rect 680 1632 696 1648
rect 504 1492 520 1508
rect 536 1492 552 1508
rect 328 1392 344 1408
rect 280 1332 296 1348
rect 312 1332 328 1348
rect 152 1312 168 1328
rect 184 1312 200 1328
rect 248 1272 264 1288
rect 248 1252 264 1268
rect 136 1172 152 1188
rect 152 1112 168 1128
rect 136 1072 152 1088
rect 8 952 24 968
rect 120 952 136 968
rect 72 932 88 948
rect 40 912 56 928
rect 8 712 24 728
rect 24 652 40 668
rect 136 912 152 928
rect 184 1152 200 1168
rect 232 1132 248 1148
rect 216 1092 232 1108
rect 328 1172 344 1188
rect 264 1112 280 1128
rect 312 1112 328 1128
rect 280 1092 296 1108
rect 184 1072 200 1088
rect 264 1032 280 1048
rect 184 992 216 1008
rect 200 972 216 988
rect 312 1052 328 1068
rect 296 992 312 1008
rect 280 952 296 968
rect 312 952 328 968
rect 216 912 232 928
rect 488 1452 504 1468
rect 392 1352 408 1368
rect 440 1332 456 1348
rect 376 1252 392 1268
rect 360 1232 376 1248
rect 376 1172 392 1188
rect 376 1152 392 1168
rect 168 892 184 908
rect 120 872 136 888
rect 232 872 248 888
rect 248 832 264 848
rect 264 772 280 788
rect 104 712 120 728
rect 152 712 168 728
rect 168 712 184 728
rect 136 692 152 708
rect 312 712 328 728
rect 344 832 360 848
rect 456 1152 472 1168
rect 440 1112 456 1128
rect 424 1092 440 1108
rect 392 1032 408 1048
rect 392 972 408 988
rect 376 932 392 948
rect 392 932 408 948
rect 440 832 456 848
rect 392 772 408 788
rect 440 732 456 748
rect 376 712 392 728
rect 200 692 216 708
rect 264 706 280 708
rect 264 692 280 706
rect 360 692 376 708
rect 184 672 200 688
rect 104 652 120 668
rect 328 592 344 608
rect 88 572 104 588
rect 280 572 296 588
rect 56 552 88 568
rect 136 552 152 568
rect 184 552 200 568
rect 40 532 56 548
rect 88 532 104 548
rect 168 532 184 548
rect 312 532 328 548
rect 8 512 24 528
rect 56 512 72 528
rect 200 512 216 528
rect 88 472 104 488
rect 8 312 24 328
rect 104 152 120 168
rect 136 152 152 168
rect 8 112 24 128
rect 136 112 152 128
rect 232 492 248 508
rect 440 692 456 708
rect 616 1492 632 1508
rect 632 1472 648 1488
rect 520 1432 536 1448
rect 568 1432 584 1448
rect 600 1432 616 1448
rect 600 1392 616 1408
rect 632 1392 648 1408
rect 616 1372 632 1388
rect 568 1132 584 1148
rect 616 1132 632 1148
rect 488 1112 520 1128
rect 472 1092 488 1108
rect 472 1012 488 1028
rect 792 1712 808 1728
rect 824 1692 840 1708
rect 776 1652 792 1668
rect 760 1632 776 1648
rect 797 1602 833 1618
rect 792 1572 808 1588
rect 744 1532 760 1548
rect 712 1512 716 1528
rect 716 1512 728 1528
rect 760 1512 776 1528
rect 680 1332 696 1348
rect 648 1052 664 1068
rect 568 992 584 1008
rect 632 992 648 1008
rect 488 932 504 948
rect 504 912 520 928
rect 520 832 536 848
rect 584 972 600 988
rect 632 932 648 948
rect 600 912 616 928
rect 824 1512 840 1528
rect 760 1472 776 1488
rect 744 1452 760 1468
rect 760 1432 776 1448
rect 776 1352 792 1368
rect 744 1292 760 1308
rect 776 1272 792 1288
rect 920 1832 936 1848
rect 1000 1792 1016 1808
rect 1128 1972 1144 1988
rect 1128 1912 1144 1928
rect 1160 2272 1176 2288
rect 1208 2272 1224 2288
rect 1208 2252 1224 2268
rect 1192 2212 1208 2228
rect 1208 2172 1224 2188
rect 1176 1992 1192 2008
rect 1096 1872 1112 1888
rect 1176 1872 1192 1888
rect 1064 1772 1080 1788
rect 1176 1752 1192 1768
rect 936 1732 952 1748
rect 968 1732 984 1748
rect 1064 1732 1080 1748
rect 904 1592 920 1608
rect 936 1592 952 1608
rect 888 1552 904 1568
rect 904 1532 920 1548
rect 968 1692 984 1708
rect 1016 1692 1036 1708
rect 1036 1692 1048 1708
rect 1080 1692 1096 1708
rect 1064 1652 1080 1668
rect 968 1632 984 1648
rect 1128 1712 1144 1728
rect 1160 1712 1176 1728
rect 1096 1612 1112 1628
rect 1096 1572 1112 1588
rect 1176 1572 1192 1588
rect 1016 1532 1032 1548
rect 1128 1532 1144 1548
rect 952 1512 984 1528
rect 840 1492 856 1508
rect 888 1492 904 1508
rect 952 1472 968 1488
rect 1048 1472 1064 1488
rect 1064 1472 1080 1488
rect 952 1432 968 1448
rect 888 1392 904 1408
rect 840 1372 856 1388
rect 856 1332 872 1348
rect 888 1312 904 1328
rect 936 1312 952 1328
rect 808 1232 824 1248
rect 797 1202 833 1218
rect 920 1292 936 1308
rect 984 1432 1000 1448
rect 968 1372 984 1388
rect 984 1312 1000 1328
rect 888 1212 904 1228
rect 840 1152 856 1168
rect 744 1132 760 1148
rect 952 1192 968 1208
rect 856 1112 872 1128
rect 920 1112 936 1128
rect 728 1092 744 1108
rect 680 912 696 928
rect 712 912 728 928
rect 584 872 600 888
rect 664 872 680 888
rect 520 732 536 748
rect 568 732 584 748
rect 760 1032 776 1048
rect 776 972 792 988
rect 792 952 808 968
rect 808 932 824 948
rect 872 932 888 948
rect 904 932 920 948
rect 728 852 760 868
rect 712 832 728 848
rect 664 732 680 748
rect 472 692 488 708
rect 584 692 600 708
rect 488 672 504 688
rect 456 652 472 668
rect 552 652 584 668
rect 408 572 424 588
rect 488 552 504 568
rect 600 592 616 608
rect 392 532 408 548
rect 472 532 488 548
rect 360 472 376 488
rect 200 432 216 448
rect 312 432 328 448
rect 360 352 376 368
rect 280 332 312 348
rect 344 332 360 348
rect 328 312 344 328
rect 312 292 328 308
rect 440 492 456 508
rect 488 492 504 508
rect 504 472 520 488
rect 568 472 584 488
rect 536 412 552 428
rect 520 372 536 388
rect 408 352 440 368
rect 408 332 424 348
rect 472 312 488 328
rect 536 352 552 368
rect 584 352 600 368
rect 568 312 584 328
rect 600 332 616 348
rect 408 272 424 288
rect 584 272 600 288
rect 248 232 264 248
rect 184 112 216 128
rect 248 112 264 128
rect 472 252 488 268
rect 680 692 696 708
rect 797 802 833 818
rect 792 732 808 748
rect 776 712 792 728
rect 632 492 648 508
rect 744 612 760 628
rect 1096 1412 1112 1428
rect 1144 1372 1160 1388
rect 1256 2472 1272 2488
rect 1272 2452 1288 2468
rect 1240 2312 1256 2328
rect 1240 2272 1256 2288
rect 1240 2132 1256 2148
rect 1304 2306 1320 2308
rect 1304 2292 1320 2306
rect 1304 2152 1320 2168
rect 1272 2112 1288 2128
rect 1304 2114 1320 2128
rect 1304 2112 1320 2114
rect 1592 2812 1608 2828
rect 1512 2772 1528 2788
rect 1464 2732 1480 2748
rect 1448 2492 1464 2508
rect 1400 2452 1416 2468
rect 1496 2632 1512 2648
rect 1496 2552 1512 2568
rect 1528 2752 1544 2768
rect 1608 2772 1624 2788
rect 1528 2712 1544 2728
rect 1592 2712 1608 2728
rect 1560 2672 1576 2688
rect 1576 2592 1592 2608
rect 1560 2572 1576 2588
rect 1480 2472 1496 2488
rect 1496 2432 1512 2448
rect 1464 2412 1480 2428
rect 1464 2392 1480 2408
rect 1432 2332 1448 2348
rect 1368 2312 1384 2328
rect 1368 2252 1384 2268
rect 1336 1952 1352 1968
rect 1256 1932 1272 1948
rect 1592 2492 1608 2508
rect 1528 2352 1544 2368
rect 1592 2352 1608 2368
rect 1512 2312 1528 2328
rect 1560 2312 1576 2328
rect 1512 2272 1528 2288
rect 1448 2232 1464 2248
rect 1544 2252 1560 2268
rect 1496 2172 1512 2188
rect 1464 2152 1480 2168
rect 1464 2132 1496 2148
rect 1512 2132 1528 2148
rect 1544 2132 1560 2148
rect 1400 2112 1416 2128
rect 1448 2032 1464 2048
rect 1480 2092 1496 2108
rect 1480 2032 1496 2048
rect 1592 2272 1608 2288
rect 1576 2232 1592 2248
rect 1736 3312 1752 3328
rect 1960 3332 1976 3348
rect 1880 3312 1896 3328
rect 1800 3292 1816 3308
rect 1896 3292 1912 3308
rect 1912 3292 1928 3308
rect 2008 3272 2024 3288
rect 1832 3152 1848 3168
rect 1912 3152 1928 3168
rect 1896 3132 1912 3148
rect 1720 3112 1736 3128
rect 1752 3112 1768 3128
rect 1832 3112 1848 3128
rect 1928 3112 1944 3128
rect 1992 3112 2008 3128
rect 1704 3092 1720 3108
rect 1800 3092 1816 3108
rect 1704 3052 1720 3068
rect 1736 3052 1752 3068
rect 1800 3052 1816 3068
rect 1880 3052 1896 3068
rect 2232 3852 2248 3868
rect 2248 3732 2264 3748
rect 2280 3852 2296 3868
rect 2312 3832 2328 3848
rect 2328 3832 2344 3848
rect 2296 3672 2312 3688
rect 2264 3572 2280 3588
rect 2280 3512 2296 3528
rect 2232 3492 2248 3508
rect 2216 3452 2232 3468
rect 2056 3292 2072 3308
rect 2120 3292 2136 3308
rect 2088 3232 2104 3248
rect 2024 3152 2056 3168
rect 2008 3092 2024 3108
rect 2056 3132 2072 3148
rect 1784 2992 1800 3008
rect 1837 3002 1873 3018
rect 1704 2972 1736 2988
rect 1688 2952 1704 2968
rect 1896 3032 1912 3048
rect 1944 3012 1960 3028
rect 1784 2952 1800 2968
rect 1928 2912 1944 2928
rect 1768 2892 1784 2908
rect 1800 2872 1816 2888
rect 1688 2832 1704 2848
rect 1656 2752 1672 2768
rect 1656 2672 1672 2688
rect 1656 2632 1672 2648
rect 1704 2632 1720 2648
rect 1624 2612 1656 2628
rect 1640 2512 1656 2528
rect 1624 2452 1640 2468
rect 1720 2592 1736 2608
rect 1704 2532 1720 2548
rect 1672 2472 1688 2488
rect 1704 2512 1720 2528
rect 1688 2432 1704 2448
rect 1656 2352 1672 2368
rect 1704 2312 1720 2328
rect 1672 2292 1704 2308
rect 1624 2272 1640 2288
rect 1640 2272 1656 2288
rect 1688 2272 1704 2288
rect 1608 2212 1624 2228
rect 1656 2192 1672 2208
rect 1576 2172 1592 2188
rect 1640 2152 1656 2168
rect 1624 2132 1640 2148
rect 1608 2112 1624 2128
rect 1560 2072 1576 2088
rect 1592 2072 1608 2088
rect 1496 2012 1528 2028
rect 1400 1952 1416 1968
rect 1464 1952 1480 1968
rect 1384 1912 1400 1928
rect 1448 1912 1464 1928
rect 1528 1912 1544 1928
rect 1560 1912 1576 1928
rect 1352 1872 1368 1888
rect 1384 1872 1400 1888
rect 1368 1832 1384 1848
rect 1320 1772 1336 1788
rect 1272 1732 1288 1748
rect 1304 1712 1320 1728
rect 1272 1692 1288 1708
rect 1240 1652 1256 1668
rect 1224 1632 1240 1648
rect 1224 1612 1240 1628
rect 1304 1532 1320 1548
rect 1288 1492 1304 1508
rect 1480 1892 1496 1908
rect 1512 1892 1528 1908
rect 1560 1892 1576 1908
rect 1592 1892 1608 1908
rect 1416 1872 1432 1888
rect 1464 1872 1480 1888
rect 1576 1872 1592 1888
rect 1448 1852 1464 1868
rect 1544 1852 1560 1868
rect 1592 1852 1608 1868
rect 1400 1832 1432 1848
rect 1400 1792 1416 1808
rect 1416 1732 1432 1748
rect 1560 1752 1592 1768
rect 1448 1732 1464 1748
rect 1528 1732 1544 1748
rect 1384 1612 1400 1628
rect 1352 1532 1368 1548
rect 1336 1492 1352 1508
rect 1208 1372 1224 1388
rect 1160 1352 1176 1368
rect 1192 1352 1208 1368
rect 1064 1332 1080 1348
rect 1144 1332 1160 1348
rect 1048 1272 1080 1288
rect 1032 1212 1048 1228
rect 968 1112 984 1128
rect 952 1052 968 1068
rect 936 1032 952 1048
rect 1016 1052 1032 1068
rect 1000 1032 1016 1048
rect 1112 1032 1128 1048
rect 1032 1012 1048 1028
rect 968 952 984 968
rect 1096 952 1112 968
rect 968 932 984 948
rect 1064 932 1080 948
rect 888 912 904 928
rect 1080 912 1096 928
rect 920 872 936 888
rect 952 872 968 888
rect 920 812 936 828
rect 872 692 888 708
rect 1064 892 1080 908
rect 984 872 1000 888
rect 968 852 984 868
rect 1016 772 1032 788
rect 1016 752 1032 768
rect 968 732 984 748
rect 936 712 952 728
rect 984 712 1016 728
rect 840 672 856 688
rect 968 592 984 608
rect 840 572 856 588
rect 920 572 936 588
rect 856 552 872 568
rect 984 572 1000 588
rect 1080 872 1096 888
rect 1064 832 1080 848
rect 1080 732 1096 748
rect 1080 692 1096 708
rect 1112 852 1128 868
rect 1128 792 1144 808
rect 1112 712 1128 728
rect 1304 1412 1320 1428
rect 1416 1532 1432 1548
rect 1672 2092 1688 2108
rect 1688 1952 1704 1968
rect 1656 1932 1672 1948
rect 1704 1912 1720 1928
rect 1672 1892 1688 1908
rect 1640 1832 1656 1848
rect 1672 1832 1688 1848
rect 1656 1752 1672 1768
rect 1784 2792 1800 2808
rect 1784 2752 1800 2768
rect 2024 2992 2040 3008
rect 1992 2952 2008 2968
rect 2040 2912 2056 2928
rect 1832 2892 1848 2908
rect 1912 2892 1928 2908
rect 1928 2892 1944 2908
rect 1880 2872 1896 2888
rect 1848 2812 1864 2828
rect 1768 2732 1784 2748
rect 1816 2732 1832 2748
rect 1752 2672 1768 2688
rect 1752 2572 1768 2588
rect 1752 2512 1768 2528
rect 1784 2692 1800 2708
rect 1832 2632 1848 2648
rect 1816 2612 1832 2628
rect 1837 2602 1873 2618
rect 1928 2812 1944 2828
rect 2264 3412 2280 3428
rect 2232 3332 2264 3348
rect 2200 3312 2216 3328
rect 2280 3372 2296 3388
rect 2536 3952 2552 3968
rect 2456 3912 2472 3928
rect 2584 4072 2600 4088
rect 2600 4052 2616 4068
rect 2632 4052 2648 4068
rect 2776 4512 2808 4528
rect 2824 4512 2840 4528
rect 2728 4452 2744 4468
rect 2792 4452 2808 4468
rect 2728 4412 2744 4428
rect 2712 4372 2728 4388
rect 2776 4352 2792 4368
rect 2744 4332 2776 4348
rect 2728 4292 2744 4308
rect 2696 4272 2712 4288
rect 2664 4252 2680 4268
rect 2680 4232 2696 4248
rect 2680 4192 2696 4208
rect 2664 4152 2680 4168
rect 2712 4172 2728 4188
rect 2664 4072 2680 4088
rect 2712 4072 2728 4088
rect 2664 4052 2680 4068
rect 2696 4052 2712 4068
rect 2648 3932 2664 3948
rect 2600 3912 2616 3928
rect 2552 3892 2568 3908
rect 2648 3892 2664 3908
rect 2456 3772 2472 3788
rect 2648 3772 2664 3788
rect 2392 3752 2408 3768
rect 2424 3752 2456 3768
rect 2488 3752 2504 3768
rect 2344 3732 2360 3748
rect 2792 4332 2808 4348
rect 2792 4312 2808 4328
rect 2792 4292 2808 4308
rect 2792 4232 2808 4248
rect 2776 4192 2792 4208
rect 2872 4532 2888 4548
rect 2968 4532 2984 4548
rect 2904 4492 2920 4508
rect 2861 4402 2897 4418
rect 2872 4372 2888 4388
rect 3000 4512 3016 4528
rect 2968 4492 2984 4508
rect 2936 4432 2952 4448
rect 2936 4392 2952 4408
rect 2920 4352 2936 4368
rect 2920 4312 2936 4328
rect 3096 4612 3112 4628
rect 3240 4612 3256 4628
rect 3096 4572 3112 4588
rect 3512 4712 3528 4728
rect 3544 4712 3560 4728
rect 3608 4712 3624 4728
rect 3400 4692 3416 4708
rect 3368 4652 3384 4668
rect 3400 4592 3432 4608
rect 3096 4532 3112 4548
rect 3080 4492 3096 4508
rect 3032 4472 3048 4488
rect 3128 4512 3144 4528
rect 3160 4512 3176 4528
rect 3208 4512 3224 4528
rect 3144 4492 3160 4508
rect 3112 4472 3128 4488
rect 3048 4432 3064 4448
rect 3176 4432 3192 4448
rect 3016 4412 3032 4428
rect 3112 4412 3128 4428
rect 3000 4352 3016 4368
rect 2952 4332 2968 4348
rect 2952 4312 2968 4328
rect 2936 4292 2952 4308
rect 3096 4372 3112 4388
rect 3032 4312 3048 4328
rect 3048 4292 3064 4308
rect 2920 4272 2936 4288
rect 2984 4272 3016 4288
rect 3064 4272 3080 4288
rect 3096 4272 3112 4288
rect 2888 4232 2904 4248
rect 2824 4212 2840 4228
rect 2872 4212 2888 4228
rect 2792 4172 2808 4188
rect 2776 4132 2792 4148
rect 2744 4032 2760 4048
rect 2744 3972 2760 3988
rect 2744 3912 2760 3928
rect 2728 3892 2744 3908
rect 2696 3872 2712 3888
rect 2744 3852 2760 3868
rect 2680 3812 2696 3828
rect 2664 3752 2680 3768
rect 2424 3732 2440 3748
rect 2504 3732 2520 3748
rect 2520 3732 2536 3748
rect 2568 3732 2584 3748
rect 2616 3732 2632 3748
rect 2344 3712 2360 3728
rect 2392 3712 2408 3728
rect 2328 3692 2344 3708
rect 2408 3692 2424 3708
rect 2360 3532 2376 3548
rect 2360 3492 2376 3508
rect 2344 3452 2360 3468
rect 2360 3412 2376 3428
rect 2344 3352 2360 3368
rect 2168 3292 2184 3308
rect 2184 3292 2200 3308
rect 2232 3292 2248 3308
rect 2152 3252 2168 3268
rect 2104 3212 2120 3228
rect 2136 3212 2152 3228
rect 2200 3212 2216 3228
rect 2328 3292 2344 3308
rect 2376 3292 2392 3308
rect 2360 3272 2392 3288
rect 2344 3252 2360 3268
rect 2296 3152 2312 3168
rect 2104 3112 2136 3128
rect 2152 3112 2168 3128
rect 2072 3072 2088 3088
rect 2088 3072 2104 3088
rect 1976 2872 1992 2888
rect 2024 2872 2040 2888
rect 2072 2772 2088 2788
rect 1960 2732 1976 2748
rect 1992 2732 2008 2748
rect 1960 2692 1976 2708
rect 1816 2572 1832 2588
rect 1800 2552 1816 2568
rect 1864 2532 1880 2548
rect 1912 2632 1928 2648
rect 1976 2652 1992 2668
rect 1944 2552 1960 2568
rect 1976 2532 1992 2548
rect 1896 2512 1912 2528
rect 1928 2512 1944 2528
rect 1960 2512 1976 2528
rect 1784 2392 1800 2408
rect 1800 2292 1816 2308
rect 1752 2272 1768 2288
rect 1768 2272 1784 2288
rect 1784 2232 1800 2248
rect 1752 2152 1768 2168
rect 1800 2092 1816 2108
rect 1800 2072 1816 2088
rect 1800 2032 1816 2048
rect 1928 2472 1944 2488
rect 2008 2672 2024 2688
rect 2008 2652 2024 2668
rect 2040 2732 2056 2748
rect 2072 2732 2088 2748
rect 2168 3092 2184 3108
rect 2200 3052 2216 3068
rect 2184 3032 2200 3048
rect 2216 2952 2232 2968
rect 2104 2872 2120 2888
rect 2136 2892 2152 2908
rect 2168 2892 2184 2908
rect 2184 2852 2200 2868
rect 2152 2832 2168 2848
rect 2120 2812 2136 2828
rect 2120 2752 2136 2768
rect 2136 2732 2152 2748
rect 2344 3092 2360 3108
rect 2296 3052 2312 3068
rect 2328 3052 2344 3068
rect 2248 3032 2264 3048
rect 2280 3032 2296 3048
rect 2312 3032 2328 3048
rect 2296 2972 2312 2988
rect 2264 2952 2280 2968
rect 2200 2832 2216 2848
rect 2200 2752 2216 2768
rect 2184 2632 2200 2648
rect 2168 2612 2184 2628
rect 2136 2592 2152 2608
rect 2104 2572 2120 2588
rect 2088 2552 2104 2568
rect 2024 2512 2040 2528
rect 2040 2472 2072 2488
rect 2104 2452 2120 2468
rect 2248 2852 2264 2868
rect 2232 2732 2248 2748
rect 2488 3672 2504 3688
rect 2632 3692 2664 3708
rect 2584 3652 2600 3668
rect 2440 3612 2456 3628
rect 2424 3472 2440 3488
rect 2424 3372 2440 3388
rect 2408 3352 2424 3368
rect 2408 3192 2424 3208
rect 2424 3172 2440 3188
rect 2424 3112 2440 3128
rect 2504 3532 2520 3548
rect 2600 3612 2616 3628
rect 2520 3492 2536 3508
rect 2584 3492 2600 3508
rect 2456 3372 2472 3388
rect 2456 3352 2472 3368
rect 2504 3472 2520 3488
rect 2472 3312 2488 3328
rect 2552 3392 2568 3408
rect 2520 3352 2536 3368
rect 2520 3312 2536 3328
rect 2536 3312 2552 3328
rect 2488 3292 2504 3308
rect 2600 3412 2616 3428
rect 2568 3252 2584 3268
rect 2616 3232 2632 3248
rect 2552 3212 2568 3228
rect 2616 3212 2632 3228
rect 2584 3172 2600 3188
rect 2552 3112 2568 3128
rect 2504 3092 2520 3108
rect 2424 3052 2440 3068
rect 2472 3052 2488 3068
rect 2408 3032 2424 3048
rect 2392 3012 2408 3028
rect 2376 2972 2392 2988
rect 2376 2952 2408 2968
rect 2296 2892 2312 2908
rect 2280 2872 2296 2888
rect 2264 2812 2280 2828
rect 2456 3032 2472 3048
rect 2312 2872 2328 2888
rect 2344 2872 2360 2888
rect 2280 2652 2296 2668
rect 2168 2512 2184 2528
rect 2168 2452 2200 2468
rect 2120 2412 2136 2428
rect 2264 2572 2280 2588
rect 2264 2512 2280 2528
rect 2248 2432 2264 2448
rect 2232 2392 2248 2408
rect 2152 2352 2168 2368
rect 1896 2332 1912 2348
rect 1976 2292 1992 2308
rect 2040 2272 2072 2288
rect 2008 2252 2040 2268
rect 1880 2232 1896 2248
rect 1837 2202 1873 2218
rect 1928 2232 1944 2248
rect 1976 2232 2008 2248
rect 1960 2212 1976 2228
rect 1928 2152 1944 2168
rect 1816 2012 1832 2028
rect 1784 1892 1800 1908
rect 1736 1872 1752 1888
rect 1784 1872 1800 1888
rect 1720 1812 1736 1828
rect 1736 1792 1752 1808
rect 1752 1752 1784 1768
rect 1592 1732 1624 1748
rect 1688 1732 1704 1748
rect 1704 1732 1720 1748
rect 1480 1712 1496 1728
rect 1512 1712 1528 1728
rect 1576 1672 1592 1688
rect 1560 1632 1576 1648
rect 1528 1612 1544 1628
rect 1480 1592 1496 1608
rect 1464 1512 1480 1528
rect 1384 1412 1400 1428
rect 1304 1392 1336 1408
rect 1288 1352 1304 1368
rect 1432 1452 1448 1468
rect 1512 1532 1528 1548
rect 1448 1412 1464 1428
rect 1480 1432 1496 1448
rect 1464 1392 1480 1408
rect 1496 1392 1512 1408
rect 1256 1332 1272 1348
rect 1336 1332 1352 1348
rect 1416 1332 1432 1348
rect 1336 1312 1352 1328
rect 1400 1312 1416 1328
rect 1464 1312 1480 1328
rect 1272 1292 1304 1308
rect 1320 1272 1336 1288
rect 1256 1252 1272 1268
rect 1192 1232 1208 1248
rect 1224 1052 1240 1068
rect 1160 1032 1176 1048
rect 1224 1012 1256 1028
rect 1208 992 1224 1008
rect 1192 912 1208 928
rect 1208 872 1224 888
rect 1192 772 1208 788
rect 1208 752 1224 768
rect 1272 1212 1288 1228
rect 1304 1212 1320 1228
rect 1288 1152 1304 1168
rect 1368 1232 1384 1248
rect 1368 1212 1384 1228
rect 1544 1492 1560 1508
rect 1592 1652 1608 1668
rect 1624 1632 1640 1648
rect 1688 1712 1704 1728
rect 1672 1572 1688 1588
rect 1656 1532 1672 1548
rect 1608 1512 1624 1528
rect 1784 1712 1800 1728
rect 1736 1572 1752 1588
rect 1608 1432 1624 1448
rect 1592 1412 1608 1428
rect 1560 1352 1576 1368
rect 1560 1332 1576 1348
rect 1512 1312 1528 1328
rect 1560 1312 1576 1328
rect 1624 1352 1640 1368
rect 1592 1292 1608 1308
rect 1832 1892 1848 1908
rect 1880 1932 1896 1948
rect 1864 1892 1880 1908
rect 1848 1872 1864 1888
rect 1912 1872 1928 1888
rect 1832 1852 1848 1868
rect 1837 1802 1873 1818
rect 1880 1752 1896 1768
rect 1928 1852 1944 1868
rect 1848 1732 1864 1748
rect 1896 1732 1912 1748
rect 1864 1672 1880 1688
rect 1976 2092 1992 2108
rect 2120 2292 2136 2308
rect 2168 2332 2184 2348
rect 2136 2272 2152 2288
rect 2200 2272 2216 2288
rect 2072 2232 2088 2248
rect 2232 2292 2248 2308
rect 2248 2292 2264 2308
rect 2200 2232 2232 2248
rect 2088 2212 2104 2228
rect 2120 2192 2136 2208
rect 2216 2192 2232 2208
rect 2136 2172 2152 2188
rect 2360 2792 2392 2808
rect 2408 2892 2424 2908
rect 2408 2752 2424 2768
rect 2328 2652 2344 2668
rect 2392 2652 2408 2668
rect 2376 2632 2392 2648
rect 2440 2852 2456 2868
rect 2440 2672 2456 2688
rect 2344 2572 2360 2588
rect 2376 2572 2408 2588
rect 2360 2552 2376 2568
rect 2472 2872 2488 2888
rect 2616 3152 2632 3168
rect 2600 3092 2616 3108
rect 2648 3512 2664 3528
rect 2648 3452 2664 3468
rect 2648 3412 2664 3428
rect 2712 3792 2728 3808
rect 2728 3752 2744 3768
rect 2696 3712 2712 3728
rect 2776 4112 2792 4128
rect 2776 3952 2792 3968
rect 3064 4232 3080 4248
rect 3048 4212 3064 4228
rect 2936 4192 2952 4208
rect 2872 4152 2888 4168
rect 2920 4152 2936 4168
rect 3032 4152 3048 4168
rect 2856 4112 2872 4128
rect 2808 4072 2824 4088
rect 2888 4052 2904 4068
rect 2861 4002 2897 4018
rect 2952 4132 2968 4148
rect 2984 4112 3000 4128
rect 2952 4072 2968 4088
rect 3016 4052 3032 4068
rect 2920 4032 2936 4048
rect 2840 3972 2856 3988
rect 2904 3972 2920 3988
rect 2840 3912 2856 3928
rect 2776 3872 2792 3888
rect 3240 4432 3256 4448
rect 3208 4372 3224 4388
rect 3240 4352 3256 4368
rect 3128 4332 3144 4348
rect 3160 4332 3176 4348
rect 3128 4272 3144 4288
rect 3320 4492 3336 4508
rect 3384 4452 3400 4468
rect 3304 4412 3320 4428
rect 3336 4412 3352 4428
rect 3576 4672 3592 4688
rect 3656 4712 3672 4728
rect 3688 4712 3704 4728
rect 3672 4672 3688 4688
rect 3720 4692 3736 4708
rect 4040 4732 4056 4748
rect 4296 4732 4312 4748
rect 4840 4732 4856 4748
rect 4904 4732 4920 4748
rect 4984 4732 5000 4748
rect 3720 4652 3736 4668
rect 3896 4652 3912 4668
rect 3640 4572 3656 4588
rect 3432 4552 3448 4568
rect 3560 4552 3576 4568
rect 3704 4552 3720 4568
rect 3496 4532 3512 4548
rect 3416 4512 3432 4528
rect 3480 4512 3496 4528
rect 3496 4512 3512 4528
rect 3464 4492 3468 4508
rect 3468 4492 3480 4508
rect 3512 4492 3528 4508
rect 3448 4452 3464 4468
rect 3576 4512 3592 4528
rect 3544 4432 3560 4448
rect 3448 4392 3464 4408
rect 3288 4352 3304 4368
rect 3336 4352 3352 4368
rect 3320 4332 3336 4348
rect 3336 4332 3352 4348
rect 3272 4312 3288 4328
rect 3256 4292 3272 4308
rect 3320 4292 3336 4308
rect 3208 4272 3224 4288
rect 3176 4252 3192 4268
rect 3192 4212 3208 4228
rect 3336 4192 3368 4208
rect 3128 4172 3144 4188
rect 3176 4172 3192 4188
rect 3320 4172 3336 4188
rect 3064 4132 3080 4148
rect 3096 4132 3112 4148
rect 3064 4052 3080 4068
rect 3080 4032 3096 4048
rect 3016 4012 3032 4028
rect 3048 4012 3064 4028
rect 3000 3952 3016 3968
rect 2968 3932 2984 3948
rect 2936 3892 2952 3908
rect 2760 3772 2776 3788
rect 2760 3752 2776 3768
rect 2744 3672 2760 3688
rect 2760 3652 2776 3668
rect 2744 3612 2760 3628
rect 2728 3532 2744 3548
rect 2696 3492 2712 3508
rect 2744 3472 2760 3488
rect 2696 3452 2712 3468
rect 2760 3412 2776 3428
rect 2760 3352 2776 3368
rect 2760 3332 2776 3348
rect 2680 3272 2696 3288
rect 2664 3132 2680 3148
rect 2696 3132 2712 3148
rect 2728 3112 2744 3128
rect 2760 3112 2776 3128
rect 2712 3092 2728 3108
rect 2760 3092 2776 3108
rect 2696 3072 2712 3088
rect 2520 3052 2552 3068
rect 2568 3052 2584 3068
rect 2648 3052 2664 3068
rect 2616 3012 2632 3028
rect 2632 2992 2648 3008
rect 2728 3052 2744 3068
rect 2680 2932 2696 2948
rect 2488 2852 2504 2868
rect 2488 2832 2504 2848
rect 2456 2652 2472 2668
rect 2472 2592 2488 2608
rect 2328 2532 2360 2548
rect 2456 2532 2488 2548
rect 2328 2472 2344 2488
rect 2312 2372 2328 2388
rect 2312 2352 2328 2368
rect 2376 2412 2392 2428
rect 2424 2412 2456 2428
rect 2344 2332 2360 2348
rect 2424 2312 2440 2328
rect 2344 2232 2360 2248
rect 2408 2272 2424 2288
rect 2392 2232 2408 2248
rect 2360 2212 2376 2228
rect 2280 2192 2296 2208
rect 2264 2152 2280 2168
rect 2328 2152 2344 2168
rect 2232 2132 2248 2148
rect 2296 2132 2312 2148
rect 2088 2112 2104 2128
rect 2008 2092 2024 2108
rect 2072 2092 2088 2108
rect 2056 2072 2072 2088
rect 2008 2052 2024 2068
rect 2040 2052 2056 2068
rect 2104 2052 2120 2068
rect 2168 2072 2184 2088
rect 1992 1972 2008 1988
rect 1960 1912 1976 1928
rect 2072 2012 2088 2028
rect 2056 1912 2072 1928
rect 2072 1912 2088 1928
rect 2040 1892 2056 1908
rect 1992 1852 2008 1868
rect 1960 1792 1976 1808
rect 1960 1732 1976 1748
rect 1944 1692 1960 1708
rect 1928 1632 1944 1648
rect 2232 2092 2248 2108
rect 2200 2072 2216 2088
rect 2072 1752 2088 1768
rect 2152 1872 2168 1888
rect 2120 1852 2136 1868
rect 2152 1852 2168 1868
rect 2120 1792 2136 1808
rect 2024 1712 2040 1728
rect 1992 1672 2008 1688
rect 1976 1652 1992 1668
rect 1976 1632 1992 1648
rect 1960 1592 1976 1608
rect 2008 1612 2024 1628
rect 2040 1612 2056 1628
rect 2008 1592 2024 1608
rect 2040 1552 2056 1568
rect 1832 1492 1848 1508
rect 2040 1492 2056 1508
rect 1704 1472 1720 1488
rect 1816 1472 1832 1488
rect 1688 1392 1704 1408
rect 2040 1472 2056 1488
rect 1992 1452 2008 1468
rect 1800 1412 1816 1428
rect 1837 1402 1873 1418
rect 1976 1412 1992 1428
rect 1736 1372 1752 1388
rect 1752 1352 1768 1368
rect 2056 1392 2072 1408
rect 2088 1712 2104 1728
rect 2072 1352 2088 1368
rect 1656 1332 1672 1348
rect 1736 1332 1752 1348
rect 1912 1332 1928 1348
rect 1992 1332 2008 1348
rect 1544 1272 1560 1288
rect 1528 1232 1544 1248
rect 1560 1232 1576 1248
rect 1480 1192 1496 1208
rect 1464 1112 1480 1128
rect 1336 1092 1352 1108
rect 1352 1092 1368 1108
rect 1544 1092 1560 1108
rect 1608 1092 1624 1108
rect 1272 992 1288 1008
rect 1368 1052 1384 1068
rect 1352 1032 1368 1048
rect 1320 1012 1336 1028
rect 1576 1072 1592 1088
rect 1464 1052 1480 1068
rect 1560 1052 1576 1068
rect 1528 1012 1544 1028
rect 1416 992 1432 1008
rect 1544 992 1576 1008
rect 1352 972 1368 988
rect 1400 972 1416 988
rect 1464 972 1480 988
rect 1544 972 1560 988
rect 1304 932 1320 948
rect 1320 912 1336 928
rect 1272 832 1288 848
rect 1336 812 1352 828
rect 1304 792 1320 808
rect 1288 772 1304 788
rect 1256 732 1272 748
rect 1160 712 1176 728
rect 1160 692 1176 708
rect 1208 692 1224 708
rect 1240 692 1256 708
rect 1272 692 1288 708
rect 1368 932 1384 948
rect 1432 932 1448 948
rect 1368 892 1384 908
rect 1432 912 1448 928
rect 1496 932 1512 948
rect 1640 1072 1656 1088
rect 1672 1092 1688 1108
rect 1672 1052 1688 1068
rect 1656 1012 1672 1028
rect 1576 952 1592 968
rect 1640 932 1656 948
rect 1544 912 1560 928
rect 1704 1092 1720 1108
rect 2024 1272 2040 1288
rect 1784 1252 1800 1268
rect 1976 1232 1992 1248
rect 2072 1172 2088 1188
rect 2024 1112 2040 1128
rect 2248 2052 2264 2068
rect 2328 2072 2344 2088
rect 2264 1992 2280 2008
rect 2328 1992 2344 2008
rect 2264 1952 2280 1968
rect 2408 2212 2424 2228
rect 2392 2112 2408 2128
rect 2408 2112 2424 2128
rect 2424 2112 2440 2128
rect 2408 1992 2424 2008
rect 2504 2812 2520 2828
rect 2504 2652 2520 2668
rect 2536 2912 2552 2928
rect 2584 2872 2600 2888
rect 2552 2852 2568 2868
rect 2568 2732 2584 2748
rect 2536 2652 2552 2668
rect 2728 2912 2744 2928
rect 2632 2672 2648 2688
rect 2696 2892 2712 2908
rect 2680 2812 2696 2828
rect 2760 2892 2776 2908
rect 2744 2792 2760 2808
rect 2728 2752 2744 2768
rect 2696 2692 2712 2708
rect 2712 2692 2728 2708
rect 3032 3952 3048 3968
rect 3112 3952 3128 3968
rect 2904 3852 2920 3868
rect 2952 3852 2968 3868
rect 2984 3852 3000 3868
rect 2888 3792 2904 3808
rect 3048 3932 3064 3948
rect 3080 3932 3096 3948
rect 3160 4112 3176 4128
rect 3192 4092 3208 4108
rect 3256 4092 3272 4108
rect 3208 4072 3224 4088
rect 3160 4052 3176 4068
rect 3256 4052 3272 4068
rect 3416 4306 3432 4308
rect 3416 4292 3432 4306
rect 3416 4192 3432 4208
rect 3480 4312 3496 4328
rect 3608 4492 3624 4508
rect 3704 4452 3720 4468
rect 3672 4432 3688 4448
rect 3656 4412 3672 4428
rect 3640 4312 3656 4328
rect 3576 4252 3592 4268
rect 3544 4232 3560 4248
rect 3624 4212 3640 4228
rect 3464 4092 3480 4108
rect 3224 3972 3240 3988
rect 3256 3972 3272 3988
rect 3272 3972 3288 3988
rect 3144 3932 3176 3948
rect 3208 3932 3224 3948
rect 3080 3912 3096 3928
rect 3128 3912 3144 3928
rect 3192 3912 3208 3928
rect 3048 3892 3064 3908
rect 3160 3892 3176 3908
rect 3128 3872 3144 3888
rect 3048 3792 3064 3808
rect 3016 3772 3032 3788
rect 3112 3772 3128 3788
rect 2824 3752 2840 3768
rect 2904 3732 2920 3748
rect 3032 3732 3048 3748
rect 2808 3712 2824 3728
rect 2840 3712 2856 3728
rect 2792 3592 2808 3608
rect 2861 3602 2897 3618
rect 2920 3592 2936 3608
rect 2952 3532 2968 3548
rect 2920 3512 2936 3528
rect 2808 3492 2824 3508
rect 2968 3492 2984 3508
rect 2936 3472 2952 3488
rect 3000 3652 3016 3668
rect 3064 3692 3080 3708
rect 3096 3692 3112 3708
rect 3208 3852 3224 3868
rect 3240 3952 3256 3968
rect 3224 3772 3240 3788
rect 3240 3772 3256 3788
rect 3208 3752 3224 3768
rect 3336 4032 3352 4048
rect 3672 4372 3688 4388
rect 3736 4632 3752 4648
rect 3832 4592 3848 4608
rect 3885 4602 3921 4618
rect 3736 4512 3752 4528
rect 3768 4492 3784 4508
rect 3752 4452 3784 4468
rect 3880 4572 3896 4588
rect 3864 4552 3880 4568
rect 3896 4532 3912 4548
rect 3816 4492 3832 4508
rect 3800 4392 3816 4408
rect 3800 4352 3816 4368
rect 3784 4332 3800 4348
rect 3720 4292 3736 4308
rect 3656 4252 3672 4268
rect 3496 4072 3512 4088
rect 3560 4072 3592 4088
rect 3480 4052 3496 4068
rect 3720 4152 3736 4168
rect 3496 4032 3512 4048
rect 3656 4032 3672 4048
rect 3464 3892 3480 3908
rect 3416 3872 3432 3888
rect 3304 3792 3320 3808
rect 3368 3792 3384 3808
rect 3288 3732 3304 3748
rect 3240 3672 3256 3688
rect 3272 3672 3288 3688
rect 3144 3632 3160 3648
rect 3096 3612 3112 3628
rect 3128 3612 3144 3628
rect 3144 3592 3160 3608
rect 3176 3552 3192 3568
rect 3240 3552 3256 3568
rect 3352 3552 3368 3568
rect 3016 3512 3032 3528
rect 3048 3512 3064 3528
rect 3080 3512 3096 3528
rect 3160 3512 3176 3528
rect 3016 3472 3032 3488
rect 3096 3472 3112 3488
rect 3064 3452 3080 3468
rect 2984 3432 3000 3448
rect 2968 3412 2984 3428
rect 2888 3392 2904 3408
rect 2856 3372 2872 3388
rect 2808 3352 2824 3368
rect 2792 3292 2808 3308
rect 2861 3202 2897 3218
rect 2840 3132 2856 3148
rect 2808 3092 2824 3108
rect 2792 2992 2808 3008
rect 2808 2952 2824 2968
rect 2776 2772 2792 2788
rect 2856 3012 2872 3028
rect 2920 3092 2936 3108
rect 3080 3412 3096 3428
rect 3128 3452 3144 3468
rect 3160 3432 3176 3448
rect 3032 3332 3048 3348
rect 3048 3312 3064 3328
rect 3016 3292 3032 3308
rect 3016 3132 3032 3148
rect 3000 3112 3016 3128
rect 3144 3332 3160 3348
rect 3128 3312 3144 3328
rect 3096 3292 3112 3308
rect 3096 3232 3112 3248
rect 3080 3152 3096 3168
rect 3064 3132 3080 3148
rect 2984 3092 3000 3108
rect 3048 3092 3064 3108
rect 3032 3072 3048 3088
rect 3064 3072 3080 3088
rect 2936 3032 2952 3048
rect 3000 3052 3016 3068
rect 3048 3052 3064 3068
rect 2952 3012 2968 3028
rect 2952 2992 2968 3008
rect 2904 2952 2920 2968
rect 2920 2872 2936 2888
rect 2861 2802 2897 2818
rect 2904 2812 2920 2828
rect 3080 3032 3096 3048
rect 3048 2992 3064 3008
rect 3128 3192 3144 3208
rect 3112 3112 3128 3128
rect 3144 3112 3160 3128
rect 3032 2972 3048 2988
rect 3096 2972 3112 2988
rect 2968 2892 2984 2908
rect 2984 2892 3000 2908
rect 3016 2892 3032 2908
rect 3080 2932 3096 2948
rect 3080 2892 3096 2908
rect 3064 2872 3080 2888
rect 2936 2852 2952 2868
rect 2952 2812 2968 2828
rect 2920 2752 2936 2768
rect 2824 2732 2840 2748
rect 3064 2792 3080 2808
rect 3096 2792 3112 2808
rect 2856 2712 2872 2728
rect 2760 2692 2776 2708
rect 2792 2692 2808 2708
rect 2680 2672 2696 2688
rect 2808 2672 2824 2688
rect 2616 2652 2632 2668
rect 2664 2652 2680 2668
rect 2776 2652 2808 2668
rect 2600 2632 2616 2648
rect 2680 2632 2696 2648
rect 2584 2612 2600 2628
rect 2520 2592 2536 2608
rect 2552 2592 2568 2608
rect 2760 2552 2776 2568
rect 2632 2532 2648 2548
rect 2520 2512 2536 2528
rect 2584 2512 2600 2528
rect 2488 2372 2504 2388
rect 2488 2272 2504 2288
rect 2456 2112 2472 2128
rect 2472 2072 2488 2088
rect 2440 1992 2456 2008
rect 2520 2472 2536 2488
rect 2552 2472 2568 2488
rect 2536 2412 2552 2428
rect 2536 2312 2552 2328
rect 2552 2272 2568 2288
rect 2824 2572 2840 2588
rect 3000 2672 3016 2688
rect 2904 2652 2920 2668
rect 2984 2652 3000 2668
rect 2952 2572 2968 2588
rect 2872 2552 2888 2568
rect 2904 2552 2920 2568
rect 2968 2552 2984 2568
rect 2792 2532 2808 2548
rect 2824 2532 2840 2548
rect 2680 2512 2696 2528
rect 2696 2512 2712 2528
rect 2616 2472 2632 2488
rect 2664 2472 2680 2488
rect 2632 2412 2648 2428
rect 2712 2452 2728 2468
rect 2696 2392 2712 2408
rect 3000 2512 3016 2528
rect 2904 2492 2920 2508
rect 2760 2472 2776 2488
rect 2792 2472 2824 2488
rect 2856 2472 2872 2488
rect 2808 2452 2824 2468
rect 2840 2452 2856 2468
rect 2776 2432 2792 2448
rect 2728 2372 2744 2388
rect 2824 2412 2840 2428
rect 2808 2352 2824 2368
rect 2664 2272 2680 2288
rect 2696 2272 2712 2288
rect 2600 2232 2616 2248
rect 2616 2132 2632 2148
rect 2744 2132 2760 2148
rect 2536 2112 2552 2128
rect 2536 2072 2552 2088
rect 2552 2052 2568 2068
rect 2328 1932 2344 1948
rect 2360 1932 2392 1948
rect 2424 1932 2440 1948
rect 2216 1872 2232 1888
rect 2200 1792 2216 1808
rect 2216 1732 2232 1748
rect 2312 1892 2328 1908
rect 2264 1832 2280 1848
rect 2312 1772 2328 1788
rect 2248 1752 2264 1768
rect 2312 1752 2328 1768
rect 2632 1932 2648 1948
rect 2616 1912 2632 1928
rect 2568 1892 2584 1908
rect 2600 1892 2616 1908
rect 2360 1852 2376 1868
rect 2344 1832 2360 1848
rect 2376 1832 2392 1848
rect 2408 1832 2424 1848
rect 2360 1772 2376 1788
rect 2184 1712 2200 1728
rect 2232 1712 2248 1728
rect 2264 1712 2280 1728
rect 2296 1712 2312 1728
rect 2328 1712 2344 1728
rect 2344 1652 2360 1668
rect 2280 1632 2296 1648
rect 2312 1632 2328 1648
rect 2104 1592 2120 1608
rect 2104 1572 2120 1588
rect 2280 1572 2296 1588
rect 2264 1552 2280 1568
rect 2248 1512 2264 1528
rect 2200 1492 2216 1508
rect 2344 1572 2360 1588
rect 2360 1532 2376 1548
rect 2520 1872 2536 1888
rect 2536 1832 2552 1848
rect 2440 1792 2456 1808
rect 2488 1792 2504 1808
rect 2456 1772 2472 1788
rect 2392 1712 2408 1728
rect 2312 1512 2328 1528
rect 2360 1512 2376 1528
rect 2216 1472 2232 1488
rect 2360 1472 2376 1488
rect 2312 1452 2328 1468
rect 2168 1412 2184 1428
rect 2104 1352 2120 1368
rect 2136 1312 2152 1328
rect 2152 1312 2168 1328
rect 2120 1252 2136 1268
rect 2104 1172 2120 1188
rect 1768 1106 1784 1108
rect 1768 1092 1784 1106
rect 1832 1092 1848 1108
rect 1864 1092 1880 1108
rect 1928 1092 1944 1108
rect 1960 1092 1976 1108
rect 2040 1092 2056 1108
rect 2088 1092 2104 1108
rect 1736 1072 1752 1088
rect 1896 1032 1912 1048
rect 1992 1032 2008 1048
rect 1688 1012 1704 1028
rect 1768 1012 1784 1028
rect 1837 1002 1873 1018
rect 2008 992 2024 1008
rect 1704 932 1720 948
rect 1768 932 1784 948
rect 1800 932 1816 948
rect 1880 932 1896 948
rect 1688 912 1704 928
rect 1400 852 1416 868
rect 1400 812 1416 828
rect 1384 792 1400 808
rect 1336 732 1352 748
rect 1064 672 1080 688
rect 1176 672 1192 688
rect 1320 672 1336 688
rect 1384 672 1400 688
rect 1032 652 1048 668
rect 1032 632 1048 648
rect 1048 572 1064 588
rect 808 492 824 508
rect 904 492 920 508
rect 936 492 952 508
rect 664 452 680 468
rect 872 452 888 468
rect 648 432 664 448
rect 632 412 648 428
rect 797 402 833 418
rect 664 372 680 388
rect 984 452 1000 468
rect 664 352 680 368
rect 936 352 952 368
rect 728 332 744 348
rect 680 312 696 328
rect 712 312 728 328
rect 712 252 728 268
rect 616 232 632 248
rect 376 112 392 128
rect 472 112 488 128
rect 504 132 520 148
rect 664 152 680 168
rect 744 312 760 328
rect 808 312 824 328
rect 856 312 872 328
rect 936 312 952 328
rect 968 312 984 328
rect 776 132 792 148
rect 872 252 888 268
rect 1000 292 1016 308
rect 920 232 936 248
rect 888 212 904 228
rect 904 172 920 188
rect 904 114 920 128
rect 904 112 920 114
rect 792 92 808 108
rect 696 72 712 88
rect 984 212 1000 228
rect 1048 392 1064 408
rect 1080 592 1096 608
rect 1112 612 1144 628
rect 1096 572 1128 588
rect 1144 552 1160 568
rect 1128 512 1144 528
rect 1240 592 1256 608
rect 1224 572 1240 588
rect 1208 552 1224 568
rect 1192 532 1208 548
rect 1080 452 1112 468
rect 1064 372 1080 388
rect 1048 312 1064 328
rect 1032 232 1048 248
rect 1032 212 1048 228
rect 984 172 1000 188
rect 1016 172 1032 188
rect 1000 152 1016 168
rect 1176 512 1192 528
rect 1304 592 1320 608
rect 1384 552 1400 568
rect 1256 532 1288 548
rect 1160 452 1176 468
rect 1256 452 1272 468
rect 1256 372 1272 388
rect 1240 352 1256 368
rect 1144 332 1160 348
rect 1176 332 1192 348
rect 1096 312 1112 328
rect 1160 312 1176 328
rect 1144 292 1160 308
rect 1064 192 1080 208
rect 1128 232 1144 248
rect 1096 192 1128 208
rect 1064 152 1080 168
rect 1080 152 1096 168
rect 1032 132 1048 148
rect 1192 312 1208 328
rect 1208 292 1224 308
rect 1336 512 1352 528
rect 1320 432 1336 448
rect 1304 392 1320 408
rect 1288 332 1304 348
rect 1288 292 1304 308
rect 1336 312 1352 328
rect 1272 272 1288 288
rect 1320 252 1336 268
rect 1416 572 1432 588
rect 1608 872 1640 888
rect 1448 852 1464 868
rect 1576 832 1592 848
rect 1448 812 1464 828
rect 1544 812 1560 828
rect 1480 692 1496 708
rect 1528 692 1544 708
rect 1608 752 1624 768
rect 1432 552 1448 568
rect 1464 552 1480 568
rect 1400 432 1416 448
rect 1384 352 1400 368
rect 1384 312 1400 328
rect 1288 232 1304 248
rect 1352 232 1368 248
rect 1176 152 1192 168
rect 1160 132 1176 148
rect 1192 132 1208 148
rect 1256 132 1272 148
rect 1272 132 1288 148
rect 968 112 984 128
rect 1016 112 1032 128
rect 1160 112 1176 128
rect 1256 112 1272 128
rect 1336 172 1352 188
rect 1384 152 1400 168
rect 1448 492 1464 508
rect 1736 912 1752 928
rect 1688 852 1704 868
rect 1848 892 1864 908
rect 1880 852 1896 868
rect 1688 812 1704 828
rect 1800 812 1816 828
rect 1720 732 1736 748
rect 1768 732 1800 748
rect 1848 732 1864 748
rect 1672 672 1688 688
rect 1752 672 1768 688
rect 1816 672 1832 688
rect 1736 652 1752 668
rect 1720 632 1736 648
rect 1800 612 1816 628
rect 1837 602 1873 618
rect 1608 572 1624 588
rect 1496 552 1512 568
rect 1800 552 1816 568
rect 1512 532 1528 548
rect 1688 532 1704 548
rect 1512 512 1528 528
rect 1480 432 1496 448
rect 1528 432 1544 448
rect 1496 372 1512 388
rect 1608 372 1624 388
rect 1464 312 1480 328
rect 1576 312 1592 328
rect 1704 312 1720 328
rect 1816 512 1832 528
rect 1928 752 1944 768
rect 2024 952 2040 968
rect 2024 732 2040 748
rect 2008 692 2024 708
rect 1960 672 1976 688
rect 1992 672 2008 688
rect 1944 632 1960 648
rect 1992 592 2008 608
rect 1928 552 1944 568
rect 1896 532 1912 548
rect 1960 532 1976 548
rect 1944 512 1960 528
rect 1976 512 1992 528
rect 2008 532 2024 548
rect 2056 532 2072 548
rect 1880 492 1896 508
rect 2008 492 2024 508
rect 1816 432 1832 448
rect 1976 352 1992 368
rect 2120 1012 2136 1028
rect 2184 1392 2200 1408
rect 2200 1352 2216 1368
rect 2296 1332 2312 1348
rect 2280 1312 2296 1328
rect 2232 1292 2248 1308
rect 2168 992 2184 1008
rect 2200 1152 2216 1168
rect 2280 1112 2296 1128
rect 2280 1092 2296 1108
rect 2216 1072 2248 1088
rect 2184 952 2200 968
rect 2104 932 2120 948
rect 2120 912 2136 928
rect 2088 892 2104 908
rect 2120 832 2136 848
rect 2104 712 2120 728
rect 2088 692 2104 708
rect 2184 912 2200 928
rect 2216 912 2232 928
rect 2168 892 2184 908
rect 2200 892 2216 908
rect 2152 812 2168 828
rect 2184 812 2200 828
rect 2136 692 2152 708
rect 2216 872 2232 888
rect 2248 1052 2264 1068
rect 2232 752 2248 768
rect 2216 732 2232 748
rect 2216 692 2232 708
rect 2152 672 2168 688
rect 2136 632 2152 648
rect 2168 632 2200 648
rect 2136 572 2152 588
rect 2104 552 2120 568
rect 2136 492 2152 508
rect 2216 592 2232 608
rect 2408 1472 2424 1488
rect 2520 1572 2536 1588
rect 2664 2114 2680 2128
rect 2664 2112 2680 2114
rect 2664 1892 2680 1908
rect 2680 1892 2696 1908
rect 2696 1872 2712 1888
rect 2728 1872 2744 1888
rect 2808 2132 2824 2148
rect 2792 2112 2808 2128
rect 2776 2092 2792 2108
rect 2776 2072 2792 2088
rect 2760 1952 2776 1968
rect 2760 1932 2776 1948
rect 2808 1932 2824 1948
rect 2744 1852 2760 1868
rect 2776 1832 2792 1848
rect 2600 1732 2616 1748
rect 2680 1732 2712 1748
rect 2616 1632 2632 1648
rect 2744 1812 2760 1828
rect 2744 1792 2760 1808
rect 2808 1792 2824 1808
rect 2861 2402 2897 2418
rect 2984 2472 3000 2488
rect 2952 2372 2968 2388
rect 2904 2312 2920 2328
rect 3080 2752 3096 2768
rect 3096 2732 3112 2748
rect 3176 3292 3192 3308
rect 3176 3132 3192 3148
rect 3192 3112 3208 3128
rect 3192 3072 3208 3088
rect 3224 3352 3240 3368
rect 3256 3532 3272 3548
rect 3352 3512 3368 3528
rect 3288 3492 3304 3508
rect 3448 3752 3464 3768
rect 3480 3752 3496 3768
rect 3464 3732 3480 3748
rect 3432 3652 3448 3668
rect 3384 3632 3400 3648
rect 3400 3532 3416 3548
rect 3336 3472 3352 3488
rect 3368 3472 3384 3488
rect 3304 3432 3320 3448
rect 3256 3412 3272 3428
rect 3288 3412 3304 3428
rect 3240 3312 3256 3328
rect 3368 3432 3384 3448
rect 3336 3372 3352 3388
rect 3304 3312 3336 3328
rect 3240 3292 3256 3308
rect 3272 3292 3288 3308
rect 3224 3272 3240 3288
rect 3224 3112 3240 3128
rect 3288 3172 3304 3188
rect 3288 3132 3304 3148
rect 3256 3112 3272 3128
rect 3240 3092 3256 3108
rect 3288 3092 3320 3108
rect 3208 3052 3224 3068
rect 3224 3032 3240 3048
rect 3192 2992 3208 3008
rect 3160 2912 3176 2928
rect 3256 2992 3272 3008
rect 3432 3492 3448 3508
rect 3416 3392 3432 3408
rect 3416 3352 3432 3368
rect 3368 3292 3384 3308
rect 3432 3272 3448 3288
rect 3464 3412 3480 3428
rect 3480 3392 3496 3408
rect 3464 3352 3480 3368
rect 3528 4012 3544 4028
rect 3528 3972 3544 3988
rect 3560 3892 3576 3908
rect 3672 3992 3688 4008
rect 3704 3992 3720 4008
rect 3720 3952 3736 3968
rect 3752 3972 3768 3988
rect 3736 3932 3752 3948
rect 3544 3872 3560 3888
rect 3624 3872 3640 3888
rect 3672 3872 3688 3888
rect 3512 3852 3528 3868
rect 3656 3852 3672 3868
rect 3624 3832 3640 3848
rect 3592 3792 3608 3808
rect 3576 3772 3592 3788
rect 3544 3752 3560 3768
rect 3512 3732 3528 3748
rect 3672 3752 3688 3768
rect 3704 3852 3720 3868
rect 3816 4332 3832 4348
rect 3816 4312 3848 4328
rect 3832 4292 3848 4308
rect 3816 4252 3832 4268
rect 3800 4212 3816 4228
rect 3784 4192 3800 4208
rect 3816 4132 3832 4148
rect 3800 4012 3816 4028
rect 3784 3912 3800 3928
rect 3768 3892 3784 3908
rect 3752 3832 3768 3848
rect 3704 3772 3720 3788
rect 3896 4512 3912 4528
rect 3928 4492 3944 4508
rect 4024 4692 4040 4708
rect 4120 4692 4136 4708
rect 4168 4692 4184 4708
rect 4104 4612 4120 4628
rect 3992 4572 4008 4588
rect 4024 4572 4040 4588
rect 4136 4672 4152 4688
rect 4104 4552 4120 4568
rect 4184 4652 4200 4668
rect 4248 4632 4264 4648
rect 4280 4612 4296 4628
rect 4312 4712 4328 4728
rect 4344 4692 4360 4708
rect 4312 4672 4328 4688
rect 4376 4712 4392 4728
rect 4328 4572 4344 4588
rect 4584 4706 4600 4708
rect 4584 4692 4600 4706
rect 4440 4672 4456 4688
rect 4696 4672 4712 4688
rect 4248 4552 4264 4568
rect 4296 4552 4312 4568
rect 4408 4552 4424 4568
rect 4136 4532 4152 4548
rect 4280 4532 4296 4548
rect 3976 4512 3992 4528
rect 4008 4472 4024 4488
rect 4024 4452 4040 4468
rect 4200 4512 4216 4528
rect 4072 4492 4088 4508
rect 3944 4432 3960 4448
rect 4024 4432 4040 4448
rect 4056 4432 4072 4448
rect 3896 4372 3912 4388
rect 3912 4312 3928 4328
rect 3960 4312 3976 4328
rect 3880 4292 3896 4308
rect 3864 4192 3880 4208
rect 3885 4202 3921 4218
rect 3976 4292 4008 4308
rect 3944 4232 3960 4248
rect 3944 4152 3960 4168
rect 3848 4012 3864 4028
rect 3896 4092 3912 4108
rect 3896 4072 3912 4088
rect 3848 3992 3880 4008
rect 3864 3972 3880 3988
rect 3848 3892 3864 3908
rect 3944 3892 3960 3908
rect 4072 4352 4088 4368
rect 4216 4492 4232 4508
rect 4264 4492 4280 4508
rect 4200 4472 4216 4488
rect 4168 4452 4184 4468
rect 4152 4372 4168 4388
rect 4088 4332 4104 4348
rect 4072 4312 4088 4328
rect 4008 4272 4024 4288
rect 4088 4272 4104 4288
rect 4008 4252 4024 4268
rect 4040 4232 4056 4248
rect 4024 4212 4040 4228
rect 4184 4232 4200 4248
rect 4120 4192 4136 4208
rect 4120 4172 4152 4188
rect 3992 4132 4008 4148
rect 4024 4132 4040 4148
rect 4072 4132 4088 4148
rect 4136 4132 4152 4148
rect 4024 4112 4040 4128
rect 4008 4092 4024 4108
rect 3976 4072 3992 4088
rect 3896 3852 3912 3868
rect 3885 3802 3921 3818
rect 3976 3852 3992 3868
rect 3960 3812 3976 3828
rect 3928 3772 3944 3788
rect 3864 3732 3880 3748
rect 4040 4092 4056 4108
rect 4072 4072 4088 4088
rect 4040 3912 4056 3928
rect 4024 3892 4040 3908
rect 3992 3832 4008 3848
rect 4168 4092 4184 4108
rect 4104 4052 4120 4068
rect 4152 3992 4168 4008
rect 4104 3972 4120 3988
rect 4056 3852 4072 3868
rect 4088 3852 4104 3868
rect 4056 3832 4072 3848
rect 4072 3752 4088 3768
rect 3688 3672 3704 3688
rect 3624 3612 3640 3628
rect 3528 3492 3544 3508
rect 3576 3492 3592 3508
rect 3592 3472 3608 3488
rect 3752 3612 3768 3628
rect 4152 3892 4168 3908
rect 4136 3852 4152 3868
rect 4152 3772 4168 3788
rect 4120 3732 4136 3748
rect 4232 4452 4248 4468
rect 4232 4432 4248 4448
rect 4216 4352 4232 4368
rect 4392 4532 4408 4548
rect 4232 4292 4248 4308
rect 4312 4312 4328 4328
rect 4232 4232 4248 4248
rect 4280 4232 4296 4248
rect 4216 4212 4232 4228
rect 4264 4092 4280 4108
rect 4232 4032 4248 4048
rect 4216 3952 4232 3968
rect 4248 3852 4264 3868
rect 4216 3792 4232 3808
rect 4040 3712 4056 3728
rect 4120 3692 4136 3708
rect 3992 3672 4008 3688
rect 4024 3672 4040 3688
rect 4056 3672 4072 3688
rect 4088 3672 4104 3688
rect 3976 3592 3992 3608
rect 3736 3552 3752 3568
rect 3688 3532 3704 3548
rect 3752 3532 3768 3548
rect 3656 3452 3672 3468
rect 4040 3552 4056 3568
rect 3800 3532 3816 3548
rect 3832 3532 3848 3548
rect 3960 3512 3976 3528
rect 3992 3512 4008 3528
rect 3768 3492 3784 3508
rect 3720 3472 3736 3488
rect 3720 3452 3736 3468
rect 3704 3432 3720 3448
rect 3640 3352 3656 3368
rect 3672 3352 3704 3368
rect 3560 3312 3576 3328
rect 3592 3312 3608 3328
rect 3448 3252 3464 3268
rect 3512 3212 3528 3228
rect 3544 3272 3560 3288
rect 3544 3232 3560 3248
rect 3400 3192 3416 3208
rect 3528 3192 3544 3208
rect 3608 3292 3624 3308
rect 3560 3172 3576 3188
rect 3368 3152 3384 3168
rect 3352 3112 3368 3128
rect 3352 3092 3368 3108
rect 3512 3132 3528 3148
rect 3416 3112 3432 3128
rect 3384 3092 3400 3108
rect 3432 3032 3448 3048
rect 3336 3012 3352 3028
rect 3400 3012 3416 3028
rect 3320 2992 3336 3008
rect 3352 2972 3368 2988
rect 3448 3012 3464 3028
rect 3464 2972 3480 2988
rect 3208 2932 3224 2948
rect 3384 2932 3400 2948
rect 3144 2892 3160 2908
rect 3176 2892 3192 2908
rect 3128 2872 3144 2888
rect 3128 2852 3144 2868
rect 3096 2672 3112 2688
rect 3048 2612 3064 2628
rect 3048 2572 3064 2588
rect 3144 2792 3160 2808
rect 3160 2752 3176 2768
rect 3144 2732 3160 2748
rect 3160 2672 3176 2688
rect 3160 2632 3176 2648
rect 3112 2552 3128 2568
rect 3144 2552 3160 2568
rect 3096 2492 3112 2508
rect 3112 2472 3128 2488
rect 3032 2452 3048 2468
rect 3080 2452 3096 2468
rect 3032 2412 3048 2428
rect 3080 2372 3096 2388
rect 3032 2312 3048 2328
rect 2840 2292 2856 2308
rect 2888 2292 2904 2308
rect 2856 2252 2872 2268
rect 2840 2112 2856 2128
rect 2904 2072 2920 2088
rect 2888 2052 2904 2068
rect 2861 2002 2897 2018
rect 2952 2292 2968 2308
rect 3016 2292 3032 2308
rect 2936 2152 2952 2168
rect 3160 2492 3176 2508
rect 3176 2372 3192 2388
rect 3144 2332 3160 2348
rect 3176 2332 3192 2348
rect 3208 2892 3224 2908
rect 3240 2892 3256 2908
rect 3224 2872 3240 2888
rect 3208 2812 3224 2828
rect 3272 2892 3288 2908
rect 3320 2852 3336 2868
rect 3368 2852 3384 2868
rect 3272 2812 3288 2828
rect 3304 2772 3320 2788
rect 3400 2752 3416 2768
rect 3448 2912 3464 2928
rect 3432 2892 3448 2908
rect 3432 2772 3448 2788
rect 3528 3072 3544 3088
rect 3528 3032 3544 3048
rect 3496 3012 3512 3028
rect 3592 3112 3608 3128
rect 3704 3332 3720 3348
rect 3656 3292 3672 3308
rect 3672 3292 3688 3308
rect 3688 3252 3704 3268
rect 3816 3472 3832 3488
rect 3848 3452 3864 3468
rect 3832 3392 3848 3408
rect 3784 3372 3800 3388
rect 3784 3332 3800 3348
rect 3816 3312 3832 3328
rect 3736 3292 3752 3308
rect 3912 3432 3928 3448
rect 3885 3402 3921 3418
rect 3944 3352 3976 3368
rect 3944 3312 3960 3328
rect 3992 3312 4008 3328
rect 3864 3292 3880 3308
rect 3896 3272 3912 3288
rect 3928 3232 3944 3248
rect 3800 3192 3816 3208
rect 3928 3172 3944 3188
rect 3896 3112 3912 3128
rect 3624 3072 3640 3088
rect 3672 3072 3688 3088
rect 3608 3052 3624 3068
rect 3624 3012 3640 3028
rect 3528 2992 3544 3008
rect 3560 2992 3576 3008
rect 3496 2912 3512 2928
rect 3480 2732 3496 2748
rect 3288 2692 3304 2708
rect 3368 2692 3384 2708
rect 3400 2692 3416 2708
rect 3480 2706 3496 2708
rect 3480 2692 3496 2706
rect 3352 2672 3368 2688
rect 3384 2672 3400 2688
rect 3256 2652 3272 2668
rect 3496 2652 3512 2668
rect 3208 2612 3224 2628
rect 3240 2592 3256 2608
rect 3208 2572 3224 2588
rect 3208 2452 3240 2468
rect 3560 2952 3576 2968
rect 3656 2932 3672 2948
rect 3592 2812 3608 2828
rect 3656 2812 3672 2828
rect 3592 2792 3608 2808
rect 3576 2712 3592 2728
rect 3544 2692 3560 2708
rect 3528 2612 3544 2628
rect 3576 2612 3592 2628
rect 3448 2572 3464 2588
rect 3528 2572 3544 2588
rect 3480 2552 3496 2568
rect 3544 2552 3560 2568
rect 3272 2532 3288 2548
rect 3320 2532 3336 2548
rect 3400 2532 3416 2548
rect 3512 2532 3528 2548
rect 3256 2392 3272 2408
rect 3208 2352 3224 2368
rect 3256 2352 3272 2368
rect 3144 2312 3176 2328
rect 3192 2312 3208 2328
rect 3048 2272 3064 2288
rect 3112 2272 3128 2288
rect 3128 2212 3144 2228
rect 3112 2172 3128 2188
rect 2936 2132 2952 2148
rect 3080 2112 3096 2128
rect 3144 2112 3160 2128
rect 2952 2092 2968 2108
rect 2984 2092 3000 2108
rect 3224 2332 3240 2348
rect 3240 2312 3256 2328
rect 3192 2292 3208 2308
rect 3320 2492 3336 2508
rect 3288 2472 3304 2488
rect 3320 2392 3336 2408
rect 3304 2312 3320 2328
rect 3272 2292 3288 2308
rect 3192 2232 3208 2248
rect 3160 2092 3176 2108
rect 3000 2072 3016 2088
rect 3080 2072 3096 2088
rect 3144 2072 3160 2088
rect 2952 2052 2968 2068
rect 3016 2052 3032 2068
rect 2936 2012 2952 2028
rect 2840 1932 2856 1948
rect 2904 1932 2920 1948
rect 2920 1932 2936 1948
rect 2840 1872 2856 1888
rect 2856 1852 2872 1868
rect 2792 1752 2808 1768
rect 2824 1752 2840 1768
rect 2776 1732 2808 1748
rect 2920 1852 2936 1868
rect 2888 1772 2904 1788
rect 2760 1712 2776 1728
rect 2696 1632 2712 1648
rect 2696 1612 2712 1628
rect 2552 1552 2568 1568
rect 2648 1552 2680 1568
rect 2520 1532 2536 1548
rect 2488 1512 2504 1528
rect 2840 1692 2856 1708
rect 2856 1692 2872 1708
rect 2856 1672 2872 1688
rect 2872 1632 2888 1648
rect 2861 1602 2897 1618
rect 2776 1552 2792 1568
rect 2856 1552 2872 1568
rect 2904 1552 2920 1568
rect 2760 1532 2776 1548
rect 2616 1512 2632 1528
rect 2696 1512 2712 1528
rect 2424 1452 2440 1468
rect 2472 1452 2488 1468
rect 2408 1432 2440 1448
rect 2344 1352 2360 1368
rect 2376 1372 2392 1388
rect 2344 1312 2360 1328
rect 2440 1312 2456 1328
rect 2344 1292 2360 1308
rect 2472 1252 2488 1268
rect 2328 1132 2344 1148
rect 2360 1112 2376 1128
rect 2456 1112 2472 1128
rect 2456 1092 2472 1108
rect 2392 1072 2408 1088
rect 2328 972 2344 988
rect 2264 932 2280 948
rect 2312 772 2328 788
rect 2440 1052 2456 1068
rect 2520 1372 2536 1388
rect 2504 1312 2520 1328
rect 2488 1212 2504 1228
rect 2632 1472 2648 1488
rect 2680 1472 2696 1488
rect 2728 1432 2744 1448
rect 2584 1412 2600 1428
rect 2584 1392 2600 1408
rect 2600 1352 2616 1368
rect 2984 2012 3000 2028
rect 2952 1852 2968 1868
rect 2936 1812 2952 1828
rect 2936 1752 2952 1768
rect 3384 2512 3400 2528
rect 3608 2772 3624 2788
rect 3688 2752 3704 2768
rect 3624 2732 3640 2748
rect 3640 2712 3644 2728
rect 3644 2712 3656 2728
rect 3672 2672 3688 2688
rect 3704 2672 3720 2688
rect 3368 2492 3384 2508
rect 3416 2492 3432 2508
rect 3496 2492 3512 2508
rect 3352 2472 3368 2488
rect 3400 2472 3416 2488
rect 3464 2472 3480 2488
rect 3432 2452 3448 2468
rect 3464 2452 3480 2468
rect 3528 2352 3544 2368
rect 3352 2312 3368 2328
rect 3368 2312 3384 2328
rect 3624 2512 3640 2528
rect 3624 2492 3640 2508
rect 3640 2472 3656 2488
rect 3784 3072 3800 3088
rect 3752 3052 3768 3068
rect 3800 3032 3816 3048
rect 3960 3152 3976 3168
rect 4008 3252 4024 3268
rect 4056 3112 4072 3128
rect 3976 3072 3992 3088
rect 4024 3072 4040 3088
rect 3885 3002 3921 3018
rect 3944 3012 3960 3028
rect 3736 2832 3752 2848
rect 3816 2912 3832 2928
rect 3944 2912 3960 2928
rect 3864 2872 3880 2888
rect 3832 2812 3848 2828
rect 3736 2652 3752 2668
rect 3720 2612 3736 2628
rect 3784 2692 3800 2708
rect 3816 2692 3832 2708
rect 3880 2732 3896 2748
rect 3928 2672 3944 2688
rect 3832 2632 3848 2648
rect 3864 2632 3880 2648
rect 3885 2602 3921 2618
rect 3768 2552 3784 2568
rect 3832 2552 3848 2568
rect 3896 2552 3912 2568
rect 3720 2512 3736 2528
rect 3688 2492 3704 2508
rect 3768 2492 3784 2508
rect 3736 2472 3752 2488
rect 3656 2452 3688 2468
rect 3656 2412 3672 2428
rect 3624 2392 3640 2408
rect 3608 2372 3624 2388
rect 3592 2312 3608 2328
rect 3624 2312 3640 2328
rect 3400 2292 3416 2308
rect 3640 2292 3656 2308
rect 3336 2252 3352 2268
rect 3304 2212 3320 2228
rect 3208 2172 3224 2188
rect 3240 2172 3256 2188
rect 3256 2152 3272 2168
rect 3208 2112 3224 2128
rect 3176 2072 3192 2088
rect 3336 2152 3352 2168
rect 3496 2272 3512 2288
rect 3416 2252 3432 2268
rect 3288 2112 3304 2128
rect 3336 2132 3352 2148
rect 3352 2112 3368 2128
rect 3336 2092 3352 2108
rect 3272 2072 3288 2088
rect 3224 2052 3240 2068
rect 3256 2052 3272 2068
rect 3096 1972 3112 1988
rect 3064 1932 3080 1948
rect 3032 1912 3048 1928
rect 3176 1952 3192 1968
rect 3208 1952 3224 1968
rect 3128 1892 3144 1908
rect 3000 1872 3016 1888
rect 3064 1872 3080 1888
rect 3000 1752 3016 1768
rect 3048 1752 3064 1768
rect 3016 1732 3032 1748
rect 2984 1712 3000 1728
rect 2968 1532 2984 1548
rect 2936 1392 2952 1408
rect 3240 1932 3256 1948
rect 3288 2032 3304 2048
rect 3320 1972 3336 1988
rect 3320 1952 3336 1968
rect 3288 1912 3304 1928
rect 3384 2112 3400 2128
rect 3448 2212 3464 2228
rect 3464 2112 3480 2128
rect 3400 2072 3416 2088
rect 3400 2032 3416 2048
rect 3368 1952 3384 1968
rect 3336 1932 3352 1948
rect 3112 1872 3128 1888
rect 3240 1872 3256 1888
rect 3192 1852 3208 1868
rect 3192 1832 3208 1848
rect 3128 1812 3144 1828
rect 3080 1792 3112 1808
rect 3112 1752 3128 1768
rect 3272 1792 3288 1808
rect 3256 1772 3272 1788
rect 3208 1712 3224 1728
rect 3112 1632 3128 1648
rect 3080 1492 3096 1508
rect 3112 1472 3128 1488
rect 3016 1392 3032 1408
rect 2984 1372 3000 1388
rect 3064 1372 3080 1388
rect 2808 1332 2824 1348
rect 2920 1332 2936 1348
rect 3096 1332 3112 1348
rect 2536 1192 2552 1208
rect 2504 1172 2520 1188
rect 2504 1092 2520 1108
rect 2536 1072 2552 1088
rect 2568 1072 2584 1088
rect 2584 1032 2600 1048
rect 2488 1012 2504 1028
rect 2344 952 2360 968
rect 2408 952 2440 968
rect 2472 952 2488 968
rect 2376 892 2392 908
rect 2344 872 2360 888
rect 2360 852 2376 868
rect 2360 832 2376 848
rect 2408 832 2424 848
rect 2248 692 2264 708
rect 2280 692 2296 708
rect 2296 692 2312 708
rect 2248 652 2264 668
rect 2248 552 2264 568
rect 2264 532 2280 548
rect 2184 512 2200 528
rect 2168 472 2184 488
rect 2152 452 2168 468
rect 2184 412 2200 428
rect 2072 352 2088 368
rect 2104 332 2120 348
rect 1464 292 1480 308
rect 1624 292 1640 308
rect 1800 292 1816 308
rect 2024 292 2040 308
rect 2120 292 2136 308
rect 1672 272 1688 288
rect 2088 276 2104 288
rect 2088 272 2104 276
rect 1656 212 1672 228
rect 1640 192 1656 208
rect 1528 152 1544 168
rect 1320 132 1336 148
rect 1384 132 1400 148
rect 1416 132 1432 148
rect 2312 672 2328 688
rect 2328 652 2344 668
rect 2344 592 2360 608
rect 2744 1312 2760 1328
rect 2792 1312 2808 1328
rect 2840 1312 2856 1328
rect 2712 1292 2728 1308
rect 2824 1292 2840 1308
rect 2760 1252 2776 1268
rect 2872 1252 2888 1268
rect 2936 1232 2952 1248
rect 2861 1202 2897 1218
rect 3000 1312 3016 1328
rect 3064 1312 3080 1328
rect 3048 1252 3064 1268
rect 3000 1232 3016 1248
rect 3016 1212 3032 1228
rect 2984 1192 3000 1208
rect 3016 1192 3032 1208
rect 2824 1152 2840 1168
rect 2968 1152 2984 1168
rect 2632 1132 2648 1148
rect 2664 1112 2680 1128
rect 2712 1112 2728 1128
rect 2760 1112 2776 1128
rect 2664 1092 2680 1108
rect 2744 1092 2760 1108
rect 2776 1092 2792 1108
rect 2552 952 2568 968
rect 2472 892 2488 908
rect 2488 852 2504 868
rect 2616 852 2632 868
rect 2520 812 2536 828
rect 2536 752 2552 768
rect 2520 732 2536 748
rect 2376 692 2392 708
rect 2424 692 2440 708
rect 2456 692 2472 708
rect 2408 672 2424 688
rect 2392 632 2408 648
rect 2312 572 2328 588
rect 2296 552 2312 568
rect 2424 592 2440 608
rect 2472 592 2488 608
rect 2504 592 2520 608
rect 2344 532 2360 548
rect 2408 532 2424 548
rect 2392 512 2408 528
rect 2248 492 2264 508
rect 2248 452 2264 468
rect 2360 452 2376 468
rect 2248 412 2264 428
rect 2232 392 2248 408
rect 2232 372 2248 388
rect 2344 352 2360 368
rect 2472 572 2488 588
rect 2456 512 2472 528
rect 2504 552 2520 568
rect 2488 532 2504 548
rect 2472 452 2488 468
rect 2456 352 2472 368
rect 2408 332 2424 348
rect 2456 332 2472 348
rect 2216 312 2232 328
rect 2248 312 2264 328
rect 2280 312 2292 328
rect 2292 312 2296 328
rect 2344 312 2360 328
rect 2376 312 2380 328
rect 2380 312 2392 328
rect 2440 312 2452 328
rect 2452 312 2456 328
rect 2184 292 2200 308
rect 2264 292 2280 308
rect 1688 252 1704 268
rect 1928 252 1944 268
rect 2024 252 2040 268
rect 2152 252 2168 268
rect 1816 232 1832 248
rect 1992 232 2008 248
rect 1688 212 1704 228
rect 1704 192 1720 208
rect 1837 202 1873 218
rect 1944 192 1960 208
rect 1752 172 1768 188
rect 1720 152 1736 168
rect 1800 152 1816 168
rect 1944 152 1960 168
rect 2120 152 2136 168
rect 2216 252 2232 268
rect 2280 232 2296 248
rect 2264 192 2280 208
rect 1992 132 2008 148
rect 2168 132 2184 148
rect 1416 112 1432 128
rect 1448 112 1464 128
rect 1512 114 1528 128
rect 1512 112 1528 114
rect 1848 112 1864 128
rect 1112 92 1128 108
rect 1224 92 1240 108
rect 1272 92 1288 108
rect 1304 92 1320 108
rect 1352 92 1368 108
rect 984 72 1000 88
rect 2392 292 2408 308
rect 2424 292 2440 308
rect 2504 412 2520 428
rect 2504 392 2520 408
rect 2488 332 2504 348
rect 3048 1192 3064 1208
rect 3080 1132 3096 1148
rect 2984 1112 3000 1128
rect 3032 1112 3048 1128
rect 2856 1092 2872 1108
rect 2840 1072 2856 1088
rect 2776 1052 2792 1068
rect 2808 992 2824 1008
rect 2680 952 2696 968
rect 2712 952 2728 968
rect 2760 912 2776 928
rect 2792 852 2808 868
rect 2936 1092 2952 1108
rect 3064 1092 3080 1108
rect 2872 1052 2888 1068
rect 2872 932 2888 948
rect 2872 912 2888 928
rect 2824 872 2840 888
rect 2808 832 2824 848
rect 2712 792 2728 808
rect 2760 792 2776 808
rect 2744 732 2760 748
rect 2584 712 2616 728
rect 2632 712 2648 728
rect 2712 712 2728 728
rect 2616 672 2632 688
rect 2680 652 2696 668
rect 2632 632 2648 648
rect 2568 572 2584 588
rect 2616 572 2632 588
rect 2600 512 2616 528
rect 2648 512 2664 528
rect 2744 612 2760 628
rect 2728 572 2744 588
rect 2616 492 2632 508
rect 2664 492 2680 508
rect 2680 492 2696 508
rect 2584 472 2600 488
rect 2616 472 2632 488
rect 2552 432 2568 448
rect 2552 392 2568 408
rect 2536 372 2552 388
rect 2584 372 2600 388
rect 2488 272 2504 288
rect 2344 252 2376 268
rect 2296 212 2312 228
rect 2424 192 2440 208
rect 2408 172 2424 188
rect 2392 152 2408 168
rect 2456 152 2472 168
rect 2312 132 2328 148
rect 2328 132 2344 148
rect 2376 132 2392 148
rect 2440 132 2456 148
rect 2520 232 2536 248
rect 2520 132 2536 148
rect 2568 312 2584 328
rect 2664 412 2680 428
rect 2840 792 2856 808
rect 2861 802 2897 818
rect 2824 772 2840 788
rect 2888 692 2904 708
rect 3048 1072 3064 1088
rect 2920 1032 2936 1048
rect 2968 1052 2984 1068
rect 3048 1052 3064 1068
rect 3000 1032 3016 1048
rect 3032 1032 3048 1048
rect 2936 992 2952 1008
rect 3000 992 3016 1008
rect 2920 952 2936 968
rect 3016 952 3032 968
rect 3112 1192 3128 1208
rect 3208 1692 3224 1708
rect 3144 1672 3176 1688
rect 3160 1592 3192 1608
rect 3160 1572 3176 1588
rect 3368 1832 3384 1848
rect 3448 2092 3464 2108
rect 3640 2232 3656 2248
rect 3592 2192 3608 2208
rect 3512 2172 3528 2188
rect 3576 2172 3592 2188
rect 3720 2392 3736 2408
rect 3816 2392 3832 2408
rect 3544 2112 3560 2128
rect 3592 2112 3608 2128
rect 3512 2092 3528 2108
rect 3560 2092 3576 2108
rect 3624 2092 3640 2108
rect 3752 2352 3768 2368
rect 3768 2332 3784 2348
rect 3800 2332 3816 2348
rect 3704 2212 3720 2228
rect 3688 2192 3704 2208
rect 3912 2532 3928 2548
rect 4184 3672 4200 3688
rect 4216 3652 4232 3668
rect 4152 3592 4168 3608
rect 4280 4012 4296 4028
rect 4312 4072 4328 4088
rect 4376 4492 4392 4508
rect 4424 4492 4436 4508
rect 4436 4492 4440 4508
rect 4392 4432 4408 4448
rect 4344 4412 4360 4428
rect 4392 4412 4408 4428
rect 4616 4652 4632 4668
rect 4568 4632 4584 4648
rect 4648 4632 4664 4648
rect 4552 4612 4568 4628
rect 4456 4592 4472 4608
rect 4456 4552 4472 4568
rect 4488 4532 4504 4548
rect 4536 4532 4552 4548
rect 4456 4492 4472 4508
rect 4488 4432 4504 4448
rect 4536 4492 4552 4508
rect 4520 4392 4536 4408
rect 4440 4352 4456 4368
rect 4424 4332 4456 4348
rect 4392 4312 4408 4328
rect 4360 4212 4376 4228
rect 4376 4132 4392 4148
rect 4536 4312 4552 4328
rect 4456 4292 4472 4308
rect 4424 4192 4440 4208
rect 4408 4132 4424 4148
rect 4456 4112 4472 4128
rect 4424 4092 4440 4108
rect 4376 4072 4408 4088
rect 4344 4052 4360 4068
rect 4584 4572 4600 4588
rect 4616 4532 4632 4548
rect 4616 4512 4632 4528
rect 4696 4592 4712 4608
rect 4680 4552 4696 4568
rect 4712 4552 4728 4568
rect 4712 4512 4728 4528
rect 4632 4432 4648 4448
rect 4664 4432 4680 4448
rect 4616 4352 4632 4368
rect 4664 4352 4680 4368
rect 4600 4312 4616 4328
rect 4632 4312 4648 4328
rect 4568 4272 4584 4288
rect 4504 4212 4520 4228
rect 4520 4192 4536 4208
rect 4536 4172 4552 4188
rect 4744 4572 4760 4588
rect 4744 4552 4760 4568
rect 4728 4492 4744 4508
rect 4696 4332 4712 4348
rect 4696 4312 4712 4328
rect 4744 4232 4760 4248
rect 4584 4212 4600 4228
rect 4680 4212 4696 4228
rect 4584 4152 4600 4168
rect 4552 4132 4568 4148
rect 4744 4132 4760 4148
rect 4520 4112 4536 4128
rect 4632 4112 4648 4128
rect 4472 4092 4488 4108
rect 4488 4092 4504 4108
rect 4328 4032 4344 4048
rect 4440 4032 4456 4048
rect 4312 3992 4328 4008
rect 4392 3992 4408 4008
rect 4296 3972 4312 3988
rect 4296 3952 4312 3968
rect 4568 4072 4584 4088
rect 4600 4052 4616 4068
rect 4632 4052 4648 4068
rect 4648 4032 4664 4048
rect 4520 3952 4536 3968
rect 4312 3912 4328 3928
rect 4376 3912 4392 3928
rect 4472 3912 4488 3928
rect 4504 3912 4520 3928
rect 4360 3892 4376 3908
rect 4456 3892 4472 3908
rect 4312 3812 4328 3828
rect 4424 3852 4440 3868
rect 4632 3932 4648 3948
rect 4584 3912 4600 3928
rect 4520 3852 4552 3868
rect 4568 3852 4584 3868
rect 4504 3832 4520 3848
rect 4344 3792 4360 3808
rect 4440 3792 4456 3808
rect 4648 3852 4664 3868
rect 4616 3832 4632 3848
rect 4648 3832 4664 3848
rect 4504 3772 4520 3788
rect 4632 3812 4648 3828
rect 4680 3812 4696 3828
rect 4728 3832 4744 3848
rect 4712 3812 4728 3828
rect 4440 3714 4456 3728
rect 4440 3712 4456 3714
rect 4328 3692 4344 3708
rect 4296 3652 4312 3668
rect 4264 3612 4280 3628
rect 4248 3592 4264 3608
rect 4216 3532 4232 3548
rect 4168 3472 4184 3488
rect 4120 3392 4136 3408
rect 4184 3452 4200 3468
rect 4168 3352 4184 3368
rect 4184 3332 4200 3348
rect 4104 3312 4120 3328
rect 4200 3312 4216 3328
rect 4088 3172 4104 3188
rect 4280 3532 4296 3548
rect 4536 3612 4552 3628
rect 4360 3512 4376 3528
rect 4392 3512 4408 3528
rect 4312 3452 4328 3468
rect 4264 3432 4280 3448
rect 4280 3392 4296 3408
rect 4248 3352 4264 3368
rect 4232 3312 4248 3328
rect 4408 3492 4424 3508
rect 4616 3732 4632 3748
rect 4664 3732 4680 3748
rect 4696 3732 4712 3748
rect 4728 3732 4744 3748
rect 4792 4692 4808 4708
rect 4840 4672 4856 4688
rect 4808 4632 4824 4648
rect 4872 4632 4888 4648
rect 4776 4612 4792 4628
rect 4856 4592 4872 4608
rect 4776 4572 4792 4588
rect 4808 4572 4824 4588
rect 4888 4592 4904 4608
rect 4888 4572 4904 4588
rect 4952 4712 4968 4728
rect 5336 4712 5352 4728
rect 4936 4692 4952 4708
rect 4968 4692 4984 4708
rect 5064 4692 5080 4708
rect 5144 4672 5160 4688
rect 5208 4672 5224 4688
rect 5304 4672 5320 4688
rect 5048 4652 5064 4668
rect 5064 4612 5080 4628
rect 5176 4612 5192 4628
rect 5240 4612 5256 4628
rect 4792 4492 4808 4508
rect 4808 4452 4824 4468
rect 4776 4432 4792 4448
rect 4856 4452 4872 4468
rect 4776 4412 4792 4428
rect 4824 4412 4840 4428
rect 4840 4392 4856 4408
rect 4968 4552 4984 4568
rect 4984 4532 5000 4548
rect 5144 4532 5160 4548
rect 4904 4512 4920 4528
rect 4968 4512 4984 4528
rect 5000 4512 5016 4528
rect 5112 4512 5128 4528
rect 5160 4512 5176 4528
rect 5032 4472 5048 4488
rect 5016 4432 5032 4448
rect 4909 4402 4945 4418
rect 4952 4312 4968 4328
rect 5032 4312 5048 4328
rect 4824 4272 4840 4288
rect 4840 4272 4856 4288
rect 4872 4272 4888 4288
rect 4840 4212 4856 4228
rect 4776 4192 4792 4208
rect 4840 4172 4856 4188
rect 4856 4132 4872 4148
rect 4808 4092 4824 4108
rect 4872 4072 4888 4088
rect 4840 4052 4856 4068
rect 4856 3992 4872 4008
rect 4776 3952 4792 3968
rect 4792 3912 4808 3928
rect 4840 3912 4856 3928
rect 4920 4172 4936 4188
rect 4936 4152 4952 4168
rect 4909 4002 4945 4018
rect 4888 3932 4904 3948
rect 4920 3932 4936 3948
rect 4936 3932 4952 3948
rect 4872 3872 4888 3888
rect 4904 3852 4920 3868
rect 4840 3832 4856 3848
rect 4760 3772 4776 3788
rect 4872 3772 4888 3788
rect 4872 3752 4904 3768
rect 4584 3712 4616 3728
rect 4648 3712 4664 3728
rect 4696 3712 4712 3728
rect 4744 3712 4760 3728
rect 4696 3692 4712 3708
rect 4648 3612 4664 3628
rect 4808 3672 4824 3688
rect 4840 3672 4856 3688
rect 4808 3532 4824 3548
rect 4760 3512 4776 3528
rect 4552 3492 4568 3508
rect 4584 3492 4600 3508
rect 4664 3492 4680 3508
rect 4728 3492 4744 3508
rect 4792 3492 4808 3508
rect 4840 3492 4856 3508
rect 4520 3432 4536 3448
rect 4936 3912 4952 3928
rect 4952 3892 4968 3908
rect 5080 4452 5096 4468
rect 5080 4392 5096 4408
rect 5096 4352 5112 4368
rect 5144 4492 5160 4508
rect 5160 4392 5176 4408
rect 5128 4332 5144 4348
rect 5096 4312 5112 4328
rect 4984 4272 5016 4288
rect 5048 4292 5064 4308
rect 5096 4292 5112 4308
rect 5064 4192 5080 4208
rect 5032 4172 5048 4188
rect 5016 4152 5032 4168
rect 5144 4192 5160 4208
rect 5064 4132 5080 4148
rect 5000 4112 5016 4128
rect 5016 4112 5032 4128
rect 5128 4112 5144 4128
rect 4984 4092 4988 4108
rect 4988 4092 5000 4108
rect 5096 4092 5112 4108
rect 5064 4072 5080 4088
rect 5080 4052 5096 4068
rect 5016 4032 5032 4048
rect 4984 3932 5000 3948
rect 4968 3752 4984 3768
rect 5112 3952 5128 3968
rect 5128 3932 5144 3948
rect 5032 3912 5048 3928
rect 5112 3912 5128 3928
rect 5000 3712 5016 3728
rect 4888 3692 4904 3708
rect 4872 3492 4888 3508
rect 4632 3472 4648 3488
rect 4760 3472 4792 3488
rect 4856 3472 4872 3488
rect 4584 3412 4600 3428
rect 4328 3352 4344 3368
rect 4520 3352 4536 3368
rect 4264 3332 4280 3348
rect 4216 3292 4248 3308
rect 4296 3312 4312 3328
rect 4280 3232 4296 3248
rect 4360 3312 4376 3328
rect 4392 3312 4408 3328
rect 4424 3312 4440 3328
rect 4488 3312 4504 3328
rect 4504 3312 4520 3328
rect 4536 3312 4552 3328
rect 4392 3292 4424 3308
rect 4456 3292 4472 3308
rect 4552 3292 4568 3308
rect 4344 3252 4360 3268
rect 4328 3192 4344 3208
rect 4376 3172 4392 3188
rect 4216 3112 4232 3128
rect 4120 3072 4136 3088
rect 4168 3072 4184 3088
rect 4168 2992 4184 3008
rect 4072 2972 4088 2988
rect 4104 2972 4136 2988
rect 4088 2952 4104 2968
rect 4072 2892 4088 2908
rect 4120 2892 4136 2908
rect 4168 2892 4184 2908
rect 4168 2812 4184 2828
rect 4072 2772 4088 2788
rect 3976 2672 3992 2688
rect 4024 2712 4040 2728
rect 4120 2752 4136 2768
rect 4136 2712 4152 2728
rect 4136 2692 4152 2708
rect 4056 2672 4072 2688
rect 4088 2672 4120 2688
rect 4008 2632 4024 2648
rect 4040 2592 4056 2608
rect 4040 2572 4056 2588
rect 3976 2552 3992 2568
rect 3960 2532 3976 2548
rect 4024 2532 4040 2548
rect 3896 2512 3912 2528
rect 3928 2512 3960 2528
rect 3976 2512 3992 2528
rect 3896 2472 3912 2488
rect 3928 2472 3944 2488
rect 3896 2372 3912 2388
rect 3800 2272 3816 2288
rect 3832 2272 3848 2288
rect 3800 2152 3816 2168
rect 3880 2292 3896 2308
rect 4200 2732 4216 2748
rect 4248 3072 4264 3088
rect 4328 3072 4344 3088
rect 4344 3052 4360 3068
rect 4584 3292 4600 3308
rect 4616 3412 4632 3428
rect 4696 3392 4712 3408
rect 4840 3452 4856 3468
rect 4744 3352 4760 3368
rect 4808 3352 4824 3368
rect 4872 3352 4888 3368
rect 4680 3332 4696 3348
rect 4712 3332 4728 3348
rect 4504 3272 4520 3288
rect 4568 3272 4584 3288
rect 4456 3252 4472 3268
rect 4440 3232 4456 3248
rect 4488 3152 4504 3168
rect 4488 3112 4504 3128
rect 4616 3252 4632 3268
rect 4600 3232 4616 3248
rect 4568 3172 4584 3188
rect 4520 3152 4552 3168
rect 4552 3092 4568 3108
rect 4440 3072 4472 3088
rect 4408 3052 4440 3068
rect 4472 3012 4488 3028
rect 4504 2992 4520 3008
rect 4280 2932 4296 2948
rect 4264 2912 4280 2928
rect 4248 2852 4264 2868
rect 4312 2792 4328 2808
rect 4632 3232 4648 3248
rect 4632 3192 4648 3208
rect 4696 3292 4712 3308
rect 4664 3212 4680 3228
rect 4744 3312 4760 3328
rect 4776 3292 4792 3308
rect 4792 3292 4808 3308
rect 4840 3312 4856 3328
rect 4728 3272 4744 3288
rect 4824 3272 4840 3288
rect 4712 3172 4728 3188
rect 4664 3152 4680 3168
rect 4712 3152 4728 3168
rect 4648 3132 4664 3148
rect 4696 3112 4712 3128
rect 4728 3112 4744 3128
rect 4760 3112 4776 3128
rect 4696 3072 4712 3088
rect 4744 3072 4760 3088
rect 4792 3072 4808 3088
rect 4568 2992 4584 3008
rect 4792 3052 4808 3068
rect 4664 3032 4680 3048
rect 4776 3032 4792 3048
rect 4648 2992 4664 3008
rect 4728 2972 4744 2988
rect 4744 2952 4760 2968
rect 4584 2932 4600 2948
rect 4712 2932 4728 2948
rect 4520 2912 4536 2928
rect 4552 2912 4568 2928
rect 4424 2892 4440 2908
rect 4456 2892 4472 2908
rect 4520 2892 4536 2908
rect 4552 2892 4568 2908
rect 4392 2812 4408 2828
rect 4376 2752 4392 2768
rect 4280 2732 4296 2748
rect 4200 2672 4216 2688
rect 4216 2672 4232 2688
rect 4200 2632 4216 2648
rect 4184 2572 4200 2588
rect 4120 2532 4136 2548
rect 4328 2712 4344 2728
rect 4248 2672 4264 2688
rect 4312 2672 4328 2688
rect 4664 2912 4680 2928
rect 4744 2912 4760 2928
rect 4664 2892 4680 2908
rect 4600 2872 4616 2888
rect 4632 2872 4648 2888
rect 4584 2812 4600 2828
rect 4440 2792 4456 2808
rect 4504 2792 4520 2808
rect 4504 2732 4520 2748
rect 4360 2672 4392 2688
rect 4344 2632 4360 2648
rect 4376 2632 4392 2648
rect 4312 2612 4328 2628
rect 4344 2592 4360 2608
rect 4264 2572 4280 2588
rect 4168 2512 4184 2528
rect 3960 2492 3976 2508
rect 4088 2492 4104 2508
rect 4200 2492 4216 2508
rect 4120 2472 4136 2488
rect 4440 2672 4456 2688
rect 4424 2632 4456 2648
rect 4408 2572 4440 2588
rect 4296 2532 4312 2548
rect 4344 2532 4360 2548
rect 4344 2512 4360 2528
rect 4376 2512 4392 2528
rect 4232 2492 4248 2508
rect 4072 2432 4088 2448
rect 4040 2392 4056 2408
rect 4072 2372 4088 2388
rect 4008 2312 4024 2328
rect 4232 2332 4248 2348
rect 3976 2252 3992 2268
rect 4024 2232 4040 2248
rect 4184 2232 4200 2248
rect 3885 2202 3921 2218
rect 3928 2192 3944 2208
rect 3960 2192 3976 2208
rect 3944 2132 3960 2148
rect 3672 2112 3688 2128
rect 3736 2112 3752 2128
rect 3656 2052 3672 2068
rect 3640 2032 3656 2048
rect 3544 2012 3560 2028
rect 3528 1992 3544 2008
rect 3592 1992 3608 2008
rect 3592 1952 3608 1968
rect 3528 1932 3544 1948
rect 3768 1992 3784 2008
rect 3640 1892 3656 1908
rect 3704 1892 3720 1908
rect 3672 1872 3688 1888
rect 3624 1852 3640 1868
rect 3560 1832 3576 1848
rect 3560 1792 3576 1808
rect 3464 1772 3480 1788
rect 3416 1752 3432 1768
rect 3352 1732 3368 1748
rect 3256 1692 3272 1708
rect 3288 1692 3304 1708
rect 3304 1692 3320 1708
rect 3272 1672 3288 1688
rect 3336 1672 3352 1688
rect 3336 1652 3352 1668
rect 3288 1612 3304 1628
rect 3288 1552 3304 1568
rect 3224 1532 3240 1548
rect 3272 1492 3288 1508
rect 3224 1472 3240 1488
rect 3176 1372 3192 1388
rect 3208 1452 3224 1468
rect 3272 1452 3288 1468
rect 3192 1312 3208 1328
rect 3144 1292 3160 1308
rect 3192 1232 3208 1248
rect 3272 1372 3288 1388
rect 3400 1712 3416 1728
rect 3560 1752 3576 1768
rect 3416 1672 3432 1688
rect 3448 1672 3480 1688
rect 3368 1632 3384 1648
rect 3304 1492 3320 1508
rect 3416 1652 3432 1668
rect 3400 1592 3416 1608
rect 3496 1692 3512 1708
rect 3528 1672 3544 1688
rect 3464 1552 3480 1568
rect 3416 1532 3432 1548
rect 3352 1472 3368 1488
rect 3432 1452 3448 1468
rect 3304 1352 3320 1368
rect 3368 1352 3384 1368
rect 3304 1314 3320 1328
rect 3304 1312 3320 1314
rect 3400 1312 3416 1328
rect 3432 1372 3448 1388
rect 3704 1812 3720 1828
rect 3624 1772 3640 1788
rect 3656 1772 3672 1788
rect 3768 1772 3784 1788
rect 3848 2112 3864 2128
rect 3816 2092 3832 2108
rect 3864 2092 3880 2108
rect 3864 2072 3880 2088
rect 3832 1906 3848 1908
rect 3832 1892 3848 1906
rect 3928 1872 3944 1888
rect 3944 1872 3960 1888
rect 3816 1812 3832 1828
rect 3704 1732 3720 1748
rect 3800 1732 3816 1748
rect 3576 1652 3608 1668
rect 3640 1612 3656 1628
rect 3528 1552 3544 1568
rect 3656 1552 3672 1568
rect 3560 1532 3576 1548
rect 3720 1672 3752 1688
rect 3704 1552 3720 1568
rect 3885 1802 3921 1818
rect 4008 2172 4024 2188
rect 4008 2152 4024 2168
rect 3992 2132 4008 2148
rect 3976 2112 3992 2128
rect 4008 2092 4024 2108
rect 3976 1912 3992 1928
rect 3960 1812 3976 1828
rect 3928 1792 3944 1808
rect 3832 1772 3848 1788
rect 3880 1772 3896 1788
rect 3784 1712 3800 1728
rect 3864 1712 3880 1728
rect 3976 1792 3992 1808
rect 3960 1752 3992 1768
rect 4104 2192 4120 2208
rect 4072 2152 4088 2168
rect 4088 2072 4104 2088
rect 4184 2212 4200 2228
rect 4200 2192 4216 2208
rect 4200 2172 4216 2188
rect 4168 2152 4184 2168
rect 4216 2152 4232 2168
rect 4184 2112 4200 2128
rect 4168 2092 4184 2108
rect 4088 2052 4104 2068
rect 4152 2052 4168 2068
rect 4040 1932 4056 1948
rect 4136 1992 4152 2008
rect 4136 1972 4152 1988
rect 4104 1912 4120 1928
rect 4040 1892 4056 1908
rect 4200 1892 4216 1908
rect 4072 1792 4088 1808
rect 4184 1832 4200 1848
rect 4120 1812 4136 1828
rect 4056 1772 4072 1788
rect 4104 1772 4120 1788
rect 4104 1752 4120 1768
rect 4088 1732 4104 1748
rect 4008 1712 4024 1728
rect 3816 1692 3832 1708
rect 3928 1692 3944 1708
rect 3960 1692 3976 1708
rect 3992 1692 4008 1708
rect 3960 1672 3976 1688
rect 3768 1652 3784 1668
rect 4232 2132 4248 2148
rect 4232 1912 4248 1928
rect 4328 2492 4344 2508
rect 4392 2492 4408 2508
rect 4296 2472 4312 2488
rect 4392 2472 4424 2488
rect 4360 2452 4376 2468
rect 4296 2432 4312 2448
rect 4488 2712 4504 2728
rect 4552 2672 4568 2688
rect 4504 2652 4520 2668
rect 4504 2612 4520 2628
rect 4488 2552 4504 2568
rect 4552 2532 4568 2548
rect 4456 2472 4472 2488
rect 4440 2432 4456 2448
rect 4520 2432 4536 2448
rect 4568 2412 4584 2428
rect 4616 2672 4632 2688
rect 4760 2892 4776 2908
rect 4808 3012 4824 3028
rect 4872 3072 4888 3088
rect 4872 3052 4888 3068
rect 4968 3672 4984 3688
rect 4909 3602 4945 3618
rect 4968 3592 4984 3608
rect 5096 3892 5112 3908
rect 5144 3892 5160 3908
rect 5112 3872 5128 3888
rect 5080 3852 5096 3868
rect 5064 3832 5080 3848
rect 5240 4592 5256 4608
rect 6280 4732 6296 4748
rect 6392 4732 6408 4748
rect 5512 4692 5528 4708
rect 5736 4706 5752 4708
rect 5736 4692 5752 4706
rect 5896 4692 5912 4708
rect 6152 4706 6168 4708
rect 6152 4692 6168 4706
rect 5640 4672 5656 4688
rect 5800 4672 5816 4688
rect 5640 4652 5656 4668
rect 5928 4652 5944 4668
rect 5528 4632 5544 4648
rect 5544 4612 5560 4628
rect 5352 4572 5368 4588
rect 5384 4572 5400 4588
rect 5432 4552 5448 4568
rect 5480 4552 5496 4568
rect 5560 4552 5576 4568
rect 5272 4532 5288 4548
rect 5448 4532 5464 4548
rect 5192 4512 5208 4528
rect 5208 4492 5224 4508
rect 5224 4472 5240 4488
rect 5256 4452 5272 4468
rect 5192 4432 5208 4448
rect 5368 4512 5384 4528
rect 5288 4472 5304 4488
rect 5320 4452 5336 4468
rect 5352 4292 5368 4308
rect 5272 4252 5304 4268
rect 5176 4172 5192 4188
rect 5224 4172 5240 4188
rect 5192 4112 5208 4128
rect 5208 4092 5224 4108
rect 5176 4032 5192 4048
rect 5240 4152 5256 4168
rect 5224 3972 5240 3988
rect 5176 3912 5192 3928
rect 5208 3912 5224 3928
rect 5176 3892 5192 3908
rect 5160 3832 5176 3848
rect 5144 3812 5160 3828
rect 5176 3732 5192 3748
rect 5080 3712 5096 3728
rect 5064 3672 5080 3688
rect 5160 3632 5176 3648
rect 5048 3612 5064 3628
rect 5096 3612 5112 3628
rect 5128 3612 5144 3628
rect 5016 3552 5032 3568
rect 5160 3592 5176 3608
rect 5032 3506 5048 3508
rect 5032 3492 5048 3506
rect 5112 3492 5128 3508
rect 5224 3752 5240 3768
rect 5208 3652 5224 3668
rect 5192 3532 5208 3548
rect 5176 3472 5192 3488
rect 4920 3432 4936 3448
rect 5144 3452 5160 3468
rect 5192 3452 5208 3468
rect 5128 3432 5144 3448
rect 5176 3432 5192 3448
rect 5064 3392 5080 3408
rect 5048 3352 5064 3368
rect 4952 3332 4968 3348
rect 5224 3412 5240 3428
rect 5144 3332 5160 3348
rect 4920 3312 4936 3328
rect 4920 3292 4936 3308
rect 5000 3312 5016 3328
rect 5032 3292 5048 3308
rect 4909 3202 4945 3218
rect 4968 3212 4984 3228
rect 5080 3292 5096 3308
rect 5112 3232 5128 3248
rect 4968 3172 4984 3188
rect 5048 3172 5064 3188
rect 4968 3152 4984 3168
rect 5176 3292 5192 3308
rect 5160 3232 5176 3248
rect 5144 3112 5160 3128
rect 5000 3092 5016 3108
rect 4888 3012 4904 3028
rect 4856 2972 4872 2988
rect 4920 2972 4936 2988
rect 4872 2912 4888 2928
rect 4904 2912 4920 2928
rect 4920 2912 4936 2928
rect 4808 2892 4824 2908
rect 4840 2892 4856 2908
rect 4824 2852 4840 2868
rect 5016 3072 5048 3088
rect 4984 3052 5000 3068
rect 4968 2952 4984 2968
rect 5000 2952 5016 2968
rect 4744 2772 4760 2788
rect 4744 2752 4760 2768
rect 4696 2672 4712 2688
rect 4728 2612 4744 2628
rect 4760 2612 4776 2628
rect 4696 2572 4712 2588
rect 4744 2572 4760 2588
rect 4632 2552 4648 2568
rect 4600 2472 4616 2488
rect 4584 2392 4600 2408
rect 4632 2392 4648 2408
rect 4600 2332 4616 2348
rect 4504 2312 4520 2328
rect 4856 2812 4872 2828
rect 4909 2802 4945 2818
rect 4904 2712 4916 2728
rect 4916 2712 4920 2728
rect 4952 2712 4968 2728
rect 4984 2912 5000 2928
rect 5032 2912 5048 2928
rect 5272 4132 5288 4148
rect 5256 4112 5272 4128
rect 5272 4092 5288 4108
rect 5256 3852 5272 3868
rect 5256 3792 5272 3808
rect 5256 3712 5272 3728
rect 5256 3472 5272 3488
rect 5256 3412 5272 3428
rect 5352 4272 5368 4288
rect 5320 4232 5336 4248
rect 5352 4232 5368 4248
rect 5304 4172 5336 4188
rect 5304 4052 5320 4068
rect 5288 3872 5304 3888
rect 5336 3932 5352 3948
rect 5933 4602 5969 4618
rect 6120 4672 6136 4688
rect 6008 4572 6024 4588
rect 6040 4572 6056 4588
rect 5912 4552 5928 4568
rect 5992 4552 6008 4568
rect 6248 4632 6264 4648
rect 5880 4532 5896 4548
rect 5944 4532 5960 4548
rect 5704 4514 5720 4528
rect 5704 4512 5720 4514
rect 5768 4512 5784 4528
rect 5816 4512 5832 4528
rect 5448 4492 5464 4508
rect 5480 4492 5496 4508
rect 5768 4492 5784 4508
rect 5464 4472 5480 4488
rect 5416 4452 5432 4468
rect 5400 4412 5416 4428
rect 5656 4472 5672 4488
rect 5528 4432 5544 4448
rect 5496 4392 5512 4408
rect 5416 4332 5432 4348
rect 5544 4312 5560 4328
rect 5448 4292 5464 4308
rect 5384 4252 5400 4268
rect 5416 4272 5432 4288
rect 5400 4232 5432 4248
rect 5368 4192 5400 4208
rect 5480 4252 5496 4268
rect 5512 4252 5528 4268
rect 5432 4192 5448 4208
rect 5416 4172 5432 4188
rect 5384 4112 5400 4128
rect 5400 4112 5416 4128
rect 5368 4072 5384 4088
rect 5448 4072 5464 4088
rect 5432 4052 5448 4068
rect 5400 3912 5416 3928
rect 5512 4232 5528 4248
rect 5528 4212 5544 4228
rect 5512 4192 5528 4208
rect 5832 4472 5848 4488
rect 5816 4452 5848 4468
rect 5592 4372 5608 4388
rect 5576 4292 5592 4308
rect 5704 4312 5716 4328
rect 5716 4312 5720 4328
rect 5736 4312 5752 4328
rect 5768 4312 5784 4328
rect 5800 4312 5816 4328
rect 5608 4292 5624 4308
rect 5688 4292 5704 4308
rect 5672 4272 5688 4288
rect 5528 4052 5544 4068
rect 5560 4052 5576 4068
rect 5512 3972 5528 3988
rect 5320 3892 5336 3908
rect 5448 3892 5464 3908
rect 5480 3892 5496 3908
rect 5336 3872 5352 3888
rect 5304 3772 5336 3788
rect 5288 3692 5304 3708
rect 5368 3752 5384 3768
rect 5448 3872 5464 3888
rect 5432 3832 5448 3848
rect 5432 3752 5448 3768
rect 5416 3732 5432 3748
rect 5384 3712 5400 3728
rect 5400 3712 5416 3728
rect 5304 3652 5320 3668
rect 5384 3632 5400 3648
rect 5336 3492 5352 3508
rect 5288 3372 5304 3388
rect 5272 3312 5288 3328
rect 5256 3292 5272 3308
rect 5368 3432 5384 3448
rect 5368 3392 5384 3408
rect 5336 3312 5352 3328
rect 5320 3232 5336 3248
rect 5240 3212 5272 3228
rect 5192 3192 5224 3208
rect 5080 3092 5096 3108
rect 5176 3092 5192 3108
rect 5096 3052 5112 3068
rect 5144 3032 5160 3048
rect 5112 3012 5128 3028
rect 5080 2912 5096 2928
rect 5048 2892 5064 2908
rect 5096 2892 5112 2908
rect 5032 2812 5048 2828
rect 5064 2872 5080 2888
rect 5080 2872 5096 2888
rect 5080 2852 5096 2868
rect 5176 2872 5192 2888
rect 5128 2752 5144 2768
rect 5160 2752 5176 2768
rect 5096 2732 5112 2748
rect 5048 2712 5064 2728
rect 4824 2552 4840 2568
rect 4680 2532 4696 2548
rect 4824 2532 4840 2548
rect 4696 2512 4712 2528
rect 4744 2512 4760 2528
rect 4792 2432 4808 2448
rect 4728 2412 4744 2428
rect 4760 2412 4776 2428
rect 4792 2392 4808 2408
rect 4712 2352 4728 2368
rect 4664 2332 4680 2348
rect 4648 2312 4664 2328
rect 4328 2292 4344 2308
rect 4536 2292 4552 2308
rect 4632 2292 4648 2308
rect 4680 2292 4696 2308
rect 4312 2272 4328 2288
rect 4584 2272 4600 2288
rect 4664 2272 4680 2288
rect 4712 2272 4728 2288
rect 4760 2272 4776 2288
rect 4472 2252 4488 2268
rect 4520 2252 4536 2268
rect 4280 2172 4296 2188
rect 4376 2152 4392 2168
rect 4392 2132 4408 2148
rect 4456 2132 4472 2148
rect 4264 2092 4280 2108
rect 4312 2092 4344 2108
rect 4280 2052 4296 2068
rect 4296 1932 4312 1948
rect 4328 1932 4344 1948
rect 4248 1872 4264 1888
rect 4232 1852 4248 1868
rect 4424 2112 4440 2128
rect 4376 2072 4392 2088
rect 4424 2052 4440 2068
rect 4456 2032 4472 2048
rect 4440 2012 4456 2028
rect 4408 1972 4424 1988
rect 4440 1972 4456 1988
rect 4408 1932 4424 1948
rect 4360 1912 4376 1928
rect 4408 1912 4424 1928
rect 4312 1892 4328 1908
rect 4280 1852 4296 1868
rect 4264 1792 4280 1808
rect 4248 1732 4264 1748
rect 4056 1712 4072 1728
rect 4104 1712 4120 1728
rect 3864 1652 3880 1668
rect 3944 1652 3960 1668
rect 4040 1652 4056 1668
rect 3848 1612 3864 1628
rect 3848 1592 3864 1608
rect 3768 1552 3784 1568
rect 3544 1492 3560 1508
rect 3672 1492 3688 1508
rect 3784 1492 3800 1508
rect 3800 1492 3816 1508
rect 3848 1492 3864 1508
rect 3896 1492 3912 1508
rect 3560 1452 3576 1468
rect 3592 1452 3608 1468
rect 3496 1392 3528 1408
rect 3464 1352 3480 1368
rect 3512 1372 3528 1388
rect 3544 1372 3560 1388
rect 3480 1332 3496 1348
rect 3448 1312 3464 1328
rect 3480 1312 3496 1328
rect 3384 1272 3400 1288
rect 3368 1252 3384 1268
rect 3208 1192 3224 1208
rect 3144 1152 3160 1168
rect 3176 1152 3192 1168
rect 3288 1152 3304 1168
rect 3144 1132 3160 1148
rect 3128 1092 3144 1108
rect 3112 1052 3128 1068
rect 3112 1012 3128 1028
rect 3176 1092 3192 1108
rect 3160 1072 3176 1088
rect 3160 1032 3176 1048
rect 3048 932 3064 948
rect 2920 892 2936 908
rect 2968 892 2984 908
rect 3080 892 3096 908
rect 3080 872 3096 888
rect 3016 792 3032 808
rect 3064 752 3080 768
rect 3208 1032 3224 1048
rect 3336 1032 3352 1048
rect 3272 1012 3288 1028
rect 3336 992 3352 1008
rect 3320 952 3352 968
rect 3160 912 3176 928
rect 3160 852 3176 868
rect 3144 752 3160 768
rect 3064 732 3080 748
rect 3096 732 3112 748
rect 3128 732 3160 748
rect 2936 712 2952 728
rect 3080 712 3096 728
rect 2920 692 2936 708
rect 2904 672 2920 688
rect 2776 632 2792 648
rect 2904 632 2920 648
rect 2792 612 2808 628
rect 2968 692 2984 708
rect 3032 692 3048 708
rect 3000 632 3016 648
rect 3000 612 3016 628
rect 3032 612 3048 628
rect 3032 572 3048 588
rect 2920 552 2936 568
rect 2760 514 2776 528
rect 2760 512 2776 514
rect 2904 452 2920 468
rect 2861 402 2897 418
rect 2728 372 2744 388
rect 2696 312 2712 328
rect 2616 252 2632 268
rect 2552 152 2568 168
rect 2328 112 2344 128
rect 2440 112 2456 128
rect 2488 112 2504 128
rect 2536 112 2552 128
rect 2632 232 2648 248
rect 2744 332 2760 348
rect 2792 332 2808 348
rect 2696 272 2712 288
rect 2856 312 2872 328
rect 2920 432 2936 448
rect 2952 372 2968 388
rect 3272 912 3288 928
rect 3224 872 3240 888
rect 3224 832 3240 848
rect 3192 732 3208 748
rect 3176 712 3192 728
rect 3208 712 3224 728
rect 3416 1172 3432 1188
rect 3432 1172 3448 1188
rect 3400 992 3416 1008
rect 3400 952 3416 968
rect 3304 912 3320 928
rect 3336 912 3352 928
rect 3368 892 3384 908
rect 3400 892 3416 908
rect 3384 792 3400 808
rect 3352 772 3368 788
rect 3240 712 3256 728
rect 3320 712 3336 728
rect 3272 692 3288 708
rect 3160 672 3176 688
rect 3224 672 3240 688
rect 3128 652 3144 668
rect 3160 652 3176 668
rect 3096 632 3112 648
rect 3208 632 3224 648
rect 3064 572 3080 588
rect 3112 572 3128 588
rect 3144 572 3160 588
rect 3192 572 3208 588
rect 3096 552 3112 568
rect 3192 532 3208 548
rect 3336 552 3352 568
rect 3272 532 3288 548
rect 3304 532 3320 548
rect 3048 492 3064 508
rect 3128 512 3144 528
rect 3064 452 3080 468
rect 3080 412 3096 428
rect 2984 332 3000 348
rect 3032 332 3048 348
rect 3016 312 3032 328
rect 3096 372 3112 388
rect 3112 352 3128 368
rect 3144 492 3176 508
rect 3288 492 3300 508
rect 3300 492 3304 508
rect 3304 492 3320 508
rect 3144 452 3160 468
rect 3288 452 3304 468
rect 3256 332 3272 348
rect 3432 1052 3448 1068
rect 3448 1032 3464 1048
rect 3432 752 3448 768
rect 3416 692 3432 708
rect 3576 1392 3592 1408
rect 3592 1352 3608 1368
rect 3576 1272 3592 1288
rect 3528 1192 3544 1208
rect 3512 1152 3528 1168
rect 3512 1112 3528 1128
rect 3496 972 3512 988
rect 3464 952 3480 968
rect 3464 912 3480 928
rect 3560 1032 3576 1048
rect 3784 1472 3800 1488
rect 3688 1452 3704 1468
rect 3736 1452 3752 1468
rect 3688 1432 3704 1448
rect 3672 1412 3688 1428
rect 3624 1352 3640 1368
rect 3752 1372 3768 1388
rect 3688 1332 3704 1348
rect 3672 1312 3688 1328
rect 3656 1292 3672 1308
rect 3688 1292 3704 1308
rect 3720 1292 3736 1308
rect 3608 1232 3624 1248
rect 3624 1212 3640 1228
rect 3736 1152 3752 1168
rect 3656 1092 3672 1108
rect 3608 1032 3624 1048
rect 3496 892 3512 908
rect 3624 952 3640 968
rect 3992 1612 4008 1628
rect 3960 1572 3976 1588
rect 4040 1552 4056 1568
rect 3960 1512 3976 1528
rect 4008 1512 4040 1528
rect 4072 1532 4088 1548
rect 4120 1692 4136 1708
rect 4120 1632 4136 1648
rect 4152 1692 4168 1708
rect 4136 1612 4152 1628
rect 4216 1652 4232 1668
rect 4232 1592 4248 1608
rect 4136 1512 4152 1528
rect 4168 1512 4184 1528
rect 4216 1512 4232 1528
rect 4232 1512 4248 1528
rect 3896 1472 3912 1488
rect 3992 1472 4008 1488
rect 4056 1472 4072 1488
rect 4088 1472 4104 1488
rect 4152 1472 4168 1488
rect 3864 1452 3880 1468
rect 3800 1432 3816 1448
rect 3784 1352 3800 1368
rect 3848 1272 3864 1288
rect 3768 1112 3784 1128
rect 3752 1072 3768 1088
rect 3672 1052 3704 1068
rect 3608 912 3624 928
rect 3656 912 3672 928
rect 3592 892 3608 908
rect 3736 992 3752 1008
rect 3720 952 3736 968
rect 3688 912 3704 928
rect 3704 892 3720 908
rect 3640 872 3656 888
rect 3576 832 3592 848
rect 3544 792 3560 808
rect 3832 1132 3848 1148
rect 3816 912 3832 928
rect 3832 772 3848 788
rect 3800 752 3816 768
rect 3736 732 3752 748
rect 3768 732 3784 748
rect 3544 712 3560 728
rect 3624 692 3640 708
rect 3688 692 3720 708
rect 3752 692 3768 708
rect 3768 692 3784 708
rect 3784 692 3800 708
rect 3528 672 3544 688
rect 3672 672 3688 688
rect 3400 632 3432 648
rect 3608 652 3624 668
rect 3528 632 3560 648
rect 3464 612 3480 628
rect 3416 532 3432 548
rect 3384 432 3400 448
rect 3304 372 3320 388
rect 3288 292 3304 308
rect 2808 272 2824 288
rect 2840 272 2856 288
rect 2952 272 2968 288
rect 3096 272 3112 288
rect 3192 272 3208 288
rect 2712 232 2728 248
rect 2776 232 2792 248
rect 2856 232 2872 248
rect 2712 212 2728 228
rect 2696 132 2712 148
rect 2744 132 2760 148
rect 2648 112 2664 128
rect 2232 92 2248 108
rect 2552 92 2568 108
rect 2600 92 2616 108
rect 2824 212 2840 228
rect 2776 192 2792 208
rect 2824 132 2840 148
rect 2888 152 2904 168
rect 3016 252 3032 268
rect 3048 252 3064 268
rect 3256 272 3272 288
rect 3288 272 3304 288
rect 3000 232 3016 248
rect 3224 232 3240 248
rect 2984 212 3000 228
rect 2968 132 2984 148
rect 3048 192 3064 208
rect 2968 112 2984 128
rect 3032 112 3048 128
rect 2824 92 2840 108
rect 3176 172 3192 188
rect 3288 212 3304 228
rect 3368 332 3384 348
rect 3320 292 3336 308
rect 3384 292 3400 308
rect 3416 292 3432 308
rect 3448 292 3464 308
rect 3400 272 3416 288
rect 3336 252 3352 268
rect 3304 192 3320 208
rect 3128 112 3144 128
rect 2760 72 2776 88
rect 3032 72 3048 88
rect 3064 72 3080 88
rect 472 52 488 68
rect 600 52 616 68
rect 936 52 952 68
rect 1432 52 1448 68
rect 2104 52 2120 68
rect 2264 52 2280 68
rect 797 2 833 18
rect 2861 2 2897 18
rect 3480 552 3496 568
rect 3496 492 3512 508
rect 3544 592 3560 608
rect 3656 592 3672 608
rect 3624 572 3640 588
rect 3576 532 3592 548
rect 3672 572 3688 588
rect 3720 572 3736 588
rect 3640 512 3656 528
rect 3704 512 3720 528
rect 3560 492 3576 508
rect 3544 472 3560 488
rect 3512 432 3544 448
rect 3528 372 3544 388
rect 3496 312 3512 328
rect 3800 552 3816 568
rect 3736 532 3752 548
rect 3768 532 3784 548
rect 3992 1452 4008 1468
rect 3944 1432 3960 1448
rect 3885 1402 3921 1418
rect 3944 1352 3960 1368
rect 3912 1314 3928 1328
rect 3912 1312 3928 1314
rect 3976 1312 3992 1328
rect 4040 1432 4056 1448
rect 4296 1732 4312 1748
rect 4296 1712 4312 1728
rect 4280 1692 4296 1708
rect 4264 1612 4280 1628
rect 4296 1592 4312 1608
rect 4264 1532 4280 1548
rect 4392 1892 4408 1908
rect 4360 1832 4376 1848
rect 4344 1692 4360 1708
rect 4360 1632 4376 1648
rect 4360 1612 4376 1628
rect 4696 2212 4712 2228
rect 4536 2192 4552 2208
rect 4648 2172 4664 2188
rect 4520 2072 4536 2088
rect 4488 2052 4504 2068
rect 4472 1992 4488 2008
rect 4600 2112 4616 2128
rect 4568 2092 4584 2108
rect 4616 2092 4632 2108
rect 4744 2112 4760 2128
rect 4664 2072 4680 2088
rect 4552 2052 4568 2068
rect 4584 2052 4600 2068
rect 4632 2052 4648 2068
rect 4648 2052 4664 2068
rect 4536 1972 4552 1988
rect 4728 1972 4744 1988
rect 4712 1912 4728 1928
rect 4552 1872 4568 1888
rect 4600 1872 4616 1888
rect 4568 1852 4584 1868
rect 4424 1792 4440 1808
rect 4392 1712 4408 1728
rect 4584 1812 4600 1828
rect 4920 2692 4936 2708
rect 4872 2672 4888 2688
rect 4888 2672 4904 2688
rect 4856 2632 4872 2648
rect 4856 2612 4872 2628
rect 4856 2552 4872 2568
rect 4840 2392 4856 2408
rect 4840 2372 4856 2388
rect 4808 2312 4824 2328
rect 4808 2272 4824 2288
rect 4824 2112 4840 2128
rect 4776 2072 4792 2088
rect 4776 2032 4792 2048
rect 4760 1932 4776 1948
rect 4824 1992 4840 2008
rect 4776 1912 4792 1928
rect 4808 1892 4824 1908
rect 4680 1872 4696 1888
rect 4616 1792 4648 1808
rect 4552 1772 4568 1788
rect 4584 1772 4600 1788
rect 4488 1752 4504 1768
rect 4520 1732 4536 1748
rect 4456 1712 4472 1728
rect 4488 1712 4504 1728
rect 4504 1692 4520 1708
rect 4472 1672 4488 1688
rect 4520 1672 4536 1688
rect 4520 1632 4536 1648
rect 4472 1612 4488 1628
rect 4376 1592 4392 1608
rect 4312 1572 4328 1588
rect 4344 1532 4360 1548
rect 4312 1512 4328 1528
rect 4248 1452 4264 1468
rect 4264 1432 4280 1448
rect 4104 1412 4120 1428
rect 4168 1412 4184 1428
rect 4072 1392 4088 1408
rect 4120 1392 4136 1408
rect 4040 1372 4056 1388
rect 4056 1332 4072 1348
rect 4232 1372 4248 1388
rect 4104 1312 4120 1328
rect 4008 1292 4024 1308
rect 4088 1292 4104 1308
rect 3992 1252 4008 1268
rect 4024 1252 4040 1268
rect 3864 1212 3880 1228
rect 3944 1172 3960 1188
rect 3864 1112 3880 1128
rect 4136 1332 4152 1348
rect 4168 1332 4184 1348
rect 4168 1292 4184 1308
rect 4120 1232 4136 1248
rect 4216 1272 4232 1288
rect 4040 1152 4056 1168
rect 4120 1152 4136 1168
rect 4200 1152 4216 1168
rect 4056 1132 4072 1148
rect 3885 1002 3921 1018
rect 3976 932 3992 948
rect 4008 932 4024 948
rect 4040 1052 4056 1068
rect 3928 912 3944 928
rect 4024 912 4040 928
rect 4088 1072 4104 1088
rect 4120 1072 4136 1088
rect 4152 992 4168 1008
rect 4120 972 4136 988
rect 4072 952 4088 968
rect 4088 952 4104 968
rect 4104 932 4120 948
rect 3976 872 3992 888
rect 4152 912 4168 928
rect 4232 1112 4248 1128
rect 4216 1052 4232 1068
rect 4248 1032 4264 1048
rect 4264 992 4280 1008
rect 4264 952 4280 968
rect 4184 932 4200 948
rect 4232 932 4248 948
rect 4136 872 4152 888
rect 4216 892 4232 908
rect 4248 912 4264 928
rect 4232 852 4248 868
rect 4264 832 4280 848
rect 4184 792 4200 808
rect 4264 792 4280 808
rect 4136 772 4152 788
rect 4056 732 4072 748
rect 4104 732 4120 748
rect 4120 732 4136 748
rect 3896 712 3912 728
rect 4008 712 4024 728
rect 4168 712 4184 728
rect 3880 672 3896 688
rect 4088 672 4104 688
rect 4104 672 4120 688
rect 4136 672 4152 688
rect 3880 652 3896 668
rect 3848 612 3864 628
rect 3864 592 3880 608
rect 3885 602 3921 618
rect 3864 572 3880 588
rect 3928 552 3944 568
rect 3960 552 3976 568
rect 3864 532 3880 548
rect 3752 512 3768 528
rect 3832 512 3848 528
rect 3752 472 3768 488
rect 3688 372 3704 388
rect 3736 372 3752 388
rect 3656 332 3672 348
rect 3640 312 3656 328
rect 3576 292 3608 308
rect 3544 272 3560 288
rect 3608 272 3624 288
rect 3432 232 3448 248
rect 3416 172 3432 188
rect 3288 132 3304 148
rect 3400 132 3416 148
rect 3256 112 3272 128
rect 3288 92 3304 108
rect 3384 92 3400 108
rect 3480 212 3496 228
rect 3496 152 3512 168
rect 3528 114 3544 128
rect 3528 112 3544 114
rect 3784 452 3800 468
rect 3976 512 3992 528
rect 3944 492 3960 508
rect 3896 472 3912 488
rect 4072 652 4088 668
rect 4264 772 4280 788
rect 4216 712 4232 728
rect 4248 692 4264 708
rect 4168 672 4184 688
rect 4152 652 4168 668
rect 4088 592 4104 608
rect 4104 552 4120 568
rect 4024 532 4040 548
rect 4056 532 4072 548
rect 4392 1492 4408 1508
rect 4504 1492 4520 1508
rect 4344 1472 4360 1488
rect 4376 1472 4392 1488
rect 4456 1472 4472 1488
rect 4424 1452 4440 1468
rect 4312 1412 4328 1428
rect 4600 1752 4616 1768
rect 4648 1632 4664 1648
rect 4552 1612 4568 1628
rect 4552 1592 4568 1608
rect 4584 1592 4600 1608
rect 4616 1592 4632 1608
rect 4680 1592 4696 1608
rect 4584 1572 4600 1588
rect 4536 1512 4552 1528
rect 4648 1512 4680 1528
rect 4632 1492 4648 1508
rect 4488 1452 4504 1468
rect 4472 1372 4488 1388
rect 4392 1292 4408 1308
rect 4472 1292 4488 1308
rect 4296 1192 4312 1208
rect 4536 1412 4552 1428
rect 4296 1172 4312 1188
rect 4488 1172 4504 1188
rect 4296 1152 4312 1168
rect 4392 1132 4408 1148
rect 4328 1112 4344 1128
rect 4360 1112 4376 1128
rect 4600 1472 4616 1488
rect 4664 1472 4680 1488
rect 4680 1472 4696 1488
rect 4840 1812 4856 1828
rect 4776 1792 4792 1808
rect 4808 1792 4824 1808
rect 4744 1772 4760 1788
rect 4776 1772 4792 1788
rect 4728 1752 4744 1768
rect 4712 1712 4728 1728
rect 4776 1712 4792 1728
rect 4744 1552 4760 1568
rect 4744 1532 4760 1548
rect 4712 1512 4728 1528
rect 4904 2452 4920 2468
rect 5096 2672 5112 2688
rect 5128 2672 5144 2688
rect 5016 2632 5032 2648
rect 5016 2612 5032 2628
rect 4968 2552 4984 2568
rect 4984 2532 5000 2548
rect 5016 2532 5032 2548
rect 4888 2392 4904 2408
rect 4909 2402 4945 2418
rect 4952 2412 4968 2428
rect 4872 2352 4888 2368
rect 4904 2132 4920 2148
rect 4904 2092 4920 2108
rect 4952 2092 4968 2108
rect 4952 2072 4968 2088
rect 4909 2002 4945 2018
rect 5112 2632 5128 2648
rect 5064 2552 5080 2568
rect 5064 2532 5080 2548
rect 5192 2852 5208 2868
rect 5192 2832 5208 2848
rect 5288 3172 5304 3188
rect 5352 3152 5368 3168
rect 5352 3132 5368 3148
rect 5336 3112 5352 3128
rect 5256 3092 5272 3108
rect 5224 3052 5240 3068
rect 5288 3052 5304 3068
rect 5352 3052 5368 3068
rect 5224 2912 5240 2928
rect 5304 3032 5320 3048
rect 5400 3412 5416 3428
rect 5464 3712 5480 3728
rect 5576 4012 5608 4028
rect 5640 4192 5656 4208
rect 5672 4172 5688 4188
rect 5656 4132 5672 4148
rect 5704 4272 5720 4288
rect 5720 4252 5736 4268
rect 6008 4512 6024 4528
rect 5896 4432 5912 4448
rect 5864 4392 5880 4408
rect 5848 4332 5864 4348
rect 5832 4312 5848 4328
rect 5816 4292 5832 4308
rect 5816 4272 5832 4288
rect 5752 4232 5768 4248
rect 5736 4212 5768 4228
rect 5704 4072 5720 4088
rect 5656 4012 5672 4028
rect 5672 3932 5688 3948
rect 5608 3912 5624 3928
rect 5688 3912 5704 3928
rect 5800 4192 5816 4208
rect 6040 4492 6056 4508
rect 5992 4472 6008 4488
rect 6056 4452 6072 4468
rect 6024 4372 6040 4388
rect 5928 4352 5944 4368
rect 5880 4332 5896 4348
rect 5848 4272 5864 4288
rect 5816 4152 5832 4168
rect 5736 4072 5752 4088
rect 5800 4072 5816 4088
rect 5880 4112 5896 4128
rect 5752 4052 5768 4068
rect 5848 4052 5864 4068
rect 5720 4012 5736 4028
rect 5640 3892 5656 3908
rect 5688 3892 5720 3908
rect 5576 3872 5592 3888
rect 5624 3872 5640 3888
rect 5672 3872 5688 3888
rect 5528 3832 5544 3848
rect 5512 3772 5528 3788
rect 5560 3772 5576 3788
rect 5640 3712 5656 3728
rect 5448 3692 5464 3708
rect 5448 3612 5464 3628
rect 6088 4492 6104 4508
rect 6136 4472 6152 4488
rect 6168 4452 6184 4468
rect 6120 4392 6136 4408
rect 6104 4352 6120 4368
rect 6024 4312 6040 4328
rect 6072 4312 6088 4328
rect 5933 4202 5969 4218
rect 5960 4152 5976 4168
rect 5912 4092 5928 4108
rect 5896 4072 5912 4088
rect 5944 4052 5960 4068
rect 5912 4032 5928 4048
rect 5912 4012 5928 4028
rect 5864 3992 5880 4008
rect 5768 3872 5784 3888
rect 5880 3872 5896 3888
rect 6056 4272 6072 4288
rect 6680 4692 6696 4708
rect 6488 4572 6504 4588
rect 6584 4572 6600 4588
rect 6376 4512 6392 4528
rect 6504 4512 6520 4528
rect 6344 4492 6360 4508
rect 6456 4492 6472 4508
rect 6648 4492 6664 4508
rect 6184 4352 6200 4368
rect 6808 4312 6824 4328
rect 6120 4252 6136 4268
rect 6184 4252 6200 4268
rect 5992 4232 6008 4248
rect 6120 4152 6136 4168
rect 5976 4112 5992 4128
rect 6040 4112 6056 4128
rect 5976 4012 5992 4028
rect 6008 4092 6024 4108
rect 6040 4092 6056 4108
rect 6088 4112 6104 4128
rect 6280 4272 6296 4288
rect 6312 4232 6328 4248
rect 6424 4272 6440 4288
rect 6200 4152 6216 4168
rect 6280 4152 6296 4168
rect 6328 4152 6344 4168
rect 6408 4152 6424 4168
rect 6296 4132 6312 4148
rect 6168 4112 6184 4128
rect 6072 4092 6088 4108
rect 6056 4072 6072 4088
rect 6040 4032 6056 4048
rect 6024 3992 6040 4008
rect 5976 3972 5992 3988
rect 5992 3972 6008 3988
rect 5960 3852 5976 3868
rect 6024 3892 6040 3908
rect 6008 3872 6024 3888
rect 6152 4092 6168 4108
rect 6120 4012 6136 4028
rect 6088 3932 6104 3948
rect 6152 3892 6168 3908
rect 6104 3872 6120 3888
rect 6136 3872 6152 3888
rect 6152 3872 6168 3888
rect 6104 3852 6120 3868
rect 5992 3832 6008 3848
rect 5933 3802 5969 3818
rect 6024 3792 6040 3808
rect 5688 3692 5704 3708
rect 5496 3592 5512 3608
rect 5608 3592 5624 3608
rect 5720 3512 5736 3528
rect 5976 3632 5992 3648
rect 5976 3552 5992 3568
rect 6008 3552 6024 3568
rect 5752 3532 5768 3548
rect 5864 3532 5880 3548
rect 5640 3492 5656 3508
rect 5448 3412 5464 3428
rect 5416 3372 5432 3388
rect 5784 3492 5800 3508
rect 5688 3472 5704 3488
rect 5480 3452 5496 3468
rect 5688 3432 5704 3448
rect 5464 3392 5480 3408
rect 5576 3392 5592 3408
rect 5464 3372 5480 3388
rect 5528 3352 5544 3368
rect 5608 3332 5640 3348
rect 5464 3312 5480 3328
rect 5496 3312 5512 3328
rect 5560 3312 5576 3328
rect 5640 3312 5656 3328
rect 5416 3272 5432 3288
rect 5544 3292 5560 3308
rect 5464 3252 5480 3268
rect 5608 3292 5624 3308
rect 5560 3132 5576 3148
rect 5416 3112 5432 3128
rect 5448 3112 5464 3128
rect 5496 3112 5512 3128
rect 5608 3192 5624 3208
rect 5384 3092 5400 3108
rect 5480 3092 5496 3108
rect 5512 3092 5528 3108
rect 5592 3092 5608 3108
rect 5400 3072 5416 3088
rect 5272 2912 5288 2928
rect 5240 2892 5256 2908
rect 5272 2892 5288 2908
rect 5208 2792 5224 2808
rect 5208 2672 5224 2688
rect 5192 2632 5208 2648
rect 5192 2612 5208 2628
rect 5192 2552 5208 2568
rect 5240 2752 5256 2768
rect 5256 2692 5272 2708
rect 5304 2792 5320 2808
rect 5240 2672 5256 2688
rect 5272 2652 5304 2668
rect 5240 2632 5256 2648
rect 5224 2532 5240 2548
rect 5192 2492 5208 2508
rect 5096 2472 5112 2488
rect 5176 2412 5192 2428
rect 5064 2352 5080 2368
rect 5096 2352 5112 2368
rect 5160 2312 5176 2328
rect 5128 2292 5144 2308
rect 5080 2272 5096 2288
rect 5096 2272 5112 2288
rect 5048 2252 5064 2268
rect 5048 2192 5064 2208
rect 5080 2132 5096 2148
rect 5208 2312 5224 2328
rect 5160 2192 5176 2208
rect 5144 2112 5160 2128
rect 5064 2092 5080 2108
rect 5144 2092 5160 2108
rect 5032 2052 5048 2068
rect 5064 2032 5080 2048
rect 5000 1992 5016 2008
rect 5112 1992 5128 2008
rect 5048 1952 5064 1968
rect 4904 1912 4920 1928
rect 5000 1912 5016 1928
rect 4968 1892 4984 1908
rect 5176 2112 5192 2128
rect 5224 2252 5240 2268
rect 5672 3272 5688 3288
rect 5656 3172 5672 3188
rect 5624 3132 5640 3148
rect 5640 3072 5656 3088
rect 5528 3052 5544 3068
rect 5416 2992 5432 3008
rect 5384 2892 5400 2908
rect 5496 2912 5512 2928
rect 5480 2892 5496 2908
rect 5480 2872 5496 2888
rect 5416 2852 5432 2868
rect 5496 2852 5512 2868
rect 5544 3032 5560 3048
rect 5544 3012 5560 3028
rect 5560 2992 5576 3008
rect 5624 3032 5640 3048
rect 5592 2972 5624 2988
rect 5656 2992 5672 3008
rect 5640 2972 5656 2988
rect 5704 3352 5720 3368
rect 5704 3332 5720 3348
rect 5784 3452 5800 3468
rect 5704 3312 5720 3328
rect 5752 3312 5768 3328
rect 5720 3272 5736 3288
rect 5704 3192 5720 3208
rect 5784 3272 5800 3288
rect 5768 3192 5784 3208
rect 5736 3132 5752 3148
rect 5816 3492 5832 3508
rect 5880 3492 5896 3508
rect 5832 3352 5848 3368
rect 5992 3492 6008 3508
rect 5960 3472 5976 3488
rect 5976 3472 5992 3488
rect 5864 3432 5880 3448
rect 5928 3432 5944 3448
rect 5933 3402 5969 3418
rect 5896 3352 5912 3368
rect 5944 3352 5960 3368
rect 5896 3332 5912 3348
rect 5832 3272 5848 3288
rect 5800 3112 5816 3128
rect 5816 3112 5832 3128
rect 5704 3092 5720 3108
rect 5704 3012 5720 3028
rect 5784 2972 5816 2988
rect 5992 3392 6008 3408
rect 6232 4092 6248 4108
rect 6216 4052 6232 4068
rect 6344 4072 6360 4088
rect 6312 3972 6328 3988
rect 6264 3912 6280 3928
rect 6280 3892 6296 3908
rect 6280 3852 6296 3868
rect 6184 3792 6200 3808
rect 6232 3792 6248 3808
rect 6056 3752 6072 3768
rect 6120 3752 6136 3768
rect 6040 3732 6056 3748
rect 6136 3732 6152 3748
rect 6088 3712 6104 3728
rect 6056 3692 6072 3708
rect 6360 3932 6376 3948
rect 6552 4192 6568 4208
rect 6552 4172 6568 4188
rect 6744 4192 6760 4208
rect 6696 4172 6712 4188
rect 6728 4172 6744 4188
rect 6472 4132 6488 4148
rect 6616 4132 6632 4148
rect 6440 4112 6456 4128
rect 6664 4112 6680 4128
rect 6536 4092 6552 4108
rect 6600 4092 6616 4108
rect 6632 4072 6648 4088
rect 6616 4052 6632 4068
rect 6440 3952 6456 3968
rect 6584 3912 6600 3928
rect 6424 3892 6440 3908
rect 6488 3906 6504 3908
rect 6488 3892 6504 3906
rect 6344 3852 6360 3868
rect 6312 3812 6328 3828
rect 6296 3752 6312 3768
rect 6280 3732 6296 3748
rect 6184 3712 6200 3728
rect 6216 3712 6232 3728
rect 6152 3632 6168 3648
rect 6152 3612 6168 3628
rect 6184 3692 6200 3708
rect 6168 3592 6184 3608
rect 6168 3572 6184 3588
rect 6152 3532 6168 3548
rect 6024 3452 6040 3468
rect 5928 3292 5944 3308
rect 5880 3212 5896 3228
rect 5864 3192 5880 3208
rect 5896 3172 5912 3188
rect 5912 3152 5928 3168
rect 5896 3132 5912 3148
rect 5848 3072 5864 3088
rect 5880 3052 5896 3068
rect 5944 3172 5960 3188
rect 5944 3052 5960 3068
rect 5928 3032 5944 3048
rect 5848 3012 5864 3028
rect 5592 2932 5608 2948
rect 5624 2932 5640 2948
rect 5720 2932 5736 2948
rect 5576 2892 5592 2908
rect 5544 2832 5560 2848
rect 5528 2792 5544 2808
rect 5576 2792 5592 2808
rect 5352 2772 5368 2788
rect 5544 2772 5560 2788
rect 5400 2752 5416 2768
rect 5432 2752 5448 2768
rect 5528 2752 5544 2768
rect 5352 2692 5368 2708
rect 5384 2692 5400 2708
rect 5352 2672 5368 2688
rect 5320 2632 5336 2648
rect 5336 2592 5352 2608
rect 5416 2692 5432 2708
rect 5512 2652 5528 2668
rect 5432 2632 5448 2648
rect 5480 2632 5496 2648
rect 5400 2612 5416 2628
rect 5464 2592 5480 2608
rect 5496 2592 5512 2608
rect 5432 2572 5448 2588
rect 5416 2552 5432 2568
rect 5272 2472 5288 2488
rect 5256 2312 5272 2328
rect 5304 2452 5320 2468
rect 5288 2312 5304 2328
rect 5272 2272 5288 2288
rect 5240 2212 5256 2228
rect 5288 2152 5304 2168
rect 5320 2272 5336 2288
rect 5400 2512 5416 2528
rect 5384 2452 5400 2468
rect 5352 2412 5368 2428
rect 5416 2312 5432 2328
rect 5656 2912 5672 2928
rect 5672 2892 5688 2908
rect 5640 2872 5656 2888
rect 5560 2692 5576 2708
rect 5608 2632 5624 2648
rect 5576 2592 5592 2608
rect 5448 2532 5464 2548
rect 5528 2532 5544 2548
rect 5480 2492 5496 2508
rect 5496 2412 5528 2428
rect 5528 2392 5544 2408
rect 5448 2312 5464 2328
rect 5368 2292 5384 2308
rect 5400 2292 5416 2308
rect 5560 2312 5576 2328
rect 5768 2892 5784 2908
rect 5752 2752 5768 2768
rect 5880 2992 5896 3008
rect 5933 3002 5969 3018
rect 5912 2932 5928 2948
rect 5880 2912 5896 2928
rect 5928 2912 5944 2928
rect 5928 2832 5944 2848
rect 5960 2772 5976 2788
rect 5832 2732 5848 2748
rect 5752 2712 5768 2728
rect 5880 2712 5896 2728
rect 5720 2692 5736 2708
rect 5800 2692 5816 2708
rect 6072 3412 6088 3428
rect 6056 3352 6072 3368
rect 6088 3352 6104 3368
rect 6040 3272 6056 3288
rect 6008 3232 6024 3248
rect 6024 3232 6040 3248
rect 6008 3212 6024 3228
rect 6104 3212 6120 3228
rect 6056 3192 6072 3208
rect 6088 3172 6104 3188
rect 6072 3152 6088 3168
rect 6008 3112 6024 3128
rect 6040 3112 6056 3128
rect 6056 3012 6072 3028
rect 6008 2952 6024 2968
rect 6104 3052 6120 3068
rect 6088 2952 6104 2968
rect 6008 2932 6024 2948
rect 6072 2892 6088 2908
rect 6264 3712 6280 3728
rect 6216 3532 6232 3548
rect 6248 3532 6264 3548
rect 6296 3712 6312 3728
rect 6296 3552 6312 3568
rect 6248 3512 6264 3528
rect 6280 3512 6296 3528
rect 6440 3792 6456 3808
rect 6408 3772 6424 3788
rect 6424 3752 6440 3768
rect 6376 3732 6392 3748
rect 6376 3712 6392 3728
rect 6456 3692 6472 3708
rect 6344 3632 6360 3648
rect 6472 3612 6488 3628
rect 6376 3592 6392 3608
rect 6328 3552 6360 3568
rect 6200 3492 6216 3508
rect 6296 3472 6312 3488
rect 6152 3452 6168 3468
rect 6184 3432 6200 3448
rect 6328 3472 6344 3488
rect 6312 3392 6328 3408
rect 6168 3352 6184 3368
rect 6312 3352 6328 3368
rect 6408 3572 6424 3588
rect 6376 3452 6392 3468
rect 6536 3812 6552 3828
rect 6504 3752 6520 3768
rect 6520 3732 6536 3748
rect 6504 3492 6520 3508
rect 6424 3432 6440 3448
rect 6344 3412 6360 3428
rect 6264 3332 6280 3348
rect 6360 3392 6376 3408
rect 6392 3392 6408 3408
rect 6504 3432 6520 3448
rect 6456 3372 6472 3388
rect 6360 3352 6376 3368
rect 6376 3352 6392 3368
rect 6488 3352 6504 3368
rect 6568 3892 6584 3908
rect 6568 3872 6584 3888
rect 6600 3872 6616 3888
rect 6552 3772 6568 3788
rect 6616 3712 6648 3728
rect 6584 3672 6600 3688
rect 6600 3632 6616 3648
rect 6632 3632 6648 3648
rect 6680 3792 6696 3808
rect 6664 3732 6680 3748
rect 6680 3712 6696 3728
rect 6664 3472 6680 3488
rect 6200 3312 6216 3328
rect 6520 3312 6536 3328
rect 6184 3292 6200 3308
rect 6216 3292 6232 3308
rect 6248 3292 6264 3308
rect 6168 3252 6184 3268
rect 6136 3192 6152 3208
rect 6024 2872 6040 2888
rect 6120 2872 6136 2888
rect 6168 2992 6184 3008
rect 6168 2972 6184 2988
rect 6152 2892 6168 2908
rect 6136 2852 6152 2868
rect 6344 3292 6360 3308
rect 6424 3292 6440 3308
rect 6264 3152 6280 3168
rect 6280 3112 6296 3128
rect 6312 3112 6328 3128
rect 6248 3092 6264 3108
rect 6280 3072 6296 3088
rect 6360 3072 6376 3088
rect 6232 3052 6248 3068
rect 6280 3052 6296 3068
rect 6200 2972 6216 2988
rect 6264 2952 6280 2968
rect 6264 2932 6280 2948
rect 6248 2892 6264 2908
rect 6184 2752 6200 2768
rect 6024 2732 6056 2748
rect 6152 2732 6168 2748
rect 5976 2692 5992 2708
rect 5992 2692 6008 2708
rect 5704 2672 5720 2688
rect 5816 2672 5832 2688
rect 5864 2672 5880 2688
rect 5704 2612 5720 2628
rect 5864 2612 5880 2628
rect 5688 2592 5704 2608
rect 5832 2572 5864 2588
rect 5640 2552 5656 2568
rect 5768 2532 5784 2548
rect 5656 2512 5672 2528
rect 5624 2352 5640 2368
rect 5608 2332 5624 2348
rect 5656 2312 5672 2328
rect 5512 2292 5528 2308
rect 5416 2272 5432 2288
rect 5496 2272 5512 2288
rect 5336 2232 5352 2248
rect 5352 2152 5368 2168
rect 5320 2112 5336 2128
rect 5208 2092 5224 2108
rect 5256 2092 5272 2108
rect 5272 2072 5288 2088
rect 5224 2052 5240 2068
rect 5208 2032 5224 2048
rect 5304 2032 5320 2048
rect 5192 2012 5208 2028
rect 5224 2012 5240 2028
rect 5240 1892 5256 1908
rect 4888 1872 4904 1888
rect 4952 1832 4968 1848
rect 4904 1732 4920 1748
rect 4840 1712 4856 1728
rect 4984 1752 5000 1768
rect 4824 1672 4840 1688
rect 4872 1672 4888 1688
rect 4909 1602 4945 1618
rect 4952 1572 4968 1588
rect 4920 1552 4936 1568
rect 4776 1512 4792 1528
rect 4728 1492 4744 1508
rect 4904 1492 4920 1508
rect 4696 1452 4712 1468
rect 5048 1872 5064 1888
rect 5096 1872 5112 1888
rect 5160 1872 5176 1888
rect 5192 1872 5208 1888
rect 5032 1852 5048 1868
rect 5080 1832 5096 1848
rect 5096 1792 5112 1808
rect 5112 1752 5128 1768
rect 5016 1732 5032 1748
rect 5064 1712 5080 1728
rect 4792 1412 4808 1428
rect 4984 1412 5000 1428
rect 4600 1372 4616 1388
rect 5080 1652 5096 1668
rect 5096 1632 5112 1648
rect 5064 1512 5080 1528
rect 5144 1772 5160 1788
rect 5208 1752 5224 1768
rect 5144 1712 5160 1728
rect 5176 1692 5192 1708
rect 5272 1832 5288 1848
rect 5272 1792 5288 1808
rect 5256 1712 5272 1728
rect 5224 1612 5240 1628
rect 5112 1512 5128 1528
rect 5128 1512 5144 1528
rect 5176 1512 5192 1528
rect 5128 1492 5144 1508
rect 5016 1372 5048 1388
rect 5128 1432 5144 1448
rect 4680 1352 4696 1368
rect 4952 1352 4968 1368
rect 4632 1332 4648 1348
rect 4712 1332 4728 1348
rect 4776 1332 4792 1348
rect 4616 1312 4632 1328
rect 4664 1312 4680 1328
rect 4728 1312 4744 1328
rect 4600 1172 4616 1188
rect 4424 1112 4440 1128
rect 4584 1112 4600 1128
rect 4568 1092 4584 1108
rect 4600 1052 4616 1068
rect 4296 1012 4312 1028
rect 4328 1012 4344 1028
rect 4456 1012 4472 1028
rect 4488 1012 4504 1028
rect 4456 992 4472 1008
rect 4488 992 4504 1008
rect 4536 992 4552 1008
rect 4312 952 4328 968
rect 4376 952 4392 968
rect 4440 952 4456 968
rect 4520 952 4536 968
rect 4296 912 4312 928
rect 4328 912 4344 928
rect 4360 892 4376 908
rect 4408 892 4424 908
rect 4632 1252 4648 1268
rect 4632 1072 4648 1088
rect 4616 1012 4632 1028
rect 4600 952 4616 968
rect 4536 872 4552 888
rect 4488 852 4504 868
rect 4472 812 4488 828
rect 4552 792 4568 808
rect 4440 772 4456 788
rect 4296 712 4312 728
rect 4392 712 4408 728
rect 4616 892 4632 908
rect 4600 792 4616 808
rect 4584 752 4600 768
rect 4504 732 4536 748
rect 4568 732 4584 748
rect 4536 712 4552 728
rect 4344 692 4360 708
rect 4376 692 4392 708
rect 4488 692 4504 708
rect 4328 672 4344 688
rect 4408 672 4424 688
rect 4456 672 4472 688
rect 4520 672 4536 688
rect 4312 652 4328 668
rect 4392 652 4408 668
rect 4248 632 4264 648
rect 4344 632 4360 648
rect 4440 632 4456 648
rect 4248 612 4264 628
rect 4408 592 4424 608
rect 4248 572 4264 588
rect 4296 572 4312 588
rect 4392 572 4408 588
rect 4120 532 4136 548
rect 4024 512 4040 528
rect 4088 512 4104 528
rect 4120 512 4136 528
rect 4040 472 4056 488
rect 3992 432 4024 448
rect 4072 432 4088 448
rect 3800 392 3816 408
rect 4008 392 4024 408
rect 3688 292 3704 308
rect 3720 292 3752 308
rect 3800 292 3816 308
rect 3832 292 3848 308
rect 3976 292 3992 308
rect 3672 272 3688 288
rect 3752 272 3768 288
rect 3832 272 3848 288
rect 3960 272 3976 288
rect 3864 232 3880 248
rect 3848 192 3864 208
rect 3885 202 3921 218
rect 3656 172 3672 188
rect 3848 172 3864 188
rect 3688 152 3704 168
rect 4024 372 4040 388
rect 4280 552 4296 568
rect 4264 532 4280 548
rect 4328 532 4344 548
rect 4424 572 4440 588
rect 4504 632 4520 648
rect 4472 592 4504 608
rect 4472 572 4488 588
rect 4472 552 4488 568
rect 4312 512 4328 528
rect 4232 492 4248 508
rect 4200 472 4216 488
rect 4184 452 4200 468
rect 4456 432 4472 448
rect 4232 372 4248 388
rect 4232 352 4248 368
rect 4168 332 4184 348
rect 4280 332 4296 348
rect 4328 332 4344 348
rect 4152 312 4168 328
rect 4120 272 4136 288
rect 4200 272 4216 288
rect 4040 252 4056 268
rect 4136 232 4152 248
rect 4040 212 4056 228
rect 4008 192 4024 208
rect 3992 152 4008 168
rect 4072 152 4088 168
rect 4120 152 4136 168
rect 3976 132 3992 148
rect 4104 132 4120 148
rect 4264 252 4280 268
rect 4168 132 4184 148
rect 4248 132 4264 148
rect 3720 114 3736 128
rect 3720 112 3736 114
rect 4088 112 4104 128
rect 3416 92 3432 108
rect 3448 92 3460 108
rect 3460 92 3464 108
rect 3592 92 3608 108
rect 3464 72 3480 88
rect 3400 52 3416 68
rect 4168 92 4184 108
rect 4312 252 4328 268
rect 4472 412 4488 428
rect 4440 352 4456 368
rect 4408 332 4424 348
rect 4392 272 4408 288
rect 4360 232 4376 248
rect 4360 192 4392 208
rect 4392 132 4408 148
rect 4584 672 4600 688
rect 4536 612 4552 628
rect 4584 552 4600 568
rect 4632 712 4648 728
rect 4808 1212 4824 1228
rect 4696 1192 4712 1208
rect 4680 1032 4696 1048
rect 4760 1132 4776 1148
rect 5144 1392 5160 1408
rect 5016 1332 5032 1348
rect 5128 1332 5144 1348
rect 5032 1312 5048 1328
rect 5144 1312 5160 1328
rect 5000 1292 5016 1308
rect 5080 1292 5096 1308
rect 4856 1272 4872 1288
rect 5000 1272 5016 1288
rect 4840 1172 4856 1188
rect 5144 1292 5160 1308
rect 5112 1232 5128 1248
rect 4909 1202 4945 1218
rect 4808 1112 4824 1128
rect 4856 1092 4872 1108
rect 5064 1172 5080 1188
rect 5128 1152 5144 1168
rect 4984 1132 5000 1148
rect 5080 1132 5096 1148
rect 4968 1072 4984 1088
rect 4776 1052 4792 1068
rect 4840 1052 4856 1068
rect 4936 1052 4952 1068
rect 5016 1052 5032 1068
rect 4904 1032 4920 1048
rect 4712 992 4728 1008
rect 4760 992 4776 1008
rect 4680 792 4696 808
rect 4664 712 4680 728
rect 4760 892 4776 908
rect 4728 812 4744 828
rect 4792 1012 4808 1028
rect 5016 952 5032 968
rect 4776 792 4792 808
rect 4696 732 4712 748
rect 4712 732 4728 748
rect 4664 672 4696 688
rect 4648 652 4664 668
rect 4680 652 4696 668
rect 4664 612 4680 628
rect 4616 532 4632 548
rect 4520 512 4536 528
rect 4760 692 4776 708
rect 4824 872 4840 888
rect 4824 832 4840 848
rect 4808 732 4824 748
rect 4872 932 4888 948
rect 4968 932 4984 948
rect 4920 912 4936 928
rect 4872 892 4888 908
rect 4984 892 5000 908
rect 4909 802 4945 818
rect 4920 712 4936 728
rect 4744 652 4760 668
rect 4840 652 4856 668
rect 4888 652 4904 668
rect 5032 932 5048 948
rect 5064 952 5080 968
rect 5048 892 5064 908
rect 5128 892 5144 908
rect 5112 872 5128 888
rect 5000 792 5016 808
rect 5000 772 5016 788
rect 5064 732 5080 748
rect 5032 712 5048 728
rect 5016 652 5032 668
rect 4984 632 5000 648
rect 4808 592 4824 608
rect 4840 592 4856 608
rect 4712 532 4728 548
rect 4744 534 4760 548
rect 4744 532 4760 534
rect 4776 532 4792 548
rect 4808 532 4824 548
rect 4568 492 4584 508
rect 4552 452 4568 468
rect 4520 432 4536 448
rect 4552 392 4568 408
rect 4632 492 4648 508
rect 4616 472 4632 488
rect 4648 472 4664 488
rect 4680 472 4696 488
rect 4728 452 4744 468
rect 4648 412 4664 428
rect 4632 312 4648 328
rect 4536 272 4552 288
rect 4520 252 4536 268
rect 4680 392 4696 408
rect 4600 272 4616 288
rect 4616 272 4632 288
rect 4712 252 4728 268
rect 4968 612 4984 628
rect 4904 532 4920 548
rect 4808 492 4824 508
rect 4840 432 4856 448
rect 4776 412 4792 428
rect 4840 412 4856 428
rect 4760 392 4792 408
rect 4728 212 4760 228
rect 4904 472 4920 488
rect 4909 402 4945 418
rect 4872 352 4888 368
rect 4904 352 4920 368
rect 4952 352 4968 368
rect 4824 292 4840 308
rect 4920 292 4936 308
rect 5000 552 5016 568
rect 5256 1512 5272 1528
rect 5240 1492 5256 1508
rect 5208 1472 5224 1488
rect 5192 1392 5208 1408
rect 5192 1352 5208 1368
rect 5240 1352 5256 1368
rect 5176 1172 5192 1188
rect 5176 1112 5192 1128
rect 5160 1072 5176 1088
rect 5160 972 5176 988
rect 5176 952 5192 968
rect 5256 1332 5272 1348
rect 5448 2212 5464 2228
rect 5432 2172 5448 2188
rect 5416 2112 5432 2128
rect 5432 2072 5448 2088
rect 5416 1992 5432 2008
rect 5352 1912 5368 1928
rect 5336 1872 5352 1888
rect 5336 1792 5352 1808
rect 5304 1732 5320 1748
rect 5288 1432 5304 1448
rect 5272 1312 5288 1328
rect 5208 1272 5224 1288
rect 5320 1652 5336 1668
rect 5384 1872 5400 1888
rect 5368 1832 5384 1848
rect 5400 1792 5416 1808
rect 5384 1752 5400 1768
rect 5608 2272 5624 2288
rect 5560 2252 5576 2268
rect 5560 2232 5576 2248
rect 5512 2192 5528 2208
rect 5480 2112 5496 2128
rect 5544 1992 5560 2008
rect 5624 2192 5640 2208
rect 5656 2252 5672 2268
rect 5704 2492 5720 2508
rect 5752 2492 5768 2508
rect 5688 2352 5704 2368
rect 5832 2532 5848 2548
rect 5800 2512 5816 2528
rect 5933 2602 5969 2618
rect 5944 2552 5960 2568
rect 5784 2432 5800 2448
rect 5736 2412 5752 2428
rect 5752 2312 5768 2328
rect 5912 2492 5928 2508
rect 5912 2472 5928 2488
rect 5896 2392 5912 2408
rect 5880 2372 5896 2388
rect 6008 2512 6024 2528
rect 5976 2412 5992 2428
rect 5944 2352 5960 2368
rect 5928 2312 5944 2328
rect 5720 2292 5736 2308
rect 5928 2292 5944 2308
rect 5960 2292 5976 2308
rect 5704 2272 5720 2288
rect 5768 2272 5784 2288
rect 5864 2252 5880 2268
rect 5640 2172 5656 2188
rect 5784 2192 5800 2208
rect 5720 2172 5736 2188
rect 5848 2232 5864 2248
rect 5960 2252 5976 2268
rect 5933 2202 5969 2218
rect 6088 2712 6104 2728
rect 6072 2632 6088 2648
rect 6120 2692 6136 2708
rect 6168 2692 6184 2708
rect 6200 2692 6216 2708
rect 6056 2612 6072 2628
rect 6104 2612 6120 2628
rect 6056 2592 6072 2608
rect 6104 2592 6120 2608
rect 6040 2572 6056 2588
rect 6040 2552 6056 2568
rect 6072 2512 6088 2528
rect 6104 2512 6120 2528
rect 6200 2672 6216 2688
rect 6168 2652 6184 2668
rect 6536 3192 6552 3208
rect 6632 3432 6648 3448
rect 6648 3432 6664 3448
rect 6568 3372 6584 3388
rect 6632 3352 6648 3368
rect 6664 3412 6680 3428
rect 6584 3332 6600 3348
rect 6552 3172 6568 3188
rect 6712 3392 6728 3408
rect 6808 3912 6824 3928
rect 6808 3712 6824 3728
rect 6776 3452 6792 3468
rect 6696 3372 6712 3388
rect 6744 3372 6760 3388
rect 6744 3352 6760 3368
rect 6712 3332 6728 3348
rect 6776 3332 6792 3348
rect 6712 3292 6728 3308
rect 6648 3132 6664 3148
rect 6536 3112 6552 3128
rect 6632 3112 6648 3128
rect 6504 3092 6536 3108
rect 6600 3106 6616 3108
rect 6600 3092 6616 3106
rect 6408 3072 6424 3088
rect 6408 3032 6424 3048
rect 6408 3012 6424 3028
rect 6376 2952 6392 2968
rect 6360 2932 6376 2948
rect 6344 2912 6360 2928
rect 6312 2892 6328 2908
rect 6248 2692 6264 2708
rect 6296 2692 6312 2708
rect 6344 2692 6360 2708
rect 6248 2672 6264 2688
rect 6280 2652 6296 2668
rect 6216 2632 6248 2648
rect 6200 2592 6216 2608
rect 6200 2572 6216 2588
rect 6264 2612 6280 2628
rect 6248 2592 6264 2608
rect 6232 2572 6248 2588
rect 6200 2512 6216 2528
rect 6056 2472 6072 2488
rect 6104 2472 6120 2488
rect 6136 2472 6152 2488
rect 6152 2472 6168 2488
rect 6040 2352 6056 2368
rect 6120 2452 6136 2468
rect 6088 2432 6104 2448
rect 6200 2472 6216 2488
rect 6056 2272 6072 2288
rect 6072 2252 6088 2268
rect 6088 2252 6104 2268
rect 6088 2232 6104 2248
rect 6056 2212 6072 2228
rect 6168 2192 6184 2208
rect 6136 2172 6152 2188
rect 6344 2672 6360 2688
rect 6472 2952 6488 2968
rect 6424 2932 6440 2948
rect 6440 2912 6456 2928
rect 6472 2892 6488 2908
rect 6568 3072 6584 3088
rect 6536 3012 6552 3028
rect 6632 3012 6648 3028
rect 6664 2972 6680 2988
rect 6552 2952 6568 2968
rect 6632 2952 6648 2968
rect 6520 2912 6536 2928
rect 6616 2912 6632 2928
rect 6520 2892 6536 2908
rect 6472 2872 6488 2888
rect 6504 2872 6520 2888
rect 6408 2792 6424 2808
rect 6424 2732 6440 2748
rect 6392 2706 6408 2708
rect 6392 2692 6408 2706
rect 6360 2652 6376 2668
rect 6328 2552 6344 2568
rect 6328 2512 6344 2528
rect 6296 2472 6312 2488
rect 6280 2432 6296 2448
rect 6392 2612 6408 2628
rect 6600 2892 6616 2908
rect 6552 2832 6568 2848
rect 6536 2712 6552 2728
rect 6488 2692 6504 2708
rect 6456 2672 6472 2688
rect 6504 2672 6520 2688
rect 6488 2572 6504 2588
rect 6520 2572 6536 2588
rect 6472 2552 6488 2568
rect 6536 2552 6552 2568
rect 6456 2532 6472 2548
rect 6392 2512 6408 2528
rect 6440 2492 6456 2508
rect 6440 2472 6456 2488
rect 6424 2432 6440 2448
rect 6376 2412 6392 2428
rect 6264 2292 6280 2308
rect 6232 2232 6248 2248
rect 6296 2232 6312 2248
rect 6264 2192 6280 2208
rect 5640 2132 5656 2148
rect 5816 2132 5832 2148
rect 5928 2132 5944 2148
rect 5976 2132 5992 2148
rect 6024 2132 6040 2148
rect 5592 2114 5608 2128
rect 5592 2112 5608 2114
rect 5496 1892 5512 1908
rect 5560 1892 5576 1908
rect 5656 2012 5672 2028
rect 5880 2092 5896 2108
rect 6232 2152 6248 2168
rect 6056 2132 6072 2148
rect 6104 2132 6120 2148
rect 6072 2112 6088 2128
rect 5816 2072 5832 2088
rect 5912 2072 5928 2088
rect 5992 2072 6008 2088
rect 6024 2072 6040 2088
rect 5768 2032 5784 2048
rect 5688 1992 5704 2008
rect 5704 1972 5720 1988
rect 5864 1972 5880 1988
rect 5464 1852 5480 1868
rect 5496 1832 5512 1848
rect 5448 1792 5464 1808
rect 5464 1772 5480 1788
rect 5480 1752 5496 1768
rect 5512 1752 5528 1768
rect 5608 1752 5624 1768
rect 5720 1932 5736 1948
rect 5736 1892 5752 1908
rect 5752 1892 5768 1908
rect 5800 1892 5816 1908
rect 5656 1772 5672 1788
rect 5704 1812 5720 1828
rect 5416 1732 5432 1748
rect 5496 1712 5512 1728
rect 5528 1712 5544 1728
rect 5624 1732 5640 1748
rect 5688 1732 5704 1748
rect 5416 1672 5432 1688
rect 5400 1652 5416 1668
rect 5352 1632 5384 1648
rect 5352 1512 5368 1528
rect 5448 1612 5464 1628
rect 5544 1672 5560 1688
rect 5624 1572 5640 1588
rect 5608 1532 5624 1548
rect 5448 1512 5464 1528
rect 5464 1512 5480 1528
rect 5512 1512 5516 1528
rect 5516 1512 5528 1528
rect 5304 1272 5320 1288
rect 5416 1472 5432 1488
rect 5464 1472 5480 1488
rect 5384 1452 5400 1468
rect 5368 1412 5384 1428
rect 5416 1392 5432 1408
rect 5352 1372 5368 1388
rect 5336 1312 5352 1328
rect 5208 1232 5224 1248
rect 5240 1232 5272 1248
rect 5320 1232 5336 1248
rect 5240 1192 5256 1208
rect 5208 932 5224 948
rect 5304 1112 5320 1128
rect 5304 1072 5320 1088
rect 5192 812 5208 828
rect 5080 712 5096 728
rect 5144 712 5176 728
rect 5240 912 5256 928
rect 5256 872 5272 888
rect 5256 812 5272 828
rect 5368 1232 5384 1248
rect 5656 1692 5672 1708
rect 5784 1852 5800 1868
rect 5800 1832 5816 1848
rect 5880 1932 5896 1948
rect 5848 1872 5864 1888
rect 5832 1812 5848 1828
rect 5720 1772 5736 1788
rect 5832 1772 5848 1788
rect 5768 1752 5784 1768
rect 5864 1752 5880 1768
rect 5800 1732 5816 1748
rect 5816 1732 5832 1748
rect 5864 1732 5880 1748
rect 5688 1552 5704 1568
rect 5656 1512 5672 1528
rect 5592 1472 5608 1488
rect 5640 1472 5656 1488
rect 5528 1432 5544 1448
rect 5480 1392 5496 1408
rect 5528 1372 5544 1388
rect 5576 1372 5592 1388
rect 5480 1352 5496 1368
rect 5528 1352 5544 1368
rect 5496 1332 5512 1348
rect 5448 1312 5464 1328
rect 5480 1292 5496 1308
rect 5480 1152 5496 1168
rect 5400 1132 5416 1148
rect 5448 1132 5464 1148
rect 5384 1112 5400 1128
rect 5368 1052 5384 1068
rect 5352 1012 5368 1028
rect 5336 992 5352 1008
rect 5320 972 5336 988
rect 5304 952 5320 968
rect 5352 972 5368 988
rect 5368 912 5384 928
rect 5400 912 5416 928
rect 5288 892 5304 908
rect 5320 852 5336 868
rect 5272 772 5288 788
rect 5272 732 5288 748
rect 5304 732 5320 748
rect 5224 692 5240 708
rect 5256 692 5272 708
rect 5288 692 5304 708
rect 5208 672 5224 688
rect 5224 672 5240 688
rect 5144 612 5160 628
rect 5144 592 5160 608
rect 5192 552 5208 568
rect 5240 652 5256 668
rect 5224 632 5240 648
rect 5240 552 5256 568
rect 5048 532 5064 548
rect 5064 532 5080 548
rect 5096 532 5112 548
rect 5112 532 5128 548
rect 5208 532 5224 548
rect 5032 512 5048 528
rect 5080 512 5096 528
rect 5000 472 5016 488
rect 4984 352 5000 368
rect 5176 512 5192 528
rect 5144 452 5160 468
rect 5128 392 5144 408
rect 5192 392 5208 408
rect 5032 352 5048 368
rect 5128 352 5144 368
rect 5048 292 5064 308
rect 5080 292 5096 308
rect 4888 272 4904 288
rect 4952 272 4968 288
rect 4968 272 4984 288
rect 4808 212 4824 228
rect 4664 192 4680 208
rect 4760 192 4776 208
rect 4584 152 4600 168
rect 4632 152 4648 168
rect 4856 172 4872 188
rect 4696 132 4712 148
rect 4824 132 4840 148
rect 4472 112 4488 128
rect 4296 32 4312 48
rect 3944 12 3960 28
rect 3976 12 3992 28
rect 4472 92 4488 108
rect 4456 32 4472 48
rect 4568 92 4584 108
rect 4920 252 4936 268
rect 5128 252 5144 268
rect 5000 172 5016 188
rect 4968 152 4984 168
rect 5096 232 5112 248
rect 5160 232 5176 248
rect 5160 212 5176 228
rect 5368 892 5384 908
rect 5336 752 5352 768
rect 5400 752 5416 768
rect 5432 892 5448 908
rect 5416 712 5432 728
rect 5336 692 5352 708
rect 5336 672 5352 688
rect 5400 652 5416 668
rect 5640 1412 5656 1428
rect 5688 1392 5704 1408
rect 5608 1372 5624 1388
rect 5736 1692 5752 1708
rect 5848 1712 5864 1728
rect 5832 1672 5848 1688
rect 5800 1652 5816 1668
rect 5896 1692 5912 1708
rect 5880 1632 5896 1648
rect 5848 1552 5864 1568
rect 5848 1532 5864 1548
rect 5752 1512 5784 1528
rect 5800 1512 5816 1528
rect 5864 1512 5880 1528
rect 6008 1972 6024 1988
rect 5928 1952 5944 1968
rect 5976 1892 5992 1908
rect 6120 2112 6136 2128
rect 6136 2092 6152 2108
rect 6088 2052 6104 2068
rect 6088 1972 6104 1988
rect 6088 1952 6104 1968
rect 6088 1932 6104 1948
rect 6024 1912 6040 1928
rect 6072 1912 6088 1928
rect 6040 1892 6056 1908
rect 5992 1872 6008 1888
rect 5928 1852 5944 1868
rect 5933 1802 5969 1818
rect 6008 1772 6024 1788
rect 5928 1712 5944 1728
rect 5912 1592 5928 1608
rect 5912 1572 5928 1588
rect 5848 1492 5864 1508
rect 5736 1472 5752 1488
rect 5800 1472 5816 1488
rect 5816 1432 5832 1448
rect 5768 1392 5784 1408
rect 5704 1352 5736 1368
rect 5576 1312 5592 1328
rect 5528 1292 5544 1308
rect 5576 1292 5592 1308
rect 5784 1372 5800 1388
rect 5656 1292 5672 1308
rect 5688 1292 5704 1308
rect 5832 1292 5848 1308
rect 5592 1252 5608 1268
rect 5624 1232 5640 1248
rect 5544 1132 5560 1148
rect 5592 1132 5608 1148
rect 5656 1132 5672 1148
rect 5672 1112 5688 1128
rect 5528 1072 5544 1088
rect 5512 992 5528 1008
rect 5496 972 5512 988
rect 5528 972 5544 988
rect 5576 972 5592 988
rect 5496 952 5512 968
rect 5512 952 5528 968
rect 5576 952 5592 968
rect 5656 1072 5672 1088
rect 5752 1232 5768 1248
rect 5848 1152 5864 1168
rect 5768 1132 5784 1148
rect 5800 1132 5816 1148
rect 5896 1372 5912 1388
rect 5944 1672 5960 1688
rect 6168 1932 6184 1948
rect 6152 1912 6168 1928
rect 6152 1892 6168 1908
rect 6120 1872 6136 1888
rect 6504 2532 6520 2548
rect 6488 2512 6504 2528
rect 6632 2772 6648 2788
rect 6632 2732 6648 2748
rect 6600 2692 6616 2708
rect 6632 2692 6648 2708
rect 6648 2672 6664 2688
rect 6680 2892 6696 2908
rect 6696 2752 6712 2768
rect 6696 2712 6712 2728
rect 6744 3032 6760 3048
rect 6728 2952 6744 2968
rect 6776 2952 6792 2968
rect 6808 2912 6824 2928
rect 6712 2692 6728 2708
rect 6680 2652 6696 2668
rect 6728 2652 6744 2668
rect 6664 2552 6680 2568
rect 6712 2552 6728 2568
rect 6696 2532 6712 2548
rect 6632 2512 6648 2528
rect 6664 2512 6680 2528
rect 6712 2512 6728 2528
rect 6504 2372 6520 2388
rect 6472 2332 6488 2348
rect 6472 2292 6488 2308
rect 6392 2272 6408 2288
rect 6376 2212 6392 2228
rect 6344 2172 6360 2188
rect 6344 2132 6360 2148
rect 6280 2112 6296 2128
rect 6184 1852 6200 1868
rect 6104 1832 6120 1848
rect 6088 1812 6104 1828
rect 6120 1792 6136 1808
rect 6104 1752 6120 1768
rect 6056 1732 6088 1748
rect 6040 1712 6056 1728
rect 6040 1692 6056 1708
rect 6024 1672 6040 1688
rect 6008 1572 6024 1588
rect 6024 1552 6056 1568
rect 5960 1472 5976 1488
rect 5928 1452 5944 1468
rect 5933 1402 5969 1418
rect 6008 1372 6024 1388
rect 5928 1352 5944 1368
rect 6024 1332 6040 1348
rect 6168 1692 6184 1708
rect 6152 1652 6168 1668
rect 6312 2112 6328 2128
rect 6296 2092 6312 2108
rect 6344 2072 6360 2088
rect 6232 1992 6248 2008
rect 6248 1892 6264 1908
rect 6424 2152 6440 2168
rect 6424 2132 6440 2148
rect 6424 2112 6440 2128
rect 6408 2092 6424 2108
rect 6392 1912 6408 1928
rect 6424 1912 6440 1928
rect 6408 1852 6424 1868
rect 6376 1812 6392 1828
rect 6488 2252 6504 2268
rect 6680 2492 6696 2508
rect 6632 2412 6648 2428
rect 6600 2372 6616 2388
rect 6568 2352 6584 2368
rect 6568 2332 6584 2348
rect 6520 2292 6536 2308
rect 6552 2292 6568 2308
rect 6584 2292 6600 2308
rect 6456 2132 6472 2148
rect 6472 2052 6488 2068
rect 6504 1952 6520 1968
rect 6504 1932 6520 1948
rect 6712 2392 6728 2408
rect 6664 2306 6680 2308
rect 6664 2292 6680 2306
rect 6536 2272 6552 2288
rect 6552 2252 6568 2268
rect 6536 2192 6552 2208
rect 6552 2172 6568 2188
rect 6600 2152 6616 2168
rect 6616 2112 6632 2128
rect 6552 2092 6568 2108
rect 6520 1912 6536 1928
rect 6648 2212 6664 2228
rect 6632 1992 6648 2008
rect 6664 2152 6680 2168
rect 6680 2132 6696 2148
rect 6696 2132 6712 2148
rect 6696 1932 6712 1948
rect 6712 1912 6728 1928
rect 6456 1892 6472 1908
rect 6600 1892 6616 1908
rect 6600 1872 6616 1888
rect 6536 1852 6552 1868
rect 6472 1832 6488 1848
rect 6456 1792 6472 1808
rect 6360 1752 6376 1768
rect 6440 1752 6456 1768
rect 6680 1892 6696 1908
rect 6744 2372 6760 2388
rect 6792 2532 6808 2548
rect 6776 2272 6792 2288
rect 6760 2212 6776 2228
rect 6744 2132 6760 2148
rect 6792 2052 6808 2068
rect 6648 1872 6664 1888
rect 6712 1872 6744 1888
rect 6616 1832 6648 1848
rect 6696 1832 6712 1848
rect 6584 1812 6600 1828
rect 6664 1792 6680 1808
rect 6328 1732 6344 1748
rect 6440 1732 6456 1748
rect 6568 1732 6584 1748
rect 6616 1732 6632 1748
rect 6408 1712 6424 1728
rect 6248 1672 6264 1688
rect 6168 1592 6184 1608
rect 6200 1592 6216 1608
rect 6104 1512 6120 1528
rect 6136 1512 6152 1528
rect 6072 1492 6088 1508
rect 6632 1712 6648 1728
rect 6488 1652 6504 1668
rect 6600 1652 6616 1668
rect 6312 1572 6328 1588
rect 6424 1572 6440 1588
rect 6472 1572 6488 1588
rect 6232 1532 6248 1548
rect 6184 1512 6200 1528
rect 6200 1512 6216 1528
rect 6216 1492 6232 1508
rect 6120 1432 6136 1448
rect 6264 1512 6280 1528
rect 6280 1492 6296 1508
rect 6408 1552 6424 1568
rect 6424 1512 6440 1528
rect 6296 1472 6312 1488
rect 6184 1432 6200 1448
rect 6248 1432 6264 1448
rect 6216 1412 6232 1428
rect 6168 1392 6184 1408
rect 6104 1372 6120 1388
rect 6168 1372 6184 1388
rect 6152 1352 6168 1368
rect 6136 1332 6152 1348
rect 5896 1292 5928 1308
rect 5928 1212 5944 1228
rect 5928 1172 5944 1188
rect 5736 1112 5752 1128
rect 5864 1112 5880 1128
rect 5880 1092 5896 1108
rect 5752 1072 5768 1088
rect 5784 1072 5800 1088
rect 5720 1052 5736 1068
rect 5704 992 5720 1008
rect 5688 932 5704 948
rect 5544 912 5560 928
rect 5624 912 5640 928
rect 5640 912 5656 928
rect 5688 912 5704 928
rect 5464 792 5480 808
rect 5528 752 5544 768
rect 5528 732 5544 748
rect 5272 632 5288 648
rect 5352 632 5368 648
rect 5336 592 5352 608
rect 5384 612 5400 628
rect 5512 652 5528 668
rect 5464 632 5480 648
rect 5384 572 5400 588
rect 5256 492 5272 508
rect 5304 392 5320 408
rect 5208 352 5224 368
rect 5240 352 5256 368
rect 5288 312 5304 328
rect 5192 212 5208 228
rect 5256 212 5272 228
rect 5192 192 5208 208
rect 5240 192 5256 208
rect 5432 512 5448 528
rect 5416 472 5432 488
rect 5384 352 5416 368
rect 5288 172 5304 188
rect 5112 152 5128 168
rect 5320 252 5336 268
rect 5368 232 5384 248
rect 5336 212 5352 228
rect 5384 212 5400 228
rect 5352 192 5368 208
rect 5384 192 5400 208
rect 5320 152 5336 168
rect 4824 112 4840 128
rect 4952 112 4968 128
rect 5096 112 5112 128
rect 5304 112 5320 128
rect 5448 372 5464 388
rect 5512 572 5528 588
rect 5528 552 5544 568
rect 5560 852 5576 868
rect 5576 732 5592 748
rect 5576 652 5592 668
rect 5624 892 5640 908
rect 5656 892 5672 908
rect 5624 872 5640 888
rect 5608 712 5624 728
rect 5640 832 5656 848
rect 5592 632 5608 648
rect 5608 612 5624 628
rect 5640 672 5656 688
rect 5688 812 5704 828
rect 5688 712 5704 728
rect 5832 1072 5848 1088
rect 5880 1052 5896 1068
rect 6072 1312 6088 1328
rect 6152 1312 6168 1328
rect 6072 1252 6088 1268
rect 6120 1252 6136 1268
rect 6056 1092 6072 1108
rect 6024 1072 6040 1088
rect 5800 1032 5832 1048
rect 5848 1012 5864 1028
rect 5736 912 5752 928
rect 5720 892 5736 908
rect 5752 852 5768 868
rect 5848 892 5864 908
rect 5848 872 5864 888
rect 5816 752 5832 768
rect 5752 732 5768 748
rect 5784 712 5800 728
rect 5736 692 5752 708
rect 5672 652 5688 668
rect 5656 592 5672 608
rect 5624 572 5640 588
rect 5688 632 5704 648
rect 5656 532 5672 548
rect 5768 652 5784 668
rect 5768 632 5784 648
rect 5816 632 5832 648
rect 5528 492 5544 508
rect 5480 472 5496 488
rect 5528 452 5544 468
rect 5480 412 5496 428
rect 5640 512 5656 528
rect 5688 512 5704 528
rect 5784 512 5800 528
rect 5576 492 5592 508
rect 5656 492 5672 508
rect 5688 492 5704 508
rect 5752 492 5768 508
rect 5800 492 5816 508
rect 5704 472 5720 488
rect 5736 472 5752 488
rect 5592 452 5608 468
rect 5576 432 5592 448
rect 5528 392 5560 408
rect 5512 312 5528 328
rect 5432 192 5448 208
rect 5464 252 5480 268
rect 5464 212 5480 228
rect 5512 192 5528 208
rect 5896 912 5912 928
rect 5896 892 5912 908
rect 5976 1032 5992 1048
rect 5933 1002 5969 1018
rect 5944 952 5960 968
rect 6008 952 6024 968
rect 5928 932 5944 948
rect 5944 932 5960 948
rect 5976 944 5992 948
rect 5976 932 5992 944
rect 5912 812 5928 828
rect 5912 772 5928 788
rect 6008 872 6024 888
rect 6056 1012 6072 1028
rect 6040 992 6056 1008
rect 6200 1272 6216 1288
rect 6168 1192 6200 1208
rect 6568 1492 6584 1508
rect 6520 1472 6536 1488
rect 6696 1472 6712 1488
rect 6376 1452 6392 1468
rect 6456 1452 6472 1468
rect 6344 1392 6360 1408
rect 6328 1332 6344 1348
rect 6280 1312 6296 1328
rect 6296 1312 6312 1328
rect 6248 1292 6264 1308
rect 6504 1392 6520 1408
rect 6472 1352 6488 1368
rect 6392 1332 6408 1348
rect 6440 1332 6456 1348
rect 6520 1332 6536 1348
rect 6248 1272 6264 1288
rect 6360 1212 6376 1228
rect 6216 1152 6232 1168
rect 6264 1152 6280 1168
rect 6200 1132 6216 1148
rect 6232 1132 6248 1148
rect 6216 1112 6232 1128
rect 6328 1112 6344 1128
rect 6280 1092 6296 1108
rect 6200 1052 6216 1068
rect 6248 1052 6264 1068
rect 6248 1012 6264 1028
rect 6264 992 6280 1008
rect 6104 912 6120 928
rect 6136 912 6152 928
rect 6184 912 6200 928
rect 6232 912 6248 928
rect 6072 892 6088 908
rect 5896 672 5912 688
rect 5896 652 5912 668
rect 5880 632 5896 648
rect 5912 592 5928 608
rect 5933 602 5969 618
rect 5992 572 6008 588
rect 5672 412 5688 428
rect 5816 412 5832 428
rect 5768 352 5784 368
rect 5736 332 5752 348
rect 5576 312 5592 328
rect 5624 312 5640 328
rect 5688 312 5704 328
rect 5640 292 5656 308
rect 5576 272 5592 288
rect 5704 272 5720 288
rect 5816 272 5832 288
rect 5608 252 5624 268
rect 5688 252 5704 268
rect 6056 852 6072 868
rect 6200 872 6216 888
rect 6264 832 6280 848
rect 6264 812 6280 828
rect 6136 792 6152 808
rect 6104 772 6120 788
rect 6168 752 6184 768
rect 6040 732 6056 748
rect 6024 692 6040 708
rect 6136 712 6152 728
rect 6120 692 6136 708
rect 6184 672 6200 688
rect 6248 672 6264 688
rect 6232 552 6248 568
rect 6344 1092 6360 1108
rect 6328 1072 6344 1088
rect 6312 1052 6328 1068
rect 6312 952 6328 968
rect 6328 932 6344 948
rect 6296 912 6312 928
rect 6328 852 6344 868
rect 6312 772 6328 788
rect 6296 732 6312 748
rect 6296 672 6312 688
rect 6328 652 6344 668
rect 6296 572 6312 588
rect 6008 532 6024 548
rect 6136 532 6152 548
rect 6168 532 6184 548
rect 6216 532 6232 548
rect 6248 532 6264 548
rect 6280 532 6296 548
rect 5992 512 6008 528
rect 6008 492 6024 508
rect 5880 472 5896 488
rect 5864 432 5880 448
rect 5848 372 5864 388
rect 6312 552 6328 568
rect 6280 492 6296 508
rect 6248 472 6264 488
rect 6232 432 6248 448
rect 6136 392 6152 408
rect 6088 372 6104 388
rect 5864 352 5880 368
rect 6024 352 6040 368
rect 5832 252 5848 268
rect 5768 152 5784 168
rect 5832 152 5848 168
rect 6024 332 6040 348
rect 5896 292 5912 308
rect 5560 132 5576 148
rect 5624 132 5640 148
rect 5624 112 5640 128
rect 5704 112 5720 128
rect 5800 114 5816 128
rect 5800 112 5816 114
rect 6168 332 6184 348
rect 6328 412 6344 428
rect 6312 312 6328 328
rect 6104 292 6120 308
rect 6152 292 6168 308
rect 6184 292 6200 308
rect 5992 272 6008 288
rect 6136 272 6152 288
rect 6152 252 6168 268
rect 5944 232 5960 248
rect 6024 232 6040 248
rect 5933 202 5969 218
rect 5944 172 5960 188
rect 5928 152 5944 168
rect 6056 132 6072 148
rect 6488 1312 6504 1328
rect 6552 1312 6568 1328
rect 6456 1292 6472 1308
rect 6424 1252 6440 1268
rect 6552 1272 6568 1288
rect 6488 1172 6504 1188
rect 6552 1172 6568 1188
rect 6488 1152 6504 1168
rect 6472 1132 6488 1148
rect 6392 1112 6408 1128
rect 6440 1112 6456 1128
rect 6696 1452 6712 1468
rect 6616 1372 6632 1388
rect 6744 1852 6760 1868
rect 6760 1812 6776 1828
rect 6744 1532 6760 1548
rect 6760 1492 6776 1508
rect 6728 1452 6744 1468
rect 6728 1352 6744 1368
rect 6584 1332 6600 1348
rect 6632 1332 6648 1348
rect 6600 1312 6616 1328
rect 6648 1312 6664 1328
rect 6680 1292 6696 1308
rect 6600 1252 6616 1268
rect 6712 1332 6728 1348
rect 6696 1172 6712 1188
rect 6568 1092 6584 1108
rect 6632 1092 6648 1108
rect 6456 1072 6472 1088
rect 6536 1072 6552 1088
rect 6376 1032 6392 1048
rect 6456 1032 6472 1048
rect 6408 972 6424 988
rect 6376 952 6392 968
rect 6424 932 6440 948
rect 6360 912 6376 928
rect 6424 912 6440 928
rect 6472 932 6488 948
rect 6408 892 6424 908
rect 6456 892 6472 908
rect 6472 872 6488 888
rect 6632 972 6648 988
rect 6600 952 6616 968
rect 6552 932 6568 948
rect 6584 932 6600 948
rect 6520 912 6536 928
rect 6584 912 6600 928
rect 6520 892 6536 908
rect 6536 872 6552 888
rect 6488 852 6504 868
rect 6520 852 6536 868
rect 6440 732 6456 748
rect 6504 732 6520 748
rect 6408 712 6424 728
rect 6376 692 6392 708
rect 6392 672 6408 688
rect 6424 632 6440 648
rect 6504 632 6520 648
rect 6472 552 6488 568
rect 6360 532 6376 548
rect 6504 532 6520 548
rect 6376 512 6392 528
rect 6360 492 6376 508
rect 6264 272 6280 288
rect 4760 92 4776 108
rect 4840 92 4844 108
rect 4844 92 4856 108
rect 4984 92 5000 108
rect 5320 92 5336 108
rect 5400 92 5432 108
rect 5592 92 5608 108
rect 5624 92 5640 108
rect 5672 92 5688 108
rect 5912 92 5928 108
rect 5960 92 5976 108
rect 4909 2 4945 18
rect 5944 12 5960 28
rect 6072 92 6088 108
rect 6024 12 6040 28
rect 6056 12 6072 28
rect 6184 132 6200 148
rect 6168 112 6184 128
rect 6200 112 6216 128
rect 6456 492 6472 508
rect 6440 292 6456 308
rect 6424 232 6440 248
rect 6440 172 6456 188
rect 6504 132 6520 148
rect 6552 832 6568 848
rect 6600 832 6616 848
rect 6568 712 6584 728
rect 6680 932 6696 948
rect 6648 712 6664 728
rect 6696 712 6712 728
rect 6744 1312 6760 1328
rect 6776 1292 6792 1308
rect 6760 1152 6776 1168
rect 6776 872 6792 888
rect 6808 872 6824 888
rect 6712 692 6728 708
rect 6616 672 6632 688
rect 6568 632 6584 648
rect 6616 632 6632 648
rect 6568 552 6584 568
rect 6632 572 6648 588
rect 6664 672 6680 688
rect 6696 672 6712 688
rect 6648 492 6664 508
rect 6728 572 6744 588
rect 6712 412 6728 428
rect 6584 352 6600 368
rect 6552 292 6568 308
rect 6680 332 6696 348
rect 6696 272 6712 288
rect 6344 112 6360 128
rect 6632 172 6648 188
rect 6760 392 6776 408
rect 6744 352 6760 368
rect 6744 312 6760 328
rect 6728 292 6744 308
rect 6808 552 6824 568
rect 6776 272 6792 288
rect 6664 112 6696 128
<< metal3 >>
rect 200 4817 216 4823
rect 376 4817 392 4823
rect 6600 4817 6616 4823
rect 808 4777 840 4783
rect 3752 4777 5176 4783
rect 5192 4777 5224 4783
rect 5240 4777 5624 4783
rect 3880 4757 4024 4763
rect 1128 4737 1160 4743
rect 2744 4737 2776 4743
rect 4056 4737 4296 4743
rect 4856 4737 4904 4743
rect 4920 4737 4984 4743
rect 6296 4737 6392 4743
rect -51 4717 8 4723
rect 2184 4717 2232 4723
rect 3352 4717 3512 4723
rect 3560 4717 3608 4723
rect 3672 4717 3688 4723
rect 4328 4717 4376 4723
rect 4968 4717 5336 4723
rect 152 4697 168 4703
rect 184 4697 248 4703
rect 264 4697 424 4703
rect 440 4697 632 4703
rect 648 4697 936 4703
rect 1160 4697 1256 4703
rect 1336 4697 1464 4703
rect 2232 4697 2360 4703
rect 2376 4697 2504 4703
rect 2776 4697 2904 4703
rect 3240 4697 3288 4703
rect 3416 4697 3720 4703
rect 4040 4697 4120 4703
rect 4184 4697 4344 4703
rect 4600 4697 4712 4703
rect 4808 4697 4936 4703
rect 4984 4697 5064 4703
rect 5144 4697 5512 4703
rect 5528 4697 5736 4703
rect 5912 4697 6152 4703
rect 6584 4697 6680 4703
rect 552 4677 584 4683
rect 904 4677 920 4683
rect 968 4677 984 4683
rect 1672 4677 1880 4683
rect 1896 4677 2200 4683
rect 2216 4677 2392 4683
rect 2408 4677 2472 4683
rect 2488 4677 2632 4683
rect 2648 4677 2968 4683
rect 2984 4677 3256 4683
rect 3272 4677 3480 4683
rect 3496 4677 3576 4683
rect 3592 4677 3672 4683
rect 4152 4677 4312 4683
rect 4456 4677 4696 4683
rect 4712 4677 4840 4683
rect 5160 4677 5208 4683
rect 5224 4677 5304 4683
rect 5320 4677 5512 4683
rect 5528 4677 5640 4683
rect 5816 4677 6120 4683
rect 120 4657 136 4663
rect 1320 4657 1384 4663
rect 1400 4657 1432 4663
rect 1512 4657 1720 4663
rect 1736 4657 2264 4663
rect 2456 4657 3368 4663
rect 3736 4657 3896 4663
rect 3912 4657 4184 4663
rect 4200 4657 4616 4663
rect 4632 4657 4664 4663
rect 4680 4657 5048 4663
rect 5656 4657 5928 4663
rect 1416 4637 1560 4643
rect 1848 4637 1992 4643
rect 2584 4637 2712 4643
rect 2824 4637 3016 4643
rect 4264 4637 4568 4643
rect 4584 4637 4648 4643
rect 4717 4637 4808 4643
rect 1080 4617 1592 4623
rect 1608 4617 1752 4623
rect 1192 4597 1384 4603
rect 2760 4617 2936 4623
rect 3112 4617 3240 4623
rect 2248 4597 2792 4603
rect 3432 4597 3832 4603
rect 4120 4617 4280 4623
rect 4296 4617 4552 4623
rect 4717 4623 4723 4637
rect 4824 4637 4872 4643
rect 5352 4637 5528 4643
rect 5544 4637 6248 4643
rect 4568 4617 4723 4623
rect 4792 4617 5064 4623
rect 5192 4617 5240 4623
rect 5256 4617 5544 4623
rect 4440 4597 4456 4603
rect 4472 4597 4696 4603
rect 4712 4597 4856 4603
rect 4904 4597 5240 4603
rect 584 4577 632 4583
rect 760 4577 936 4583
rect 1144 4577 1240 4583
rect 1528 4577 1592 4583
rect 1992 4577 2216 4583
rect 2296 4577 2648 4583
rect 2856 4577 3096 4583
rect 3656 4577 3880 4583
rect 4008 4577 4024 4583
rect 4344 4577 4584 4583
rect 4760 4577 4776 4583
rect 4824 4577 4888 4583
rect 5368 4577 5384 4583
rect 6024 4577 6040 4583
rect 6504 4577 6584 4583
rect 1144 4557 1272 4563
rect 1304 4557 2584 4563
rect 2077 4548 2083 4557
rect 3000 4557 3432 4563
rect 3880 4557 4104 4563
rect 4264 4557 4296 4563
rect 4424 4557 4456 4563
rect 4696 4557 4712 4563
rect 4760 4557 4968 4563
rect 5448 4557 5480 4563
rect 5576 4557 5640 4563
rect 5928 4557 5992 4563
rect 3565 4548 3571 4552
rect 472 4537 696 4543
rect 712 4537 1000 4543
rect 1112 4537 1288 4543
rect 1400 4537 1608 4543
rect 1704 4537 1784 4543
rect 1848 4537 1859 4543
rect 2104 4537 2136 4543
rect 2296 4537 2472 4543
rect 2632 4537 2680 4543
rect 2840 4537 2872 4543
rect 3112 4537 3496 4543
rect 3912 4537 4136 4543
rect 4264 4537 4280 4543
rect 4296 4537 4392 4543
rect 4632 4537 4984 4543
rect 5160 4537 5272 4543
rect 5464 4537 5880 4543
rect 5896 4537 5944 4543
rect -51 4517 8 4523
rect 280 4517 360 4523
rect 440 4517 968 4523
rect 984 4517 1048 4523
rect 1144 4517 1320 4523
rect 1336 4517 2152 4523
rect 2408 4517 2536 4523
rect 2557 4517 2563 4532
rect 2760 4517 2776 4523
rect 2808 4517 2824 4523
rect 2840 4517 3000 4523
rect 3144 4517 3160 4523
rect 3224 4517 3416 4523
rect 3432 4517 3480 4523
rect 3512 4517 3560 4523
rect 3592 4517 3736 4523
rect 3880 4517 3896 4523
rect 4008 4517 4200 4523
rect 4216 4517 4616 4523
rect 4984 4517 5000 4523
rect 5128 4517 5160 4523
rect 5208 4517 5368 4523
rect 5720 4517 5768 4523
rect 5832 4517 6008 4523
rect 6392 4517 6504 4523
rect 1069 4508 1075 4512
rect 1128 4497 1144 4503
rect 1160 4497 1272 4503
rect 1592 4497 1720 4503
rect 1928 4497 2488 4503
rect 2504 4497 2776 4503
rect 2792 4497 2904 4503
rect 2920 4497 2968 4503
rect 2984 4497 3080 4503
rect 3096 4497 3144 4503
rect 3208 4497 3320 4503
rect 3480 4497 3512 4503
rect 3624 4497 3768 4503
rect 3784 4497 3816 4503
rect 3832 4497 3928 4503
rect 4088 4497 4216 4503
rect 4232 4497 4264 4503
rect 4392 4497 4424 4503
rect 4472 4497 4536 4503
rect 4744 4497 4792 4503
rect 4856 4497 5144 4503
rect 5496 4497 5768 4503
rect 6056 4497 6088 4503
rect 6360 4497 6456 4503
rect 6472 4497 6648 4503
rect 248 4477 296 4483
rect 600 4477 760 4483
rect 776 4477 1096 4483
rect 1192 4477 1240 4483
rect 1464 4477 1896 4483
rect 2008 4477 2040 4483
rect 2072 4477 2104 4483
rect 2184 4477 3032 4483
rect 3048 4477 3112 4483
rect 3336 4477 4008 4483
rect 4024 4477 4200 4483
rect 4216 4477 5032 4483
rect 5048 4477 5224 4483
rect 5240 4477 5288 4483
rect 5304 4477 5464 4483
rect 5672 4477 5832 4483
rect 6008 4477 6136 4483
rect 472 4457 1816 4463
rect 1976 4457 2520 4463
rect 2536 4457 2728 4463
rect 2808 4457 3384 4463
rect 3400 4457 3448 4463
rect 3720 4457 3752 4463
rect 3784 4457 4024 4463
rect 4040 4457 4168 4463
rect 4184 4457 4232 4463
rect 4728 4457 4808 4463
rect 4872 4457 5080 4463
rect 5096 4457 5256 4463
rect 5272 4457 5320 4463
rect 5432 4457 5816 4463
rect 5848 4457 6056 4463
rect 1064 4437 1640 4443
rect 1656 4437 1752 4443
rect 1912 4437 2120 4443
rect 2136 4437 2184 4443
rect 2280 4437 2936 4443
rect 2952 4437 3048 4443
rect 3256 4437 3544 4443
rect 3560 4437 3672 4443
rect 3960 4437 4024 4443
rect 4072 4437 4120 4443
rect 4248 4437 4392 4443
rect 4408 4437 4488 4443
rect 4504 4437 4632 4443
rect 4680 4437 4696 4443
rect 4792 4437 5016 4443
rect 5112 4437 5192 4443
rect 5544 4437 5896 4443
rect 1112 4417 1224 4423
rect 1272 4417 1352 4423
rect 1432 4417 1576 4423
rect 1720 4417 1896 4423
rect 1912 4417 2024 4423
rect 2152 4417 2264 4423
rect 2744 4417 2824 4423
rect 1096 4397 1560 4403
rect 2040 4397 2568 4403
rect 3032 4417 3112 4423
rect 3128 4417 3304 4423
rect 3352 4417 3656 4423
rect 4360 4417 4376 4423
rect 4408 4417 4776 4423
rect 2952 4397 3448 4403
rect 3464 4397 3800 4403
rect 3816 4397 4520 4403
rect 4536 4397 4840 4403
rect 5416 4417 6168 4423
rect 5096 4397 5160 4403
rect 5512 4397 5864 4403
rect 5880 4397 6120 4403
rect 680 4377 856 4383
rect 1048 4377 1128 4383
rect 1240 4377 1464 4383
rect 1672 4377 1736 4383
rect 2008 4377 2248 4383
rect 2264 4377 2280 4383
rect 2616 4377 2712 4383
rect 2728 4377 2872 4383
rect 2888 4377 3096 4383
rect 3112 4377 3208 4383
rect 3688 4377 3896 4383
rect 4168 4377 5528 4383
rect 5608 4377 6024 4383
rect 520 4357 600 4363
rect 632 4357 712 4363
rect 760 4357 840 4363
rect 920 4357 936 4363
rect 984 4357 1672 4363
rect 1816 4357 2088 4363
rect 2152 4357 2776 4363
rect 2888 4357 2920 4363
rect 3016 4357 3048 4363
rect 3064 4357 3240 4363
rect 3304 4357 3336 4363
rect 3816 4357 4072 4363
rect 4232 4357 4440 4363
rect 4808 4357 5096 4363
rect 5544 4357 5928 4363
rect 5944 4357 6104 4363
rect 6120 4357 6184 4363
rect 600 4337 664 4343
rect 696 4337 824 4343
rect 840 4337 888 4343
rect 904 4337 968 4343
rect 1224 4337 1800 4343
rect 2248 4337 2312 4343
rect 2408 4337 2632 4343
rect 2648 4337 2680 4343
rect 2776 4337 2792 4343
rect 2968 4337 3128 4343
rect 3176 4337 3320 4343
rect 3352 4337 3784 4343
rect 3832 4337 4088 4343
rect 4456 4337 4696 4343
rect 4712 4337 5128 4343
rect 5432 4337 5848 4343
rect -51 4317 40 4323
rect 424 4317 456 4323
rect 664 4317 979 4323
rect 1005 4317 1011 4332
rect 4429 4328 4435 4332
rect 173 4308 179 4312
rect 296 4297 488 4303
rect 536 4297 632 4303
rect 680 4297 744 4303
rect 765 4297 904 4303
rect 392 4277 536 4283
rect 765 4283 771 4297
rect 920 4297 952 4303
rect 973 4303 979 4317
rect 1032 4317 1048 4323
rect 1112 4317 1128 4323
rect 1160 4317 1208 4323
rect 1512 4317 1720 4323
rect 1752 4317 1992 4323
rect 2008 4317 2200 4323
rect 2216 4317 2248 4323
rect 2264 4317 2408 4323
rect 2456 4317 2536 4323
rect 2616 4317 2744 4323
rect 2760 4317 2792 4323
rect 2936 4317 2952 4323
rect 3048 4317 3272 4323
rect 3656 4317 3720 4323
rect 3736 4317 3816 4323
rect 3848 4317 3912 4323
rect 3976 4317 4072 4323
rect 4328 4317 4392 4323
rect 4552 4317 4600 4323
rect 4648 4317 4696 4323
rect 4968 4317 5032 4323
rect 5560 4317 5704 4323
rect 5816 4317 5832 4323
rect 5885 4323 5891 4332
rect 5880 4317 5891 4323
rect 6040 4317 6072 4323
rect 6824 4317 6867 4323
rect 3485 4308 3491 4312
rect 973 4297 1112 4303
rect 1128 4297 1144 4303
rect 1160 4297 1384 4303
rect 1464 4297 1544 4303
rect 1560 4297 1960 4303
rect 2312 4297 2728 4303
rect 2808 4297 2936 4303
rect 3064 4297 3256 4303
rect 3336 4297 3416 4303
rect 3736 4297 3832 4303
rect 3896 4297 3976 4303
rect 4008 4297 4232 4303
rect 4472 4297 5048 4303
rect 5112 4297 5352 4303
rect 5368 4297 5448 4303
rect 5464 4297 5576 4303
rect 5592 4297 5608 4303
rect 5704 4297 5816 4303
rect 616 4277 771 4283
rect 808 4277 920 4283
rect 952 4277 1048 4283
rect 1208 4277 1272 4283
rect 1448 4277 1560 4283
rect 1784 4277 1912 4283
rect 2248 4277 2472 4283
rect 2488 4277 2696 4283
rect 2712 4277 2824 4283
rect 2936 4277 2984 4283
rect 3016 4277 3064 4283
rect 3085 4277 3096 4283
rect 3085 4268 3091 4277
rect 3144 4277 3208 4283
rect 3304 4277 3816 4283
rect 3832 4277 4008 4283
rect 4104 4277 4520 4283
rect 4552 4277 4568 4283
rect 4584 4277 4824 4283
rect 4856 4277 4872 4283
rect 5016 4277 5352 4283
rect 5688 4277 5704 4283
rect 5736 4277 5816 4283
rect 5864 4277 6056 4283
rect 6296 4277 6424 4283
rect -51 4257 8 4263
rect 40 4257 136 4263
rect 200 4257 424 4263
rect 456 4257 1112 4263
rect 1208 4257 1224 4263
rect 1256 4257 1288 4263
rect 1357 4257 1416 4263
rect 376 4237 600 4243
rect 669 4237 968 4243
rect 669 4223 675 4237
rect 984 4237 1064 4243
rect 1357 4243 1363 4257
rect 1960 4257 2120 4263
rect 2136 4257 2152 4263
rect 2424 4257 2664 4263
rect 3192 4257 3576 4263
rect 3672 4257 3816 4263
rect 4024 4257 4952 4263
rect 4968 4257 5272 4263
rect 5400 4257 5480 4263
rect 5528 4257 5720 4263
rect 6136 4257 6184 4263
rect 1112 4237 1363 4243
rect 1672 4237 1944 4243
rect 2120 4237 2456 4243
rect 2472 4237 2627 4243
rect 440 4217 675 4223
rect 696 4217 856 4223
rect 888 4217 1000 4223
rect 1144 4217 1416 4223
rect 1544 4217 1704 4223
rect 1453 4208 1459 4212
rect 504 4197 952 4203
rect 968 4197 1032 4203
rect 1048 4197 1432 4203
rect 1528 4197 1592 4203
rect 2072 4217 2120 4223
rect 2136 4217 2280 4223
rect 2621 4223 2627 4237
rect 2696 4237 2792 4243
rect 2904 4237 2920 4243
rect 3080 4237 3544 4243
rect 3560 4237 3928 4243
rect 3960 4237 4040 4243
rect 4200 4237 4232 4243
rect 4296 4237 4744 4243
rect 4760 4237 4872 4243
rect 5032 4237 5320 4243
rect 5368 4237 5400 4243
rect 5432 4237 5512 4243
rect 5768 4237 5992 4243
rect 6168 4237 6312 4243
rect 2621 4217 2824 4223
rect 2888 4217 3048 4223
rect 3640 4217 3800 4223
rect 2040 4197 2072 4203
rect 2088 4197 2344 4203
rect 2360 4197 2472 4203
rect 2488 4197 2568 4203
rect 2584 4197 2680 4203
rect 2792 4197 2936 4203
rect 2952 4197 3336 4203
rect 3432 4197 3768 4203
rect 3800 4197 3864 4203
rect 4040 4217 4216 4223
rect 4344 4217 4360 4223
rect 4520 4217 4584 4223
rect 4696 4217 4808 4223
rect 4856 4217 5528 4223
rect 5544 4217 5736 4223
rect 4136 4197 4280 4203
rect 4296 4197 4424 4203
rect 4440 4197 4504 4203
rect 4536 4197 4776 4203
rect 4792 4197 4888 4203
rect 5160 4197 5368 4203
rect 5400 4197 5432 4203
rect 5656 4197 5800 4203
rect 6568 4197 6744 4203
rect 488 4177 504 4183
rect 760 4177 904 4183
rect 920 4177 1512 4183
rect 1528 4177 1576 4183
rect 1624 4177 1736 4183
rect 1752 4177 1784 4183
rect 1800 4177 2136 4183
rect 2152 4177 2232 4183
rect 2568 4177 2712 4183
rect 2808 4177 3128 4183
rect 3144 4177 3176 4183
rect 3480 4177 4120 4183
rect 4152 4177 4536 4183
rect 4552 4177 4840 4183
rect 4936 4177 5032 4183
rect 5048 4177 5176 4183
rect 5240 4177 5304 4183
rect 5336 4177 5416 4183
rect 5544 4177 5672 4183
rect 5832 4177 6552 4183
rect 6712 4177 6728 4183
rect 632 4157 920 4163
rect 936 4157 1080 4163
rect 1117 4157 1208 4163
rect 568 4137 760 4143
rect 840 4137 856 4143
rect 888 4137 936 4143
rect 1016 4137 1080 4143
rect 1117 4143 1123 4157
rect 1272 4157 1368 4163
rect 1432 4157 1608 4163
rect 1832 4157 1992 4163
rect 2008 4157 2280 4163
rect 2328 4157 2600 4163
rect 2680 4157 2872 4163
rect 2936 4157 3032 4163
rect 3048 4157 3336 4163
rect 3736 4157 3864 4163
rect 3880 4157 3944 4163
rect 3981 4157 4472 4163
rect 1213 4148 1219 4152
rect 1096 4137 1123 4143
rect 1368 4137 1384 4143
rect 1416 4137 1528 4143
rect 1576 4137 1656 4143
rect 1704 4137 1816 4143
rect 1832 4137 2760 4143
rect 2792 4137 2952 4143
rect 3112 4137 3816 4143
rect 3981 4143 3987 4157
rect 4488 4157 4584 4163
rect 4952 4157 5016 4163
rect 5032 4157 5192 4163
rect 5256 4157 5816 4163
rect 5832 4157 5960 4163
rect 6136 4157 6200 4163
rect 6296 4157 6328 4163
rect 3832 4137 3987 4143
rect 4008 4137 4024 4143
rect 4088 4137 4136 4143
rect 4424 4137 4536 4143
rect 4568 4137 4744 4143
rect 4872 4137 5016 4143
rect 5288 4137 5416 4143
rect 5672 4137 6280 4143
rect 6440 4137 6472 4143
rect 6488 4137 6616 4143
rect 600 4117 728 4123
rect 744 4117 1416 4123
rect 1432 4117 1608 4123
rect 1624 4117 2008 4123
rect 2216 4117 2280 4123
rect 2360 4117 2376 4123
rect 2472 4117 2776 4123
rect 2792 4117 2840 4123
rect 2872 4117 2888 4123
rect 2920 4117 2984 4123
rect 3000 4117 3160 4123
rect 3192 4117 4024 4123
rect 4040 4117 4456 4123
rect 4536 4117 4632 4123
rect 4728 4117 5000 4123
rect 5037 4117 5128 4123
rect 2429 4108 2435 4112
rect 424 4097 584 4103
rect 776 4097 792 4103
rect 840 4097 883 4103
rect 440 4077 520 4083
rect 680 4077 840 4083
rect 877 4083 883 4097
rect 984 4097 1032 4103
rect 1064 4097 1160 4103
rect 1176 4097 1192 4103
rect 1352 4097 1432 4103
rect 1448 4097 1496 4103
rect 1512 4097 2024 4103
rect 2088 4097 2296 4103
rect 2328 4097 2344 4103
rect 2376 4097 2408 4103
rect 2568 4097 3176 4103
rect 3272 4097 3464 4103
rect 3912 4097 4008 4103
rect 4024 4097 4040 4103
rect 4280 4097 4408 4103
rect 4440 4097 4472 4103
rect 4504 4097 4792 4103
rect 4824 4097 4968 4103
rect 5037 4103 5043 4117
rect 5272 4117 5384 4123
rect 6120 4117 6168 4123
rect 6456 4117 6664 4123
rect 5000 4097 5043 4103
rect 5112 4097 5208 4103
rect 5288 4097 5912 4103
rect 5928 4097 6008 4103
rect 6056 4097 6072 4103
rect 6168 4097 6232 4103
rect 6552 4097 6600 4103
rect 877 4077 1016 4083
rect 1080 4077 1320 4083
rect 1400 4077 1448 4083
rect 1464 4077 1640 4083
rect 1672 4077 1736 4083
rect 1816 4077 1832 4083
rect 1864 4077 1944 4083
rect 2104 4077 2216 4083
rect 2344 4077 2584 4083
rect 2680 4077 2712 4083
rect 2824 4077 2904 4083
rect 2968 4077 3208 4083
rect 3240 4077 3496 4083
rect 3512 4077 3560 4083
rect 3592 4077 3896 4083
rect 3992 4077 4072 4083
rect 4328 4077 4376 4083
rect 4408 4077 4568 4083
rect 4584 4077 4872 4083
rect 4888 4077 4984 4083
rect 5384 4077 5448 4083
rect 5464 4077 5688 4083
rect 5720 4077 5736 4083
rect 5816 4077 5896 4083
rect 6360 4077 6632 4083
rect 312 4057 408 4063
rect 968 4057 1272 4063
rect 1288 4057 1464 4063
rect 1480 4057 1672 4063
rect 1720 4057 1896 4063
rect 2536 4057 2600 4063
rect 2648 4057 2664 4063
rect 2712 4057 2888 4063
rect 3032 4057 3064 4063
rect 3176 4057 3256 4063
rect 3496 4057 4088 4063
rect 4424 4057 4600 4063
rect 4648 4057 4840 4063
rect 4856 4057 5080 4063
rect 5320 4057 5432 4063
rect 5448 4057 5528 4063
rect 5576 4057 5752 4063
rect 5960 4057 6216 4063
rect 6232 4057 6616 4063
rect 328 4037 680 4043
rect 968 4037 1240 4043
rect 1624 4037 1672 4043
rect 1896 4037 1928 4043
rect 2280 4037 2392 4043
rect 2456 4037 2744 4043
rect 2760 4037 2920 4043
rect 3096 4037 3336 4043
rect 3672 4037 4232 4043
rect 4248 4037 4328 4043
rect 4664 4037 5016 4043
rect 5192 4037 5896 4043
rect 5928 4037 6040 4043
rect 24 4017 216 4023
rect 232 4017 360 4023
rect 392 4017 648 4023
rect 936 4017 1192 4023
rect 1240 4017 1416 4023
rect 1496 4017 2072 4023
rect 2296 4017 2520 4023
rect 920 3997 1096 4003
rect 1112 3997 1544 4003
rect 1640 3997 2424 4003
rect 3032 4017 3048 4023
rect 3544 4017 3784 4023
rect 3864 4017 4280 4023
rect 2936 3997 3672 4003
rect 3720 3997 3848 4003
rect 3880 3997 4152 4003
rect 4328 3997 4392 4003
rect 4472 3997 4856 4003
rect 4984 4017 5576 4023
rect 5608 4017 5656 4023
rect 5736 4017 5912 4023
rect 5928 4017 5960 4023
rect 5992 4017 6120 4023
rect 5192 3997 5864 4003
rect 5880 3997 6024 4003
rect 152 3977 312 3983
rect 536 3977 680 3983
rect 1112 3977 1528 3983
rect 1736 3977 1928 3983
rect 1944 3977 2200 3983
rect 2760 3977 2840 3983
rect 2920 3977 3224 3983
rect 3240 3977 3256 3983
rect 3288 3977 3528 3983
rect 3544 3977 3752 3983
rect 3768 3977 3864 3983
rect 3880 3977 4104 3983
rect 4120 3977 4296 3983
rect 4312 3977 5224 3983
rect 5528 3977 5976 3983
rect 6008 3977 6312 3983
rect 696 3957 1352 3963
rect 1432 3957 1864 3963
rect 1880 3957 2024 3963
rect 2552 3957 2776 3963
rect 2792 3957 3000 3963
rect 3048 3957 3112 3963
rect 3128 3957 3240 3963
rect 3256 3957 3720 3963
rect 3944 3957 4211 3963
rect 664 3937 1096 3943
rect 1320 3937 1688 3943
rect 1752 3937 1992 3943
rect 2008 3937 2136 3943
rect 2152 3937 2328 3943
rect 2664 3937 2808 3943
rect 2984 3937 3048 3943
rect 3096 3937 3144 3943
rect 3176 3937 3208 3943
rect 3752 3937 4056 3943
rect 4205 3943 4211 3957
rect 4232 3957 4296 3963
rect 4312 3957 4520 3963
rect 4792 3957 5112 3963
rect 5336 3957 6440 3963
rect 4205 3937 4632 3943
rect 4904 3937 4920 3943
rect 4952 3937 4984 3943
rect 5048 3937 5128 3943
rect 5352 3937 5672 3943
rect 6104 3937 6360 3943
rect 1709 3928 1715 3932
rect 5693 3928 5699 3932
rect -51 3917 8 3923
rect 248 3917 296 3923
rect 376 3917 440 3923
rect 824 3917 904 3923
rect 920 3917 1016 3923
rect 1032 3917 1128 3923
rect 1192 3917 1512 3923
rect 1784 3917 2296 3923
rect 2488 3917 2600 3923
rect 2856 3917 3080 3923
rect 3144 3917 3192 3923
rect 4056 3917 4312 3923
rect 4392 3917 4472 3923
rect 4520 3917 4584 3923
rect 4808 3917 4840 3923
rect 4888 3917 4936 3923
rect 5016 3917 5032 3923
rect 5128 3917 5176 3923
rect 5224 3917 5400 3923
rect 5416 3917 5608 3923
rect 6280 3917 6584 3923
rect 6824 3917 6867 3923
rect 328 3897 392 3903
rect 520 3897 552 3903
rect 568 3897 632 3903
rect 760 3897 792 3903
rect 1208 3897 2552 3903
rect 2664 3897 2712 3903
rect 2744 3897 2920 3903
rect 3480 3897 3560 3903
rect 3576 3897 3768 3903
rect 3784 3897 3848 3903
rect 3880 3897 3944 3903
rect 4072 3897 4152 3903
rect 4488 3897 4952 3903
rect 5112 3897 5144 3903
rect 5192 3897 5320 3903
rect 5336 3897 5448 3903
rect 5464 3897 5480 3903
rect 5656 3897 5688 3903
rect 6040 3897 6152 3903
rect 6296 3897 6424 3903
rect 6504 3897 6568 3903
rect 5885 3888 5891 3892
rect 456 3877 504 3883
rect 520 3877 568 3883
rect 728 3877 760 3883
rect 861 3877 872 3883
rect 904 3877 1096 3883
rect 1112 3877 1192 3883
rect 1240 3877 1560 3883
rect 1704 3877 1752 3883
rect 1768 3877 1816 3883
rect 1896 3877 1976 3883
rect 1992 3877 2104 3883
rect 2712 3877 2776 3883
rect 2856 3877 3128 3883
rect 3432 3877 3480 3883
rect 3560 3877 3624 3883
rect 3688 3877 4376 3883
rect 4392 3877 4872 3883
rect 4888 3877 5112 3883
rect 5352 3877 5448 3883
rect 5592 3877 5624 3883
rect 5688 3877 5768 3883
rect 5992 3877 6008 3883
rect 6120 3877 6136 3883
rect 6584 3877 6600 3883
rect 1565 3868 1571 3872
rect 2125 3868 2131 3872
rect 72 3857 168 3863
rect 392 3857 616 3863
rect 728 3857 840 3863
rect 968 3857 1000 3863
rect 1016 3857 1336 3863
rect 1608 3857 1656 3863
rect 1672 3857 1736 3863
rect 1752 3857 1800 3863
rect 2248 3857 2280 3863
rect 2760 3857 2776 3863
rect 2920 3857 2952 3863
rect 3000 3857 3208 3863
rect 3672 3857 3704 3863
rect 3912 3857 3976 3863
rect 3992 3857 4056 3863
rect 4152 3857 4248 3863
rect 4472 3857 4520 3863
rect 4584 3857 4648 3863
rect 4664 3857 4888 3863
rect 5000 3857 5080 3863
rect 5096 3857 5256 3863
rect 5976 3857 6104 3863
rect 6296 3857 6344 3863
rect 664 3837 776 3843
rect 792 3837 840 3843
rect 856 3837 968 3843
rect 1000 3837 1064 3843
rect 1288 3837 1496 3843
rect 1704 3837 1992 3843
rect 2120 3837 2312 3843
rect 2344 3837 2984 3843
rect 3640 3837 3752 3843
rect 3768 3837 3992 3843
rect 4008 3837 4056 3843
rect 4301 3837 4504 3843
rect 376 3817 408 3823
rect 424 3817 536 3823
rect 552 3817 936 3823
rect 1080 3817 1112 3823
rect 1176 3817 1256 3823
rect 488 3797 552 3803
rect 1160 3797 1272 3803
rect 1528 3797 1576 3803
rect 1592 3797 1768 3803
rect 2088 3817 2680 3823
rect 2696 3817 3224 3823
rect 2728 3797 2888 3803
rect 3064 3797 3304 3803
rect 3320 3797 3368 3803
rect 3480 3797 3592 3803
rect 4301 3823 4307 3837
rect 4712 3837 4728 3843
rect 4856 3837 5064 3843
rect 5544 3837 5992 3843
rect 3976 3817 4307 3823
rect 4328 3817 4344 3823
rect 4360 3817 4632 3823
rect 4648 3817 4680 3823
rect 4728 3817 5144 3823
rect 3944 3797 4216 3803
rect 4248 3797 4344 3803
rect 4360 3797 4440 3803
rect 4456 3797 5256 3803
rect 6328 3817 6536 3823
rect 6040 3797 6184 3803
rect 6200 3797 6232 3803
rect 6248 3797 6440 3803
rect 6696 3797 6867 3803
rect 1000 3777 1112 3783
rect 1688 3777 1944 3783
rect 2024 3777 2456 3783
rect 2664 3777 2760 3783
rect 3032 3777 3112 3783
rect 3256 3777 3576 3783
rect 3720 3777 3864 3783
rect 3944 3777 4152 3783
rect 4520 3777 4760 3783
rect 4781 3777 4872 3783
rect 685 3763 691 3772
rect 536 3757 840 3763
rect 856 3757 1144 3763
rect 1624 3757 1688 3763
rect 1848 3757 1928 3763
rect 1944 3757 2088 3763
rect 2408 3757 2424 3763
rect 2456 3757 2472 3763
rect 2504 3757 2648 3763
rect 2680 3757 2728 3763
rect 2776 3757 2824 3763
rect 3464 3757 3475 3763
rect 3496 3757 3544 3763
rect 3688 3757 3928 3763
rect 4781 3763 4787 3777
rect 4904 3777 5304 3783
rect 5336 3777 5512 3783
rect 5528 3777 5560 3783
rect 6424 3777 6552 3783
rect 4088 3757 4787 3763
rect 4840 3757 4872 3763
rect 4904 3757 4968 3763
rect 4984 3757 5224 3763
rect 5384 3757 5432 3763
rect 5672 3757 6056 3763
rect 6136 3757 6296 3763
rect 6440 3757 6504 3763
rect 6808 3757 6867 3763
rect 1741 3748 1747 3752
rect 264 3737 392 3743
rect 440 3737 456 3743
rect 488 3737 888 3743
rect 1224 3737 1656 3743
rect 1688 3737 1704 3743
rect 1816 3737 1880 3743
rect 2088 3737 2147 3743
rect 413 3728 419 3732
rect 248 3717 280 3723
rect 568 3717 696 3723
rect 936 3717 984 3723
rect 1256 3717 1384 3723
rect 1544 3717 1624 3723
rect 1784 3717 1816 3723
rect 1976 3717 1992 3723
rect 2008 3717 2120 3723
rect 2141 3723 2147 3737
rect 2376 3737 2419 3743
rect 2141 3717 2200 3723
rect 2360 3717 2392 3723
rect 2413 3723 2419 3737
rect 2440 3737 2504 3743
rect 2536 3737 2568 3743
rect 2840 3737 2904 3743
rect 3048 3737 3288 3743
rect 3480 3737 3512 3743
rect 3880 3737 4120 3743
rect 4632 3737 4664 3743
rect 4712 3737 4728 3743
rect 4744 3737 5176 3743
rect 5432 3737 5448 3743
rect 5464 3737 6040 3743
rect 6152 3737 6280 3743
rect 6392 3737 6520 3743
rect 2413 3717 2696 3723
rect 2712 3717 2792 3723
rect 2824 3717 2840 3723
rect 2861 3717 4040 3723
rect 312 3697 360 3703
rect 376 3697 424 3703
rect 760 3697 904 3703
rect 1576 3697 1608 3703
rect 2024 3697 2088 3703
rect 2104 3697 2168 3703
rect 2184 3697 2328 3703
rect 2424 3697 2632 3703
rect 2861 3703 2867 3717
rect 4056 3717 4072 3723
rect 4456 3717 4584 3723
rect 4616 3717 4632 3723
rect 4664 3717 4696 3723
rect 4733 3717 4744 3723
rect 5016 3717 5080 3723
rect 5272 3717 5384 3723
rect 5480 3717 5640 3723
rect 6104 3717 6184 3723
rect 6232 3717 6264 3723
rect 6312 3717 6376 3723
rect 6584 3717 6616 3723
rect 6648 3717 6680 3723
rect 6824 3717 6867 3723
rect 2664 3697 2867 3703
rect 3112 3697 4120 3703
rect 4152 3697 4328 3703
rect 4344 3697 4696 3703
rect 4712 3697 4888 3703
rect 5464 3697 5688 3703
rect 6072 3697 6184 3703
rect 6200 3697 6456 3703
rect 408 3677 456 3683
rect 808 3677 1176 3683
rect 1224 3677 1256 3683
rect 1464 3677 1576 3683
rect 1976 3677 2040 3683
rect 2312 3677 2488 3683
rect 2760 3677 3240 3683
rect 3288 3677 3640 3683
rect 3736 3677 3800 3683
rect 3816 3677 3992 3683
rect 4040 3677 4056 3683
rect 4120 3677 4184 3683
rect 4568 3677 4808 3683
rect 4856 3677 4968 3683
rect 5032 3677 5064 3683
rect 5080 3677 5800 3683
rect 6296 3677 6584 3683
rect 280 3657 424 3663
rect 792 3657 920 3663
rect 1784 3657 2152 3663
rect 2600 3657 2760 3663
rect 2776 3657 3000 3663
rect 3016 3657 3432 3663
rect 3448 3657 4216 3663
rect 4312 3657 4968 3663
rect 5224 3657 5304 3663
rect 5320 3657 5976 3663
rect 216 3637 312 3643
rect 328 3637 616 3643
rect 744 3637 968 3643
rect 1352 3637 1448 3643
rect 1528 3637 3144 3643
rect 3160 3637 3384 3643
rect 3400 3637 5160 3643
rect 5176 3637 5384 3643
rect 5400 3637 5976 3643
rect 6168 3637 6344 3643
rect 6360 3637 6600 3643
rect 6616 3637 6632 3643
rect 376 3617 488 3623
rect 504 3617 568 3623
rect 856 3617 1112 3623
rect 1656 3617 1704 3623
rect 2456 3617 2600 3623
rect 984 3597 1080 3603
rect 1096 3597 1128 3603
rect 1608 3597 2424 3603
rect 2680 3597 2792 3603
rect 3080 3617 3096 3623
rect 3144 3617 3624 3623
rect 4280 3617 4536 3623
rect 2936 3597 3144 3603
rect 3992 3597 4152 3603
rect 4184 3597 4248 3603
rect 4264 3597 4675 3603
rect 5064 3617 5096 3623
rect 5144 3617 5448 3623
rect 6168 3617 6456 3623
rect 1368 3577 1480 3583
rect 1496 3577 1976 3583
rect 1992 3577 2232 3583
rect 2280 3577 4648 3583
rect 4669 3583 4675 3597
rect 4984 3597 5160 3603
rect 5304 3597 5496 3603
rect 5624 3597 6168 3603
rect 6184 3597 6264 3603
rect 6280 3597 6376 3603
rect 4669 3577 5224 3583
rect 5816 3577 5912 3583
rect 5928 3577 6168 3583
rect 200 3557 360 3563
rect 456 3557 872 3563
rect 920 3557 984 3563
rect 1000 3557 1112 3563
rect 1976 3557 3176 3563
rect 3256 3557 3352 3563
rect 3752 3557 4040 3563
rect 4376 3557 5016 3563
rect 5032 3557 5976 3563
rect 6024 3557 6072 3563
rect 6088 3557 6296 3563
rect 6312 3557 6328 3563
rect 232 3537 264 3543
rect 312 3537 472 3543
rect 520 3537 568 3543
rect 632 3537 664 3543
rect 680 3537 1032 3543
rect 1048 3537 2088 3543
rect 2168 3537 2360 3543
rect 2440 3537 2504 3543
rect 2584 3537 2728 3543
rect 2968 3537 3256 3543
rect 3272 3537 3400 3543
rect 3704 3537 3752 3543
rect 3816 3537 3832 3543
rect 4232 3537 4280 3543
rect 4616 3537 4808 3543
rect 5128 3537 5192 3543
rect 5768 3537 5864 3543
rect 6040 3537 6152 3543
rect 6232 3537 6248 3543
rect 120 3517 248 3523
rect 296 3517 392 3523
rect 440 3517 472 3523
rect 568 3517 648 3523
rect 664 3517 712 3523
rect 872 3517 920 3523
rect 1016 3517 1192 3523
rect 1256 3517 1464 3523
rect 1544 3517 1560 3523
rect 1592 3517 1624 3523
rect 1688 3517 1736 3523
rect 1768 3517 2008 3523
rect 2296 3517 2648 3523
rect 2824 3517 2920 3523
rect 3032 3517 3048 3523
rect 3096 3517 3112 3523
rect 3176 3517 3352 3523
rect 3448 3517 3960 3523
rect 4008 3517 4360 3523
rect 4376 3517 4392 3523
rect 4776 3517 5720 3523
rect 6264 3517 6280 3523
rect 861 3508 867 3512
rect 2237 3508 2243 3512
rect 216 3497 408 3503
rect 424 3497 584 3503
rect 600 3497 744 3503
rect 952 3497 1080 3503
rect 1656 3497 1752 3503
rect 1784 3497 1944 3503
rect 2024 3497 2040 3503
rect 2392 3497 2520 3503
rect 2600 3497 2696 3503
rect 3304 3497 3432 3503
rect 3480 3497 3528 3503
rect 3592 3497 3768 3503
rect 3864 3497 4408 3503
rect 4568 3497 4584 3503
rect 4600 3497 4664 3503
rect 4808 3497 4840 3503
rect 4856 3497 4872 3503
rect 5048 3497 5112 3503
rect 5240 3497 5336 3503
rect 5464 3497 5640 3503
rect 5800 3497 5816 3503
rect 5896 3497 5992 3503
rect 6040 3497 6168 3503
rect 6184 3497 6200 3503
rect 6232 3497 6504 3503
rect 941 3488 947 3492
rect 360 3477 504 3483
rect 568 3477 584 3483
rect 616 3477 760 3483
rect 968 3477 1032 3483
rect 1480 3477 1720 3483
rect 1960 3477 2424 3483
rect 2440 3477 2504 3483
rect 2520 3477 2744 3483
rect 2760 3477 2936 3483
rect 2952 3477 3016 3483
rect 3112 3477 3336 3483
rect 3384 3477 3592 3483
rect 3608 3477 3720 3483
rect 4184 3477 4328 3483
rect 4648 3477 4760 3483
rect 4792 3477 4856 3483
rect 4872 3477 5176 3483
rect 5192 3477 5256 3483
rect 5704 3477 5960 3483
rect 5992 3477 6296 3483
rect 6312 3477 6328 3483
rect 6456 3477 6664 3483
rect 248 3457 568 3463
rect 760 3457 1048 3463
rect 1064 3457 1096 3463
rect 1608 3457 1704 3463
rect 1752 3457 2104 3463
rect 2232 3457 2312 3463
rect 2360 3457 2648 3463
rect 2712 3457 3064 3463
rect 3576 3457 3656 3463
rect 3864 3457 4184 3463
rect 4232 3457 4312 3463
rect 4333 3463 4339 3472
rect 4333 3457 4488 3463
rect 4504 3457 4840 3463
rect 4856 3457 5048 3463
rect 5064 3457 5096 3463
rect 5160 3457 5192 3463
rect 5213 3457 5480 3463
rect 488 3437 648 3443
rect 680 3437 888 3443
rect 984 3437 1016 3443
rect 1352 3437 1560 3443
rect 1640 3437 1688 3443
rect 1816 3437 2984 3443
rect 3176 3437 3304 3443
rect 3384 3437 3704 3443
rect 3720 3437 3912 3443
rect 4072 3437 4264 3443
rect 4360 3437 4520 3443
rect 4936 3437 5128 3443
rect 5213 3443 5219 3457
rect 5800 3457 6024 3463
rect 6168 3457 6376 3463
rect 6760 3457 6776 3463
rect 5192 3437 5219 3443
rect 5384 3437 5688 3443
rect 5880 3437 5928 3443
rect 6333 3437 6424 3443
rect 248 3417 280 3423
rect 536 3417 680 3423
rect 696 3417 824 3423
rect 888 3417 904 3423
rect 1048 3417 1112 3423
rect 1128 3417 1528 3423
rect 1544 3417 1800 3423
rect 280 3397 456 3403
rect 520 3397 600 3403
rect 648 3397 984 3403
rect 1016 3397 1064 3403
rect 1560 3397 1816 3403
rect 2104 3417 2264 3423
rect 2376 3417 2600 3423
rect 2776 3417 2968 3423
rect 3096 3417 3256 3423
rect 3304 3417 3464 3423
rect 1944 3397 2056 3403
rect 2088 3397 2552 3403
rect 2568 3397 2888 3403
rect 2920 3397 3416 3403
rect 3496 3397 3816 3403
rect 4312 3417 4584 3423
rect 4632 3417 5224 3423
rect 5304 3417 5400 3423
rect 5464 3417 5880 3423
rect 3944 3397 4120 3403
rect 4296 3397 4552 3403
rect 4712 3397 4776 3403
rect 5080 3397 5160 3403
rect 5176 3397 5368 3403
rect 5384 3397 5464 3403
rect 5592 3397 5688 3403
rect 6333 3423 6339 3437
rect 6520 3437 6632 3443
rect 6088 3417 6339 3423
rect 6360 3417 6664 3423
rect 6008 3397 6312 3403
rect 6376 3397 6392 3403
rect 152 3377 248 3383
rect 296 3377 568 3383
rect 584 3377 696 3383
rect 712 3377 824 3383
rect 840 3377 1208 3383
rect 1256 3377 1496 3383
rect 1816 3377 2008 3383
rect 2024 3377 2200 3383
rect 2216 3377 2248 3383
rect 2264 3377 2280 3383
rect 2472 3377 2568 3383
rect 2632 3377 2856 3383
rect 3352 3377 3784 3383
rect 3816 3377 5288 3383
rect 5480 3377 6456 3383
rect 6584 3377 6696 3383
rect 6712 3377 6744 3383
rect 56 3357 104 3363
rect 184 3357 344 3363
rect 456 3357 520 3363
rect 1592 3357 1800 3363
rect 1880 3357 2088 3363
rect 2333 3357 2344 3363
rect 2424 3357 2456 3363
rect 2536 3357 2760 3363
rect 2824 3357 2952 3363
rect 3176 3357 3224 3363
rect 3432 3357 3464 3363
rect 3480 3357 3640 3363
rect 3656 3357 3672 3363
rect 3704 3357 3944 3363
rect 3976 3357 4168 3363
rect 4413 3357 4520 3363
rect 589 3348 595 3352
rect 893 3348 899 3352
rect 104 3337 328 3343
rect 344 3337 376 3343
rect 1544 3337 1672 3343
rect 1688 3337 1960 3343
rect 1976 3337 2040 3343
rect 2056 3337 2232 3343
rect 2600 3337 2760 3343
rect 2776 3337 2968 3343
rect 2984 3337 3032 3343
rect 3192 3337 3704 3343
rect 3800 3337 4008 3343
rect 4200 3337 4264 3343
rect 4413 3343 4419 3357
rect 4536 3357 4744 3363
rect 4824 3357 4872 3363
rect 4888 3357 5048 3363
rect 5064 3357 5288 3363
rect 5320 3357 5528 3363
rect 5720 3357 5832 3363
rect 5880 3357 5896 3363
rect 5960 3357 6056 3363
rect 6072 3357 6088 3363
rect 6104 3357 6152 3363
rect 6184 3357 6280 3363
rect 6328 3357 6360 3363
rect 6392 3357 6488 3363
rect 6648 3357 6744 3363
rect 4280 3337 4419 3343
rect 4696 3337 4707 3343
rect 4728 3337 4952 3343
rect 5080 3337 5144 3343
rect 5160 3337 5608 3343
rect 5912 3337 6104 3343
rect 6280 3337 6584 3343
rect 6728 3337 6776 3343
rect 72 3317 88 3323
rect 136 3317 328 3323
rect 424 3317 440 3323
rect 456 3317 595 3323
rect 605 3317 611 3332
rect 4429 3328 4435 3332
rect 4509 3328 4515 3332
rect 88 3297 152 3303
rect 168 3297 184 3303
rect 232 3297 248 3303
rect 376 3297 488 3303
rect 589 3303 595 3317
rect 808 3317 867 3323
rect 589 3297 632 3303
rect 808 3297 840 3303
rect 861 3303 867 3317
rect 920 3317 1064 3323
rect 1640 3317 1736 3323
rect 1896 3317 2072 3323
rect 2088 3317 2200 3323
rect 2216 3317 2472 3323
rect 2488 3317 2520 3323
rect 2552 3317 2840 3323
rect 2856 3317 3048 3323
rect 3144 3317 3240 3323
rect 3336 3317 3560 3323
rect 3608 3317 3816 3323
rect 4008 3317 4072 3323
rect 4120 3317 4200 3323
rect 4248 3317 4296 3323
rect 4568 3317 4744 3323
rect 4760 3317 4840 3323
rect 4936 3317 4995 3323
rect 1181 3308 1187 3312
rect 861 3297 952 3303
rect 1576 3297 1624 3303
rect 1672 3297 1800 3303
rect 1816 3297 1896 3303
rect 1928 3297 1992 3303
rect 2072 3297 2120 3303
rect 2136 3297 2168 3303
rect 2248 3297 2328 3303
rect 2344 3297 2376 3303
rect 2504 3297 2792 3303
rect 3032 3297 3096 3303
rect 3117 3297 3176 3303
rect 40 3277 216 3283
rect 296 3277 584 3283
rect 856 3277 936 3283
rect 952 3277 1000 3283
rect 2024 3277 2360 3283
rect 2392 3277 2664 3283
rect 3117 3283 3123 3297
rect 3208 3297 3240 3303
rect 3288 3297 3368 3303
rect 3624 3297 3656 3303
rect 3688 3297 3736 3303
rect 3752 3297 3864 3303
rect 3880 3297 4216 3303
rect 4376 3297 4392 3303
rect 4472 3297 4552 3303
rect 4712 3297 4776 3303
rect 4808 3297 4920 3303
rect 4989 3303 4995 3317
rect 5032 3317 5272 3323
rect 5352 3317 5432 3323
rect 5448 3317 5464 3323
rect 5512 3317 5560 3323
rect 5629 3317 5635 3332
rect 5720 3317 5752 3323
rect 5848 3317 6200 3323
rect 6216 3317 6520 3323
rect 4989 3297 5032 3303
rect 5096 3297 5176 3303
rect 5208 3297 5256 3303
rect 5560 3297 5608 3303
rect 5656 3297 5928 3303
rect 5944 3297 6184 3303
rect 6264 3297 6344 3303
rect 6440 3297 6712 3303
rect 2696 3277 3123 3283
rect 3144 3277 3224 3283
rect 3240 3277 3432 3283
rect 3448 3277 3528 3283
rect 3560 3277 3896 3283
rect 3912 3277 4344 3283
rect 4520 3277 4568 3283
rect 4584 3277 4728 3283
rect 4744 3277 4824 3283
rect 4840 3277 5416 3283
rect 5432 3277 5672 3283
rect 5736 3277 5784 3283
rect 5848 3277 5896 3283
rect 5912 3277 6040 3283
rect 328 3257 520 3263
rect 712 3257 904 3263
rect 1128 3257 1144 3263
rect 1160 3257 1432 3263
rect 1704 3257 2152 3263
rect 2168 3257 2344 3263
rect 2360 3257 2568 3263
rect 2728 3257 3448 3263
rect 3464 3257 3496 3263
rect 3704 3257 3832 3263
rect 4024 3257 4344 3263
rect 4360 3257 4456 3263
rect 4632 3257 5080 3263
rect 5480 3257 6168 3263
rect 88 3237 328 3243
rect 584 3237 1064 3243
rect 1496 3237 1672 3243
rect 2104 3237 2616 3243
rect 3112 3237 3544 3243
rect 3944 3237 4168 3243
rect 4184 3237 4280 3243
rect 4456 3237 4600 3243
rect 4648 3237 5096 3243
rect 5176 3237 5320 3243
rect 5336 3237 6008 3243
rect 6040 3237 6216 3243
rect 328 3197 424 3203
rect 2120 3217 2136 3223
rect 2568 3217 2616 3223
rect 2168 3197 2232 3203
rect 2248 3197 2408 3203
rect 2952 3217 3512 3223
rect 3528 3217 3992 3223
rect 4344 3217 4664 3223
rect 2936 3197 3128 3203
rect 3144 3197 3400 3203
rect 3752 3197 3800 3203
rect 4024 3197 4328 3203
rect 4360 3197 4632 3203
rect 5096 3217 5240 3223
rect 5272 3217 5352 3223
rect 5597 3217 5880 3223
rect 5597 3203 5603 3217
rect 5896 3217 5992 3223
rect 6024 3217 6104 3223
rect 5224 3197 5603 3203
rect 5624 3197 5704 3203
rect 5784 3197 5864 3203
rect 5896 3197 6056 3203
rect 6152 3197 6536 3203
rect 632 3177 1608 3183
rect 1992 3177 2424 3183
rect 2600 3177 3272 3183
rect 3576 3177 3928 3183
rect 4408 3177 4504 3183
rect 4520 3177 4568 3183
rect 4584 3177 4712 3183
rect 4984 3177 5048 3183
rect 5304 3177 5320 3183
rect 5496 3177 5656 3183
rect 5672 3177 5896 3183
rect 5960 3177 6088 3183
rect 6104 3177 6552 3183
rect 296 3157 408 3163
rect 712 3157 920 3163
rect 1192 3157 1240 3163
rect 1848 3157 1912 3163
rect 1928 3157 2024 3163
rect 2312 3157 2568 3163
rect 2632 3157 3080 3163
rect 3208 3157 3368 3163
rect 3976 3157 4136 3163
rect 4504 3157 4520 3163
rect 4552 3157 4664 3163
rect 4728 3157 4968 3163
rect 5368 3157 5688 3163
rect 5704 3157 5912 3163
rect 6088 3157 6264 3163
rect 312 3137 472 3143
rect 536 3137 600 3143
rect 616 3137 1160 3143
rect 1256 3137 1400 3143
rect 1416 3137 1592 3143
rect 1608 3137 1656 3143
rect 1832 3137 1896 3143
rect 2072 3137 2664 3143
rect 2712 3137 2840 3143
rect 2856 3137 3016 3143
rect 3080 3137 3176 3143
rect 3304 3137 3512 3143
rect 3528 3137 4648 3143
rect 4680 3137 4808 3143
rect 4824 3137 5352 3143
rect 5576 3137 5624 3143
rect 5640 3137 5736 3143
rect 5912 3137 6040 3143
rect 6056 3137 6552 3143
rect 6568 3137 6648 3143
rect 264 3117 360 3123
rect 616 3117 712 3123
rect 824 3117 1272 3123
rect 1288 3117 1336 3123
rect 1448 3117 1480 3123
rect 1496 3117 1720 3123
rect 1736 3117 1752 3123
rect 1768 3117 1832 3123
rect 1944 3117 1992 3123
rect 2008 3117 2104 3123
rect 2168 3117 2424 3123
rect 2568 3117 2728 3123
rect 2776 3117 3000 3123
rect 3016 3117 3112 3123
rect 3160 3117 3192 3123
rect 3240 3117 3256 3123
rect 3368 3117 3384 3123
rect 3912 3117 3928 3123
rect 4072 3117 4216 3123
rect 4232 3117 4488 3123
rect 4504 3117 4552 3123
rect 4712 3117 4728 3123
rect 4776 3117 5144 3123
rect 5352 3117 5416 3123
rect 5528 3117 5800 3123
rect 5832 3117 6008 3123
rect 6056 3117 6067 3123
rect 6296 3117 6312 3123
rect 6552 3117 6632 3123
rect 408 3097 424 3103
rect 440 3097 648 3103
rect 728 3097 776 3103
rect 920 3097 1080 3103
rect 1160 3097 1208 3103
rect 1224 3097 1256 3103
rect 1304 3097 1704 3103
rect 1816 3097 2008 3103
rect 2120 3097 2168 3103
rect 2184 3097 2344 3103
rect 2520 3097 2600 3103
rect 2728 3097 2760 3103
rect 2824 3097 2920 3103
rect 3000 3097 3032 3103
rect 3064 3097 3219 3103
rect 3037 3088 3043 3092
rect 312 3077 408 3083
rect 424 3077 728 3083
rect 904 3077 1256 3083
rect 1336 3077 2072 3083
rect 2104 3077 2184 3083
rect 2200 3077 2616 3083
rect 2712 3077 2723 3083
rect 3080 3077 3144 3083
rect 3213 3083 3219 3097
rect 3256 3097 3288 3103
rect 3400 3097 4552 3103
rect 4568 3097 4712 3103
rect 5016 3097 5080 3103
rect 5096 3097 5176 3103
rect 5192 3097 5256 3103
rect 5272 3097 5336 3103
rect 5496 3097 5512 3103
rect 5544 3097 5592 3103
rect 5720 3097 5795 3103
rect 3213 3077 3528 3083
rect 3560 3077 3624 3083
rect 3800 3077 3848 3083
rect 3864 3077 3976 3083
rect 4136 3077 4168 3083
rect 4264 3077 4312 3083
rect 4344 3077 4440 3083
rect 4472 3077 4696 3083
rect 4733 3083 4739 3092
rect 4733 3077 4744 3083
rect 4808 3077 4872 3083
rect 4888 3077 5016 3083
rect 5048 3077 5256 3083
rect 5272 3077 5400 3083
rect 5416 3077 5640 3083
rect 5656 3077 5720 3083
rect 5789 3083 5795 3097
rect 6264 3097 6504 3103
rect 6536 3097 6600 3103
rect 5789 3077 5848 3083
rect 6296 3077 6360 3083
rect 6424 3077 6568 3083
rect 248 3057 520 3063
rect 552 3057 632 3063
rect 744 3057 1192 3063
rect 1416 3057 1624 3063
rect 1720 3057 1736 3063
rect 1752 3057 1800 3063
rect 1896 3057 2184 3063
rect 2216 3057 2296 3063
rect 2344 3057 2360 3063
rect 2408 3057 2424 3063
rect 2552 3057 2568 3063
rect 2600 3057 2648 3063
rect 2744 3057 3000 3063
rect 3016 3057 3048 3063
rect 3160 3057 3208 3063
rect 3368 3057 3608 3063
rect 3624 3057 3736 3063
rect 3768 3057 4344 3063
rect 4440 3057 4792 3063
rect 4888 3057 4984 3063
rect 5000 3057 5096 3063
rect 5112 3057 5224 3063
rect 5304 3057 5352 3063
rect 5368 3057 5528 3063
rect 5896 3057 5944 3063
rect 5960 3057 6104 3063
rect 6248 3057 6280 3063
rect 136 3037 440 3043
rect 872 3037 920 3043
rect 1032 3037 1144 3043
rect 1192 3037 1224 3043
rect 1336 3037 1416 3043
rect 1480 3037 1560 3043
rect 1640 3037 1656 3043
rect 1720 3037 1896 3043
rect 2200 3037 2248 3043
rect 2264 3037 2280 3043
rect 2328 3037 2408 3043
rect 2472 3037 2904 3043
rect 2952 3037 3080 3043
rect 3240 3037 3368 3043
rect 3448 3037 3528 3043
rect 3816 3037 3976 3043
rect 4680 3037 4776 3043
rect 5160 3037 5304 3043
rect 5320 3037 5480 3043
rect 5560 3037 5624 3043
rect 5816 3037 5928 3043
rect 6424 3037 6744 3043
rect 856 3017 888 3023
rect 984 3017 1048 3023
rect 1512 3017 1800 3023
rect 408 2997 424 3003
rect 440 2997 904 3003
rect 1144 2997 1176 3003
rect 1656 2997 1784 3003
rect 1800 2997 1816 3003
rect 1960 3017 2392 3023
rect 2632 3017 2856 3023
rect 2968 3017 3336 3023
rect 3352 3017 3400 3023
rect 3416 3017 3448 3023
rect 3512 3017 3624 3023
rect 2040 2997 2200 3003
rect 2648 2997 2792 3003
rect 2968 2997 3048 3003
rect 3208 2997 3256 3003
rect 3272 2997 3320 3003
rect 3544 2997 3560 3003
rect 3960 3017 4472 3023
rect 4488 3017 4664 3023
rect 4824 3017 4888 3023
rect 5560 3017 5704 3023
rect 5720 3017 5848 3023
rect 4184 2997 4200 3003
rect 4520 2997 4568 3003
rect 4664 2997 4888 3003
rect 5432 2997 5560 3003
rect 5672 2997 5880 3003
rect 6072 3017 6408 3023
rect 6552 3017 6632 3023
rect 6184 2997 6808 3003
rect 392 2977 616 2983
rect 984 2977 1032 2983
rect 1352 2977 1416 2983
rect 1464 2977 1704 2983
rect 1768 2977 2296 2983
rect 2392 2977 2600 2983
rect 3048 2977 3096 2983
rect 3368 2977 3384 2983
rect 3400 2977 3464 2983
rect 4088 2977 4104 2983
rect 4136 2977 4232 2983
rect 4264 2977 4728 2983
rect 4744 2977 4856 2983
rect 4936 2977 4952 2983
rect 5624 2977 5640 2983
rect 5816 2977 6168 2983
rect 6216 2977 6664 2983
rect 221 2968 227 2972
rect 1725 2968 1731 2972
rect 552 2957 664 2963
rect 936 2957 1192 2963
rect 1336 2957 1448 2963
rect 1464 2957 1688 2963
rect 2008 2957 2088 2963
rect 2280 2957 2376 2963
rect 2408 2957 2808 2963
rect 2920 2957 3560 2963
rect 4104 2957 4744 2963
rect 4792 2957 4968 2963
rect 5016 2957 5896 2963
rect 6024 2957 6088 2963
rect 6280 2957 6376 2963
rect 6392 2957 6472 2963
rect 6648 2957 6728 2963
rect 6744 2957 6776 2963
rect 6824 2957 6867 2963
rect 6557 2948 6563 2952
rect -51 2937 216 2943
rect 360 2937 456 2943
rect 584 2937 616 2943
rect 664 2937 984 2943
rect 1160 2937 1272 2943
rect 1304 2937 1560 2943
rect 1576 2937 2280 2943
rect 2696 2937 3080 2943
rect 3224 2937 3384 2943
rect 3416 2937 3656 2943
rect 3672 2937 4280 2943
rect 4552 2937 4584 2943
rect 4648 2937 4712 2943
rect 4728 2937 5416 2943
rect 5608 2937 5624 2943
rect 5640 2937 5720 2943
rect 5928 2937 6008 2943
rect 6376 2937 6424 2943
rect 333 2928 339 2932
rect 200 2917 280 2923
rect 456 2917 584 2923
rect 664 2917 712 2923
rect 1048 2917 1112 2923
rect 1128 2917 1272 2923
rect 1576 2917 1592 2923
rect 1752 2917 1928 2923
rect 2120 2917 2536 2923
rect 2744 2917 3160 2923
rect 3464 2917 3496 2923
rect 3832 2917 3944 2923
rect 3960 2917 4264 2923
rect 4536 2917 4552 2923
rect 4760 2917 4872 2923
rect 4888 2917 4904 2923
rect 4936 2917 4984 2923
rect 5048 2917 5080 2923
rect 5240 2917 5272 2923
rect 5512 2917 5656 2923
rect 5896 2917 5928 2923
rect 5944 2917 5976 2923
rect 5992 2917 6339 2923
rect 4429 2908 4435 2912
rect 40 2897 200 2903
rect 344 2897 392 2903
rect 536 2897 552 2903
rect 600 2897 680 2903
rect 696 2897 712 2903
rect 1096 2897 1160 2903
rect 1320 2897 1400 2903
rect 1544 2897 1624 2903
rect 1672 2897 1768 2903
rect 1848 2897 1912 2903
rect 1944 2897 2136 2903
rect 2312 2897 2408 2903
rect 2712 2897 2760 2903
rect 3000 2897 3016 2903
rect 3101 2897 3144 2903
rect 269 2888 275 2892
rect 296 2877 488 2883
rect 504 2877 1096 2883
rect 1480 2877 1496 2883
rect 1816 2877 1880 2883
rect 1992 2877 2024 2883
rect 2120 2877 2280 2883
rect 2328 2877 2344 2883
rect 2488 2877 2584 2883
rect 2600 2877 2920 2883
rect 3101 2883 3107 2897
rect 3224 2897 3240 2903
rect 3288 2897 3432 2903
rect 3768 2897 4072 2903
rect 4088 2897 4120 2903
rect 4472 2897 4520 2903
rect 4568 2897 4664 2903
rect 4776 2897 4808 2903
rect 4856 2897 5048 2903
rect 5112 2897 5128 2903
rect 5256 2897 5272 2903
rect 5400 2897 5480 2903
rect 5592 2897 5672 2903
rect 5688 2897 5768 2903
rect 5992 2897 6072 2903
rect 6168 2897 6248 2903
rect 6264 2897 6312 2903
rect 6333 2903 6339 2917
rect 6360 2917 6440 2923
rect 6536 2917 6616 2923
rect 6632 2917 6712 2923
rect 6824 2917 6867 2923
rect 6333 2897 6472 2903
rect 6488 2897 6520 2903
rect 6616 2897 6680 2903
rect 6696 2897 6712 2903
rect 3080 2877 3107 2883
rect 3144 2877 3224 2883
rect 3240 2877 3864 2883
rect 3880 2877 4600 2883
rect 4616 2877 4632 2883
rect 4664 2877 5064 2883
rect 5096 2877 5176 2883
rect 5432 2877 5480 2883
rect 5656 2877 6024 2883
rect 6040 2877 6120 2883
rect 6488 2877 6504 2883
rect 120 2857 360 2863
rect 712 2857 1032 2863
rect 1816 2857 2184 2863
rect 2200 2857 2248 2863
rect 2456 2857 2488 2863
rect 2504 2857 2552 2863
rect 2568 2857 2936 2863
rect 2952 2857 3128 2863
rect 3144 2857 3320 2863
rect 3384 2857 4248 2863
rect 4840 2857 5080 2863
rect 5432 2857 5496 2863
rect 5560 2857 6136 2863
rect 136 2837 280 2843
rect 312 2837 376 2843
rect 664 2837 1624 2843
rect 1832 2837 2152 2843
rect 2216 2837 2488 2843
rect 2584 2837 3736 2843
rect 3752 2837 4328 2843
rect 4344 2837 5176 2843
rect 5208 2837 5544 2843
rect 5944 2837 6552 2843
rect 1000 2817 1192 2823
rect 1368 2817 1592 2823
rect 1709 2817 1848 2823
rect 1709 2803 1715 2817
rect 1944 2817 2088 2823
rect 2136 2817 2264 2823
rect 2520 2817 2680 2823
rect 1416 2797 1715 2803
rect 1800 2797 2360 2803
rect 2392 2797 2744 2803
rect 2920 2817 2952 2823
rect 2968 2817 3208 2823
rect 3608 2817 3656 2823
rect 3784 2817 3832 2823
rect 4184 2817 4392 2823
rect 4600 2817 4856 2823
rect 3080 2797 3096 2803
rect 3160 2797 3592 2803
rect 4328 2797 4440 2803
rect 4520 2797 4760 2803
rect 5048 2817 6584 2823
rect 5224 2797 5304 2803
rect 5544 2797 5576 2803
rect 872 2777 1288 2783
rect 1624 2777 2072 2783
rect 2088 2777 2776 2783
rect 2792 2777 3208 2783
rect 3320 2777 3427 2783
rect 600 2757 856 2763
rect 1016 2757 1048 2763
rect 1064 2757 1256 2763
rect 1320 2757 1352 2763
rect 1373 2757 1528 2763
rect 728 2737 840 2743
rect 888 2737 1064 2743
rect 1096 2737 1128 2743
rect 1192 2737 1272 2743
rect 1373 2743 1379 2757
rect 1672 2757 1784 2763
rect 2056 2757 2120 2763
rect 2136 2757 2200 2763
rect 2424 2757 2728 2763
rect 2936 2757 3080 2763
rect 3176 2757 3320 2763
rect 3336 2757 3400 2763
rect 3421 2763 3427 2777
rect 3448 2777 3608 2783
rect 4088 2777 4376 2783
rect 4392 2777 4600 2783
rect 4760 2777 5352 2783
rect 5560 2777 5960 2783
rect 6104 2777 6632 2783
rect 3421 2757 3688 2763
rect 4088 2757 4120 2763
rect 4136 2757 4344 2763
rect 4392 2757 4744 2763
rect 5016 2757 5128 2763
rect 5144 2757 5160 2763
rect 5176 2757 5240 2763
rect 5416 2757 5432 2763
rect 5768 2757 6184 2763
rect 6200 2757 6552 2763
rect 6600 2757 6696 2763
rect 1304 2737 1379 2743
rect 1784 2737 1816 2743
rect 1976 2737 1992 2743
rect 2152 2737 2232 2743
rect 2840 2737 2952 2743
rect 3112 2737 3144 2743
rect 3496 2737 3624 2743
rect 3896 2737 4200 2743
rect 4296 2737 4504 2743
rect 5256 2737 5832 2743
rect 5848 2737 6024 2743
rect 6056 2737 6152 2743
rect 6440 2737 6632 2743
rect -51 2717 8 2723
rect 168 2717 232 2723
rect 712 2717 904 2723
rect 984 2717 1528 2723
rect 1608 2717 2104 2723
rect 2152 2717 2856 2723
rect 2872 2717 3528 2723
rect 3592 2717 3640 2723
rect 4040 2717 4136 2723
rect 4344 2717 4488 2723
rect 4920 2717 4952 2723
rect 5064 2717 5752 2723
rect 5768 2717 5784 2723
rect 5896 2717 5912 2723
rect 6104 2717 6536 2723
rect 6552 2717 6696 2723
rect 136 2697 392 2703
rect 872 2697 936 2703
rect 1048 2697 1064 2703
rect 1080 2697 1128 2703
rect 1272 2697 1784 2703
rect 1800 2697 1896 2703
rect 1976 2697 2120 2703
rect 2136 2697 2696 2703
rect 2728 2697 2760 2703
rect 3096 2697 3288 2703
rect 3416 2697 3480 2703
rect 3560 2697 3784 2703
rect 4152 2697 4472 2703
rect 4488 2697 4520 2703
rect 4936 2697 4952 2703
rect 4968 2697 5240 2703
rect 5272 2697 5283 2703
rect 136 2677 328 2683
rect 344 2677 408 2683
rect 424 2677 792 2683
rect 856 2677 1032 2683
rect 1048 2677 1080 2683
rect 1112 2677 1144 2683
rect 1272 2677 1368 2683
rect 1624 2677 1656 2683
rect 1736 2677 1752 2683
rect 1768 2677 2008 2683
rect 2024 2677 2440 2683
rect 2456 2677 2632 2683
rect 2696 2677 2808 2683
rect 3112 2677 3160 2683
rect 3400 2677 3672 2683
rect 3896 2677 3928 2683
rect 3992 2677 4056 2683
rect 4120 2677 4200 2683
rect 4232 2677 4248 2683
rect 4280 2677 4312 2683
rect 4392 2677 4440 2683
rect 4632 2677 4680 2683
rect 4712 2677 4872 2683
rect 4904 2677 5048 2683
rect 5112 2677 5128 2683
rect 5160 2677 5208 2683
rect 5277 2683 5283 2697
rect 5368 2697 5384 2703
rect 5432 2697 5560 2703
rect 5576 2697 5720 2703
rect 5736 2697 5800 2703
rect 5869 2688 5875 2703
rect 5928 2697 5976 2703
rect 6008 2697 6120 2703
rect 6232 2697 6248 2703
rect 6312 2697 6344 2703
rect 6408 2697 6488 2703
rect 6616 2697 6632 2703
rect 6648 2697 6712 2703
rect 5277 2677 5352 2683
rect 5368 2677 5699 2683
rect 56 2657 136 2663
rect 728 2657 744 2663
rect 808 2657 840 2663
rect 856 2657 1160 2663
rect 1272 2657 1416 2663
rect 1448 2657 1976 2663
rect 2040 2657 2280 2663
rect 2344 2657 2392 2663
rect 2472 2657 2504 2663
rect 2552 2657 2616 2663
rect 2680 2657 2707 2663
rect 440 2637 504 2643
rect 760 2637 984 2643
rect 1000 2637 1096 2643
rect 1224 2637 1384 2643
rect 1400 2637 1496 2643
rect 1672 2637 1704 2643
rect 1725 2637 1832 2643
rect 1448 2617 1624 2623
rect 1725 2623 1731 2637
rect 1928 2637 2056 2643
rect 2200 2637 2232 2643
rect 2392 2637 2600 2643
rect 2616 2637 2680 2643
rect 2701 2643 2707 2657
rect 2808 2657 2904 2663
rect 2920 2657 2984 2663
rect 3000 2657 3256 2663
rect 3688 2657 3736 2663
rect 3752 2657 4504 2663
rect 4760 2657 5272 2663
rect 5304 2657 5512 2663
rect 5693 2663 5699 2677
rect 5720 2677 5816 2683
rect 6008 2677 6200 2683
rect 6360 2677 6456 2683
rect 6520 2677 6648 2683
rect 5693 2657 6168 2663
rect 6184 2657 6280 2663
rect 6296 2657 6360 2663
rect 6696 2657 6728 2663
rect 2701 2637 3160 2643
rect 3256 2637 3832 2643
rect 3880 2637 4008 2643
rect 4216 2637 4344 2643
rect 4392 2637 4424 2643
rect 4456 2637 4728 2643
rect 4744 2637 4856 2643
rect 5032 2637 5112 2643
rect 5208 2637 5240 2643
rect 5336 2637 5432 2643
rect 5496 2637 5528 2643
rect 5624 2637 6072 2643
rect 1656 2617 1731 2623
rect 1800 2617 1816 2623
rect 344 2597 616 2603
rect 968 2597 1176 2603
rect 1192 2597 1576 2603
rect 1640 2597 1720 2603
rect 2184 2617 2584 2623
rect 2616 2617 3048 2623
rect 3224 2617 3528 2623
rect 3544 2617 3576 2623
rect 3736 2617 3864 2623
rect 2104 2597 2136 2603
rect 2408 2597 2472 2603
rect 2536 2597 2552 2603
rect 2568 2597 2680 2603
rect 2696 2597 3144 2603
rect 3160 2597 3240 2603
rect 3256 2597 3832 2603
rect 3976 2617 4312 2623
rect 4328 2617 4499 2623
rect 4056 2597 4344 2603
rect 4493 2603 4499 2617
rect 4520 2617 4632 2623
rect 4744 2617 4760 2623
rect 4872 2617 5016 2623
rect 5208 2617 5400 2623
rect 5416 2617 5704 2623
rect 5880 2617 5912 2623
rect 4493 2597 5336 2603
rect 5592 2597 5688 2603
rect 6008 2617 6056 2623
rect 6120 2617 6264 2623
rect 6280 2617 6392 2623
rect 6072 2597 6104 2603
rect 6216 2597 6248 2603
rect 2269 2588 2275 2592
rect 152 2577 424 2583
rect 456 2577 472 2583
rect 632 2577 872 2583
rect 1208 2577 1400 2583
rect 1416 2577 1528 2583
rect 1576 2577 1752 2583
rect 1832 2577 2104 2583
rect 2360 2577 2376 2583
rect 2408 2577 2760 2583
rect 2840 2577 2936 2583
rect 2968 2577 3048 2583
rect 3064 2577 3208 2583
rect 3464 2577 3528 2583
rect 3544 2577 4040 2583
rect 4200 2577 4264 2583
rect 4280 2577 4408 2583
rect 4440 2577 4696 2583
rect 4760 2577 5432 2583
rect 5448 2577 5832 2583
rect 5864 2577 6040 2583
rect 6216 2577 6232 2583
rect 6504 2577 6520 2583
rect 488 2557 552 2563
rect 568 2557 680 2563
rect 696 2557 728 2563
rect 744 2557 1128 2563
rect 1144 2557 1240 2563
rect 1512 2557 1800 2563
rect 1816 2557 1944 2563
rect 2104 2557 2360 2563
rect 2376 2557 2760 2563
rect 2776 2557 2872 2563
rect 3128 2557 3144 2563
rect 3496 2557 3544 2563
rect 3912 2557 3976 2563
rect 4648 2557 4664 2563
rect 4840 2557 4856 2563
rect 4984 2557 5064 2563
rect 5272 2557 5416 2563
rect 5432 2557 5640 2563
rect 5960 2557 5992 2563
rect 6056 2557 6328 2563
rect 6365 2557 6472 2563
rect 1501 2548 1507 2552
rect 2973 2548 2979 2552
rect 3837 2548 3843 2552
rect 56 2537 168 2543
rect 472 2537 744 2543
rect 760 2537 1144 2543
rect 1176 2537 1208 2543
rect 1832 2537 1864 2543
rect 1992 2537 2328 2543
rect 2488 2537 2632 2543
rect 3048 2537 3272 2543
rect 3336 2537 3400 2543
rect 3528 2537 3544 2543
rect 3928 2537 3960 2543
rect 4040 2537 4120 2543
rect 4360 2537 4408 2543
rect 4424 2537 4488 2543
rect 4568 2537 4680 2543
rect 5000 2537 5016 2543
rect 5080 2537 5144 2543
rect 5240 2537 5416 2543
rect 5464 2537 5512 2543
rect 5688 2537 5768 2543
rect 6365 2543 6371 2557
rect 6552 2557 6664 2563
rect 6728 2557 6760 2563
rect 5848 2537 6371 2543
rect 6472 2537 6504 2543
rect 6728 2537 6792 2543
rect 120 2517 168 2523
rect 184 2517 440 2523
rect 584 2517 776 2523
rect 792 2517 856 2523
rect 941 2517 952 2523
rect 1256 2517 1560 2523
rect 1656 2517 1704 2523
rect 1768 2517 1896 2523
rect 1912 2517 1928 2523
rect 1976 2517 1992 2523
rect 2040 2517 2168 2523
rect 2232 2517 2264 2523
rect 2600 2517 2680 2523
rect 2712 2517 3000 2523
rect 3064 2517 3384 2523
rect 3400 2517 3560 2523
rect 3640 2517 3720 2523
rect 3736 2517 3896 2523
rect 3960 2517 3976 2523
rect 4056 2517 4168 2523
rect 4184 2517 4328 2523
rect 4360 2517 4376 2523
rect 4712 2517 4744 2523
rect 4776 2517 5400 2523
rect 5672 2517 5800 2523
rect 6024 2517 6072 2523
rect 6136 2517 6200 2523
rect 6344 2517 6392 2523
rect 6408 2517 6488 2523
rect 6504 2517 6616 2523
rect 6680 2517 6712 2523
rect 168 2497 200 2503
rect 360 2497 424 2503
rect 504 2497 680 2503
rect 856 2497 952 2503
rect 1016 2497 1336 2503
rect 1400 2497 1448 2503
rect 1608 2497 2440 2503
rect 2456 2497 2904 2503
rect 2920 2497 3096 2503
rect 3176 2497 3320 2503
rect 3384 2497 3416 2503
rect 3512 2497 3624 2503
rect 3704 2497 3768 2503
rect 3976 2497 4088 2503
rect 4216 2497 4232 2503
rect 4248 2497 4328 2503
rect 4344 2497 4392 2503
rect 4888 2497 5192 2503
rect 5208 2497 5480 2503
rect 5496 2497 5704 2503
rect 5928 2497 6040 2503
rect 6424 2497 6440 2503
rect 6456 2497 6680 2503
rect 1224 2477 1256 2483
rect 1496 2477 1672 2483
rect 1688 2477 1928 2483
rect 1976 2477 2040 2483
rect 2072 2477 2152 2483
rect 2344 2477 2360 2483
rect 2536 2477 2552 2483
rect 2632 2477 2659 2483
rect 360 2457 520 2463
rect 664 2457 760 2463
rect 840 2457 984 2463
rect 1000 2457 1144 2463
rect 1288 2457 1379 2463
rect 424 2437 712 2443
rect 728 2437 1016 2443
rect 1240 2437 1352 2443
rect 1373 2443 1379 2457
rect 1416 2457 1624 2463
rect 2120 2457 2168 2463
rect 2200 2457 2632 2463
rect 2653 2463 2659 2477
rect 2680 2477 2760 2483
rect 2776 2477 2792 2483
rect 2824 2477 2856 2483
rect 3000 2477 3112 2483
rect 3128 2477 3288 2483
rect 3304 2477 3352 2483
rect 3416 2477 3464 2483
rect 3656 2477 3736 2483
rect 3912 2477 3928 2483
rect 4136 2477 4296 2483
rect 4376 2477 4392 2483
rect 4424 2477 4456 2483
rect 4616 2477 5096 2483
rect 5288 2477 5912 2483
rect 5928 2477 6056 2483
rect 6120 2477 6136 2483
rect 6168 2477 6200 2483
rect 6216 2477 6296 2483
rect 6312 2477 6440 2483
rect 2653 2457 2712 2463
rect 2728 2457 2808 2463
rect 2856 2457 3032 2463
rect 3096 2457 3208 2463
rect 3240 2457 3432 2463
rect 3480 2457 3656 2463
rect 3688 2457 4040 2463
rect 4376 2457 4904 2463
rect 4920 2457 5304 2463
rect 5320 2457 5368 2463
rect 5416 2457 6120 2463
rect 1373 2437 1496 2443
rect 2264 2437 2776 2443
rect 2792 2437 3352 2443
rect 3528 2437 4072 2443
rect 4312 2437 4440 2443
rect 4456 2437 4520 2443
rect 4648 2437 4792 2443
rect 4808 2437 5448 2443
rect 5800 2437 6088 2443
rect 6296 2437 6424 2443
rect 5517 2428 5523 2432
rect 264 2417 488 2423
rect 504 2417 584 2423
rect 616 2417 632 2423
rect 232 2397 296 2403
rect 312 2397 408 2403
rect 920 2417 936 2423
rect 1128 2417 1224 2423
rect 1480 2417 1496 2423
rect 2136 2417 2376 2423
rect 2552 2417 2632 2423
rect 1480 2397 1544 2403
rect 1720 2397 1784 2403
rect 2205 2397 2232 2403
rect 328 2377 520 2383
rect 2205 2383 2211 2397
rect 2264 2397 2696 2403
rect 3048 2417 3656 2423
rect 4024 2417 4568 2423
rect 4744 2417 4760 2423
rect 2920 2397 3256 2403
rect 3336 2397 3624 2403
rect 3736 2397 3816 2403
rect 3832 2397 4040 2403
rect 4056 2397 4072 2403
rect 4472 2397 4584 2403
rect 4648 2397 4792 2403
rect 4808 2397 4840 2403
rect 4968 2417 5176 2423
rect 5368 2417 5496 2423
rect 5752 2417 5976 2423
rect 6392 2417 6632 2423
rect 5192 2397 5256 2403
rect 5272 2397 5528 2403
rect 5752 2397 5896 2403
rect 5912 2397 6712 2403
rect 1240 2377 2211 2383
rect 2328 2377 2488 2383
rect 2744 2377 2952 2383
rect 3096 2377 3176 2383
rect 3240 2377 3608 2383
rect 3624 2377 3656 2383
rect 3672 2377 3896 2383
rect 3912 2377 4056 2383
rect 4088 2377 4840 2383
rect 4856 2377 5432 2383
rect 5448 2377 5880 2383
rect 5912 2377 6504 2383
rect 6616 2377 6744 2383
rect 680 2357 840 2363
rect 856 2357 1080 2363
rect 1096 2357 1160 2363
rect 1176 2357 1416 2363
rect 1432 2357 1528 2363
rect 1608 2357 1656 2363
rect 2328 2357 2648 2363
rect 2824 2357 3208 2363
rect 3224 2357 3256 2363
rect 3544 2357 3752 2363
rect 4360 2357 4712 2363
rect 4888 2357 5064 2363
rect 5112 2357 5624 2363
rect 5640 2357 5688 2363
rect 5704 2357 5944 2363
rect 5960 2357 6040 2363
rect 6584 2357 6696 2363
rect 40 2337 72 2343
rect 168 2337 200 2343
rect 232 2337 312 2343
rect 792 2337 1064 2343
rect 1080 2337 1432 2343
rect 1448 2337 1896 2343
rect 2088 2337 2168 2343
rect 2360 2337 2728 2343
rect 3032 2337 3144 2343
rect 3192 2337 3224 2343
rect 3784 2337 3800 2343
rect 4248 2337 4600 2343
rect 4616 2337 4664 2343
rect 4680 2337 5608 2343
rect 6488 2337 6568 2343
rect 72 2317 296 2323
rect 328 2317 408 2323
rect 424 2317 440 2323
rect 536 2317 648 2323
rect 728 2317 776 2323
rect 952 2317 1176 2323
rect 1192 2317 1240 2323
rect 1384 2317 1432 2323
rect 1480 2317 1512 2323
rect 1576 2317 1704 2323
rect 1720 2317 2408 2323
rect 2440 2317 2536 2323
rect 2552 2317 2904 2323
rect 3048 2317 3144 2323
rect 3176 2317 3192 2323
rect 3256 2317 3304 2323
rect 3336 2317 3352 2323
rect 3384 2317 3592 2323
rect 3640 2317 3848 2323
rect 4040 2317 4392 2323
rect 4520 2317 4648 2323
rect 5176 2317 5208 2323
rect 5272 2317 5288 2323
rect 5432 2317 5448 2323
rect 5576 2317 5656 2323
rect 5768 2317 5928 2323
rect 184 2297 360 2303
rect 376 2297 472 2303
rect 664 2297 680 2303
rect 984 2297 1080 2303
rect 1144 2297 1304 2303
rect 1368 2297 1672 2303
rect 1704 2297 1800 2303
rect 1816 2297 1976 2303
rect 2136 2297 2232 2303
rect 2264 2297 2840 2303
rect 2904 2297 2952 2303
rect 2968 2297 3016 2303
rect 3112 2297 3176 2303
rect 3288 2297 3352 2303
rect 3656 2297 3704 2303
rect 3864 2297 3880 2303
rect 3944 2297 4328 2303
rect 4552 2297 4632 2303
rect 4696 2297 4712 2303
rect 5144 2297 5368 2303
rect 5528 2297 5720 2303
rect 5736 2297 5832 2303
rect 5944 2297 5960 2303
rect 6280 2297 6408 2303
rect 6488 2297 6520 2303
rect 6536 2297 6552 2303
rect 6600 2297 6664 2303
rect 104 2277 264 2283
rect 440 2277 472 2283
rect 493 2283 499 2292
rect 5421 2288 5427 2292
rect 493 2277 856 2283
rect 1048 2277 1096 2283
rect 1176 2277 1208 2283
rect 1528 2277 1592 2283
rect 1656 2277 1688 2283
rect 1784 2277 2040 2283
rect 2072 2277 2088 2283
rect 2216 2277 2408 2283
rect 2440 2277 2488 2283
rect 2568 2277 2584 2283
rect 2680 2277 2696 2283
rect 2712 2277 2792 2283
rect 2808 2277 3048 2283
rect 3064 2277 3112 2283
rect 3128 2277 3464 2283
rect 3480 2277 3496 2283
rect 3816 2277 3832 2283
rect 3880 2277 4312 2283
rect 4328 2277 4344 2283
rect 4461 2277 4584 2283
rect 56 2257 440 2263
rect 488 2257 504 2263
rect 536 2257 568 2263
rect 584 2257 728 2263
rect 1128 2257 1208 2263
rect 1384 2257 1400 2263
rect 1416 2257 1544 2263
rect 1560 2257 2008 2263
rect 2040 2257 2600 2263
rect 3096 2257 3336 2263
rect 3528 2257 3976 2263
rect 4461 2263 4467 2277
rect 4600 2277 4648 2283
rect 4680 2277 4712 2283
rect 4776 2277 4808 2283
rect 4824 2277 5080 2283
rect 5112 2277 5272 2283
rect 5288 2277 5320 2283
rect 5512 2277 5608 2283
rect 5784 2277 5896 2283
rect 5912 2277 5976 2283
rect 6408 2277 6424 2283
rect 6552 2277 6776 2283
rect 4040 2257 4467 2263
rect 4488 2257 4520 2263
rect 5064 2257 5224 2263
rect 5240 2257 5560 2263
rect 5672 2257 5864 2263
rect 5976 2257 6072 2263
rect 6104 2257 6440 2263
rect 6504 2257 6552 2263
rect 472 2237 488 2243
rect 504 2237 568 2243
rect 632 2237 776 2243
rect 920 2237 952 2243
rect 968 2237 1032 2243
rect 1464 2237 1576 2243
rect 1592 2237 1784 2243
rect 1800 2237 1880 2243
rect 1944 2237 1976 2243
rect 2056 2237 2072 2243
rect 2088 2237 2200 2243
rect 2232 2237 2344 2243
rect 2408 2237 2600 2243
rect 2616 2237 2632 2243
rect 3208 2237 3640 2243
rect 3656 2237 4024 2243
rect 4200 2237 5336 2243
rect 5352 2237 5560 2243
rect 5576 2237 5736 2243
rect 5864 2237 6088 2243
rect 6120 2237 6232 2243
rect 6248 2237 6296 2243
rect 264 2217 392 2223
rect 408 2217 680 2223
rect 728 2217 904 2223
rect 920 2217 1064 2223
rect 1208 2217 1480 2223
rect 1496 2217 1608 2223
rect 680 2197 712 2203
rect 728 2197 1560 2203
rect 1608 2197 1656 2203
rect 1976 2217 2088 2223
rect 2376 2217 2408 2223
rect 3144 2217 3224 2223
rect 3320 2217 3448 2223
rect 3560 2217 3704 2223
rect 2136 2197 2216 2203
rect 2232 2197 2280 2203
rect 2296 2197 3592 2203
rect 3608 2197 3688 2203
rect 4200 2217 4264 2223
rect 4296 2217 4552 2223
rect 5256 2217 5448 2223
rect 3944 2197 3960 2203
rect 3976 2197 4104 2203
rect 4216 2197 4280 2203
rect 4504 2197 4536 2203
rect 4552 2197 5048 2203
rect 5176 2197 5384 2203
rect 5640 2197 5784 2203
rect 6072 2217 6376 2223
rect 6664 2217 6760 2223
rect 6184 2197 6264 2203
rect 6280 2197 6536 2203
rect 6552 2197 6632 2203
rect 200 2177 216 2183
rect 232 2177 360 2183
rect 504 2177 600 2183
rect 776 2177 856 2183
rect 984 2177 1144 2183
rect 1160 2177 1208 2183
rect 1464 2177 1496 2183
rect 1592 2177 2072 2183
rect 2104 2177 2136 2183
rect 2152 2177 2824 2183
rect 3128 2177 3208 2183
rect 3256 2177 3320 2183
rect 3832 2177 4008 2183
rect 4296 2177 4536 2183
rect 4552 2177 4648 2183
rect 5448 2177 5640 2183
rect 5656 2177 5720 2183
rect 5736 2177 6136 2183
rect 6360 2177 6552 2183
rect 136 2157 280 2163
rect 936 2157 1112 2163
rect 1128 2157 1304 2163
rect 1448 2157 1464 2163
rect 1656 2157 1752 2163
rect 1768 2157 1928 2163
rect 2280 2157 2328 2163
rect 2952 2157 3256 2163
rect 3352 2157 3800 2163
rect 4024 2157 4072 2163
rect 4104 2157 4168 2163
rect 4232 2157 4376 2163
rect 5304 2157 5352 2163
rect 5544 2157 5624 2163
rect 5640 2157 6232 2163
rect 6616 2157 6664 2163
rect 541 2148 547 2152
rect 280 2137 296 2143
rect 328 2137 392 2143
rect 440 2137 520 2143
rect 600 2137 648 2143
rect 776 2137 840 2143
rect 856 2137 1016 2143
rect 1288 2137 1464 2143
rect 1496 2137 1512 2143
rect 1560 2137 1624 2143
rect 1768 2137 2232 2143
rect 2312 2137 2504 2143
rect 2552 2137 2616 2143
rect 2952 2137 3336 2143
rect 3384 2137 3944 2143
rect 3960 2137 3992 2143
rect 4008 2137 4232 2143
rect 4248 2137 4392 2143
rect 4408 2137 4456 2143
rect 4840 2137 4904 2143
rect 5096 2137 5240 2143
rect 5256 2137 5640 2143
rect 5832 2137 5928 2143
rect 5992 2137 6024 2143
rect 6072 2137 6104 2143
rect 6360 2137 6424 2143
rect 6568 2137 6680 2143
rect 6712 2137 6744 2143
rect 248 2117 467 2123
rect 248 2097 280 2103
rect 376 2097 440 2103
rect 461 2103 467 2117
rect 568 2117 616 2123
rect 1245 2123 1251 2132
rect 4829 2128 4835 2132
rect 1245 2117 1256 2123
rect 1288 2117 1304 2123
rect 1416 2117 1608 2123
rect 1656 2117 2088 2123
rect 2104 2117 2392 2123
rect 2440 2117 2456 2123
rect 2680 2117 2776 2123
rect 2808 2117 2840 2123
rect 2856 2117 3080 2123
rect 3160 2117 3208 2123
rect 3304 2117 3352 2123
rect 3400 2117 3464 2123
rect 3565 2117 3576 2123
rect 3517 2108 3523 2112
rect 3565 2108 3571 2117
rect 3688 2117 3736 2123
rect 3752 2117 3848 2123
rect 3992 2117 4072 2123
rect 4173 2117 4184 2123
rect 4440 2117 4595 2123
rect 461 2097 1480 2103
rect 1688 2097 1784 2103
rect 1816 2097 1976 2103
rect 2088 2097 2232 2103
rect 2792 2097 2952 2103
rect 3048 2097 3160 2103
rect 3352 2097 3448 2103
rect 3640 2097 3816 2103
rect 3880 2097 4008 2103
rect 4184 2097 4264 2103
rect 4344 2097 4568 2103
rect 4589 2103 4595 2117
rect 4616 2117 4744 2123
rect 5160 2117 5176 2123
rect 5336 2117 5416 2123
rect 5496 2117 5592 2123
rect 5880 2117 6072 2123
rect 6136 2117 6280 2123
rect 6328 2117 6376 2123
rect 6440 2117 6616 2123
rect 6648 2117 6867 2123
rect 4589 2097 4616 2103
rect 4920 2097 4952 2103
rect 5080 2097 5144 2103
rect 5224 2097 5256 2103
rect 5432 2097 5880 2103
rect 5896 2097 6136 2103
rect 6312 2097 6408 2103
rect 6520 2097 6552 2103
rect 232 2077 248 2083
rect 520 2077 616 2083
rect 632 2077 648 2083
rect 664 2077 1080 2083
rect 1096 2077 1560 2083
rect 1608 2077 1720 2083
rect 1736 2077 1800 2083
rect 2072 2077 2168 2083
rect 2344 2077 2472 2083
rect 2488 2077 2536 2083
rect 2552 2077 2776 2083
rect 2920 2077 3000 2083
rect 3096 2077 3144 2083
rect 3192 2077 3272 2083
rect 3416 2077 3864 2083
rect 4104 2077 4376 2083
rect 4392 2077 4520 2083
rect 4536 2077 4664 2083
rect 4792 2077 4952 2083
rect 5288 2077 5432 2083
rect 5832 2077 5912 2083
rect 6040 2077 6344 2083
rect 1240 2057 2008 2063
rect 2056 2057 2104 2063
rect 2216 2057 2248 2063
rect 2264 2057 2552 2063
rect 2904 2057 2952 2063
rect 3032 2057 3224 2063
rect 3272 2057 3656 2063
rect 3672 2057 4088 2063
rect 4104 2057 4152 2063
rect 4296 2057 4424 2063
rect 4440 2057 4488 2063
rect 4504 2057 4552 2063
rect 4600 2057 4632 2063
rect 4664 2057 5032 2063
rect 5048 2057 5224 2063
rect 5240 2057 5384 2063
rect 6104 2057 6472 2063
rect 6488 2057 6792 2063
rect 285 2037 296 2043
rect 285 2028 291 2037
rect 1000 2037 1016 2043
rect 1032 2037 1096 2043
rect 1112 2037 1448 2043
rect 1496 2037 1800 2043
rect 1816 2037 2472 2043
rect 3304 2037 3400 2043
rect 3656 2037 4424 2043
rect 4440 2037 4456 2043
rect 4792 2037 5064 2043
rect 5080 2037 5192 2043
rect 5224 2037 5304 2043
rect 5320 2037 5768 2043
rect 1416 2017 1496 2023
rect 1528 2017 1816 2023
rect 2088 2017 2392 2023
rect 1160 1997 1176 2003
rect 1192 1997 2264 2003
rect 2424 1997 2440 2003
rect 2952 2017 2984 2023
rect 3080 2017 3544 2023
rect 4136 2017 4248 2023
rect 4264 2017 4440 2023
rect 3416 1997 3528 2003
rect 3608 1997 3768 2003
rect 4152 1997 4472 2003
rect 4536 1997 4824 2003
rect 5208 2017 5224 2023
rect 5368 2017 5656 2023
rect 5128 1997 5416 2003
rect 5560 1997 5576 2003
rect 5704 1997 6232 2003
rect 6248 1997 6632 2003
rect 440 1977 584 1983
rect 744 1977 936 1983
rect 952 1977 1128 1983
rect 2008 1977 3096 1983
rect 3336 1977 4136 1983
rect 4456 1977 4536 1983
rect 4744 1977 5704 1983
rect 5720 1977 5864 1983
rect 6024 1977 6088 1983
rect 120 1957 264 1963
rect 760 1957 824 1963
rect 1016 1957 1064 1963
rect 1352 1957 1400 1963
rect 1480 1957 1592 1963
rect 1704 1957 2056 1963
rect 2088 1957 2264 1963
rect 2776 1957 3176 1963
rect 3224 1957 3320 1963
rect 3384 1957 3592 1963
rect 4248 1957 5048 1963
rect 5064 1957 5880 1963
rect 5944 1957 6088 1963
rect 408 1937 456 1943
rect 504 1937 552 1943
rect 664 1937 744 1943
rect 776 1937 856 1943
rect 888 1937 1032 1943
rect 1272 1937 1656 1943
rect 1896 1937 2328 1943
rect 2344 1937 2360 1943
rect 2440 1937 2632 1943
rect 2648 1937 2760 1943
rect 2776 1937 2808 1943
rect 2856 1937 2904 1943
rect 2936 1937 2968 1943
rect 2984 1937 3064 1943
rect 3144 1937 3240 1943
rect 3352 1937 3528 1943
rect 4056 1937 4296 1943
rect 4344 1937 4408 1943
rect 4776 1937 5720 1943
rect 5736 1937 5880 1943
rect 5896 1937 6040 1943
rect 6104 1937 6168 1943
rect 6520 1937 6696 1943
rect 6712 1937 6728 1943
rect 216 1917 312 1923
rect 440 1917 536 1923
rect 568 1917 632 1923
rect 680 1917 840 1923
rect 856 1917 1128 1923
rect 1144 1917 1288 1923
rect 1400 1917 1448 1923
rect 1464 1917 1528 1923
rect 1576 1917 1704 1923
rect 1976 1917 2056 1923
rect 2408 1917 2616 1923
rect 2632 1917 3032 1923
rect 3080 1917 3288 1923
rect 4008 1917 4104 1923
rect 4248 1917 4264 1923
rect 4376 1917 4408 1923
rect 4728 1917 4776 1923
rect 4920 1917 5000 1923
rect 5368 1917 6024 1923
rect 6088 1917 6152 1923
rect 6536 1917 6712 1923
rect 2077 1908 2083 1912
rect 3981 1908 3987 1912
rect 248 1897 328 1903
rect 360 1897 376 1903
rect 424 1897 520 1903
rect 552 1897 600 1903
rect 696 1897 888 1903
rect 920 1897 1192 1903
rect 1208 1897 1480 1903
rect 1528 1897 1560 1903
rect 1608 1897 1672 1903
rect 1848 1897 1864 1903
rect 1896 1897 2040 1903
rect 2301 1897 2312 1903
rect 2344 1897 2456 1903
rect 2472 1897 2568 1903
rect 2616 1897 2664 1903
rect 2712 1897 3128 1903
rect 3144 1897 3208 1903
rect 3528 1897 3640 1903
rect 4024 1897 4040 1903
rect 4216 1897 4312 1903
rect 4824 1897 4968 1903
rect 5256 1897 5464 1903
rect 5576 1897 5736 1903
rect 5768 1897 5800 1903
rect 5992 1897 6040 1903
rect 6168 1897 6248 1903
rect 6616 1897 6632 1903
rect 2685 1888 2691 1892
rect 4605 1888 4611 1892
rect 280 1877 344 1883
rect 536 1877 552 1883
rect 744 1877 776 1883
rect 856 1877 968 1883
rect 1064 1877 1096 1883
rect 1192 1877 1352 1883
rect 1368 1877 1384 1883
rect 1432 1877 1464 1883
rect 1752 1877 1784 1883
rect 1864 1877 1896 1883
rect 1928 1877 2152 1883
rect 2184 1877 2216 1883
rect 2712 1877 2728 1883
rect 2744 1877 2840 1883
rect 3016 1877 3064 1883
rect 3128 1877 3160 1883
rect 3176 1877 3240 1883
rect 3256 1877 3672 1883
rect 3688 1877 3928 1883
rect 3960 1877 4120 1883
rect 4264 1877 4552 1883
rect 4696 1877 4888 1883
rect 5112 1877 5160 1883
rect 5176 1877 5192 1883
rect 5352 1877 5384 1883
rect 5496 1877 5848 1883
rect 6136 1877 6600 1883
rect 6664 1877 6712 1883
rect 205 1868 211 1872
rect 669 1868 675 1872
rect 4237 1868 4243 1872
rect 328 1857 392 1863
rect 408 1857 616 1863
rect 920 1857 952 1863
rect 968 1857 1048 1863
rect 1064 1857 1448 1863
rect 1560 1857 1592 1863
rect 1848 1857 1928 1863
rect 2008 1857 2120 1863
rect 2168 1857 2360 1863
rect 2760 1857 2856 1863
rect 2936 1857 2952 1863
rect 2968 1857 3192 1863
rect 3256 1857 3624 1863
rect 3640 1857 4056 1863
rect 4264 1857 4280 1863
rect 4584 1857 5032 1863
rect 5064 1857 5464 1863
rect 5800 1857 5928 1863
rect 6424 1857 6536 1863
rect 6552 1857 6744 1863
rect 296 1837 456 1843
rect 648 1837 664 1843
rect 1384 1837 1400 1843
rect 1432 1837 1640 1843
rect 1688 1837 2264 1843
rect 2280 1837 2328 1843
rect 2360 1837 2376 1843
rect 2392 1837 2408 1843
rect 2424 1837 2536 1843
rect 2792 1837 3080 1843
rect 3208 1837 3368 1843
rect 3576 1837 3784 1843
rect 4056 1837 4088 1843
rect 4104 1837 4184 1843
rect 4376 1837 4952 1843
rect 5096 1837 5272 1843
rect 5288 1837 5368 1843
rect 5384 1837 5496 1843
rect 5816 1837 6104 1843
rect 6456 1837 6472 1843
rect 6568 1837 6616 1843
rect 6648 1837 6696 1843
rect 296 1817 360 1823
rect 616 1817 1720 1823
rect 424 1797 632 1803
rect 648 1797 968 1803
rect 1016 1797 1400 1803
rect 1416 1797 1432 1803
rect 1592 1797 1736 1803
rect 2760 1817 2936 1823
rect 3144 1817 3496 1823
rect 3720 1817 3816 1823
rect 1896 1797 1960 1803
rect 2136 1797 2200 1803
rect 2504 1797 2744 1803
rect 2824 1797 3016 1803
rect 3032 1797 3080 1803
rect 3112 1797 3272 1803
rect 3288 1797 3560 1803
rect 3976 1817 4120 1823
rect 4600 1817 4840 1823
rect 5720 1817 5832 1823
rect 5101 1808 5107 1812
rect 3944 1797 3976 1803
rect 4088 1797 4264 1803
rect 4280 1797 4424 1803
rect 4440 1797 4616 1803
rect 4648 1797 4776 1803
rect 4792 1797 4808 1803
rect 5112 1797 5224 1803
rect 5240 1797 5272 1803
rect 5352 1797 5400 1803
rect 5464 1797 5688 1803
rect 6104 1817 6376 1823
rect 6600 1817 6760 1823
rect 6056 1797 6120 1803
rect 6136 1797 6232 1803
rect 6472 1797 6664 1803
rect 2445 1788 2451 1792
rect 600 1777 648 1783
rect 760 1777 1064 1783
rect 1309 1777 1320 1783
rect 1640 1777 2312 1783
rect 2376 1777 2440 1783
rect 2472 1777 2728 1783
rect 2744 1777 2888 1783
rect 2904 1777 3048 1783
rect 3272 1777 3384 1783
rect 3480 1777 3624 1783
rect 3640 1777 3656 1783
rect 3672 1777 3768 1783
rect 3896 1777 4056 1783
rect 4120 1777 4552 1783
rect 4600 1777 4744 1783
rect 4792 1777 5000 1783
rect 5016 1777 5144 1783
rect 5224 1777 5464 1783
rect 5672 1777 5720 1783
rect 5848 1777 6008 1783
rect 6024 1777 6216 1783
rect 216 1757 232 1763
rect 376 1757 424 1763
rect 872 1757 1176 1763
rect 1320 1757 1560 1763
rect 1592 1757 1640 1763
rect 1672 1757 1752 1763
rect 1784 1757 1880 1763
rect 2088 1757 2248 1763
rect 2328 1757 2792 1763
rect 2952 1757 3000 1763
rect 3064 1757 3112 1763
rect 3240 1757 3416 1763
rect 3576 1757 3960 1763
rect 3992 1757 4104 1763
rect 4120 1757 4296 1763
rect 4504 1757 4600 1763
rect 4616 1757 4728 1763
rect 4904 1757 4984 1763
rect 5000 1757 5112 1763
rect 5224 1757 5384 1763
rect 5496 1757 5512 1763
rect 5624 1757 5768 1763
rect 5880 1757 6104 1763
rect 6120 1757 6360 1763
rect 6456 1757 6712 1763
rect 253 1748 259 1752
rect 1048 1737 1064 1743
rect 1432 1737 1448 1743
rect 1544 1737 1592 1743
rect 1624 1737 1688 1743
rect 1864 1737 1896 1743
rect 1976 1737 2088 1743
rect 2200 1737 2216 1743
rect 2616 1737 2680 1743
rect 2712 1737 2776 1743
rect 2808 1737 3016 1743
rect 3816 1737 4083 1743
rect 456 1717 760 1723
rect 904 1717 1112 1723
rect 1288 1717 1304 1723
rect 1501 1723 1507 1732
rect 3357 1728 3363 1732
rect 1496 1717 1507 1723
rect 1528 1717 1688 1723
rect 1704 1717 1752 1723
rect 2040 1717 2088 1723
rect 2200 1717 2232 1723
rect 2312 1717 2328 1723
rect 2408 1717 2760 1723
rect 3224 1717 3336 1723
rect 3421 1723 3427 1732
rect 3709 1728 3715 1732
rect 3416 1717 3427 1723
rect 3800 1717 3864 1723
rect 4024 1717 4056 1723
rect 4077 1723 4083 1737
rect 4264 1737 4296 1743
rect 4552 1737 4904 1743
rect 5032 1737 5304 1743
rect 5432 1737 5624 1743
rect 5704 1737 5800 1743
rect 5832 1737 5864 1743
rect 5896 1737 6056 1743
rect 6344 1737 6440 1743
rect 6456 1737 6504 1743
rect 6584 1737 6616 1743
rect 4077 1717 4104 1723
rect 4312 1717 4371 1723
rect 248 1697 376 1703
rect 408 1697 488 1703
rect 552 1697 584 1703
rect 600 1697 696 1703
rect 728 1697 824 1703
rect 840 1697 968 1703
rect 1005 1697 1016 1703
rect 1048 1697 1080 1703
rect 1288 1697 1384 1703
rect 1400 1697 1896 1703
rect 1960 1697 2840 1703
rect 2872 1697 3208 1703
rect 3272 1697 3288 1703
rect 3320 1697 3496 1703
rect 3832 1697 3928 1703
rect 3976 1697 3992 1703
rect 4136 1697 4152 1703
rect 4168 1697 4200 1703
rect 4296 1697 4344 1703
rect 4365 1703 4371 1717
rect 4408 1717 4456 1723
rect 4504 1717 4712 1723
rect 4792 1717 4840 1723
rect 5080 1717 5112 1723
rect 5160 1717 5256 1723
rect 5400 1717 5496 1723
rect 5512 1717 5528 1723
rect 5544 1717 5848 1723
rect 5944 1717 5992 1723
rect 6424 1717 6632 1723
rect 4365 1697 4504 1703
rect 4760 1697 5176 1703
rect 5192 1697 5656 1703
rect 5752 1697 5896 1703
rect 5912 1697 6040 1703
rect 6056 1697 6168 1703
rect 344 1677 888 1683
rect 1128 1677 1576 1683
rect 1592 1677 1688 1683
rect 1704 1677 1864 1683
rect 1880 1677 1992 1683
rect 2680 1677 2856 1683
rect 3176 1677 3272 1683
rect 3352 1677 3416 1683
rect 3480 1677 3528 1683
rect 3752 1677 3960 1683
rect 4488 1677 4520 1683
rect 4840 1677 4872 1683
rect 5432 1677 5544 1683
rect 5848 1677 5944 1683
rect 6040 1677 6248 1683
rect 376 1657 456 1663
rect 472 1657 680 1663
rect 696 1657 776 1663
rect 792 1657 1064 1663
rect 1080 1657 1240 1663
rect 1608 1657 1976 1663
rect 1992 1657 2200 1663
rect 2360 1657 3336 1663
rect 3352 1657 3400 1663
rect 3432 1657 3576 1663
rect 3608 1657 3768 1663
rect 3880 1657 3928 1663
rect 3960 1657 4040 1663
rect 4056 1657 4216 1663
rect 4280 1657 5080 1663
rect 5336 1657 5400 1663
rect 5816 1657 6152 1663
rect 6168 1657 6488 1663
rect 6504 1657 6600 1663
rect 488 1637 520 1643
rect 616 1637 680 1643
rect 776 1637 968 1643
rect 1240 1637 1352 1643
rect 1576 1637 1624 1643
rect 1640 1637 1928 1643
rect 1944 1637 1976 1643
rect 2296 1637 2312 1643
rect 2632 1637 2696 1643
rect 2888 1637 2936 1643
rect 3128 1637 3368 1643
rect 3400 1637 4120 1643
rect 4376 1637 4520 1643
rect 4536 1637 4648 1643
rect 4664 1637 5096 1643
rect 5112 1637 5352 1643
rect 5896 1637 6040 1643
rect 360 1597 424 1603
rect 1112 1617 1224 1623
rect 1400 1617 1528 1623
rect 1624 1617 2008 1623
rect 2056 1617 2696 1623
rect 952 1597 1064 1603
rect 1080 1597 1480 1603
rect 1496 1597 1960 1603
rect 2024 1597 2104 1603
rect 3304 1617 3544 1623
rect 3656 1617 3848 1623
rect 3869 1617 3992 1623
rect 3016 1597 3160 1603
rect 3192 1597 3400 1603
rect 3869 1603 3875 1617
rect 4008 1617 4136 1623
rect 4280 1617 4312 1623
rect 4328 1617 4360 1623
rect 4488 1617 4552 1623
rect 3864 1597 3875 1603
rect 3885 1597 4232 1603
rect 120 1577 200 1583
rect 296 1577 792 1583
rect 808 1577 1096 1583
rect 1192 1577 1672 1583
rect 1752 1577 2104 1583
rect 2296 1577 2344 1583
rect 2536 1577 3144 1583
rect 3885 1583 3891 1597
rect 4312 1597 4376 1603
rect 4568 1597 4584 1603
rect 4600 1597 4616 1603
rect 4632 1597 4680 1603
rect 5240 1617 5448 1623
rect 5928 1597 6168 1603
rect 6216 1597 6376 1603
rect 3176 1577 3891 1583
rect 3976 1577 4312 1583
rect 4344 1577 4584 1583
rect 4888 1577 4952 1583
rect 5640 1577 5800 1583
rect 5816 1577 5912 1583
rect 6024 1577 6312 1583
rect 6440 1577 6472 1583
rect 136 1557 216 1563
rect 904 1557 2040 1563
rect 2280 1557 2392 1563
rect 2680 1557 2776 1563
rect 2872 1557 2904 1563
rect 3304 1557 3464 1563
rect 3480 1557 3528 1563
rect 3672 1557 3704 1563
rect 3784 1557 4040 1563
rect 4061 1557 4744 1563
rect -51 1537 120 1543
rect 248 1537 376 1543
rect 552 1537 744 1543
rect 920 1537 1016 1543
rect 1032 1537 1128 1543
rect 1368 1537 1416 1543
rect 1432 1537 1512 1543
rect 1528 1537 1656 1543
rect 2776 1537 2968 1543
rect 2984 1537 3224 1543
rect 3432 1537 3560 1543
rect 4061 1543 4067 1557
rect 4840 1557 4920 1563
rect 4936 1557 5336 1563
rect 5352 1557 5688 1563
rect 5864 1557 6024 1563
rect 6056 1557 6408 1563
rect 3576 1537 4067 1543
rect 4088 1537 4264 1543
rect 4360 1537 4680 1543
rect 4760 1537 5608 1543
rect 5864 1537 6200 1543
rect 6424 1537 6600 1543
rect 6616 1537 6744 1543
rect 328 1517 408 1523
rect 600 1517 632 1523
rect 728 1517 760 1523
rect 840 1517 952 1523
rect 984 1517 1464 1523
rect 1544 1517 1608 1523
rect 1624 1517 2168 1523
rect 2264 1517 2312 1523
rect 2328 1517 2360 1523
rect 2504 1517 2616 1523
rect 2712 1517 2808 1523
rect 2840 1517 3960 1523
rect 3992 1517 4008 1523
rect 4040 1517 4136 1523
rect 4184 1517 4216 1523
rect 4248 1517 4312 1523
rect 4328 1517 4536 1523
rect 4568 1517 4648 1523
rect 4680 1517 4712 1523
rect 4728 1517 4776 1523
rect 5080 1517 5112 1523
rect 5144 1517 5176 1523
rect 5368 1517 5448 1523
rect 5480 1517 5512 1523
rect 5672 1517 5752 1523
rect 5784 1517 5800 1523
rect 6120 1517 6136 1523
rect 6152 1517 6184 1523
rect 6216 1517 6243 1523
rect -51 1497 8 1503
rect 248 1497 264 1503
rect 392 1497 440 1503
rect 552 1497 616 1503
rect 856 1497 888 1503
rect 1304 1497 1336 1503
rect 1464 1497 1544 1503
rect 1848 1497 2040 1503
rect 2216 1497 2408 1503
rect 2424 1497 3080 1503
rect 3288 1497 3304 1503
rect 3528 1497 3544 1503
rect 3704 1497 3784 1503
rect 3837 1497 3848 1503
rect 3912 1497 4248 1503
rect 4264 1497 4376 1503
rect 4408 1497 4504 1503
rect 4589 1497 4632 1503
rect 477 1477 632 1483
rect -51 1457 88 1463
rect 216 1457 264 1463
rect 280 1457 312 1463
rect 477 1463 483 1477
rect 749 1477 760 1483
rect 968 1477 1048 1483
rect 1080 1477 1160 1483
rect 1176 1477 1704 1483
rect 1832 1477 2040 1483
rect 2344 1477 2360 1483
rect 2424 1477 2632 1483
rect 2648 1477 2664 1483
rect 2936 1477 3096 1483
rect 3368 1477 3672 1483
rect 3688 1477 3752 1483
rect 3800 1477 3896 1483
rect 4008 1477 4056 1483
rect 4104 1477 4152 1483
rect 4360 1477 4376 1483
rect 4589 1483 4595 1497
rect 4920 1497 5128 1503
rect 5256 1497 5848 1503
rect 5885 1497 6072 1503
rect 4685 1488 4691 1492
rect 4733 1488 4739 1492
rect 4472 1477 4595 1483
rect 4616 1477 4664 1483
rect 4776 1477 5208 1483
rect 5432 1477 5464 1483
rect 5608 1477 5640 1483
rect 5656 1477 5736 1483
rect 5885 1483 5891 1497
rect 6237 1503 6243 1517
rect 6280 1517 6424 1523
rect 6237 1497 6280 1503
rect 6712 1497 6728 1503
rect 6744 1497 6760 1503
rect 5816 1477 5891 1483
rect 5912 1477 5960 1483
rect 5976 1477 6296 1483
rect 6408 1477 6520 1483
rect 6600 1477 6696 1483
rect 4429 1468 4435 1472
rect 328 1457 483 1463
rect 504 1457 744 1463
rect 1448 1457 1528 1463
rect 2008 1457 2312 1463
rect 2328 1457 2424 1463
rect 2456 1457 2472 1463
rect 2488 1457 3208 1463
rect 3288 1457 3432 1463
rect 3448 1457 3560 1463
rect 3608 1457 3688 1463
rect 3752 1457 3864 1463
rect 4008 1457 4248 1463
rect 4504 1457 4696 1463
rect 4712 1457 5384 1463
rect 5400 1457 5928 1463
rect 5944 1457 6376 1463
rect 6392 1457 6456 1463
rect 6712 1457 6728 1463
rect 536 1437 568 1443
rect 616 1437 760 1443
rect 968 1437 984 1443
rect 1560 1437 1608 1443
rect 1736 1437 2408 1443
rect 2440 1437 2728 1443
rect 2760 1437 3208 1443
rect 3704 1437 3800 1443
rect 3816 1437 3944 1443
rect 4056 1437 4264 1443
rect 4664 1437 5128 1443
rect 5304 1437 5528 1443
rect 5832 1437 6120 1443
rect 6200 1437 6248 1443
rect 184 1417 696 1423
rect 712 1417 1096 1423
rect 1112 1417 1304 1423
rect 1400 1417 1448 1423
rect 1464 1417 1592 1423
rect 1608 1417 1800 1423
rect 136 1397 328 1403
rect 648 1397 888 1403
rect 1128 1397 1304 1403
rect 1336 1397 1464 1403
rect 1480 1397 1496 1403
rect 1512 1397 1688 1403
rect 1992 1417 2168 1423
rect 2344 1417 2584 1423
rect 3208 1417 3672 1423
rect 2072 1397 2120 1403
rect 2200 1397 2584 1403
rect 2952 1397 3016 1403
rect 3032 1397 3496 1403
rect 3528 1397 3576 1403
rect 3992 1417 4104 1423
rect 4184 1417 4312 1423
rect 4552 1417 4792 1423
rect 4840 1417 4984 1423
rect 5384 1417 5640 1423
rect 3944 1397 4072 1403
rect 4136 1397 4952 1403
rect 4968 1397 4984 1403
rect 5000 1397 5144 1403
rect 5208 1397 5416 1403
rect 5496 1397 5635 1403
rect 605 1388 611 1392
rect 632 1377 840 1383
rect 984 1377 1144 1383
rect 1224 1377 1736 1383
rect 2392 1377 2520 1383
rect 3000 1377 3064 1383
rect 3192 1377 3272 1383
rect 3448 1377 3512 1383
rect 3560 1377 3752 1383
rect 4056 1377 4088 1383
rect 4104 1377 4168 1383
rect 4216 1377 4232 1383
rect 4488 1377 4600 1383
rect 4712 1377 5016 1383
rect 5048 1377 5352 1383
rect 5544 1377 5576 1383
rect 5592 1377 5608 1383
rect 5629 1383 5635 1397
rect 5704 1397 5768 1403
rect 6232 1417 6440 1423
rect 6184 1397 6344 1403
rect 6440 1397 6504 1403
rect 6520 1397 6728 1403
rect 5629 1377 5784 1383
rect 5912 1377 6008 1383
rect 6120 1377 6168 1383
rect 6344 1377 6616 1383
rect -51 1357 136 1363
rect 376 1357 392 1363
rect 792 1357 1160 1363
rect 1304 1357 1544 1363
rect 1576 1357 1624 1363
rect 2088 1357 2104 1363
rect 2184 1357 2200 1363
rect 2360 1357 2600 1363
rect 3320 1357 3368 1363
rect 3480 1357 3592 1363
rect 3640 1357 3784 1363
rect 3800 1357 3928 1363
rect 4696 1357 4952 1363
rect 5208 1357 5240 1363
rect 5496 1357 5523 1363
rect 120 1337 280 1343
rect 328 1337 440 1343
rect 696 1337 856 1343
rect 872 1337 888 1343
rect 936 1337 1064 1343
rect 1160 1337 1256 1343
rect 1272 1337 1336 1343
rect 1432 1337 1560 1343
rect 1688 1337 1736 1343
rect 1768 1337 1912 1343
rect 2008 1337 2296 1343
rect 2824 1337 2920 1343
rect 2936 1337 3096 1343
rect 3448 1337 3480 1343
rect 3496 1337 3688 1343
rect 3704 1337 3928 1343
rect 3949 1343 3955 1352
rect 3949 1337 3960 1343
rect 4072 1337 4136 1343
rect 4184 1337 4632 1343
rect 4696 1337 4712 1343
rect 4728 1337 4776 1343
rect 5032 1337 5123 1343
rect -51 1317 8 1323
rect 200 1317 264 1323
rect 904 1317 936 1323
rect 1352 1317 1400 1323
rect 1480 1317 1512 1323
rect 1592 1317 1912 1323
rect 2168 1317 2264 1323
rect 2456 1317 2504 1323
rect 2648 1317 2744 1323
rect 2808 1317 2819 1323
rect 2872 1317 3000 1323
rect 3048 1317 3064 1323
rect 3080 1317 3192 1323
rect 3320 1317 3400 1323
rect 3464 1317 3480 1323
rect 3688 1317 3768 1323
rect 3928 1317 3976 1323
rect 4120 1317 4616 1323
rect 4680 1317 4696 1323
rect 5048 1317 5064 1323
rect 5117 1323 5123 1337
rect 5144 1337 5256 1343
rect 5272 1337 5496 1343
rect 5517 1343 5523 1357
rect 5544 1357 5704 1363
rect 5736 1357 5928 1363
rect 6168 1357 6472 1363
rect 6664 1357 6728 1363
rect 5517 1337 6024 1343
rect 6152 1337 6328 1343
rect 6408 1337 6440 1343
rect 6600 1337 6632 1343
rect 6525 1328 6531 1332
rect 5117 1317 5144 1323
rect 5288 1317 5336 1323
rect 5432 1317 5448 1323
rect 5464 1317 5576 1323
rect 6088 1317 6152 1323
rect 6168 1317 6280 1323
rect 6312 1317 6488 1323
rect 6568 1317 6600 1323
rect 6728 1317 6744 1323
rect 760 1297 920 1303
rect 1304 1297 1592 1303
rect 1608 1297 1928 1303
rect 2248 1297 2344 1303
rect 2728 1297 2824 1303
rect 2840 1297 3144 1303
rect 3672 1297 3688 1303
rect 3736 1297 4008 1303
rect 4104 1297 4168 1303
rect 4408 1297 4472 1303
rect 5016 1297 5080 1303
rect 5160 1297 5400 1303
rect 5496 1297 5528 1303
rect 5592 1297 5656 1303
rect 5704 1297 5832 1303
rect 5848 1297 5896 1303
rect 5928 1297 6248 1303
rect 6472 1297 6680 1303
rect 6712 1297 6776 1303
rect 56 1277 248 1283
rect 792 1277 1048 1283
rect 1336 1277 1544 1283
rect 1565 1277 2024 1283
rect 264 1257 376 1263
rect 1565 1263 1571 1277
rect 2072 1277 3384 1283
rect 3400 1277 3560 1283
rect 3592 1277 3848 1283
rect 3864 1277 4216 1283
rect 4360 1277 4856 1283
rect 5016 1277 5208 1283
rect 5320 1277 5896 1283
rect 6264 1277 6552 1283
rect 1272 1257 1571 1263
rect 2136 1257 2472 1263
rect 2776 1257 2872 1263
rect 2888 1257 3048 1263
rect 3384 1257 3992 1263
rect 4040 1257 4632 1263
rect 4872 1257 5592 1263
rect 6088 1257 6120 1263
rect 6136 1257 6424 1263
rect 6440 1257 6600 1263
rect 376 1237 808 1243
rect 1208 1237 1368 1243
rect 1544 1237 1560 1243
rect 1992 1237 2040 1243
rect 2952 1237 3000 1243
rect 3208 1237 3320 1243
rect 3336 1237 3608 1243
rect 3672 1237 4120 1243
rect 5128 1237 5208 1243
rect 5224 1237 5240 1243
rect 5272 1237 5320 1243
rect 5336 1237 5368 1243
rect 904 1217 1032 1223
rect 1048 1217 1272 1223
rect 1288 1217 1304 1223
rect 1384 1217 1507 1223
rect 968 1197 1480 1203
rect 1501 1203 1507 1217
rect 1800 1217 2488 1223
rect 1501 1197 2536 1203
rect 3032 1217 3112 1223
rect 3128 1217 3624 1223
rect 3880 1217 4264 1223
rect 4296 1217 4808 1223
rect 3000 1197 3016 1203
rect 3064 1197 3112 1203
rect 3224 1197 3528 1203
rect 3544 1197 4296 1203
rect 4312 1197 4696 1203
rect 5944 1217 6360 1223
rect 4984 1197 5240 1203
rect 5480 1197 6168 1203
rect 152 1177 328 1183
rect 344 1177 376 1183
rect 392 1177 2072 1183
rect 2520 1177 3416 1183
rect 3960 1177 3976 1183
rect 3992 1177 4296 1183
rect 4504 1177 4600 1183
rect 4856 1177 5064 1183
rect 5192 1177 5928 1183
rect 6504 1177 6552 1183
rect 6568 1177 6696 1183
rect 40 1157 184 1163
rect 392 1157 424 1163
rect 440 1157 456 1163
rect 472 1157 840 1163
rect 856 1157 1288 1163
rect 1304 1157 1608 1163
rect 2168 1157 2200 1163
rect 2216 1157 2680 1163
rect 2760 1157 2824 1163
rect 2984 1157 3144 1163
rect 3192 1157 3288 1163
rect 3528 1157 3736 1163
rect 3800 1157 4040 1163
rect 4136 1157 4200 1163
rect 4312 1157 4888 1163
rect 4904 1157 5128 1163
rect 5144 1157 5480 1163
rect 5496 1157 5528 1163
rect 5544 1157 5848 1163
rect 6248 1157 6264 1163
rect 6504 1157 6760 1163
rect 56 1137 232 1143
rect 584 1137 616 1143
rect 632 1137 744 1143
rect 760 1137 2328 1143
rect 2344 1137 2632 1143
rect 2648 1137 3080 1143
rect 3160 1137 3832 1143
rect 3848 1137 4056 1143
rect 4136 1137 4392 1143
rect 4488 1137 4760 1143
rect 4776 1137 4968 1143
rect 5000 1137 5080 1143
rect 5416 1137 5448 1143
rect 5464 1137 5544 1143
rect 5560 1137 5592 1143
rect 5608 1137 5656 1143
rect 5784 1137 5800 1143
rect 6216 1137 6232 1143
rect 6317 1137 6472 1143
rect 168 1117 264 1123
rect 280 1117 312 1123
rect 456 1117 488 1123
rect 520 1117 856 1123
rect 872 1117 920 1123
rect 984 1117 1048 1123
rect 1080 1117 1464 1123
rect 2040 1117 2280 1123
rect 2472 1117 2664 1123
rect 2680 1117 2712 1123
rect 2776 1117 2984 1123
rect 3048 1117 3512 1123
rect 3592 1117 3768 1123
rect 4248 1117 4328 1123
rect 4376 1117 4424 1123
rect 4824 1117 5176 1123
rect 5320 1117 5384 1123
rect 5688 1117 5736 1123
rect 5880 1117 6216 1123
rect 6317 1123 6323 1137
rect 6232 1117 6323 1123
rect 6344 1117 6392 1123
rect 6408 1117 6440 1123
rect 3869 1108 3875 1112
rect 56 1097 88 1103
rect 232 1097 280 1103
rect 440 1097 472 1103
rect 744 1097 1336 1103
rect 1368 1097 1544 1103
rect 1624 1097 1672 1103
rect 1720 1097 1768 1103
rect 1816 1097 1832 1103
rect 1848 1097 1864 1103
rect 1944 1097 1955 1103
rect 1976 1097 2040 1103
rect 2104 1097 2120 1103
rect 2296 1097 2456 1103
rect 2520 1097 2664 1103
rect 2760 1097 2776 1103
rect 2829 1097 2856 1103
rect 88 1077 136 1083
rect 200 1077 1032 1083
rect 1048 1077 1224 1083
rect 1240 1077 1576 1083
rect 1656 1077 1736 1083
rect 1752 1077 2216 1083
rect 2248 1077 2392 1083
rect 2408 1077 2536 1083
rect 2829 1083 2835 1097
rect 3144 1097 3176 1103
rect 3272 1097 3352 1103
rect 3368 1097 3656 1103
rect 3880 1097 4568 1103
rect 4893 1097 5512 1103
rect 2584 1077 2835 1083
rect 2856 1077 3048 1083
rect 3544 1077 3752 1083
rect 3944 1077 4088 1083
rect 4136 1077 4627 1083
rect 328 1057 648 1063
rect 664 1057 952 1063
rect 989 1057 1016 1063
rect 280 1037 392 1043
rect 477 1037 488 1043
rect 477 1028 483 1037
rect 776 1037 920 1043
rect 989 1043 995 1057
rect 1064 1057 1208 1063
rect 1256 1057 1368 1063
rect 1400 1057 1464 1063
rect 1480 1057 1560 1063
rect 1688 1057 1704 1063
rect 1725 1057 2099 1063
rect 952 1037 995 1043
rect 1016 1037 1112 1043
rect 1176 1037 1288 1043
rect 1725 1043 1731 1057
rect 1368 1037 1731 1043
rect 1832 1037 1896 1043
rect 2093 1043 2099 1057
rect 2264 1057 2424 1063
rect 2456 1057 2776 1063
rect 2792 1057 2872 1063
rect 2984 1057 3000 1063
rect 3064 1057 3112 1063
rect 3144 1057 3432 1063
rect 3704 1057 4040 1063
rect 4232 1057 4600 1063
rect 4621 1063 4627 1077
rect 4893 1083 4899 1097
rect 5528 1097 5880 1103
rect 6072 1097 6280 1103
rect 6360 1097 6568 1103
rect 6584 1097 6632 1103
rect 4648 1077 4899 1083
rect 4984 1077 5160 1083
rect 5176 1077 5304 1083
rect 5400 1077 5528 1083
rect 5544 1077 5656 1083
rect 5768 1077 5784 1083
rect 5848 1077 6019 1083
rect 5373 1068 5379 1072
rect 4621 1057 4776 1063
rect 4952 1057 5016 1063
rect 5736 1057 5880 1063
rect 6013 1063 6019 1077
rect 6040 1077 6216 1083
rect 6232 1077 6328 1083
rect 6472 1077 6536 1083
rect 6013 1057 6200 1063
rect 6264 1057 6312 1063
rect 2093 1037 2584 1043
rect 2600 1037 2920 1043
rect 2936 1037 3000 1043
rect 3016 1037 3032 1043
rect 3176 1037 3208 1043
rect 3352 1037 3448 1043
rect 3576 1037 3608 1043
rect 3624 1037 4248 1043
rect 4264 1037 4680 1043
rect 4696 1037 4904 1043
rect 4936 1037 5800 1043
rect 5832 1037 5976 1043
rect 6392 1037 6456 1043
rect 1048 1017 1224 1023
rect 1256 1017 1320 1023
rect 1544 1017 1656 1023
rect 1704 1017 1768 1023
rect 216 997 296 1003
rect 312 997 568 1003
rect 600 997 632 1003
rect 648 997 1208 1003
rect 1288 997 1416 1003
rect 1432 997 1544 1003
rect 1576 997 1816 1003
rect 1976 1017 2120 1023
rect 2136 1017 2216 1023
rect 2328 1017 2408 1023
rect 2424 1017 2488 1023
rect 3128 1017 3272 1023
rect 2024 997 2168 1003
rect 2184 997 2808 1003
rect 2893 997 2936 1003
rect 216 977 392 983
rect 600 977 776 983
rect 792 977 1080 983
rect 1368 977 1400 983
rect 1560 977 2312 983
rect 2893 983 2899 997
rect 3016 997 3160 1003
rect 3352 997 3400 1003
rect 3752 997 3864 1003
rect 4312 1017 4328 1023
rect 4472 1017 4488 1023
rect 4632 1017 4792 1023
rect 5368 1017 5848 1023
rect 4168 997 4264 1003
rect 4280 997 4456 1003
rect 4552 997 4712 1003
rect 4776 997 4920 1003
rect 5352 997 5512 1003
rect 5992 1017 6056 1023
rect 6136 1017 6248 1023
rect 6264 1017 6424 1023
rect 6056 997 6136 1003
rect 6152 997 6264 1003
rect 6280 997 6520 1003
rect 2344 977 2899 983
rect 2909 977 3480 983
rect -51 957 8 963
rect 136 957 280 963
rect 808 957 968 963
rect 984 957 1096 963
rect 1112 957 1576 963
rect 1592 957 1960 963
rect 2040 957 2184 963
rect 2360 957 2408 963
rect 2440 957 2472 963
rect 2568 957 2680 963
rect 2909 963 2915 977
rect 3528 977 4120 983
rect 4136 977 5160 983
rect 5240 977 5320 983
rect 5336 977 5352 983
rect 5512 977 5528 983
rect 5560 977 5576 983
rect 6392 977 6408 983
rect 6424 977 6632 983
rect 2728 957 2915 963
rect 3192 957 3320 963
rect 3352 957 3400 963
rect 3736 957 4072 963
rect 4104 957 4264 963
rect 4328 957 4376 963
rect 4456 957 4520 963
rect 4616 957 4696 963
rect 5032 957 5064 963
rect 5320 957 5496 963
rect 5528 957 5576 963
rect 5960 957 6008 963
rect 6328 957 6376 963
rect 6392 957 6600 963
rect 317 948 323 952
rect 2925 948 2931 952
rect 88 937 312 943
rect 408 937 488 943
rect 648 937 808 943
rect 888 937 904 943
rect 984 937 1064 943
rect 1080 937 1112 943
rect 1448 937 1496 943
rect 1512 937 1640 943
rect 1656 937 1704 943
rect 1816 937 1880 943
rect 2120 937 2264 943
rect 2296 937 2872 943
rect 3064 937 3976 943
rect 4024 937 4104 943
rect 4248 937 4856 943
rect 4984 937 5032 943
rect 5181 943 5187 952
rect 5176 937 5187 943
rect 5229 937 5688 943
rect 381 928 387 932
rect 1373 928 1379 932
rect 2109 928 2115 932
rect 56 917 136 923
rect 200 917 216 923
rect 232 917 360 923
rect 520 917 600 923
rect 696 917 712 923
rect 728 917 888 923
rect 904 917 1080 923
rect 1448 917 1544 923
rect 1704 917 1736 923
rect 2168 917 2184 923
rect 2232 917 2760 923
rect 2888 917 3160 923
rect 3320 917 3336 923
rect 3624 917 3656 923
rect 3704 917 3816 923
rect 3944 917 4024 923
rect 4168 917 4248 923
rect 4344 917 4376 923
rect 4392 917 4920 923
rect 5229 923 5235 937
rect 5960 937 5976 943
rect 6344 937 6408 943
rect 6440 937 6472 943
rect 6536 937 6552 943
rect 6600 937 6680 943
rect 4936 917 5235 923
rect 5256 917 5368 923
rect 5384 917 5400 923
rect 5560 917 5624 923
rect 5704 917 5736 923
rect 5912 917 6104 923
rect 6152 917 6184 923
rect 6200 917 6232 923
rect 6312 917 6360 923
rect 6440 917 6515 923
rect 184 897 776 903
rect 792 897 1064 903
rect 1384 897 1848 903
rect 2104 897 2168 903
rect 2184 897 2200 903
rect 2392 897 2472 903
rect 2936 897 2968 903
rect 2984 897 3080 903
rect 3112 897 3368 903
rect 3416 897 3496 903
rect 3512 897 3576 903
rect 3608 897 3704 903
rect 3736 897 4216 903
rect 4232 897 4360 903
rect 4376 897 4408 903
rect 4424 897 4552 903
rect 4632 897 4760 903
rect 4888 897 4984 903
rect 5064 897 5128 903
rect 5144 897 5288 903
rect 5400 897 5432 903
rect 5640 897 5656 903
rect 5672 897 5720 903
rect 5864 897 5896 903
rect 6088 897 6408 903
rect 6424 897 6456 903
rect 6509 903 6515 917
rect 6536 917 6584 923
rect 6509 897 6520 903
rect 1085 888 1091 892
rect 136 877 232 883
rect 600 877 664 883
rect 680 877 920 883
rect 968 877 984 883
rect 1224 877 1608 883
rect 1640 877 1896 883
rect 1912 877 2216 883
rect 2360 877 2824 883
rect 3096 877 3224 883
rect 3656 877 3976 883
rect 3992 877 4136 883
rect 4152 877 4536 883
rect 4840 877 5112 883
rect 5128 877 5256 883
rect 5272 877 5624 883
rect 5864 877 6008 883
rect 6024 877 6200 883
rect 6216 877 6472 883
rect 6488 877 6536 883
rect 6792 877 6808 883
rect 760 857 968 863
rect 1128 857 1256 863
rect 1272 857 1400 863
rect 1464 857 1688 863
rect 1896 857 2360 863
rect 2504 857 2616 863
rect 2808 857 3160 863
rect 3176 857 3432 863
rect 3464 857 4232 863
rect 4312 857 4488 863
rect 4504 857 4995 863
rect 264 837 344 843
rect 360 837 440 843
rect 536 837 712 843
rect 1080 837 1272 843
rect 1592 837 2120 843
rect 2136 837 2200 843
rect 2376 837 2408 843
rect 2824 837 3224 843
rect 3240 837 3576 843
rect 4280 837 4424 843
rect 4440 837 4824 843
rect 4989 843 4995 857
rect 5336 857 5544 863
rect 5576 857 5752 863
rect 5768 857 6056 863
rect 6216 857 6328 863
rect 6344 857 6488 863
rect 6536 857 6552 863
rect 4989 837 5640 843
rect 6280 837 6552 843
rect 6568 837 6600 843
rect 6616 837 6632 843
rect 936 817 984 823
rect 1000 817 1336 823
rect 1416 817 1448 823
rect 1560 817 1608 823
rect 1704 817 1800 823
rect 2200 817 2520 823
rect 1144 797 1304 803
rect 1320 797 1384 803
rect 1400 797 2328 803
rect 2728 797 2760 803
rect 3000 817 4472 823
rect 3032 797 3384 803
rect 3576 797 3720 803
rect 3736 797 4184 803
rect 4280 797 4552 803
rect 4568 797 4600 803
rect 4696 797 4776 803
rect 5208 817 5256 823
rect 5272 817 5688 823
rect 5928 817 6264 823
rect 5016 797 5464 803
rect 5480 797 6136 803
rect 280 777 392 783
rect 1032 777 1192 783
rect 1208 777 1288 783
rect 2024 777 2312 783
rect 2840 777 3352 783
rect 3368 777 3832 783
rect 4152 777 4264 783
rect 4456 777 5000 783
rect 5304 777 5912 783
rect 6120 777 6312 783
rect 1032 757 1208 763
rect 1624 757 1928 763
rect 1944 757 2232 763
rect 2552 757 2984 763
rect 3080 757 3144 763
rect 3208 757 3432 763
rect 3816 757 4584 763
rect 4600 757 5336 763
rect 5416 757 5528 763
rect 5640 757 5816 763
rect 5832 757 6168 763
rect 456 737 520 743
rect 584 737 664 743
rect 808 737 968 743
rect 1096 737 1256 743
rect 1352 737 1384 743
rect 1736 737 1768 743
rect 1800 737 1848 743
rect 1864 737 2024 743
rect 2232 737 2312 743
rect 2536 737 2744 743
rect 2760 737 3064 743
rect 3112 737 3128 743
rect 3160 737 3192 743
rect 3752 737 3768 743
rect 4072 737 4104 743
rect 4136 737 4360 743
rect 4381 737 4504 743
rect -51 717 8 723
rect 120 717 152 723
rect 184 717 312 723
rect 392 717 776 723
rect 952 717 984 723
rect 1016 717 1112 723
rect 1208 717 2104 723
rect 2376 717 2584 723
rect 2728 717 2936 723
rect 3096 717 3176 723
rect 3224 717 3240 723
rect 3304 717 3320 723
rect 3336 717 3528 723
rect 3560 717 3896 723
rect 4024 717 4168 723
rect 4232 717 4280 723
rect 4381 723 4387 737
rect 4536 737 4568 743
rect 4728 737 4808 743
rect 4824 737 5064 743
rect 5288 737 5304 743
rect 5592 737 5752 743
rect 6056 737 6296 743
rect 6456 737 6504 743
rect 5533 728 5539 732
rect 4312 717 4387 723
rect 4408 717 4419 723
rect 4552 717 4632 723
rect 4680 717 4776 723
rect 4904 717 4920 723
rect 5048 717 5080 723
rect 5128 717 5144 723
rect 5261 717 5416 723
rect 2221 708 2227 712
rect 152 697 168 703
rect 216 697 264 703
rect 376 697 440 703
rect 488 697 584 703
rect 888 697 1080 703
rect 1176 697 1208 703
rect 1368 697 1480 703
rect 1496 697 1512 703
rect 1544 697 2008 703
rect 2104 697 2136 703
rect 2264 697 2280 703
rect 2312 697 2376 703
rect 2392 697 2424 703
rect 2637 703 2643 712
rect 5261 708 5267 717
rect 5624 717 5688 723
rect 5704 717 5784 723
rect 5805 717 6136 723
rect 2472 697 2888 703
rect 2952 697 2968 703
rect 3048 697 3272 703
rect 3432 697 3624 703
rect 3640 697 3672 703
rect 3800 697 4179 703
rect 685 688 691 692
rect 3693 688 3699 692
rect 3757 688 3763 692
rect 4173 688 4179 697
rect 4264 697 4344 703
rect 4392 697 4424 703
rect 4504 697 4760 703
rect 4776 697 5224 703
rect 5805 703 5811 717
rect 6424 717 6568 723
rect 6664 717 6696 723
rect 5752 697 5811 703
rect 6040 697 6120 703
rect 6136 697 6376 703
rect 200 677 488 683
rect 856 677 1064 683
rect 1192 677 1320 683
rect 1400 677 1496 683
rect 1512 677 1672 683
rect 1688 677 1752 683
rect 1768 677 1816 683
rect 2040 677 2152 683
rect 2328 677 2408 683
rect 2440 677 2616 683
rect 2632 677 2904 683
rect 2920 677 3160 683
rect 3544 677 3672 683
rect 3768 677 3864 683
rect 3896 677 4088 683
rect 4120 677 4136 683
rect 4184 677 4200 683
rect 4344 677 4408 683
rect 4472 677 4520 683
rect 4600 677 4664 683
rect 4696 677 5208 683
rect 5240 677 5336 683
rect 5352 677 5496 683
rect 5512 677 5640 683
rect 5656 677 5896 683
rect 6200 677 6248 683
rect 6312 677 6392 683
rect 6632 677 6664 683
rect 6712 677 6792 683
rect 573 668 579 672
rect 40 657 104 663
rect 472 657 552 663
rect 1048 657 1736 663
rect 1752 657 2088 663
rect 2264 657 2328 663
rect 2696 657 3128 663
rect 3176 657 3512 663
rect 3624 657 3880 663
rect 3912 657 4072 663
rect 4168 657 4312 663
rect 4408 657 4536 663
rect 4664 657 4680 663
rect 4760 657 4840 663
rect 4856 657 4888 663
rect 4904 657 5016 663
rect 5256 657 5400 663
rect 5528 657 5576 663
rect 5688 657 5768 663
rect 5912 657 6328 663
rect 696 637 1032 643
rect 1736 637 1944 643
rect 2152 637 2168 643
rect 2200 637 2392 643
rect 2648 637 2771 643
rect 760 617 1112 623
rect 1144 617 1560 623
rect 1576 617 1800 623
rect 344 597 600 603
rect 984 597 1080 603
rect 1128 597 1240 603
rect 1256 597 1304 603
rect 2712 617 2744 623
rect 2765 623 2771 637
rect 2792 637 2904 643
rect 2920 637 3000 643
rect 3112 637 3192 643
rect 3224 637 3400 643
rect 3432 637 3528 643
rect 3560 637 4248 643
rect 4296 637 4344 643
rect 4456 637 4504 643
rect 4520 637 4984 643
rect 5000 637 5224 643
rect 5288 637 5352 643
rect 5480 637 5592 643
rect 5704 637 5768 643
rect 5832 637 5880 643
rect 6440 637 6504 643
rect 6584 637 6616 643
rect 2765 617 2792 623
rect 3016 617 3032 623
rect 3480 617 3848 623
rect 2008 597 2216 603
rect 2360 597 2424 603
rect 2440 597 2472 603
rect 2520 597 3544 603
rect 3672 597 3864 603
rect 4264 617 4536 623
rect 4680 617 4840 623
rect 5000 617 5144 623
rect 5160 617 5256 623
rect 5400 617 5608 623
rect 4104 597 4408 603
rect 4504 597 4568 603
rect 4600 597 4808 603
rect 4856 597 5144 603
rect 5672 597 5912 603
rect 104 577 280 583
rect 424 577 840 583
rect 936 577 984 583
rect 1064 577 1096 583
rect 1128 577 1224 583
rect 1240 577 1400 583
rect 1432 577 1608 583
rect 1928 577 2136 583
rect 2152 577 2280 583
rect 2344 577 2472 583
rect 2584 577 2616 583
rect 2744 577 3032 583
rect 3048 577 3064 583
rect 3128 577 3144 583
rect 3208 577 3448 583
rect 3640 577 3672 583
rect 3736 577 3827 583
rect -51 557 56 563
rect 88 557 136 563
rect 200 557 488 563
rect 872 557 1128 563
rect 1160 557 1208 563
rect 1224 557 1384 563
rect 1400 557 1432 563
rect 1480 557 1496 563
rect 1944 557 2104 563
rect 2120 557 2248 563
rect 2312 557 2424 563
rect 2520 557 2920 563
rect 3112 557 3176 563
rect 3192 557 3336 563
rect 3496 557 3688 563
rect 3704 557 3800 563
rect 3821 563 3827 577
rect 3880 577 4248 583
rect 4264 577 4296 583
rect 4312 577 4392 583
rect 4440 577 4456 583
rect 4488 577 5384 583
rect 5640 577 5768 583
rect 5784 577 5992 583
rect 6312 577 6632 583
rect 6648 577 6728 583
rect 3821 557 3928 563
rect 3976 557 4104 563
rect 4120 557 4147 563
rect 56 537 88 543
rect 328 537 392 543
rect 488 537 1192 543
rect 1288 537 1512 543
rect 1704 537 1896 543
rect 1976 537 2008 543
rect 2072 537 2264 543
rect 2424 537 2488 543
rect 2504 537 3192 543
rect 3288 537 3304 543
rect 3432 537 3560 543
rect 3592 537 3736 543
rect 1197 528 1203 532
rect 1261 528 1267 532
rect 2349 528 2355 532
rect 3757 528 3763 543
rect 3800 537 3864 543
rect 4072 537 4120 543
rect 4141 543 4147 557
rect 4296 557 4472 563
rect 4600 557 5000 563
rect 5016 557 5160 563
rect 5208 557 5240 563
rect 5272 557 5528 563
rect 5544 557 5640 563
rect 5656 557 6120 563
rect 6248 557 6312 563
rect 6488 557 6568 563
rect 6824 557 6867 563
rect 4141 537 4264 543
rect 4344 537 4616 543
rect 4728 537 4744 543
rect 4920 537 5048 543
rect 5080 537 5096 543
rect 5128 537 5208 543
rect 5224 537 5368 543
rect 5384 537 5656 543
rect 5672 537 5960 543
rect 5976 537 6008 543
rect 6184 537 6216 543
rect 6264 537 6280 543
rect 6376 537 6504 543
rect 3773 528 3779 532
rect -51 517 8 523
rect 72 517 200 523
rect 216 517 1128 523
rect 1352 517 1496 523
rect 1832 517 1944 523
rect 1992 517 2184 523
rect 2408 517 2456 523
rect 2664 517 2760 523
rect 3144 517 3640 523
rect 3688 517 3704 523
rect 3848 517 3976 523
rect 4040 517 4088 523
rect 4264 517 4312 523
rect 4328 517 4520 523
rect 4536 517 5000 523
rect 5048 517 5080 523
rect 5208 517 5432 523
rect 5448 517 5624 523
rect 5656 517 5688 523
rect 6008 517 6376 523
rect 2605 508 2611 512
rect 248 497 440 503
rect 456 497 488 503
rect 504 497 632 503
rect 824 497 904 503
rect 952 497 1448 503
rect 1464 497 1880 503
rect 1896 497 2008 503
rect 2152 497 2248 503
rect 2632 497 2664 503
rect 3064 497 3144 503
rect 3176 497 3288 503
rect 3512 497 3560 503
rect 3576 497 3944 503
rect 3960 497 4232 503
rect 4664 497 4808 503
rect 4968 497 5256 503
rect 5544 497 5576 503
rect 5592 497 5656 503
rect 5672 497 5688 503
rect 5768 497 5800 503
rect 5821 497 6008 503
rect 104 477 360 483
rect 376 477 504 483
rect 520 477 552 483
rect 584 477 1384 483
rect 2184 477 2584 483
rect 2632 477 2904 483
rect 3560 477 3752 483
rect 3768 477 3896 483
rect 3912 477 4040 483
rect 4216 477 4616 483
rect 4664 477 4680 483
rect 4920 477 5000 483
rect 5016 477 5304 483
rect 5320 477 5416 483
rect 5432 477 5480 483
rect 5496 477 5704 483
rect 5821 483 5827 497
rect 6296 497 6360 503
rect 6488 497 6648 503
rect 5752 477 5827 483
rect 5896 477 6248 483
rect 680 457 872 463
rect 1000 457 1080 463
rect 1112 457 1160 463
rect 1176 457 1256 463
rect 1277 457 1912 463
rect 216 437 312 443
rect 1277 443 1283 457
rect 2168 457 2248 463
rect 2349 457 2360 463
rect 2488 457 2904 463
rect 3080 457 3144 463
rect 3304 457 3768 463
rect 3944 457 4184 463
rect 4376 457 4552 463
rect 4744 457 5144 463
rect 5160 457 5528 463
rect 5560 457 5592 463
rect 664 437 1283 443
rect 1336 437 1400 443
rect 1416 437 1480 443
rect 1496 437 1528 443
rect 1832 437 2488 443
rect 2568 437 2920 443
rect 2936 437 3384 443
rect 3400 437 3512 443
rect 3544 437 3992 443
rect 4024 437 4072 443
rect 4296 437 4456 443
rect 4536 437 4728 443
rect 4856 437 5576 443
rect 5661 437 5864 443
rect 552 417 632 423
rect 648 417 760 423
rect 856 417 2184 423
rect 2264 417 2504 423
rect 2680 417 2808 423
rect 1064 397 1304 403
rect 2248 397 2392 403
rect 2520 397 2552 403
rect 2920 417 3080 423
rect 3096 417 4472 423
rect 4664 417 4776 423
rect 4792 417 4840 423
rect 3672 397 3800 403
rect 3816 397 4008 403
rect 4568 397 4680 403
rect 4696 397 4760 403
rect 4792 397 4888 403
rect 5224 417 5480 423
rect 5661 423 5667 437
rect 5880 437 6232 443
rect 5496 417 5667 423
rect 5688 417 5816 423
rect 6344 417 6712 423
rect 4989 397 5128 403
rect 536 377 664 383
rect 1080 377 1256 383
rect 1512 377 1608 383
rect 2248 377 2536 383
rect 2600 377 2728 383
rect 2968 377 3096 383
rect 3112 377 3304 383
rect 3544 377 3592 383
rect 3752 377 4024 383
rect 4040 377 4232 383
rect 4989 383 4995 397
rect 5208 397 5224 403
rect 5320 397 5528 403
rect 5560 397 6136 403
rect 6765 388 6771 392
rect 4248 377 4995 383
rect 5016 377 5448 383
rect 5464 377 5848 383
rect 5864 377 6088 383
rect 376 357 408 363
rect 440 357 536 363
rect 552 357 584 363
rect 680 357 936 363
rect 1256 357 1384 363
rect 1992 357 2072 363
rect 2088 357 2344 363
rect 2472 357 3112 363
rect 3128 357 3928 363
rect 4248 357 4259 363
rect 4456 357 4872 363
rect 4920 357 4952 363
rect 5048 357 5128 363
rect 5256 357 5384 363
rect 5416 357 5768 363
rect 5880 357 6024 363
rect 6600 357 6744 363
rect 285 348 291 352
rect 312 337 344 343
rect 424 337 600 343
rect 616 337 728 343
rect 744 337 1144 343
rect 1192 337 1288 343
rect 2120 337 2408 343
rect 2472 337 2488 343
rect 2520 337 2744 343
rect 2808 337 2968 343
rect 3000 337 3032 343
rect 3272 337 3368 343
rect 3672 337 4168 343
rect 4248 337 4280 343
rect 4344 337 4408 343
rect 4424 337 4872 343
rect 4888 337 5736 343
rect 6040 337 6168 343
rect 6696 337 6867 343
rect -51 317 8 323
rect 344 317 472 323
rect 488 317 568 323
rect 696 317 707 323
rect 824 317 840 323
rect 952 317 968 323
rect 1064 317 1096 323
rect 1208 317 1336 323
rect 1400 317 1464 323
rect 1592 317 1704 323
rect 2232 317 2248 323
rect 2296 317 2344 323
rect 2365 317 2376 323
rect 2456 317 2568 323
rect 2712 317 2856 323
rect 2872 317 2952 323
rect 3032 317 3480 323
rect 3512 317 3640 323
rect 3656 317 4152 323
rect 4168 317 4632 323
rect 4648 317 5288 323
rect 5528 317 5544 323
rect 5592 317 5624 323
rect 5640 317 5688 323
rect 5704 317 6312 323
rect 6632 317 6744 323
rect 6861 317 6867 337
rect 328 297 376 303
rect 392 297 1000 303
rect 1016 297 1144 303
rect 1160 297 1208 303
rect 1304 297 1464 303
rect 1640 297 1800 303
rect 2040 297 2120 303
rect 2200 297 2264 303
rect 2328 297 2392 303
rect 2440 297 3288 303
rect 3400 297 3416 303
rect 3437 297 3448 303
rect 3608 297 3656 303
rect 3752 297 3800 303
rect 3880 297 3976 303
rect 3992 297 4824 303
rect 5096 297 5640 303
rect 5656 297 5896 303
rect 6120 297 6152 303
rect 6200 297 6440 303
rect 6456 297 6552 303
rect 3693 288 3699 292
rect 4957 288 4963 292
rect 376 277 408 283
rect 424 277 584 283
rect 600 277 1272 283
rect 1608 277 1672 283
rect 1688 277 2088 283
rect 2104 277 2488 283
rect 2504 277 2696 283
rect 2728 277 2808 283
rect 2856 277 2952 283
rect 2968 277 3096 283
rect 3208 277 3240 283
rect 3453 277 3544 283
rect 488 257 568 263
rect 584 257 712 263
rect 728 257 872 263
rect 888 257 1320 263
rect 1944 257 2024 263
rect 2168 257 2216 263
rect 2333 257 2344 263
rect 2376 257 2424 263
rect 2632 257 2824 263
rect 2840 257 3016 263
rect 3064 257 3336 263
rect 3453 263 3459 277
rect 3720 277 3752 283
rect 3848 277 3864 283
rect 3992 277 4120 283
rect 4216 277 4392 283
rect 4440 277 4536 283
rect 4552 277 4584 283
rect 4632 277 4888 283
rect 4984 277 5576 283
rect 5640 277 5704 283
rect 5720 277 5816 283
rect 5832 277 5992 283
rect 6152 277 6264 283
rect 6712 277 6776 283
rect 6792 277 6867 283
rect 3352 257 3459 263
rect 3480 257 4040 263
rect 4280 257 4312 263
rect 4392 257 4520 263
rect 4760 257 4920 263
rect 4936 257 5128 263
rect 5144 257 5320 263
rect 5624 257 5688 263
rect 5704 257 5832 263
rect 264 237 616 243
rect 936 237 1032 243
rect 1048 237 1128 243
rect 1144 237 1288 243
rect 1368 237 1816 243
rect 2008 237 2280 243
rect 2536 237 2632 243
rect 2728 237 2776 243
rect 2872 237 3000 243
rect 3016 237 3224 243
rect 3240 237 3432 243
rect 3448 237 3672 243
rect 3688 237 3864 243
rect 3880 237 4136 243
rect 4152 237 4360 243
rect 4968 237 5096 243
rect 5176 237 5368 243
rect 5928 237 5944 243
rect 5976 237 6024 243
rect 6040 237 6424 243
rect 904 217 984 223
rect 1048 217 1656 223
rect 1704 217 1784 223
rect 1080 197 1096 203
rect 1128 197 1640 203
rect 1656 197 1704 203
rect 2312 217 2712 223
rect 2840 217 2984 223
rect 3304 217 3480 223
rect 3496 217 3768 223
rect 1960 197 2184 203
rect 2280 197 2424 203
rect 2792 197 3048 203
rect 3320 197 3848 203
rect 4056 217 4728 223
rect 4760 217 4808 223
rect 4824 217 5160 223
rect 5181 217 5192 223
rect 4024 197 4360 203
rect 4680 197 4760 203
rect 5181 203 5187 217
rect 5272 217 5336 223
rect 5400 217 5464 223
rect 4776 197 5187 203
rect 5208 197 5240 203
rect 5368 197 5384 203
rect 5448 197 5512 203
rect 1000 177 1016 183
rect 1032 177 1336 183
rect 1352 177 1752 183
rect 1768 177 2408 183
rect 2424 177 3128 183
rect 3432 177 3656 183
rect 3864 177 4280 183
rect 4381 183 4387 192
rect 4376 177 4387 183
rect 4872 177 5000 183
rect 5304 177 5944 183
rect 5960 177 6008 183
rect 6456 177 6584 183
rect 6616 177 6632 183
rect 120 157 136 163
rect 909 163 915 172
rect 3181 168 3187 172
rect 680 157 920 163
rect 1016 157 1064 163
rect 1096 157 1160 163
rect 1192 157 1384 163
rect 1416 157 1528 163
rect 1736 157 1800 163
rect 1816 157 1944 163
rect 2136 157 2152 163
rect 2568 157 2888 163
rect 3192 157 3496 163
rect 3512 157 3688 163
rect 3944 157 3992 163
rect 4088 157 4120 163
rect 4600 157 4632 163
rect 4648 157 4968 163
rect 5128 157 5320 163
rect 5352 157 5768 163
rect 5848 157 5928 163
rect 2397 148 2403 152
rect 2461 148 2467 152
rect 6509 148 6515 152
rect 520 137 584 143
rect 792 137 1032 143
rect 1288 137 1320 143
rect 1400 137 1416 143
rect 1704 137 1992 143
rect 2184 137 2312 143
rect 2344 137 2376 143
rect 2429 137 2440 143
rect 2504 137 2520 143
rect 2760 137 2824 143
rect 2984 137 3288 143
rect 3416 137 3976 143
rect 3992 137 4104 143
rect 4184 137 4248 143
rect 4408 137 4696 143
rect 4840 137 5560 143
rect 5640 137 5731 143
rect -51 117 8 123
rect 152 117 184 123
rect 216 117 248 123
rect 392 117 472 123
rect 920 117 968 123
rect 1176 117 1256 123
rect 1272 117 1320 123
rect 1352 117 1416 123
rect 1464 117 1512 123
rect 1864 117 2259 123
rect 808 97 1112 103
rect 1128 97 1224 103
rect 1320 97 1352 103
rect 2253 103 2259 117
rect 2424 117 2440 123
rect 2504 117 2536 123
rect 2568 117 2648 123
rect 2664 117 2968 123
rect 3048 117 3128 123
rect 3272 117 3528 123
rect 3549 117 3720 123
rect 2253 97 2552 103
rect 2616 97 2824 103
rect 3277 97 3288 103
rect 3400 97 3416 103
rect 3549 103 3555 117
rect 3784 117 4088 123
rect 4104 117 4472 123
rect 4840 117 4952 123
rect 4989 117 5000 123
rect 4989 108 4995 117
rect 5112 117 5304 123
rect 5336 117 5624 123
rect 5656 117 5704 123
rect 5725 123 5731 137
rect 6072 137 6184 143
rect 5725 117 5800 123
rect 6184 117 6200 123
rect 6696 117 6867 123
rect 3464 97 3555 103
rect 3608 97 4168 103
rect 4200 97 4472 103
rect 4488 97 4568 103
rect 4584 97 4696 103
rect 4776 97 4840 103
rect 5336 97 5400 103
rect 5432 97 5592 103
rect 5640 97 5672 103
rect 5928 97 5960 103
rect 5976 97 6072 103
rect 712 77 984 83
rect 2776 77 3032 83
rect 3080 77 3464 83
rect 488 57 600 63
rect 952 57 1432 63
rect 2120 57 2264 63
rect 3144 57 3400 63
rect 4312 37 4456 43
rect 4472 37 4824 43
rect 4840 37 5624 43
rect 3960 17 3976 23
rect 5928 17 5944 23
rect 6040 17 6056 23
<< m4contact >>
rect 798 4802 826 4818
rect 2862 4802 2890 4818
rect 3496 4812 3512 4828
rect 4910 4802 4938 4818
rect 3736 4772 3752 4788
rect 168 4692 184 4708
rect 936 4692 952 4708
rect 2216 4692 2232 4708
rect 2568 4692 2584 4708
rect 3064 4692 3080 4708
rect 3736 4692 3752 4708
rect 4712 4692 4728 4708
rect 5128 4692 5144 4708
rect 6568 4692 6584 4708
rect 1656 4672 1672 4688
rect 2472 4672 2488 4688
rect 3480 4672 3496 4688
rect 5512 4672 5528 4688
rect 1304 4652 1320 4668
rect 1496 4652 1512 4668
rect 4664 4652 4680 4668
rect 3720 4632 3736 4648
rect 1064 4612 1080 4628
rect 1752 4612 1768 4628
rect 1838 4602 1866 4618
rect 2680 4612 2696 4628
rect 3886 4602 3914 4618
rect 5336 4632 5352 4648
rect 4424 4592 4440 4608
rect 5934 4602 5962 4618
rect 1704 4572 1720 4588
rect 1272 4552 1288 4568
rect 2584 4552 2600 4568
rect 2984 4552 3000 4568
rect 3432 4552 3448 4568
rect 3704 4552 3720 4568
rect 5640 4552 5656 4568
rect 1096 4532 1112 4548
rect 1672 4532 1688 4548
rect 1832 4532 1848 4548
rect 1944 4532 1960 4548
rect 2280 4532 2296 4548
rect 2552 4532 2568 4548
rect 2776 4532 2808 4548
rect 2824 4532 2840 4548
rect 2984 4532 3000 4548
rect 3560 4532 3576 4548
rect 4248 4532 4264 4548
rect 4504 4532 4536 4548
rect 1048 4512 1080 4528
rect 1128 4512 1144 4528
rect 2536 4512 2552 4528
rect 2584 4512 2600 4528
rect 2616 4512 2632 4528
rect 2744 4512 2760 4528
rect 3560 4512 3576 4528
rect 3864 4512 3880 4528
rect 3992 4512 4008 4528
rect 4696 4512 4712 4528
rect 4888 4512 4904 4528
rect 1112 4492 1128 4508
rect 1544 4492 1560 4508
rect 1560 4492 1576 4508
rect 1576 4492 1592 4508
rect 2776 4492 2792 4508
rect 3192 4492 3208 4508
rect 4840 4492 4856 4508
rect 5192 4492 5208 4508
rect 5448 4492 5464 4508
rect 3320 4472 3336 4488
rect 456 4452 472 4468
rect 4712 4452 4728 4468
rect 6168 4452 6184 4468
rect 3160 4432 3176 4448
rect 4120 4432 4136 4448
rect 4696 4432 4712 4448
rect 5096 4432 5112 4448
rect 798 4402 826 4418
rect 1224 4412 1240 4428
rect 1256 4412 1272 4428
rect 2632 4412 2648 4428
rect 2824 4412 2840 4428
rect 1560 4392 1576 4408
rect 2862 4402 2890 4418
rect 3336 4412 3352 4428
rect 4376 4412 4392 4428
rect 4808 4412 4824 4428
rect 4910 4402 4938 4418
rect 6168 4412 6184 4428
rect 1032 4372 1048 4388
rect 1480 4372 1496 4388
rect 2248 4372 2264 4388
rect 2568 4372 2584 4388
rect 5528 4372 5544 4388
rect 856 4352 872 4368
rect 888 4352 920 4368
rect 1672 4352 1688 4368
rect 2872 4352 2888 4368
rect 3048 4352 3064 4368
rect 4632 4352 4648 4368
rect 4664 4352 4680 4368
rect 4792 4352 4808 4368
rect 5528 4352 5544 4368
rect 664 4332 680 4348
rect 1000 4332 1016 4348
rect 1192 4332 1224 4348
rect 2232 4332 2248 4348
rect 2680 4332 2696 4348
rect 2728 4332 2744 4348
rect 168 4292 184 4308
rect 664 4292 680 4308
rect 952 4292 968 4308
rect 1240 4312 1256 4328
rect 1272 4312 1288 4328
rect 1496 4312 1512 4328
rect 1720 4312 1736 4328
rect 1992 4312 2008 4328
rect 2744 4312 2760 4328
rect 3720 4312 3736 4328
rect 4424 4312 4440 4328
rect 5080 4312 5096 4328
rect 5720 4312 5736 4328
rect 5784 4312 5800 4328
rect 5864 4312 5880 4328
rect 1960 4292 1976 4308
rect 3480 4292 3496 4308
rect 920 4272 936 4288
rect 1176 4272 1192 4288
rect 1272 4272 1288 4288
rect 2824 4272 2840 4288
rect 3288 4272 3304 4288
rect 3816 4272 3832 4288
rect 4520 4272 4552 4288
rect 4824 4272 4840 4288
rect 4968 4272 4984 4288
rect 5416 4272 5432 4288
rect 5720 4272 5736 4288
rect 184 4252 200 4268
rect 1112 4252 1128 4268
rect 1192 4252 1208 4268
rect 1240 4252 1256 4268
rect 1064 4232 1080 4248
rect 1656 4252 1672 4268
rect 2328 4252 2344 4268
rect 2376 4252 2392 4268
rect 3080 4252 3096 4268
rect 4952 4252 4968 4268
rect 5288 4252 5304 4268
rect 856 4212 872 4228
rect 1000 4212 1016 4228
rect 1448 4212 1464 4228
rect 1592 4192 1608 4208
rect 1838 4202 1866 4218
rect 2920 4232 2936 4248
rect 3928 4232 3944 4248
rect 4872 4232 4888 4248
rect 5016 4232 5032 4248
rect 6152 4232 6168 4248
rect 3192 4212 3208 4228
rect 2776 4192 2792 4208
rect 3368 4192 3384 4208
rect 3768 4192 3784 4208
rect 3886 4202 3914 4218
rect 4328 4212 4344 4228
rect 4808 4212 4824 4228
rect 4280 4192 4296 4208
rect 4504 4192 4520 4208
rect 4888 4192 4904 4208
rect 5064 4192 5080 4208
rect 5512 4192 5528 4208
rect 5934 4202 5962 4218
rect 1736 4172 1752 4188
rect 3320 4172 3336 4188
rect 3464 4172 3480 4188
rect 5528 4172 5544 4188
rect 5816 4172 5832 4188
rect 1080 4152 1096 4168
rect 456 4132 472 4148
rect 1224 4152 1240 4168
rect 1800 4152 1816 4168
rect 2280 4152 2296 4168
rect 3336 4152 3352 4168
rect 3864 4152 3880 4168
rect 1144 4132 1160 4148
rect 1208 4132 1224 4148
rect 1320 4132 1336 4148
rect 1352 4132 1368 4148
rect 1400 4132 1416 4148
rect 1688 4132 1704 4148
rect 2760 4132 2776 4148
rect 3080 4132 3096 4148
rect 4472 4152 4488 4168
rect 5192 4152 5208 4168
rect 6392 4152 6408 4168
rect 4360 4132 4376 4148
rect 4536 4132 4552 4148
rect 5016 4132 5032 4148
rect 5048 4132 5064 4148
rect 5256 4132 5272 4148
rect 5416 4132 5432 4148
rect 6280 4132 6296 4148
rect 6424 4132 6440 4148
rect 584 4112 600 4128
rect 1608 4112 1624 4128
rect 2392 4112 2408 4128
rect 2440 4112 2456 4128
rect 2840 4112 2856 4128
rect 2888 4112 2920 4128
rect 3176 4112 3192 4128
rect 4712 4112 4728 4128
rect 5016 4112 5032 4128
rect 904 4092 920 4108
rect 1192 4092 1208 4108
rect 1320 4092 1336 4108
rect 1496 4092 1512 4108
rect 2424 4092 2440 4108
rect 3176 4092 3192 4108
rect 4152 4092 4168 4108
rect 4408 4092 4424 4108
rect 4792 4092 4808 4108
rect 4968 4092 4984 4108
rect 5176 4112 5192 4128
rect 5400 4112 5416 4128
rect 5880 4112 5896 4128
rect 5960 4112 5976 4128
rect 6056 4112 6088 4128
rect 6104 4112 6120 4128
rect 6024 4092 6040 4108
rect 1320 4072 1336 4088
rect 2264 4072 2280 4088
rect 2584 4072 2600 4088
rect 2904 4072 2920 4088
rect 3224 4072 3240 4088
rect 4984 4072 5000 4088
rect 5080 4072 5096 4088
rect 5688 4072 5704 4088
rect 6040 4072 6056 4088
rect 936 4052 952 4068
rect 4088 4052 4104 4068
rect 4344 4052 4360 4068
rect 4408 4052 4424 4068
rect 4616 4052 4632 4068
rect 5848 4052 5864 4068
rect 952 4032 968 4048
rect 1256 4032 1272 4048
rect 1560 4032 1576 4048
rect 1672 4032 1688 4048
rect 1832 4032 1848 4048
rect 1928 4032 1944 4048
rect 3496 4032 3512 4048
rect 4456 4032 4472 4048
rect 5896 4032 5912 4048
rect 216 4012 232 4028
rect 798 4002 826 4018
rect 920 4012 936 4028
rect 904 3992 920 4008
rect 1544 3992 1560 4008
rect 2862 4002 2890 4018
rect 3784 4012 3800 4028
rect 3816 4012 3832 4028
rect 2920 3992 2936 4008
rect 4456 3992 4472 4008
rect 4910 4002 4938 4018
rect 4968 4012 4984 4028
rect 5960 4012 5976 4028
rect 5176 3992 5192 4008
rect 520 3972 536 3988
rect 680 3972 696 3988
rect 968 3972 984 3988
rect 1080 3972 1096 3988
rect 3928 3952 3944 3968
rect 1304 3932 1320 3948
rect 1688 3932 1704 3948
rect 2808 3932 2824 3948
rect 4056 3932 4072 3948
rect 5320 3952 5336 3968
rect 5032 3932 5048 3948
rect 5688 3932 5704 3948
rect 1560 3912 1576 3928
rect 1704 3912 1720 3928
rect 1768 3912 1784 3928
rect 2472 3912 2488 3928
rect 2744 3912 2760 3928
rect 3784 3912 3800 3928
rect 4024 3912 4040 3928
rect 4312 3912 4328 3928
rect 4872 3912 4888 3928
rect 5000 3912 5016 3928
rect 6264 3912 6280 3928
rect 1000 3892 1016 3908
rect 1160 3892 1176 3908
rect 2712 3892 2728 3908
rect 2920 3892 2936 3908
rect 2952 3892 2968 3908
rect 3048 3892 3064 3908
rect 3176 3892 3192 3908
rect 3848 3892 3864 3908
rect 3864 3892 3880 3908
rect 4040 3892 4072 3908
rect 4376 3892 4392 3908
rect 4472 3892 4488 3908
rect 5880 3892 5896 3908
rect 712 3872 728 3888
rect 872 3872 888 3888
rect 1560 3872 1576 3888
rect 1816 3872 1832 3888
rect 2120 3872 2136 3888
rect 2184 3872 2200 3888
rect 2248 3872 2264 3888
rect 2840 3872 2856 3888
rect 3480 3872 3496 3888
rect 4376 3872 4392 3888
rect 5272 3872 5288 3888
rect 5976 3872 5992 3888
rect 840 3852 856 3868
rect 1000 3852 1016 3868
rect 1400 3852 1416 3868
rect 1480 3852 1496 3868
rect 1592 3852 1608 3868
rect 2776 3852 2792 3868
rect 3512 3852 3528 3868
rect 4072 3852 4088 3868
rect 4440 3852 4472 3868
rect 4552 3852 4568 3868
rect 4888 3852 4904 3868
rect 4984 3852 5000 3868
rect 984 3832 1000 3848
rect 1688 3832 1704 3848
rect 2984 3832 3000 3848
rect 360 3812 376 3828
rect 936 3812 952 3828
rect 1112 3812 1128 3828
rect 1768 3792 1784 3808
rect 1838 3802 1866 3818
rect 3224 3812 3240 3828
rect 3464 3792 3480 3808
rect 3886 3802 3914 3818
rect 4632 3832 4648 3848
rect 4664 3832 4680 3848
rect 4696 3832 4712 3848
rect 5160 3832 5176 3848
rect 5432 3832 5448 3848
rect 4344 3812 4360 3828
rect 3928 3792 3944 3808
rect 4232 3792 4248 3808
rect 5934 3802 5962 3818
rect 1944 3772 1960 3788
rect 3864 3772 3880 3788
rect 1784 3752 1800 3768
rect 2472 3752 2488 3768
rect 2648 3752 2664 3768
rect 3224 3752 3240 3768
rect 3448 3752 3464 3768
rect 3928 3752 3944 3768
rect 4888 3772 4904 3788
rect 4824 3752 4840 3768
rect 5656 3752 5672 3768
rect 6792 3752 6808 3768
rect 232 3732 248 3748
rect 408 3732 424 3748
rect 888 3732 904 3748
rect 1656 3732 1672 3748
rect 1736 3732 1752 3748
rect 1800 3732 1816 3748
rect 1992 3732 2024 3748
rect 72 3712 88 3728
rect 984 3712 1000 3728
rect 1992 3712 2008 3728
rect 2232 3732 2248 3748
rect 2360 3732 2376 3748
rect 2600 3732 2616 3748
rect 2824 3732 2840 3748
rect 5448 3732 5464 3748
rect 6664 3732 6680 3748
rect 2792 3712 2808 3728
rect 2168 3692 2184 3708
rect 4072 3712 4088 3728
rect 4632 3712 4648 3728
rect 4648 3712 4664 3728
rect 4744 3712 4760 3728
rect 6568 3712 6584 3728
rect 3080 3692 3096 3708
rect 4136 3692 4152 3708
rect 5288 3692 5304 3708
rect 3640 3672 3656 3688
rect 3704 3672 3736 3688
rect 3800 3672 3816 3688
rect 4072 3672 4088 3688
rect 4104 3672 4120 3688
rect 4552 3672 4568 3688
rect 5016 3672 5032 3688
rect 5800 3672 5816 3688
rect 6280 3672 6296 3688
rect 424 3652 440 3668
rect 1016 3652 1032 3668
rect 1768 3652 1784 3668
rect 4968 3652 4984 3668
rect 5976 3652 5992 3668
rect 200 3632 216 3648
rect 616 3632 632 3648
rect 968 3632 984 3648
rect 1512 3632 1528 3648
rect 568 3612 584 3628
rect 798 3602 826 3618
rect 840 3612 856 3628
rect 1704 3612 1720 3628
rect 2744 3612 2760 3628
rect 2424 3592 2440 3608
rect 2664 3592 2680 3608
rect 2862 3602 2890 3618
rect 3064 3612 3080 3628
rect 3768 3612 3784 3628
rect 4664 3612 4680 3628
rect 4168 3592 4184 3608
rect 4910 3602 4938 3618
rect 5112 3612 5128 3628
rect 6456 3612 6472 3628
rect 2232 3572 2248 3588
rect 4648 3572 4664 3588
rect 5288 3592 5304 3608
rect 6264 3592 6280 3608
rect 5224 3572 5240 3588
rect 5800 3572 5816 3588
rect 5912 3572 5928 3588
rect 6392 3572 6408 3588
rect 1960 3552 1976 3568
rect 3192 3552 3208 3568
rect 4360 3552 4376 3568
rect 6072 3552 6088 3568
rect 2424 3532 2440 3548
rect 2568 3532 2584 3548
rect 4600 3532 4616 3548
rect 5112 3532 5128 3548
rect 6024 3532 6040 3548
rect 920 3512 936 3528
rect 1240 3512 1256 3528
rect 1736 3512 1752 3528
rect 2232 3512 2248 3528
rect 2808 3512 2824 3528
rect 3112 3512 3128 3528
rect 3432 3512 3448 3528
rect 3976 3512 3992 3528
rect 6232 3512 6248 3528
rect 856 3492 872 3508
rect 2008 3492 2024 3508
rect 2344 3492 2360 3508
rect 2376 3492 2392 3508
rect 2824 3492 2840 3508
rect 2952 3492 2968 3508
rect 3464 3492 3480 3508
rect 3848 3492 3864 3508
rect 4744 3492 4760 3508
rect 5224 3492 5240 3508
rect 5448 3492 5464 3508
rect 6024 3492 6040 3508
rect 6168 3492 6184 3508
rect 6216 3492 6232 3508
rect 200 3472 216 3488
rect 328 3472 344 3488
rect 536 3472 552 3488
rect 584 3472 616 3488
rect 936 3472 952 3488
rect 1912 3472 1928 3488
rect 3832 3472 3848 3488
rect 4328 3472 4344 3488
rect 6440 3472 6456 3488
rect 2312 3452 2328 3468
rect 3144 3452 3160 3468
rect 3560 3452 3576 3468
rect 3704 3452 3720 3468
rect 4216 3452 4232 3468
rect 4488 3452 4504 3468
rect 5048 3452 5064 3468
rect 5096 3452 5112 3468
rect 664 3432 680 3448
rect 4056 3432 4072 3448
rect 4344 3432 4360 3448
rect 6744 3452 6760 3468
rect 6200 3432 6216 3448
rect 280 3412 296 3428
rect 440 3412 456 3428
rect 1112 3412 1128 3428
rect 1528 3412 1544 3428
rect 600 3392 632 3408
rect 1838 3402 1866 3418
rect 2648 3412 2664 3428
rect 1896 3392 1912 3408
rect 1928 3392 1944 3408
rect 2072 3392 2088 3408
rect 2904 3392 2920 3408
rect 3816 3392 3832 3408
rect 3848 3392 3864 3408
rect 3886 3402 3914 3418
rect 4296 3412 4312 3428
rect 5272 3412 5304 3428
rect 5880 3412 5896 3428
rect 3928 3392 3944 3408
rect 4552 3392 4568 3408
rect 4776 3392 4792 3408
rect 5160 3392 5176 3408
rect 5688 3392 5704 3408
rect 5934 3402 5962 3418
rect 6664 3432 6680 3448
rect 6712 3392 6728 3408
rect 280 3372 296 3388
rect 1512 3372 1528 3388
rect 2200 3372 2216 3388
rect 2248 3372 2264 3388
rect 2408 3372 2424 3388
rect 2568 3372 2584 3388
rect 2616 3372 2632 3388
rect 3800 3372 3816 3388
rect 5416 3372 5432 3388
rect 344 3352 360 3368
rect 360 3352 376 3368
rect 2344 3352 2360 3368
rect 2952 3352 2968 3368
rect 3160 3352 3176 3368
rect 4264 3352 4280 3368
rect 4328 3352 4344 3368
rect 392 3332 408 3348
rect 584 3332 600 3348
rect 600 3332 632 3348
rect 664 3332 680 3348
rect 888 3332 904 3348
rect 1000 3332 1016 3348
rect 2040 3332 2056 3348
rect 2584 3332 2600 3348
rect 2968 3332 2984 3348
rect 3160 3332 3192 3348
rect 3704 3332 3720 3348
rect 4008 3332 4024 3348
rect 5288 3352 5320 3368
rect 5864 3352 5880 3368
rect 6152 3352 6168 3368
rect 6280 3352 6296 3368
rect 4424 3332 4440 3348
rect 4504 3332 4520 3348
rect 4680 3332 4696 3348
rect 5064 3332 5080 3348
rect 5624 3332 5640 3348
rect 5720 3332 5736 3348
rect 6104 3332 6120 3348
rect 328 3312 344 3328
rect 440 3312 456 3328
rect 1064 3312 1080 3328
rect 1176 3312 1192 3328
rect 2072 3312 2088 3328
rect 2840 3312 2856 3328
rect 3944 3312 3960 3328
rect 4072 3312 4088 3328
rect 4376 3312 4392 3328
rect 4392 3312 4408 3328
rect 4472 3312 4488 3328
rect 4552 3312 4568 3328
rect 1992 3292 2008 3308
rect 2200 3292 2216 3308
rect 2472 3292 2488 3308
rect 2664 3272 2680 3288
rect 3192 3292 3208 3308
rect 4248 3292 4264 3308
rect 4360 3292 4376 3308
rect 4408 3292 4424 3308
rect 4584 3292 4600 3308
rect 5016 3312 5032 3328
rect 5432 3312 5448 3328
rect 5656 3312 5672 3328
rect 5832 3312 5848 3328
rect 5192 3292 5208 3308
rect 5640 3292 5656 3308
rect 6200 3292 6216 3308
rect 3128 3272 3144 3288
rect 3528 3272 3544 3288
rect 4344 3272 4360 3288
rect 5896 3272 5912 3288
rect 1016 3252 1032 3268
rect 1432 3252 1448 3268
rect 2712 3252 2728 3268
rect 3496 3252 3512 3268
rect 3832 3252 3848 3268
rect 5080 3252 5096 3268
rect 568 3232 584 3248
rect 1480 3232 1496 3248
rect 1672 3232 1688 3248
rect 4168 3232 4184 3248
rect 5096 3232 5112 3248
rect 6216 3232 6232 3248
rect 798 3202 826 3218
rect 2216 3212 2232 3228
rect 2152 3192 2168 3208
rect 2232 3192 2248 3208
rect 2862 3202 2890 3218
rect 2936 3212 2952 3228
rect 3992 3212 4008 3228
rect 4328 3212 4344 3228
rect 2920 3192 2936 3208
rect 3528 3192 3544 3208
rect 3736 3192 3752 3208
rect 4008 3192 4024 3208
rect 4344 3192 4360 3208
rect 4910 3202 4938 3218
rect 4984 3212 5000 3228
rect 5080 3212 5096 3228
rect 5352 3212 5368 3228
rect 5192 3192 5208 3208
rect 5992 3212 6008 3228
rect 5880 3192 5896 3208
rect 1976 3172 1992 3188
rect 3272 3172 3288 3188
rect 4088 3172 4104 3188
rect 4392 3172 4408 3188
rect 4504 3172 4520 3188
rect 5320 3172 5336 3188
rect 5480 3172 5496 3188
rect 2568 3152 2584 3168
rect 3192 3152 3208 3168
rect 4136 3152 4152 3168
rect 5688 3152 5704 3168
rect 1208 3132 1224 3148
rect 1688 3132 1704 3148
rect 1816 3132 1832 3148
rect 4664 3132 4680 3148
rect 4808 3132 4824 3148
rect 6040 3132 6056 3148
rect 6552 3132 6568 3148
rect 2136 3112 2152 3128
rect 3192 3112 3208 3128
rect 3384 3112 3416 3128
rect 3608 3112 3624 3128
rect 3928 3112 3944 3128
rect 4552 3112 4568 3128
rect 5432 3112 5448 3128
rect 5512 3112 5528 3128
rect 6040 3112 6056 3128
rect 424 3092 440 3108
rect 648 3092 664 3108
rect 1080 3092 1096 3108
rect 1112 3092 1128 3108
rect 1288 3092 1304 3108
rect 2104 3092 2120 3108
rect 3032 3092 3048 3108
rect 408 3072 424 3088
rect 888 3072 904 3088
rect 1320 3072 1336 3088
rect 2184 3072 2200 3088
rect 2616 3072 2632 3088
rect 2696 3072 2712 3088
rect 3144 3072 3160 3088
rect 3176 3072 3192 3088
rect 3368 3092 3384 3108
rect 4712 3092 4744 3108
rect 5336 3092 5352 3108
rect 5368 3092 5384 3108
rect 5528 3092 5544 3108
rect 3544 3072 3560 3088
rect 3688 3072 3704 3088
rect 3848 3072 3864 3088
rect 4008 3072 4024 3088
rect 4312 3072 4328 3088
rect 5256 3072 5272 3088
rect 5720 3072 5736 3088
rect 72 3052 88 3068
rect 1192 3052 1208 3068
rect 1640 3052 1656 3068
rect 2184 3052 2200 3068
rect 2360 3052 2408 3068
rect 2456 3052 2472 3068
rect 2504 3052 2520 3068
rect 2584 3052 2600 3068
rect 3144 3052 3160 3068
rect 3352 3052 3368 3068
rect 3736 3052 3752 3068
rect 3752 3052 3768 3068
rect 4360 3052 4376 3068
rect 4392 3052 4408 3068
rect 1176 3032 1192 3048
rect 1416 3032 1432 3048
rect 1576 3032 1592 3048
rect 1656 3032 1672 3048
rect 1704 3032 1720 3048
rect 1912 3032 1928 3048
rect 2904 3032 2920 3048
rect 3368 3032 3384 3048
rect 3976 3032 3992 3048
rect 5480 3032 5496 3048
rect 5800 3032 5816 3048
rect 840 3012 856 3028
rect 1800 3012 1832 3028
rect 392 2992 408 3008
rect 904 2992 920 3008
rect 1816 2992 1832 3008
rect 1838 3002 1866 3018
rect 2200 2992 2216 3008
rect 3886 3002 3914 3018
rect 4664 3012 4680 3028
rect 5112 3012 5128 3028
rect 4200 2992 4216 3008
rect 4888 2992 4904 3008
rect 5934 3002 5962 3018
rect 6808 2992 6824 3008
rect 1752 2972 1768 2988
rect 2600 2972 2616 2988
rect 3384 2972 3400 2988
rect 4232 2972 4264 2988
rect 4952 2972 4968 2988
rect 5576 2972 5592 2988
rect 216 2952 232 2968
rect 296 2952 312 2968
rect 1720 2952 1736 2968
rect 1784 2952 1800 2968
rect 2088 2952 2104 2968
rect 2216 2952 2232 2968
rect 2392 2952 2408 2968
rect 4776 2952 4792 2968
rect 5896 2952 5912 2968
rect 6808 2952 6824 2968
rect 328 2932 344 2948
rect 648 2932 664 2948
rect 1272 2932 1288 2948
rect 1560 2932 1576 2948
rect 2280 2932 2296 2948
rect 3400 2932 3416 2948
rect 4536 2932 4552 2948
rect 4632 2932 4648 2948
rect 5416 2932 5432 2948
rect 6248 2932 6264 2948
rect 6552 2932 6568 2948
rect 1272 2912 1288 2928
rect 1320 2912 1336 2928
rect 1368 2912 1384 2928
rect 1384 2912 1400 2928
rect 1736 2912 1752 2928
rect 2024 2912 2040 2928
rect 2104 2912 2120 2928
rect 2536 2912 2552 2928
rect 3176 2912 3192 2928
rect 4424 2912 4440 2928
rect 4648 2912 4664 2928
rect 5976 2912 5992 2928
rect 264 2892 280 2908
rect 1064 2892 1080 2908
rect 1160 2892 1176 2908
rect 1400 2892 1416 2908
rect 1656 2892 1672 2908
rect 2184 2892 2200 2908
rect 2952 2892 2968 2908
rect 3080 2892 3096 2908
rect 3192 2892 3208 2908
rect 3752 2892 3768 2908
rect 4168 2892 4184 2908
rect 4440 2892 4456 2908
rect 4840 2892 4856 2908
rect 5128 2892 5144 2908
rect 5976 2892 5992 2908
rect 6712 2912 6728 2928
rect 6712 2892 6728 2908
rect 4648 2872 4664 2888
rect 5416 2872 5432 2888
rect 5624 2872 5640 2888
rect 1032 2852 1048 2868
rect 1800 2852 1816 2868
rect 5208 2852 5224 2868
rect 5544 2852 5560 2868
rect 1704 2832 1720 2848
rect 1816 2832 1832 2848
rect 2152 2832 2168 2848
rect 2568 2832 2584 2848
rect 4328 2832 4344 2848
rect 5176 2832 5192 2848
rect 798 2802 826 2818
rect 2088 2812 2104 2828
rect 2862 2802 2890 2818
rect 3272 2812 3288 2828
rect 3768 2812 3784 2828
rect 4760 2792 4776 2808
rect 4910 2802 4938 2818
rect 6584 2812 6600 2828
rect 6408 2792 6424 2808
rect 200 2772 216 2788
rect 1528 2772 1544 2788
rect 3208 2772 3224 2788
rect 1000 2752 1016 2768
rect 1256 2752 1272 2768
rect 1080 2732 1096 2748
rect 2040 2752 2056 2768
rect 3320 2752 3336 2768
rect 4376 2772 4392 2788
rect 4600 2772 4616 2788
rect 6088 2772 6104 2788
rect 4072 2752 4088 2768
rect 4344 2752 4360 2768
rect 5000 2752 5016 2768
rect 5528 2752 5544 2768
rect 5752 2752 5768 2768
rect 6552 2752 6568 2768
rect 6584 2752 6600 2768
rect 1464 2732 1480 2748
rect 2040 2732 2056 2748
rect 2072 2732 2088 2748
rect 2248 2732 2264 2748
rect 2568 2732 2584 2748
rect 2952 2732 2968 2748
rect 5096 2732 5112 2748
rect 5240 2732 5256 2748
rect 696 2712 712 2728
rect 920 2712 936 2728
rect 2104 2712 2120 2728
rect 2136 2712 2152 2728
rect 3528 2712 3544 2728
rect 5784 2712 5800 2728
rect 5912 2712 5928 2728
rect 1064 2692 1080 2708
rect 1128 2692 1144 2708
rect 1224 2692 1240 2708
rect 1896 2692 1912 2708
rect 1944 2692 1960 2708
rect 2120 2692 2136 2708
rect 2792 2692 2808 2708
rect 3080 2692 3096 2708
rect 3304 2692 3320 2708
rect 3352 2692 3368 2708
rect 3800 2692 3816 2708
rect 4472 2692 4488 2708
rect 4520 2692 4536 2708
rect 4952 2692 4968 2708
rect 5240 2692 5256 2708
rect 328 2672 344 2688
rect 1080 2672 1112 2688
rect 1160 2672 1176 2688
rect 1256 2672 1272 2688
rect 1448 2672 1464 2688
rect 1544 2672 1560 2688
rect 1608 2672 1624 2688
rect 1720 2672 1736 2688
rect 2984 2672 3000 2688
rect 3368 2672 3384 2688
rect 3704 2672 3720 2688
rect 3880 2672 3896 2688
rect 4264 2672 4280 2688
rect 4344 2672 4360 2688
rect 4536 2672 4552 2688
rect 4680 2672 4696 2688
rect 4872 2672 4888 2688
rect 5048 2672 5064 2688
rect 5144 2672 5160 2688
rect 5240 2672 5256 2688
rect 5256 2672 5272 2688
rect 5816 2692 5832 2708
rect 5912 2692 5928 2708
rect 6184 2692 6200 2708
rect 6200 2692 6216 2708
rect 6216 2692 6232 2708
rect 472 2652 488 2668
rect 840 2652 856 2668
rect 1432 2652 1448 2668
rect 1976 2652 1992 2668
rect 1992 2652 2008 2668
rect 2024 2652 2040 2668
rect 2328 2652 2344 2668
rect 1432 2612 1448 2628
rect 2056 2632 2072 2648
rect 2232 2632 2248 2648
rect 2760 2652 2776 2668
rect 3480 2652 3496 2668
rect 3672 2652 3688 2668
rect 4744 2652 4760 2668
rect 5864 2672 5880 2688
rect 5992 2672 6008 2688
rect 6232 2672 6248 2688
rect 3240 2632 3256 2648
rect 4728 2632 4744 2648
rect 5528 2632 5544 2648
rect 6200 2632 6216 2648
rect 6248 2632 6264 2648
rect 1784 2612 1800 2628
rect 1592 2592 1608 2608
rect 1624 2592 1640 2608
rect 1838 2602 1866 2618
rect 2600 2612 2616 2628
rect 3864 2612 3880 2628
rect 2088 2592 2104 2608
rect 2264 2592 2280 2608
rect 2392 2592 2408 2608
rect 2680 2592 2696 2608
rect 3144 2592 3160 2608
rect 3832 2592 3848 2608
rect 3886 2602 3914 2618
rect 3960 2612 3976 2628
rect 4632 2612 4648 2628
rect 5912 2612 5928 2628
rect 5480 2592 5496 2608
rect 5512 2592 5528 2608
rect 5934 2602 5962 2618
rect 5992 2612 6008 2628
rect 424 2572 456 2588
rect 1528 2572 1544 2588
rect 2760 2572 2776 2588
rect 2936 2572 2952 2588
rect 2952 2572 2968 2588
rect 1240 2552 1256 2568
rect 2888 2552 2904 2568
rect 3784 2552 3800 2568
rect 4488 2552 4504 2568
rect 4664 2552 4680 2568
rect 5208 2552 5224 2568
rect 5256 2552 5272 2568
rect 5992 2552 6008 2568
rect 6040 2552 6056 2568
rect 1144 2532 1160 2548
rect 1304 2532 1320 2548
rect 1496 2532 1512 2548
rect 1720 2532 1736 2548
rect 1816 2532 1832 2548
rect 2344 2532 2360 2548
rect 2456 2532 2472 2548
rect 2776 2532 2792 2548
rect 2824 2532 2840 2548
rect 2968 2532 2984 2548
rect 3032 2532 3048 2548
rect 3544 2532 3560 2548
rect 3832 2532 3848 2548
rect 4280 2532 4296 2548
rect 4408 2532 4424 2548
rect 4488 2532 4504 2548
rect 4808 2532 4824 2548
rect 5144 2532 5160 2548
rect 5416 2532 5432 2548
rect 5512 2532 5528 2548
rect 5544 2532 5560 2548
rect 5672 2532 5688 2548
rect 6760 2552 6776 2568
rect 6440 2532 6456 2548
rect 6712 2532 6728 2548
rect 776 2512 792 2528
rect 856 2512 872 2528
rect 952 2512 968 2528
rect 1144 2512 1160 2528
rect 1560 2512 1576 2528
rect 1992 2512 2008 2528
rect 2216 2512 2232 2528
rect 2504 2512 2520 2528
rect 3000 2512 3016 2528
rect 3048 2512 3064 2528
rect 3560 2512 3576 2528
rect 4040 2512 4056 2528
rect 4328 2512 4344 2528
rect 4760 2512 4776 2528
rect 6088 2512 6104 2528
rect 6120 2512 6136 2528
rect 6216 2512 6232 2528
rect 6616 2512 6632 2528
rect 6648 2512 6664 2528
rect 680 2492 712 2508
rect 1336 2492 1352 2508
rect 1384 2492 1400 2508
rect 2440 2492 2456 2508
rect 4872 2492 4888 2508
rect 5752 2492 5768 2508
rect 6040 2492 6056 2508
rect 6408 2492 6424 2508
rect 1960 2472 1976 2488
rect 2152 2472 2168 2488
rect 2360 2472 2376 2488
rect 520 2452 536 2468
rect 1048 2432 1064 2448
rect 1352 2432 1368 2448
rect 2632 2452 2648 2468
rect 4360 2472 4376 2488
rect 4040 2452 4056 2468
rect 5368 2452 5384 2468
rect 5400 2452 5416 2468
rect 1688 2432 1704 2448
rect 3352 2432 3368 2448
rect 3512 2432 3528 2448
rect 4632 2432 4648 2448
rect 5448 2432 5464 2448
rect 5512 2432 5528 2448
rect 488 2412 504 2428
rect 632 2412 648 2428
rect 296 2392 312 2408
rect 408 2392 424 2408
rect 798 2402 826 2418
rect 1496 2412 1512 2428
rect 2408 2412 2424 2428
rect 2456 2412 2472 2428
rect 2840 2412 2856 2428
rect 1544 2392 1560 2408
rect 1704 2392 1720 2408
rect 2248 2392 2264 2408
rect 2862 2402 2890 2418
rect 4008 2412 4024 2428
rect 2904 2392 2920 2408
rect 4072 2392 4088 2408
rect 4456 2392 4472 2408
rect 4888 2392 4904 2408
rect 4910 2402 4938 2418
rect 5176 2392 5192 2408
rect 5256 2392 5272 2408
rect 5736 2392 5752 2408
rect 3208 2372 3240 2388
rect 3656 2372 3672 2388
rect 4056 2372 4072 2388
rect 5432 2372 5448 2388
rect 5896 2372 5912 2388
rect 664 2352 680 2368
rect 1416 2352 1432 2368
rect 2168 2352 2184 2368
rect 2648 2352 2664 2368
rect 4344 2352 4360 2368
rect 6696 2352 6712 2368
rect 2072 2332 2088 2348
rect 2728 2332 2744 2348
rect 3016 2332 3032 2348
rect 1432 2312 1448 2328
rect 1464 2312 1480 2328
rect 2408 2312 2424 2328
rect 3144 2312 3160 2328
rect 3320 2312 3336 2328
rect 3848 2312 3864 2328
rect 4024 2312 4040 2328
rect 4392 2312 4408 2328
rect 4792 2312 4808 2328
rect 472 2292 488 2308
rect 680 2292 696 2308
rect 936 2292 952 2308
rect 1352 2292 1368 2308
rect 2120 2292 2136 2308
rect 3096 2292 3112 2308
rect 3176 2292 3192 2308
rect 3352 2292 3368 2308
rect 3416 2292 3432 2308
rect 3704 2292 3720 2308
rect 3848 2292 3864 2308
rect 3928 2292 3944 2308
rect 4712 2292 4728 2308
rect 5416 2292 5432 2308
rect 5832 2292 5848 2308
rect 6408 2292 6424 2308
rect 1256 2272 1272 2288
rect 1608 2272 1624 2288
rect 1736 2272 1752 2288
rect 2088 2272 2104 2288
rect 2136 2272 2152 2288
rect 2424 2272 2440 2288
rect 2584 2272 2600 2288
rect 2792 2272 2808 2288
rect 3464 2272 3480 2288
rect 3864 2272 3880 2288
rect 4344 2272 4360 2288
rect 1400 2252 1416 2268
rect 2600 2252 2616 2268
rect 2856 2252 2872 2268
rect 3080 2252 3096 2268
rect 3416 2252 3432 2268
rect 3512 2252 3528 2268
rect 3992 2252 4008 2268
rect 4024 2252 4040 2268
rect 4648 2272 4664 2288
rect 5688 2272 5704 2288
rect 5896 2272 5912 2288
rect 5976 2272 5992 2288
rect 6040 2272 6056 2288
rect 6392 2272 6408 2288
rect 6424 2272 6440 2288
rect 6440 2252 6456 2268
rect 184 2232 200 2248
rect 456 2232 472 2248
rect 568 2232 584 2248
rect 904 2232 920 2248
rect 1032 2232 1048 2248
rect 1928 2232 1944 2248
rect 1992 2232 2008 2248
rect 2040 2232 2056 2248
rect 2632 2232 2648 2248
rect 5736 2232 5752 2248
rect 6104 2232 6120 2248
rect 248 2212 264 2228
rect 696 2212 712 2228
rect 1480 2212 1496 2228
rect 712 2192 728 2208
rect 1560 2192 1576 2208
rect 1592 2192 1608 2208
rect 1838 2202 1866 2218
rect 3224 2212 3240 2228
rect 3544 2212 3560 2228
rect 3886 2202 3914 2218
rect 4264 2212 4296 2228
rect 4552 2212 4568 2228
rect 4680 2212 4696 2228
rect 4280 2192 4296 2208
rect 4488 2192 4504 2208
rect 5384 2192 5400 2208
rect 5496 2192 5512 2208
rect 5934 2202 5962 2218
rect 6632 2192 6648 2208
rect 360 2172 376 2188
rect 856 2172 872 2188
rect 968 2172 984 2188
rect 1144 2172 1160 2188
rect 1448 2172 1464 2188
rect 2072 2172 2104 2188
rect 2824 2172 2840 2188
rect 3208 2172 3224 2188
rect 3320 2172 3336 2188
rect 3496 2172 3512 2188
rect 3576 2172 3592 2188
rect 3816 2172 3832 2188
rect 4216 2172 4232 2188
rect 4536 2172 4552 2188
rect 1432 2152 1448 2168
rect 4088 2152 4104 2168
rect 5528 2152 5544 2168
rect 5624 2152 5640 2168
rect 6424 2152 6440 2168
rect 200 2132 216 2148
rect 296 2132 312 2148
rect 536 2132 552 2148
rect 648 2132 664 2148
rect 840 2132 856 2148
rect 1272 2132 1288 2148
rect 1752 2132 1768 2148
rect 2248 2132 2264 2148
rect 2280 2132 2296 2148
rect 2504 2132 2520 2148
rect 2536 2132 2552 2148
rect 2728 2132 2744 2148
rect 2792 2132 2808 2148
rect 3368 2132 3384 2148
rect 4824 2132 4840 2148
rect 5240 2132 5256 2148
rect 6456 2132 6472 2148
rect 6552 2132 6568 2148
rect 232 2112 248 2128
rect 1256 2112 1272 2128
rect 1640 2112 1656 2128
rect 2520 2112 2536 2128
rect 2776 2112 2792 2128
rect 3512 2112 3528 2128
rect 3544 2112 3560 2128
rect 3576 2112 3592 2128
rect 3608 2112 3624 2128
rect 4072 2112 4088 2128
rect 4184 2112 4200 2128
rect 1672 2092 1688 2108
rect 1784 2092 1800 2108
rect 2024 2092 2040 2108
rect 2968 2092 2984 2108
rect 3032 2092 3048 2108
rect 4024 2092 4040 2108
rect 4312 2092 4328 2108
rect 5864 2112 5880 2128
rect 6376 2112 6392 2128
rect 6632 2112 6648 2128
rect 5416 2092 5432 2108
rect 6504 2092 6520 2108
rect 504 2072 520 2088
rect 616 2072 632 2088
rect 1080 2072 1096 2088
rect 1720 2072 1736 2088
rect 2216 2072 2232 2088
rect 5992 2072 6008 2088
rect 1224 2052 1240 2068
rect 2200 2052 2216 2068
rect 5384 2052 5400 2068
rect 2472 2032 2488 2048
rect 4424 2032 4440 2048
rect 5192 2032 5208 2048
rect 280 2012 296 2028
rect 798 2002 826 2018
rect 1400 2012 1416 2028
rect 2392 2012 2408 2028
rect 1144 1992 1160 2008
rect 2328 1992 2344 2008
rect 2862 2002 2890 2018
rect 3064 2012 3080 2028
rect 4120 2012 4136 2028
rect 4248 2012 4264 2028
rect 3400 1992 3416 2008
rect 4520 1992 4536 2008
rect 4910 2002 4938 2018
rect 5352 2012 5368 2028
rect 5000 1992 5016 2008
rect 5576 1992 5592 2008
rect 392 1972 408 1988
rect 424 1972 440 1988
rect 4392 1972 4408 1988
rect 1592 1952 1608 1968
rect 2056 1952 2088 1968
rect 4232 1952 4248 1968
rect 5880 1952 5896 1968
rect 6520 1952 6536 1968
rect 648 1932 664 1948
rect 2968 1932 2984 1948
rect 3128 1932 3144 1948
rect 6040 1932 6056 1948
rect 6184 1932 6200 1948
rect 6728 1932 6744 1948
rect 840 1912 856 1928
rect 1288 1912 1304 1928
rect 2392 1912 2408 1928
rect 3048 1912 3080 1928
rect 3992 1912 4008 1928
rect 4264 1912 4280 1928
rect 6408 1912 6424 1928
rect 328 1892 344 1908
rect 376 1892 392 1908
rect 408 1892 424 1908
rect 1192 1892 1208 1908
rect 1496 1892 1512 1908
rect 1768 1892 1784 1908
rect 1880 1892 1896 1908
rect 2072 1892 2088 1908
rect 2312 1892 2328 1908
rect 2328 1892 2344 1908
rect 2456 1892 2472 1908
rect 2696 1892 2712 1908
rect 3208 1892 3224 1908
rect 3512 1892 3528 1908
rect 3704 1892 3720 1908
rect 3848 1892 3864 1908
rect 3976 1892 3992 1908
rect 4008 1892 4024 1908
rect 4376 1892 4392 1908
rect 4600 1892 4616 1908
rect 5464 1892 5480 1908
rect 5512 1892 5528 1908
rect 6456 1892 6472 1908
rect 6632 1892 6648 1908
rect 6696 1892 6712 1908
rect 200 1872 216 1888
rect 440 1872 456 1888
rect 520 1872 536 1888
rect 664 1872 696 1888
rect 1560 1872 1576 1888
rect 1896 1872 1912 1888
rect 2168 1872 2184 1888
rect 2504 1872 2520 1888
rect 2680 1872 2696 1888
rect 3160 1872 3176 1888
rect 4120 1872 4136 1888
rect 4232 1872 4248 1888
rect 5032 1872 5048 1888
rect 5480 1872 5496 1888
rect 6008 1872 6024 1888
rect 1048 1852 1064 1868
rect 1448 1852 1464 1868
rect 3240 1852 3256 1868
rect 4056 1852 4072 1868
rect 4248 1852 4264 1868
rect 5048 1852 5064 1868
rect 6184 1852 6200 1868
rect 632 1832 648 1848
rect 920 1832 936 1848
rect 2328 1832 2344 1848
rect 3080 1832 3096 1848
rect 3784 1832 3800 1848
rect 4040 1832 4056 1848
rect 4088 1832 4104 1848
rect 4952 1832 4968 1848
rect 6440 1832 6456 1848
rect 6552 1832 6568 1848
rect 968 1792 984 1808
rect 1432 1792 1448 1808
rect 1576 1792 1592 1808
rect 1838 1802 1866 1818
rect 3496 1812 3512 1828
rect 1880 1792 1896 1808
rect 3016 1792 3032 1808
rect 3886 1802 3914 1818
rect 5096 1812 5112 1828
rect 5224 1792 5240 1808
rect 5688 1792 5704 1808
rect 5934 1802 5962 1818
rect 6040 1792 6056 1808
rect 6232 1792 6248 1808
rect 648 1772 664 1788
rect 1320 1772 1336 1788
rect 1624 1772 1640 1788
rect 2440 1772 2456 1788
rect 2728 1772 2744 1788
rect 3048 1772 3064 1788
rect 3384 1772 3400 1788
rect 3848 1772 3864 1788
rect 5000 1772 5016 1788
rect 5208 1772 5224 1788
rect 6216 1772 6232 1788
rect 1304 1752 1320 1768
rect 1640 1752 1656 1768
rect 2840 1752 2856 1768
rect 3224 1752 3240 1768
rect 4296 1752 4312 1768
rect 4888 1752 4904 1768
rect 6712 1752 6728 1768
rect 248 1732 264 1748
rect 504 1732 520 1748
rect 952 1732 968 1748
rect 968 1732 984 1748
rect 1032 1732 1048 1748
rect 1288 1732 1304 1748
rect 1496 1732 1528 1748
rect 1720 1732 1736 1748
rect 2088 1732 2104 1748
rect 2184 1732 2200 1748
rect 3416 1732 3432 1748
rect 776 1712 792 1728
rect 888 1712 904 1728
rect 1112 1712 1128 1728
rect 1144 1712 1160 1728
rect 1272 1712 1288 1728
rect 1752 1712 1784 1728
rect 2280 1712 2296 1728
rect 2968 1712 2984 1728
rect 3336 1712 3368 1728
rect 3704 1712 3720 1728
rect 4104 1732 4120 1748
rect 4536 1732 4552 1748
rect 5880 1732 5896 1748
rect 6504 1732 6520 1748
rect 392 1692 408 1708
rect 1016 1692 1032 1708
rect 1384 1692 1400 1708
rect 1896 1692 1912 1708
rect 3224 1692 3240 1708
rect 4200 1692 4216 1708
rect 5112 1712 5128 1728
rect 5384 1712 5400 1728
rect 5992 1712 6008 1728
rect 6040 1712 6056 1728
rect 6648 1712 6664 1728
rect 4744 1692 4760 1708
rect 888 1672 904 1688
rect 1112 1672 1128 1688
rect 1688 1672 1704 1688
rect 2664 1672 2680 1688
rect 2200 1652 2216 1668
rect 3400 1652 3416 1668
rect 3864 1652 3880 1668
rect 3928 1652 3944 1668
rect 4264 1652 4280 1668
rect 5080 1652 5096 1668
rect 600 1632 616 1648
rect 1352 1632 1368 1648
rect 2936 1632 2952 1648
rect 3384 1632 3400 1648
rect 6040 1632 6056 1648
rect 424 1592 440 1608
rect 798 1602 826 1618
rect 1608 1612 1624 1628
rect 904 1592 920 1608
rect 1064 1592 1080 1608
rect 2862 1602 2890 1618
rect 3544 1612 3560 1628
rect 3000 1592 3016 1608
rect 4312 1612 4328 1628
rect 3144 1572 3160 1588
rect 4910 1602 4938 1618
rect 6376 1592 6392 1608
rect 4328 1572 4344 1588
rect 4872 1572 4888 1588
rect 5800 1572 5816 1588
rect 424 1552 440 1568
rect 2392 1552 2408 1568
rect 2552 1552 2568 1568
rect 536 1532 552 1548
rect 1304 1532 1320 1548
rect 2360 1532 2376 1548
rect 2536 1532 2552 1548
rect 4824 1552 4840 1568
rect 5336 1552 5352 1568
rect 4680 1532 4696 1548
rect 6200 1532 6232 1548
rect 6408 1532 6424 1548
rect 6600 1532 6616 1548
rect 1528 1512 1544 1528
rect 2168 1512 2184 1528
rect 2616 1512 2632 1528
rect 2808 1512 2840 1528
rect 3976 1512 3992 1528
rect 4552 1512 4568 1528
rect 5256 1512 5272 1528
rect 5848 1512 5864 1528
rect 488 1492 504 1508
rect 1448 1492 1464 1508
rect 2408 1492 2424 1508
rect 3080 1492 3096 1508
rect 3512 1492 3528 1508
rect 3656 1492 3672 1508
rect 3688 1492 3704 1508
rect 3816 1492 3832 1508
rect 3848 1492 3864 1508
rect 4248 1492 4264 1508
rect 4376 1492 4392 1508
rect 200 1452 216 1468
rect 312 1452 328 1468
rect 760 1472 776 1488
rect 1160 1472 1176 1488
rect 2200 1472 2216 1488
rect 2328 1472 2344 1488
rect 2664 1472 2680 1488
rect 2696 1472 2712 1488
rect 2920 1472 2936 1488
rect 3096 1472 3112 1488
rect 3208 1472 3224 1488
rect 3672 1472 3688 1488
rect 3752 1472 3768 1488
rect 4424 1472 4440 1488
rect 4680 1492 4696 1508
rect 4728 1472 4744 1488
rect 4760 1472 4776 1488
rect 6200 1492 6216 1508
rect 6584 1492 6600 1508
rect 6696 1492 6712 1508
rect 6728 1492 6744 1508
rect 5896 1472 5912 1488
rect 6392 1472 6408 1488
rect 6584 1472 6600 1488
rect 1528 1452 1544 1468
rect 2440 1452 2456 1468
rect 3736 1452 3752 1468
rect 6456 1452 6472 1468
rect 1480 1432 1496 1448
rect 1544 1432 1560 1448
rect 1720 1432 1736 1448
rect 2744 1432 2760 1448
rect 3208 1432 3224 1448
rect 4648 1432 4664 1448
rect 696 1412 712 1428
rect 1304 1412 1320 1428
rect 904 1392 920 1408
rect 1112 1392 1128 1408
rect 1838 1402 1866 1418
rect 2328 1412 2344 1428
rect 3192 1412 3208 1428
rect 2120 1392 2136 1408
rect 3886 1402 3914 1418
rect 3976 1412 3992 1428
rect 4824 1412 4840 1428
rect 3928 1392 3944 1408
rect 4952 1392 4968 1408
rect 4984 1392 5000 1408
rect 600 1372 616 1388
rect 4088 1372 4104 1388
rect 4168 1372 4184 1388
rect 4200 1372 4216 1388
rect 4696 1372 4712 1388
rect 5934 1402 5962 1418
rect 6440 1412 6456 1428
rect 6424 1392 6440 1408
rect 6728 1392 6744 1408
rect 6328 1372 6344 1388
rect 360 1352 376 1368
rect 1208 1352 1224 1368
rect 1544 1352 1560 1368
rect 1736 1352 1752 1368
rect 2104 1352 2120 1368
rect 2168 1352 2184 1368
rect 3928 1352 3944 1368
rect 5480 1352 5496 1368
rect 888 1332 904 1348
rect 920 1332 936 1348
rect 1080 1332 1096 1348
rect 1640 1332 1656 1348
rect 1672 1332 1688 1348
rect 1752 1332 1768 1348
rect 3432 1332 3448 1348
rect 3928 1332 3944 1348
rect 3960 1332 3976 1348
rect 4680 1332 4696 1348
rect 168 1312 184 1328
rect 264 1312 280 1328
rect 984 1312 1000 1328
rect 1576 1312 1592 1328
rect 1912 1312 1928 1328
rect 2136 1312 2152 1328
rect 2264 1312 2280 1328
rect 2360 1312 2376 1328
rect 2632 1312 2648 1328
rect 2792 1312 2808 1328
rect 2824 1312 2840 1328
rect 2856 1312 2872 1328
rect 3032 1312 3048 1328
rect 3768 1312 3784 1328
rect 4088 1312 4104 1328
rect 4696 1312 4712 1328
rect 4744 1312 4760 1328
rect 5016 1312 5032 1328
rect 5064 1312 5080 1328
rect 6648 1352 6664 1368
rect 6728 1332 6744 1348
rect 5416 1312 5432 1328
rect 6520 1312 6536 1328
rect 6632 1312 6648 1328
rect 6712 1312 6728 1328
rect 1928 1292 1944 1308
rect 2824 1292 2840 1308
rect 5400 1292 5416 1308
rect 5688 1292 5704 1308
rect 6696 1292 6712 1308
rect 2056 1272 2072 1288
rect 3560 1272 3576 1288
rect 4344 1272 4360 1288
rect 5896 1272 5912 1288
rect 6200 1272 6216 1288
rect 1800 1252 1816 1268
rect 4008 1252 4024 1268
rect 4856 1252 4872 1268
rect 2040 1232 2056 1248
rect 3320 1232 3336 1248
rect 3656 1232 3672 1248
rect 5624 1232 5640 1248
rect 5752 1232 5768 1248
rect 798 1202 826 1218
rect 1784 1212 1800 1228
rect 2862 1202 2890 1218
rect 3112 1212 3128 1228
rect 4264 1212 4296 1228
rect 4910 1202 4938 1218
rect 4968 1192 4984 1208
rect 5464 1192 5480 1208
rect 2088 1172 2104 1188
rect 3448 1172 3464 1188
rect 3976 1172 3992 1188
rect 424 1152 440 1168
rect 1608 1152 1624 1168
rect 2152 1152 2168 1168
rect 2680 1152 2696 1168
rect 2744 1152 2760 1168
rect 3784 1152 3800 1168
rect 4888 1152 4904 1168
rect 5528 1152 5544 1168
rect 6216 1152 6232 1168
rect 6232 1152 6248 1168
rect 4120 1132 4136 1148
rect 4472 1132 4488 1148
rect 4968 1132 4984 1148
rect 1048 1112 1080 1128
rect 2360 1112 2376 1128
rect 3576 1112 3592 1128
rect 4568 1112 4584 1128
rect 1800 1092 1816 1108
rect 1928 1092 1944 1108
rect 2120 1092 2136 1108
rect 1032 1072 1048 1088
rect 1224 1072 1240 1088
rect 2952 1092 2968 1108
rect 3048 1092 3064 1108
rect 3256 1092 3272 1108
rect 3352 1092 3368 1108
rect 3864 1092 3880 1108
rect 4872 1092 4888 1108
rect 3160 1072 3176 1088
rect 3528 1072 3544 1088
rect 3928 1072 3944 1088
rect 488 1032 504 1048
rect 920 1032 936 1048
rect 1048 1052 1064 1068
rect 1208 1052 1224 1068
rect 1240 1052 1256 1068
rect 1384 1052 1400 1068
rect 1704 1052 1720 1068
rect 1288 1032 1304 1048
rect 1816 1032 1832 1048
rect 1976 1032 1992 1048
rect 2424 1052 2440 1068
rect 3000 1052 3016 1068
rect 3128 1052 3144 1068
rect 4632 1072 4648 1088
rect 5512 1092 5528 1108
rect 5368 1072 5400 1088
rect 4824 1052 4840 1068
rect 6216 1072 6232 1088
rect 4920 1032 4936 1048
rect 584 992 600 1008
rect 1816 992 1832 1008
rect 1838 1002 1866 1018
rect 1960 1012 1976 1028
rect 2216 1012 2232 1028
rect 2312 1012 2328 1028
rect 2408 1012 2424 1028
rect 3272 1012 3288 1028
rect 1080 972 1096 988
rect 1464 972 1480 988
rect 2312 972 2328 988
rect 3160 992 3176 1008
rect 3864 992 3880 1008
rect 3886 1002 3914 1018
rect 4504 992 4520 1008
rect 4920 992 4936 1008
rect 5688 992 5704 1008
rect 5934 1002 5962 1018
rect 5976 1012 5992 1028
rect 6120 1012 6136 1028
rect 6424 1012 6440 1028
rect 6136 992 6152 1008
rect 6520 992 6536 1008
rect 1960 952 1976 968
rect 3480 972 3496 988
rect 3512 972 3528 988
rect 5224 972 5240 988
rect 5544 972 5560 988
rect 6376 972 6392 988
rect 3032 952 3048 968
rect 3176 952 3192 968
rect 3480 952 3496 968
rect 3608 952 3624 968
rect 4696 952 4712 968
rect 312 932 328 948
rect 488 932 504 948
rect 1112 932 1128 948
rect 1288 932 1304 948
rect 1752 932 1768 948
rect 2280 932 2296 948
rect 2920 932 2936 948
rect 4168 932 4184 948
rect 4856 932 4872 948
rect 5160 932 5176 948
rect 5208 932 5224 948
rect 184 912 200 928
rect 360 912 392 928
rect 1208 912 1224 928
rect 1304 912 1320 928
rect 1368 912 1384 928
rect 2104 912 2120 928
rect 2120 912 2136 928
rect 2152 912 2168 928
rect 3256 912 3272 928
rect 3464 912 3480 928
rect 4312 912 4328 928
rect 4376 912 4392 928
rect 6408 932 6424 948
rect 6520 932 6536 948
rect 5640 912 5656 928
rect 776 892 792 908
rect 1064 892 1080 908
rect 1080 892 1096 908
rect 3096 892 3112 908
rect 3576 892 3592 908
rect 3720 892 3736 908
rect 4552 892 4568 908
rect 5384 892 5400 908
rect 1896 872 1912 888
rect 2344 872 2360 888
rect 1256 852 1272 868
rect 3432 852 3464 868
rect 4296 852 4312 868
rect 2200 832 2216 848
rect 4424 832 4440 848
rect 5544 852 5560 868
rect 6200 852 6216 868
rect 6552 852 6568 868
rect 6632 832 6648 848
rect 798 802 826 818
rect 984 812 1000 828
rect 1608 812 1624 828
rect 2152 812 2168 828
rect 2328 792 2344 808
rect 2840 792 2856 808
rect 2862 802 2890 818
rect 2984 812 3000 828
rect 4744 812 4760 828
rect 3544 792 3560 808
rect 3560 792 3576 808
rect 3720 792 3736 808
rect 4680 792 4696 808
rect 4910 802 4938 818
rect 2008 772 2024 788
rect 5288 772 5304 788
rect 2984 752 3000 768
rect 3192 752 3208 768
rect 5624 752 5640 768
rect 1384 732 1400 748
rect 2312 732 2328 748
rect 4360 732 4376 748
rect 1144 712 1160 728
rect 1192 712 1208 728
rect 2216 712 2232 728
rect 2360 712 2376 728
rect 2584 712 2616 728
rect 3288 712 3304 728
rect 3528 712 3544 728
rect 4280 712 4296 728
rect 4696 732 4712 748
rect 4392 712 4408 728
rect 4776 712 4792 728
rect 4888 712 4904 728
rect 5096 712 5128 728
rect 5160 712 5176 728
rect 168 692 184 708
rect 1224 692 1240 708
rect 1288 692 1304 708
rect 1352 692 1368 708
rect 1512 692 1528 708
rect 2456 692 2472 708
rect 5528 712 5544 728
rect 2904 692 2920 708
rect 2936 692 2952 708
rect 3672 692 3688 708
rect 3720 692 3736 708
rect 3784 692 3800 708
rect 4424 692 4440 708
rect 5304 692 5320 708
rect 5352 692 5368 708
rect 6728 692 6744 708
rect 568 672 584 688
rect 680 672 696 688
rect 1496 672 1512 688
rect 1976 672 1992 688
rect 2008 672 2040 688
rect 2424 672 2440 688
rect 3208 672 3224 688
rect 3688 672 3704 688
rect 3752 672 3768 688
rect 3864 672 3880 688
rect 4200 672 4216 688
rect 5496 672 5512 688
rect 6792 672 6808 688
rect 2088 652 2104 668
rect 3512 652 3528 668
rect 3896 652 3912 668
rect 4536 652 4552 668
rect 4728 652 4744 668
rect 680 632 696 648
rect 1560 612 1576 628
rect 1112 592 1128 608
rect 1838 602 1866 618
rect 2696 612 2712 628
rect 3192 632 3208 648
rect 3208 632 3224 648
rect 3416 632 3432 648
rect 4280 632 4296 648
rect 3886 602 3914 618
rect 4840 612 4856 628
rect 4952 612 4968 628
rect 4984 612 5000 628
rect 5256 612 5272 628
rect 4472 592 4488 608
rect 4568 592 4600 608
rect 5336 592 5352 608
rect 5934 602 5962 618
rect 1400 572 1416 588
rect 1912 572 1928 588
rect 2280 572 2296 588
rect 2328 572 2344 588
rect 3448 572 3464 588
rect 488 552 504 568
rect 1128 552 1144 568
rect 1800 552 1816 568
rect 2424 552 2440 568
rect 3176 552 3192 568
rect 3688 552 3704 568
rect 4456 572 4472 588
rect 5512 572 5528 588
rect 5768 572 5784 588
rect 168 532 184 548
rect 3560 532 3576 548
rect 3784 532 3800 548
rect 4040 532 4056 548
rect 4264 552 4280 568
rect 4584 552 4600 568
rect 5160 552 5176 568
rect 5256 552 5272 568
rect 5640 552 5656 568
rect 6120 552 6136 568
rect 4776 532 4792 548
rect 4792 532 4808 548
rect 5368 532 5384 548
rect 5960 532 5976 548
rect 6120 532 6136 548
rect 1160 512 1176 528
rect 1192 512 1208 528
rect 1256 512 1272 528
rect 1496 512 1512 528
rect 2344 512 2360 528
rect 3656 512 3688 528
rect 3752 512 3768 528
rect 3768 512 3784 528
rect 4104 512 4120 528
rect 4248 512 4264 528
rect 5000 512 5016 528
rect 5192 512 5208 528
rect 5624 512 5640 528
rect 5768 512 5784 528
rect 2600 492 2616 508
rect 2696 492 2712 508
rect 3320 492 3336 508
rect 4584 492 4600 508
rect 4616 492 4632 508
rect 4648 492 4664 508
rect 4952 492 4968 508
rect 5688 492 5704 508
rect 552 472 568 488
rect 1384 472 1400 488
rect 2904 472 2920 488
rect 3544 472 3560 488
rect 5304 472 5320 488
rect 6472 492 6488 508
rect 1912 452 1928 468
rect 2360 452 2376 468
rect 3768 452 3784 468
rect 3784 452 3800 468
rect 3928 452 3944 468
rect 4360 452 4376 468
rect 5544 452 5560 468
rect 2488 432 2504 448
rect 4280 432 4296 448
rect 4728 432 4744 448
rect 760 412 776 428
rect 798 402 826 418
rect 840 412 856 428
rect 2808 412 2824 428
rect 2392 392 2408 408
rect 2862 402 2890 418
rect 2904 412 2920 428
rect 3656 392 3672 408
rect 4680 392 4696 408
rect 4888 392 4904 408
rect 4910 402 4938 418
rect 5208 412 5224 428
rect 3592 372 3608 388
rect 3672 372 3688 388
rect 5224 392 5240 408
rect 5288 392 5304 408
rect 5000 372 5016 388
rect 6760 372 6776 388
rect 280 352 296 368
rect 424 352 440 368
rect 3928 352 3944 368
rect 4232 352 4248 368
rect 4984 352 5000 368
rect 5208 352 5224 368
rect 2504 332 2520 348
rect 2968 332 2984 348
rect 4232 332 4248 348
rect 4296 332 4312 348
rect 4872 332 4888 348
rect 680 312 696 328
rect 712 312 728 328
rect 728 312 744 328
rect 840 312 856 328
rect 872 312 888 328
rect 1176 312 1192 328
rect 2376 312 2392 328
rect 2952 312 2968 328
rect 3480 312 3496 328
rect 5544 312 5560 328
rect 6616 312 6632 328
rect 376 292 392 308
rect 2312 292 2328 308
rect 3304 292 3320 308
rect 3448 292 3464 308
rect 3576 292 3592 308
rect 3656 292 3672 308
rect 3704 292 3720 308
rect 3816 292 3832 308
rect 3864 292 3880 308
rect 4904 292 4920 308
rect 4952 292 4968 308
rect 5048 292 5064 308
rect 5064 292 5080 308
rect 6568 292 6584 308
rect 6744 292 6760 308
rect 360 272 376 288
rect 1272 272 1288 288
rect 1592 272 1608 288
rect 2712 272 2728 288
rect 3240 272 3256 288
rect 3256 272 3272 288
rect 3272 272 3288 288
rect 3416 272 3432 288
rect 568 252 584 268
rect 1688 252 1704 268
rect 2344 252 2360 268
rect 2424 252 2440 268
rect 2824 252 2840 268
rect 3624 272 3640 288
rect 3656 272 3672 288
rect 3688 272 3720 288
rect 3864 272 3880 288
rect 3960 272 3976 288
rect 3976 272 3992 288
rect 4424 272 4440 288
rect 4584 272 4600 288
rect 4600 272 4616 288
rect 5624 272 5640 288
rect 3464 252 3480 268
rect 4376 252 4392 268
rect 4728 252 4760 268
rect 5320 252 5336 268
rect 5448 252 5464 268
rect 6136 252 6152 268
rect 3672 232 3688 248
rect 4952 232 4968 248
rect 5912 232 5928 248
rect 5960 232 5976 248
rect 1784 212 1800 228
rect 1838 202 1866 218
rect 3768 212 3784 228
rect 2184 192 2200 208
rect 3886 202 3914 218
rect 4360 192 4376 208
rect 5934 202 5962 218
rect 3128 172 3144 188
rect 4280 172 4296 188
rect 4360 172 4376 188
rect 6008 172 6024 188
rect 6584 172 6616 188
rect 920 152 936 168
rect 1160 152 1176 168
rect 1400 152 1416 168
rect 2152 152 2168 168
rect 3176 152 3192 168
rect 3928 152 3944 168
rect 4984 152 5000 168
rect 5336 152 5352 168
rect 6504 152 6520 168
rect 584 132 600 148
rect 1144 132 1160 148
rect 1176 132 1192 148
rect 1272 132 1288 148
rect 1688 132 1704 148
rect 2392 132 2408 148
rect 2440 132 2456 148
rect 2456 132 2472 148
rect 2488 132 2504 148
rect 2696 132 2712 148
rect 1016 112 1032 128
rect 1320 112 1352 128
rect 1272 92 1288 108
rect 2216 92 2232 108
rect 2344 112 2360 128
rect 2408 112 2424 128
rect 2552 112 2568 128
rect 3288 92 3304 108
rect 3768 112 3784 128
rect 4472 112 4488 128
rect 5000 112 5016 128
rect 5320 112 5336 128
rect 5640 112 5656 128
rect 6328 112 6344 128
rect 6648 112 6664 128
rect 4184 92 4200 108
rect 4696 92 4712 108
rect 5960 92 5976 108
rect 3128 52 3144 68
rect 4824 32 4840 48
rect 5624 32 5640 48
rect 798 2 826 18
rect 2862 2 2890 18
rect 4910 2 4938 18
rect 5912 12 5928 28
<< metal4 >>
rect 826 4806 832 4814
rect 2890 4806 2896 4814
rect 924 4703 932 4704
rect 924 4697 936 4703
rect 924 4696 932 4697
rect 173 4308 179 4692
rect 1069 4528 1075 4612
rect 1277 4544 1283 4552
rect 1276 4536 1284 4544
rect 77 3124 83 3712
rect 76 3116 84 3124
rect 77 3068 83 3116
rect 173 1328 179 4292
rect 189 2248 195 4252
rect 461 4148 467 4452
rect 826 4406 832 4414
rect 844 4363 852 4364
rect 844 4357 856 4363
rect 844 4356 852 4357
rect 669 4308 675 4332
rect 205 3488 211 3632
rect 221 2968 227 4012
rect 173 708 179 1312
rect 189 928 195 2232
rect 205 2148 211 2772
rect 237 2128 243 3732
rect 285 3388 291 3412
rect 333 3328 339 3472
rect 365 3368 371 3812
rect 349 3324 355 3352
rect 348 3316 356 3324
rect 269 2844 275 2892
rect 268 2836 276 2844
rect 205 1468 211 1872
rect 253 1748 259 2212
rect 269 1328 275 2836
rect 301 2408 307 2952
rect 333 2948 339 3312
rect 397 3008 403 3332
rect 413 3088 419 3732
rect 429 3108 435 3652
rect 445 3328 451 3412
rect 333 2688 339 2932
rect 429 2588 435 3092
rect 284 2036 292 2044
rect 285 2028 291 2036
rect 301 1944 307 2132
rect 300 1936 308 1944
rect 333 1884 339 1892
rect 332 1876 340 1884
rect 317 948 323 1452
rect 365 1368 371 2172
rect 381 928 387 1892
rect 397 1708 403 1972
rect 413 1908 419 2392
rect 429 1988 435 2572
rect 429 1608 435 1972
rect 445 1888 451 2572
rect 461 2248 467 4132
rect 477 2308 483 2652
rect 525 2468 531 3972
rect 493 2284 499 2412
rect 492 2276 500 2284
rect 429 1168 435 1552
rect 493 1508 499 2276
rect 541 2148 547 3472
rect 573 3248 579 3612
rect 589 3488 595 4112
rect 684 4076 692 4084
rect 685 3988 691 4076
rect 826 4006 832 4014
rect 861 3884 867 4212
rect 860 3883 868 3884
rect 860 3877 872 3883
rect 860 3876 868 3877
rect 605 3408 611 3472
rect 621 3408 627 3632
rect 588 3356 596 3364
rect 589 3348 595 3356
rect 669 3348 675 3432
rect 605 3324 611 3332
rect 604 3316 612 3324
rect 509 1748 515 2072
rect 541 1548 547 2132
rect 476 1043 484 1044
rect 476 1037 488 1043
rect 476 1036 484 1037
rect 173 548 179 692
rect 285 344 291 352
rect 284 336 292 344
rect 365 288 371 912
rect 381 308 387 912
rect 493 568 499 932
rect 556 876 564 884
rect 557 488 563 876
rect 573 688 579 2232
rect 621 2088 627 3332
rect 637 1848 643 2412
rect 653 2148 659 2932
rect 701 2508 707 2712
rect 653 1948 659 2132
rect 653 1788 659 1932
rect 669 1888 675 2352
rect 685 2308 691 2492
rect 684 2196 692 2204
rect 685 1888 691 2196
rect 605 1388 611 1632
rect 429 344 435 352
rect 428 336 436 344
rect 573 268 579 672
rect 589 148 595 992
rect 685 688 691 1872
rect 701 1428 707 2212
rect 717 2208 723 3872
rect 845 3628 851 3852
rect 893 3748 899 4352
rect 1005 4324 1011 4332
rect 1004 4316 1012 4324
rect 826 3606 832 3614
rect 826 3206 832 3214
rect 845 3028 851 3612
rect 826 2806 832 2814
rect 845 2668 851 3012
rect 781 1728 787 2512
rect 826 2406 832 2414
rect 845 2148 851 2652
rect 861 2528 867 3492
rect 893 3348 899 3732
rect 893 3088 899 3332
rect 909 3008 915 3992
rect 925 3528 931 4012
rect 941 3828 947 4052
rect 957 4048 963 4292
rect 1005 3984 1011 4212
rect 1004 3976 1012 3984
rect 941 3488 947 3812
rect 973 3648 979 3972
rect 1005 3908 1011 3976
rect 989 3728 995 3832
rect 1005 3348 1011 3852
rect 909 2248 915 2992
rect 1005 2768 1011 3332
rect 1021 3268 1027 3652
rect 1037 2868 1043 4372
rect 1053 3044 1059 4512
rect 1069 4044 1075 4232
rect 1068 4036 1076 4044
rect 1085 3988 1091 4152
rect 1069 3164 1075 3312
rect 1068 3156 1076 3164
rect 1084 3136 1092 3144
rect 1085 3108 1091 3136
rect 1052 3036 1060 3044
rect 1068 2916 1076 2924
rect 1069 2908 1075 2916
rect 826 2006 832 2014
rect 748 1483 756 1484
rect 748 1477 760 1483
rect 748 1476 756 1477
rect 781 908 787 1712
rect 826 1606 832 1614
rect 826 1206 832 1214
rect 826 806 832 814
rect 685 648 691 672
rect 845 428 851 1912
rect 861 904 867 2172
rect 925 1848 931 2712
rect 940 2523 948 2524
rect 940 2517 952 2523
rect 940 2516 948 2517
rect 941 2308 947 2516
rect 1053 2304 1059 2432
rect 1052 2296 1060 2304
rect 973 1808 979 2172
rect 973 1748 979 1792
rect 1037 1748 1043 2232
rect 1053 1868 1059 2296
rect 957 1724 963 1732
rect 956 1716 964 1724
rect 893 1688 899 1712
rect 1004 1703 1012 1704
rect 1004 1697 1016 1703
rect 1004 1696 1012 1697
rect 893 1348 899 1672
rect 909 1408 915 1592
rect 925 1048 931 1332
rect 860 896 868 904
rect 989 828 995 1312
rect 1037 1088 1043 1732
rect 1069 1608 1075 2692
rect 1085 2688 1091 2732
rect 1101 2688 1107 4532
rect 1117 4268 1123 4492
rect 1117 3828 1123 4252
rect 1117 3108 1123 3412
rect 1133 2708 1139 4512
rect 1181 4204 1187 4272
rect 1197 4268 1203 4332
rect 1180 4196 1188 4204
rect 1213 4148 1219 4332
rect 1229 4168 1235 4412
rect 1245 4268 1251 4312
rect 1149 4104 1155 4132
rect 1196 4116 1204 4124
rect 1197 4108 1203 4116
rect 1148 4096 1156 4104
rect 1261 4048 1267 4412
rect 1277 4288 1283 4312
rect 1309 3948 1315 4652
rect 1485 4324 1491 4372
rect 1501 4328 1507 4652
rect 1532 4503 1540 4504
rect 1532 4497 1544 4503
rect 1532 4496 1540 4497
rect 1565 4408 1571 4492
rect 1484 4316 1492 4324
rect 1453 4204 1459 4212
rect 1452 4196 1460 4204
rect 1324 4156 1332 4164
rect 1325 4148 1331 4156
rect 1357 4104 1363 4132
rect 1405 4124 1411 4132
rect 1404 4116 1412 4124
rect 1548 4116 1556 4124
rect 1356 4096 1364 4104
rect 1165 2964 1171 3892
rect 1181 3048 1187 3312
rect 1228 3143 1236 3144
rect 1224 3137 1236 3143
rect 1228 3136 1236 3137
rect 1164 2956 1172 2964
rect 1165 2908 1171 2956
rect 1197 2704 1203 3052
rect 1196 2696 1204 2704
rect 1149 2528 1155 2532
rect 1149 2188 1155 2512
rect 1085 1348 1091 2072
rect 1149 1728 1155 1992
rect 1117 1688 1123 1712
rect 1149 1704 1155 1712
rect 1148 1696 1156 1704
rect 1117 1408 1123 1672
rect 1165 1488 1171 2672
rect 1229 2068 1235 2692
rect 1245 2568 1251 3512
rect 1277 2904 1283 2912
rect 1276 2896 1284 2904
rect 1261 2688 1267 2752
rect 1261 2288 1267 2672
rect 1277 2148 1283 2896
rect 1244 2123 1252 2124
rect 1244 2117 1256 2123
rect 1244 2116 1252 2117
rect 1293 1928 1299 3092
rect 1325 3088 1331 4072
rect 1468 3976 1476 3984
rect 1452 3876 1460 3884
rect 1388 3863 1396 3864
rect 1388 3857 1400 3863
rect 1388 3856 1396 3857
rect 1325 2928 1331 3072
rect 1389 2928 1395 3856
rect 1053 1068 1059 1112
rect 1069 908 1075 1112
rect 1084 1096 1092 1104
rect 1085 988 1091 1096
rect 1085 908 1091 972
rect 1117 608 1123 932
rect 1197 728 1203 1892
rect 1308 1783 1316 1784
rect 1308 1777 1320 1783
rect 1308 1776 1316 1777
rect 1213 1144 1219 1352
rect 1212 1136 1220 1144
rect 1213 904 1219 912
rect 1212 896 1220 904
rect 1133 524 1139 552
rect 1132 516 1140 524
rect 716 336 724 344
rect 717 328 723 336
rect 700 323 708 324
rect 696 317 708 323
rect 700 316 708 317
rect 765 324 771 412
rect 826 406 832 414
rect 845 328 851 412
rect 1149 344 1155 712
rect 1197 528 1203 712
rect 1229 708 1235 1072
rect 1245 1044 1251 1052
rect 1293 1048 1299 1732
rect 1309 1548 1315 1752
rect 1309 1428 1315 1532
rect 1244 1036 1252 1044
rect 1341 944 1347 2492
rect 1357 2308 1363 2432
rect 1308 936 1316 944
rect 1340 936 1348 944
rect 1261 528 1267 852
rect 1293 708 1299 932
rect 1309 928 1315 936
rect 1357 708 1363 1632
rect 1373 928 1379 2912
rect 1389 1708 1395 2492
rect 1405 2268 1411 2892
rect 1421 2368 1427 3032
rect 1437 2668 1443 3252
rect 1453 2688 1459 3876
rect 1469 2748 1475 3976
rect 1485 3248 1491 3852
rect 1437 2328 1443 2612
rect 1453 2204 1459 2672
rect 1501 2548 1507 4092
rect 1549 4008 1555 4116
rect 1565 4048 1571 4392
rect 1661 4268 1667 4672
rect 1677 4368 1683 4532
rect 1548 3923 1556 3924
rect 1548 3917 1560 3923
rect 1548 3916 1556 3917
rect 1517 3388 1523 3632
rect 1533 2788 1539 3412
rect 1565 2948 1571 3872
rect 1597 3868 1603 4192
rect 1452 2196 1460 2204
rect 1389 748 1395 1052
rect 1180 523 1188 524
rect 1176 517 1188 523
rect 1180 516 1188 517
rect 1148 336 1156 344
rect 748 323 756 324
rect 744 317 756 323
rect 748 316 756 317
rect 764 316 772 324
rect 860 323 868 324
rect 860 317 872 323
rect 860 316 868 317
rect 908 163 916 164
rect 908 157 920 163
rect 908 156 916 157
rect 1149 148 1155 336
rect 1164 323 1172 324
rect 1164 317 1176 323
rect 1164 316 1172 317
rect 1261 324 1267 512
rect 1389 488 1395 732
rect 1405 588 1411 2012
rect 1437 1808 1443 2152
rect 1453 1868 1459 2172
rect 1453 1508 1459 1852
rect 1469 988 1475 2312
rect 1485 1448 1491 2212
rect 1501 1908 1507 2412
rect 1516 1936 1524 1944
rect 1517 1748 1523 1936
rect 1501 1724 1507 1732
rect 1500 1716 1508 1724
rect 1533 1528 1539 2572
rect 1549 2408 1555 2672
rect 1581 2644 1587 3032
rect 1613 2864 1619 4112
rect 1677 4048 1683 4352
rect 1693 4084 1699 4132
rect 1692 4076 1700 4084
rect 1693 3848 1699 3932
rect 1709 3928 1715 4572
rect 1661 3324 1667 3732
rect 1660 3316 1668 3324
rect 1677 3144 1683 3232
rect 1676 3143 1684 3144
rect 1676 3137 1688 3143
rect 1676 3136 1684 3137
rect 1645 2884 1651 3052
rect 1709 3048 1715 3612
rect 1661 2908 1667 3032
rect 1725 2968 1731 4312
rect 1741 3748 1747 4172
rect 1757 2988 1763 4612
rect 1866 4606 1872 4614
rect 1852 4543 1860 4544
rect 1848 4537 1860 4543
rect 1852 4536 1860 4537
rect 1866 4206 1872 4214
rect 1773 3668 1779 3792
rect 1789 3744 1795 3752
rect 1805 3748 1811 4152
rect 1852 4043 1860 4044
rect 1848 4037 1860 4043
rect 1852 4036 1860 4037
rect 1788 3736 1796 3744
rect 1821 3304 1827 3872
rect 1866 3806 1872 3814
rect 1916 3496 1924 3504
rect 1917 3488 1923 3496
rect 1933 3484 1939 4032
rect 1949 3788 1955 4532
rect 1965 3568 1971 4292
rect 1997 3748 2003 4312
rect 2028 3743 2036 3744
rect 2024 3737 2036 3743
rect 2028 3736 2036 3737
rect 1932 3476 1940 3484
rect 1866 3406 1872 3414
rect 1933 3408 1939 3476
rect 1820 3296 1828 3304
rect 1821 3028 1827 3132
rect 1901 3084 1907 3392
rect 1997 3308 2003 3712
rect 2077 3364 2083 3392
rect 2076 3356 2084 3364
rect 1900 3076 1908 3084
rect 1788 2976 1796 2984
rect 1789 2968 1795 2976
rect 1644 2876 1652 2884
rect 1805 2868 1811 3012
rect 1866 3006 1872 3014
rect 1612 2856 1620 2864
rect 1613 2688 1619 2856
rect 1821 2848 1827 2992
rect 1580 2636 1588 2644
rect 1565 2208 1571 2512
rect 1597 2208 1603 2592
rect 1629 2544 1635 2592
rect 1628 2536 1636 2544
rect 1709 2444 1715 2832
rect 1901 2708 1907 3076
rect 1725 2548 1731 2672
rect 1708 2436 1716 2444
rect 1628 2283 1636 2284
rect 1624 2277 1636 2283
rect 1628 2276 1636 2277
rect 1565 1888 1571 2192
rect 1533 1468 1539 1512
rect 1549 1368 1555 1432
rect 1516 716 1524 724
rect 1517 708 1523 716
rect 1501 528 1507 672
rect 1565 628 1571 1872
rect 1581 1328 1587 1792
rect 1260 316 1268 324
rect 1597 288 1603 1952
rect 1629 1788 1635 2276
rect 1645 1768 1651 2112
rect 1613 1168 1619 1612
rect 1677 1348 1683 2092
rect 1693 1688 1699 2432
rect 1660 1343 1668 1344
rect 1656 1337 1668 1343
rect 1660 1336 1668 1337
rect 1613 828 1619 1152
rect 1709 1068 1715 2392
rect 1725 1748 1731 2072
rect 1725 1448 1731 1732
rect 1741 1484 1747 2272
rect 1757 1728 1763 2132
rect 1789 2108 1795 2612
rect 1866 2606 1872 2614
rect 1772 1916 1780 1924
rect 1773 1908 1779 1916
rect 1788 1723 1796 1724
rect 1784 1717 1796 1723
rect 1788 1716 1796 1717
rect 1740 1476 1748 1484
rect 1741 1368 1747 1476
rect 1788 1263 1796 1264
rect 1788 1257 1800 1263
rect 1788 1256 1796 1257
rect 1756 956 1764 964
rect 1757 948 1763 956
rect 1020 136 1028 144
rect 1021 128 1027 136
rect 1165 124 1171 152
rect 1277 148 1283 272
rect 1693 148 1699 252
rect 1789 228 1795 1212
rect 1805 568 1811 1092
rect 1821 1048 1827 2532
rect 1917 2464 1923 3032
rect 1981 2904 1987 3172
rect 1980 2896 1988 2904
rect 1964 2703 1972 2704
rect 1960 2697 1972 2703
rect 1964 2696 1972 2697
rect 1997 2668 2003 3292
rect 2028 2936 2036 2944
rect 2029 2928 2035 2936
rect 2028 2876 2036 2884
rect 2029 2668 2035 2876
rect 2045 2768 2051 3332
rect 2060 3256 2068 3264
rect 2045 2748 2051 2752
rect 1964 2636 1972 2644
rect 1965 2488 1971 2636
rect 1916 2456 1924 2464
rect 1884 2436 1892 2444
rect 1866 2206 1872 2214
rect 1885 1908 1891 2436
rect 1866 1806 1872 1814
rect 1885 1784 1891 1792
rect 1884 1776 1892 1784
rect 1901 1708 1907 1872
rect 1866 1406 1872 1414
rect 1821 1008 1827 1032
rect 1866 1006 1872 1014
rect 1901 888 1907 1692
rect 1866 606 1872 614
rect 1917 588 1923 1312
rect 1933 1308 1939 2232
rect 1965 1924 1971 2472
rect 1964 1916 1972 1924
rect 1981 1144 1987 2652
rect 1997 2564 2003 2652
rect 2061 2648 2067 3256
rect 2077 2748 2083 3312
rect 2108 3116 2116 3124
rect 2109 3108 2115 3116
rect 2093 2904 2099 2952
rect 2092 2896 2100 2904
rect 2109 2864 2115 2912
rect 2108 2856 2116 2864
rect 2093 2608 2099 2812
rect 1996 2556 2004 2564
rect 1997 2248 2003 2512
rect 2012 2103 2020 2104
rect 2012 2097 2024 2103
rect 2012 2096 2020 2097
rect 2045 1248 2051 2232
rect 2077 2188 2083 2332
rect 2076 2036 2084 2044
rect 2077 1968 2083 2036
rect 2061 1288 2067 1952
rect 2076 1936 2084 1944
rect 2077 1908 2083 1936
rect 2093 1748 2099 2172
rect 2109 1584 2115 2712
rect 2125 2708 2131 3872
rect 2141 2844 2147 3112
rect 2157 2848 2163 3192
rect 2140 2836 2148 2844
rect 2141 2728 2147 2836
rect 2173 2523 2179 3692
rect 2189 3088 2195 3872
rect 2205 3308 2211 3372
rect 2221 3228 2227 4692
rect 2237 3748 2243 4332
rect 2253 3888 2259 4372
rect 2285 4304 2291 4532
rect 2396 4376 2404 4384
rect 2284 4296 2292 4304
rect 2285 4168 2291 4296
rect 2316 4263 2324 4264
rect 2316 4257 2328 4263
rect 2316 4256 2324 4257
rect 2237 3588 2243 3732
rect 2237 3564 2243 3572
rect 2236 3556 2244 3564
rect 2348 3516 2356 3524
rect 2237 3208 2243 3512
rect 2349 3508 2355 3516
rect 2188 2936 2196 2944
rect 2189 2908 2195 2936
rect 2173 2517 2195 2523
rect 2108 1576 2116 1584
rect 2125 1408 2131 2292
rect 1980 1136 1988 1144
rect 1948 1103 1956 1104
rect 1944 1097 1956 1103
rect 1948 1096 1956 1097
rect 1980 1056 1988 1064
rect 1981 1048 1987 1056
rect 1965 968 1971 1012
rect 2013 688 2019 772
rect 1964 683 1972 684
rect 1964 677 1976 683
rect 1964 676 1972 677
rect 2093 668 2099 1172
rect 2109 928 2115 1352
rect 2141 1328 2147 2272
rect 2157 2124 2163 2472
rect 2156 2116 2164 2124
rect 2157 1168 2163 2116
rect 2173 1528 2179 1872
rect 2189 1748 2195 2517
rect 2205 2068 2211 2992
rect 2221 2528 2227 2952
rect 2253 2748 2259 3372
rect 2237 2524 2243 2632
rect 2269 2584 2275 2592
rect 2268 2576 2276 2584
rect 2236 2516 2244 2524
rect 2220 2176 2228 2184
rect 2221 2088 2227 2176
rect 2173 1368 2179 1512
rect 2205 1488 2211 1652
rect 2205 984 2211 1472
rect 2237 1264 2243 2516
rect 2253 2148 2259 2392
rect 2285 2148 2291 2932
rect 2317 2184 2323 3452
rect 2332 3363 2340 3364
rect 2332 3357 2344 3363
rect 2332 3356 2340 3357
rect 2365 3264 2371 3732
rect 2381 3644 2387 4252
rect 2397 4164 2403 4376
rect 2396 4156 2404 4164
rect 2397 4128 2403 4156
rect 2460 4123 2468 4124
rect 2456 4117 2468 4123
rect 2460 4116 2468 4117
rect 2380 3636 2388 3644
rect 2364 3256 2372 3264
rect 2381 3068 2387 3492
rect 2397 3068 2403 4112
rect 2429 4084 2435 4092
rect 2428 4076 2436 4084
rect 2460 4076 2468 4084
rect 2429 3548 2435 3592
rect 2461 3068 2467 4076
rect 2477 3928 2483 4672
rect 2557 4524 2563 4532
rect 2556 4516 2564 4524
rect 2541 4504 2547 4512
rect 2540 4496 2548 4504
rect 2573 4388 2579 4692
rect 2636 4523 2644 4524
rect 2632 4517 2644 4523
rect 2636 4516 2644 4517
rect 2589 4504 2595 4512
rect 2588 4496 2596 4504
rect 2620 4423 2628 4424
rect 2620 4417 2632 4423
rect 2620 4416 2628 4417
rect 2685 4348 2691 4612
rect 2989 4548 2995 4552
rect 2764 4523 2772 4524
rect 2760 4517 2772 4523
rect 2764 4516 2772 4517
rect 2748 4343 2756 4344
rect 2744 4337 2756 4343
rect 2748 4336 2756 4337
rect 2477 3744 2483 3752
rect 2476 3736 2484 3744
rect 2492 3456 2500 3464
rect 2316 2176 2324 2184
rect 2333 2008 2339 2652
rect 2349 2484 2355 2532
rect 2365 2488 2371 3052
rect 2396 3036 2404 3044
rect 2397 2968 2403 3036
rect 2348 2476 2356 2484
rect 2397 2028 2403 2592
rect 2461 2548 2467 3052
rect 2413 2328 2419 2412
rect 2300 1903 2308 1904
rect 2300 1897 2312 1903
rect 2300 1896 2308 1897
rect 2333 1848 2339 1892
rect 2268 1576 2276 1584
rect 2269 1328 2275 1576
rect 2236 1256 2244 1264
rect 2204 976 2212 984
rect 2125 884 2131 912
rect 2157 904 2163 912
rect 2156 896 2164 904
rect 2124 876 2132 884
rect 2205 848 2211 976
rect 2157 664 2163 812
rect 2221 728 2227 1012
rect 2285 948 2291 1712
rect 2333 1488 2339 1832
rect 2397 1568 2403 1912
rect 2317 988 2323 1012
rect 2333 808 2339 1412
rect 2365 1328 2371 1532
rect 2413 1508 2419 2312
rect 2445 1788 2451 2492
rect 2461 1908 2467 2412
rect 2477 2048 2483 3292
rect 2364 1136 2372 1144
rect 2365 1128 2371 1136
rect 2428 1076 2436 1084
rect 2429 1068 2435 1076
rect 2156 656 2164 664
rect 1917 468 1923 572
rect 1866 206 1872 214
rect 1324 136 1332 144
rect 1164 116 1172 124
rect 1277 108 1283 132
rect 1325 128 1331 136
rect 2189 124 2195 192
rect 2188 116 2196 124
rect 2221 108 2227 712
rect 2284 616 2292 624
rect 2285 588 2291 616
rect 2317 344 2323 732
rect 2333 588 2339 792
rect 2349 528 2355 872
rect 2348 463 2356 464
rect 2348 457 2360 463
rect 2348 456 2356 457
rect 2316 336 2324 344
rect 2317 308 2323 336
rect 2364 323 2372 324
rect 2364 317 2376 323
rect 2364 316 2372 317
rect 2332 263 2340 264
rect 2332 257 2344 263
rect 2332 256 2340 257
rect 2397 148 2403 392
rect 2348 136 2356 144
rect 2349 128 2355 136
rect 2413 128 2419 1012
rect 2445 944 2451 1452
rect 2444 936 2452 944
rect 2429 568 2435 672
rect 2429 268 2435 552
rect 2461 148 2467 692
rect 2493 448 2499 3456
rect 2573 3388 2579 3532
rect 2589 3348 2595 4072
rect 2749 3928 2755 4312
rect 2765 4148 2771 4516
rect 2781 4508 2787 4532
rect 2797 4424 2803 4532
rect 2829 4428 2835 4532
rect 2796 4416 2804 4424
rect 2890 4406 2896 4414
rect 2989 4384 2995 4532
rect 2988 4376 2996 4384
rect 2781 3868 2787 4192
rect 2812 4096 2820 4104
rect 2813 3948 2819 4096
rect 2620 3743 2628 3744
rect 2616 3737 2628 3743
rect 2620 3736 2628 3737
rect 2796 3736 2804 3744
rect 2797 3728 2803 3736
rect 2748 3636 2756 3644
rect 2749 3628 2755 3636
rect 2620 3556 2628 3564
rect 2621 3388 2627 3556
rect 2524 3063 2532 3064
rect 2520 3057 2532 3063
rect 2524 3056 2532 3057
rect 2508 2536 2516 2544
rect 2509 2528 2515 2536
rect 2524 2456 2532 2464
rect 2509 1888 2515 2132
rect 2525 2128 2531 2456
rect 2541 2148 2547 2912
rect 2573 2848 2579 3152
rect 2653 3104 2659 3412
rect 2669 3288 2675 3592
rect 2813 3528 2819 3932
rect 2829 3748 2835 4272
rect 2845 3888 2851 4112
rect 2877 4044 2883 4352
rect 2892 4136 2900 4144
rect 2893 4128 2899 4136
rect 2909 4088 2915 4112
rect 2876 4036 2884 4044
rect 2890 4006 2896 4014
rect 2925 4008 2931 4232
rect 2925 3984 2931 3992
rect 2924 3976 2932 3984
rect 3053 3908 3059 4352
rect 2940 3903 2948 3904
rect 2940 3897 2952 3903
rect 2940 3896 2948 3897
rect 2890 3606 2896 3614
rect 2828 3556 2836 3564
rect 2813 3384 2819 3512
rect 2829 3508 2835 3556
rect 2829 3484 2835 3492
rect 2828 3476 2836 3484
rect 2812 3376 2820 3384
rect 2652 3096 2660 3104
rect 2589 2984 2595 3052
rect 2588 2976 2596 2984
rect 2573 2724 2579 2732
rect 2572 2716 2580 2724
rect 2605 2584 2611 2612
rect 2604 2576 2612 2584
rect 2572 2283 2580 2284
rect 2572 2277 2584 2283
rect 2572 2276 2580 2277
rect 2525 2084 2531 2112
rect 2524 2076 2532 2084
rect 2509 1464 2515 1872
rect 2524 1543 2532 1544
rect 2524 1537 2536 1543
rect 2524 1536 2532 1537
rect 2508 1456 2516 1464
rect 2557 664 2563 1552
rect 2605 784 2611 2252
rect 2621 1664 2627 3072
rect 2636 2936 2644 2944
rect 2637 2468 2643 2936
rect 2653 2368 2659 3096
rect 2717 3084 2723 3252
rect 2716 3083 2724 3084
rect 2712 3077 2724 3083
rect 2716 3076 2724 3077
rect 2620 1656 2628 1664
rect 2621 1528 2627 1656
rect 2637 1524 2643 2232
rect 2685 1888 2691 2592
rect 2765 2588 2771 2652
rect 2765 2524 2771 2572
rect 2780 2556 2788 2564
rect 2781 2548 2787 2556
rect 2764 2516 2772 2524
rect 2733 2148 2739 2332
rect 2797 2288 2803 2692
rect 2829 2188 2835 2532
rect 2845 2428 2851 3312
rect 2890 3206 2896 3214
rect 2909 3048 2915 3392
rect 2925 3208 2931 3892
rect 2989 3684 2995 3832
rect 2988 3676 2996 3684
rect 3069 3628 3075 4692
rect 3180 4516 3188 4524
rect 3084 4276 3092 4284
rect 3085 4268 3091 4276
rect 3165 4084 3171 4432
rect 3181 4128 3187 4516
rect 3197 4344 3203 4492
rect 3196 4336 3204 4344
rect 3292 4296 3300 4304
rect 3293 4288 3299 4296
rect 3197 4164 3203 4212
rect 3325 4188 3331 4472
rect 3341 4168 3347 4412
rect 3373 4184 3379 4192
rect 3372 4176 3380 4184
rect 3196 4156 3204 4164
rect 3164 4076 3172 4084
rect 3181 3908 3187 4092
rect 3084 3716 3092 3724
rect 3085 3708 3091 3716
rect 2957 3484 2963 3492
rect 2956 3476 2964 3484
rect 2957 3368 2963 3476
rect 2890 2806 2896 2814
rect 2941 2588 2947 3212
rect 2957 2588 2963 2732
rect 2893 2544 2899 2552
rect 2973 2548 2979 3332
rect 2988 2716 2996 2724
rect 2989 2688 2995 2716
rect 3037 2548 3043 3092
rect 3085 2708 3091 2892
rect 2892 2536 2900 2544
rect 2890 2406 2896 2414
rect 2909 2284 2915 2392
rect 2908 2276 2916 2284
rect 2861 2184 2867 2252
rect 2860 2176 2868 2184
rect 2796 2156 2804 2164
rect 2797 2148 2803 2156
rect 2700 1916 2708 1924
rect 2701 1908 2707 1916
rect 2733 1788 2739 2132
rect 2636 1516 2644 1524
rect 2637 1328 2643 1516
rect 2669 1488 2675 1672
rect 2829 1528 2835 2172
rect 2972 2116 2980 2124
rect 2973 2108 2979 2116
rect 2890 2006 2896 2014
rect 2813 1504 2819 1512
rect 2812 1496 2820 1504
rect 2684 1483 2692 1484
rect 2684 1477 2696 1483
rect 2684 1476 2692 1477
rect 2685 1168 2691 1476
rect 2749 1168 2755 1432
rect 2829 1328 2835 1512
rect 2812 1323 2820 1324
rect 2808 1317 2820 1323
rect 2812 1316 2820 1317
rect 2829 944 2835 1292
rect 2828 936 2836 944
rect 2604 776 2612 784
rect 2605 728 2611 776
rect 2556 656 2564 664
rect 2604 516 2612 524
rect 2605 508 2611 516
rect 2701 508 2707 612
rect 2812 496 2820 504
rect 2813 428 2819 496
rect 2509 324 2515 332
rect 2508 316 2516 324
rect 2717 264 2723 272
rect 2829 268 2835 936
rect 2845 808 2851 1752
rect 2973 1728 2979 1932
rect 2890 1606 2896 1614
rect 2890 1206 2896 1214
rect 2925 964 2931 1472
rect 2924 956 2932 964
rect 2925 948 2931 956
rect 2908 896 2916 904
rect 2890 806 2896 814
rect 2845 324 2851 792
rect 2909 708 2915 896
rect 2941 708 2947 1632
rect 3005 1608 3011 2512
rect 3021 1808 3027 2332
rect 3053 1928 3059 2512
rect 3068 2476 3076 2484
rect 3069 2028 3075 2476
rect 3069 1904 3075 1912
rect 3068 1896 3076 1904
rect 3085 1848 3091 2252
rect 2957 1084 2963 1092
rect 2956 1076 2964 1084
rect 2957 804 2963 1076
rect 2988 1063 2996 1064
rect 2988 1057 3000 1063
rect 2988 1056 2996 1057
rect 3037 968 3043 1312
rect 3053 1108 3059 1772
rect 3085 1508 3091 1832
rect 3101 1488 3107 2292
rect 3117 1228 3123 3512
rect 3132 3463 3140 3464
rect 3132 3457 3144 3463
rect 3132 3456 3140 3457
rect 3132 3356 3140 3364
rect 3133 3288 3139 3356
rect 3165 3348 3171 3352
rect 3181 3348 3187 3892
rect 3197 3884 3203 4156
rect 3196 3876 3204 3884
rect 3229 3828 3235 4072
rect 3229 3768 3235 3812
rect 3149 3068 3155 3072
rect 3149 2608 3155 3052
rect 3149 2328 3155 2592
rect 3165 1888 3171 3332
rect 3197 3308 3203 3552
rect 3437 3528 3443 4552
rect 3485 4308 3491 4672
rect 3469 4044 3475 4172
rect 3468 4036 3476 4044
rect 3469 3808 3475 4036
rect 3485 3888 3491 4292
rect 3501 4048 3507 4812
rect 4938 4806 4944 4814
rect 3741 4708 3747 4772
rect 3564 4556 3572 4564
rect 3565 4548 3571 4556
rect 3709 4524 3715 4552
rect 3708 4516 3716 4524
rect 3468 3763 3476 3764
rect 3464 3757 3476 3763
rect 3468 3756 3476 3757
rect 3485 3584 3491 3872
rect 3484 3576 3492 3584
rect 3356 3296 3364 3304
rect 3197 3128 3203 3152
rect 3181 3064 3187 3072
rect 3180 3056 3188 3064
rect 3181 2308 3187 2912
rect 3148 1636 3156 1644
rect 3149 1588 3155 1636
rect 3197 1428 3203 2892
rect 3277 2828 3283 3172
rect 3357 3068 3363 3296
rect 3372 3116 3380 3124
rect 3373 3108 3379 3116
rect 3213 2388 3219 2772
rect 3229 2228 3235 2372
rect 3245 2364 3251 2632
rect 3244 2356 3252 2364
rect 3325 2328 3331 2752
rect 3357 2684 3363 2692
rect 3373 2688 3379 3032
rect 3389 2988 3395 3112
rect 3404 2956 3412 2964
rect 3405 2948 3411 2956
rect 3356 2676 3364 2684
rect 3357 2448 3363 2676
rect 3325 2188 3331 2312
rect 3213 2144 3219 2172
rect 3212 2136 3220 2144
rect 3229 1708 3235 1752
rect 3213 1448 3219 1472
rect 3053 1084 3059 1092
rect 3052 1076 3060 1084
rect 3165 1008 3171 1072
rect 3180 976 3188 984
rect 3181 968 3187 976
rect 2956 796 2964 804
rect 2989 768 2995 812
rect 3101 784 3107 892
rect 3100 776 3108 784
rect 2941 584 2947 692
rect 3197 648 3203 752
rect 3213 688 3219 1432
rect 3245 1144 3251 1852
rect 3357 1728 3363 2292
rect 3421 2268 3427 2292
rect 3469 2288 3475 3492
rect 3517 3484 3523 3852
rect 3516 3476 3524 3484
rect 3244 1136 3252 1144
rect 3261 928 3267 1092
rect 3212 656 3220 664
rect 3213 648 3219 656
rect 2940 576 2948 584
rect 2909 428 2915 472
rect 2890 406 2896 414
rect 2972 356 2980 364
rect 2973 348 2979 356
rect 2844 316 2852 324
rect 2716 256 2724 264
rect 2957 264 2963 312
rect 2956 256 2964 264
rect 2700 156 2708 164
rect 2701 148 2707 156
rect 2428 143 2436 144
rect 2428 137 2440 143
rect 2428 136 2436 137
rect 2508 143 2516 144
rect 2504 137 2516 143
rect 2508 136 2516 137
rect 3133 68 3139 172
rect 3181 168 3187 552
rect 3244 296 3252 304
rect 3245 288 3251 296
rect 3261 288 3267 912
rect 3277 288 3283 1012
rect 3325 524 3331 1232
rect 3357 1108 3363 1712
rect 3389 1648 3395 1772
rect 3405 1668 3411 1992
rect 3421 1724 3427 1732
rect 3420 1716 3428 1724
rect 3437 868 3443 1332
rect 3485 988 3491 2652
rect 3501 2188 3507 3252
rect 3517 2448 3523 3476
rect 3565 3468 3571 4512
rect 3725 4328 3731 4632
rect 3708 3856 3716 3864
rect 3709 3688 3715 3856
rect 3724 3736 3732 3744
rect 3725 3688 3731 3736
rect 3645 3604 3651 3672
rect 3692 3656 3700 3664
rect 3644 3596 3652 3604
rect 3532 3376 3540 3384
rect 3533 3288 3539 3376
rect 3533 3044 3539 3192
rect 3532 3036 3540 3044
rect 3533 2728 3539 3036
rect 3549 2548 3555 3072
rect 3501 1828 3507 2172
rect 3517 2128 3523 2252
rect 3549 2228 3555 2532
rect 3565 2528 3571 3452
rect 3596 3136 3604 3144
rect 3597 3124 3603 3136
rect 3596 3123 3604 3124
rect 3596 3117 3608 3123
rect 3596 3116 3604 3117
rect 3693 3088 3699 3656
rect 3709 3544 3715 3672
rect 3708 3536 3716 3544
rect 3709 3468 3715 3536
rect 3580 2276 3588 2284
rect 3549 2164 3555 2212
rect 3581 2188 3587 2276
rect 3548 2156 3556 2164
rect 3612 2156 3620 2164
rect 3613 2128 3619 2156
rect 3564 2123 3572 2124
rect 3564 2117 3576 2123
rect 3564 2116 3572 2117
rect 3517 1508 3523 1892
rect 3549 1628 3555 2112
rect 3661 1508 3667 2372
rect 3677 1488 3683 2652
rect 3693 1508 3699 3072
rect 3709 2688 3715 3332
rect 3741 3208 3747 4692
rect 3914 4606 3920 4614
rect 4252 4556 4260 4564
rect 4253 4548 4259 4556
rect 4124 4516 4132 4524
rect 3772 4436 3780 4444
rect 3773 4208 3779 4436
rect 3821 4028 3827 4272
rect 3869 4168 3875 4512
rect 3914 4206 3920 4214
rect 3789 3928 3795 4012
rect 3933 3968 3939 4232
rect 3853 3864 3859 3892
rect 3852 3856 3860 3864
rect 3869 3788 3875 3892
rect 3914 3806 3920 3814
rect 3933 3768 3939 3792
rect 3756 3096 3764 3104
rect 3757 3068 3763 3096
rect 3709 2308 3715 2672
rect 3709 1728 3715 1892
rect 3741 1468 3747 3052
rect 3757 1644 3763 2892
rect 3773 2828 3779 3612
rect 3805 3388 3811 3672
rect 3980 3576 3988 3584
rect 3981 3528 3987 3576
rect 3805 2708 3811 3372
rect 3772 2563 3780 2564
rect 3772 2557 3784 2563
rect 3772 2556 3780 2557
rect 3821 2188 3827 3392
rect 3837 3268 3843 3472
rect 3853 3408 3859 3492
rect 3964 3456 3972 3464
rect 3914 3406 3920 3414
rect 3837 2608 3843 3252
rect 3933 3128 3939 3392
rect 3948 3336 3956 3344
rect 3949 3328 3955 3336
rect 3837 2548 3843 2592
rect 3853 2328 3859 3072
rect 3914 3006 3920 3014
rect 3853 2308 3859 2312
rect 3869 2288 3875 2612
rect 3914 2606 3920 2614
rect 3933 2308 3939 3112
rect 3965 2628 3971 3456
rect 3997 3228 4003 4512
rect 4125 4448 4131 4516
rect 4044 3923 4052 3924
rect 4040 3917 4052 3923
rect 4044 3916 4052 3917
rect 4061 3908 4067 3932
rect 4028 3716 4036 3724
rect 4013 3208 4019 3332
rect 3914 2206 3920 2214
rect 3756 1636 3764 1644
rect 3724 1456 3732 1464
rect 3469 904 3475 912
rect 3468 896 3476 904
rect 3421 624 3427 632
rect 3420 616 3428 624
rect 3453 588 3459 852
rect 3324 516 3332 524
rect 3325 508 3331 516
rect 3485 328 3491 952
rect 3517 668 3523 972
rect 3533 728 3539 1072
rect 3565 808 3571 1272
rect 3581 908 3587 1112
rect 3628 963 3636 964
rect 3624 957 3636 963
rect 3628 956 3636 957
rect 3549 488 3555 792
rect 3581 784 3587 892
rect 3580 776 3588 784
rect 3565 524 3571 532
rect 3661 528 3667 1232
rect 3725 908 3731 1456
rect 3676 736 3684 744
rect 3677 708 3683 736
rect 3725 708 3731 792
rect 3692 696 3700 704
rect 3693 688 3699 696
rect 3757 688 3763 1472
rect 3564 516 3572 524
rect 3596 416 3604 424
rect 3597 388 3603 416
rect 3628 336 3636 344
rect 3324 303 3332 304
rect 3320 297 3332 303
rect 3324 296 3332 297
rect 3436 303 3444 304
rect 3436 297 3448 303
rect 3436 296 3444 297
rect 3581 284 3587 292
rect 3629 288 3635 336
rect 3661 308 3667 392
rect 3580 276 3588 284
rect 3581 184 3587 276
rect 3677 248 3683 372
rect 3693 288 3699 552
rect 3756 536 3764 544
rect 3757 528 3763 536
rect 3773 528 3779 1312
rect 3789 1168 3795 1832
rect 3853 1788 3859 1892
rect 3914 1806 3920 1814
rect 3933 1668 3939 2292
rect 3981 1908 3987 3032
rect 4013 2428 4019 3072
rect 3997 2224 4003 2252
rect 3996 2216 4004 2224
rect 3820 1516 3828 1524
rect 3821 1508 3827 1516
rect 3836 1503 3844 1504
rect 3836 1497 3848 1503
rect 3836 1496 3844 1497
rect 3869 1108 3875 1652
rect 3981 1584 3987 1892
rect 3980 1576 3988 1584
rect 3997 1544 4003 1912
rect 4013 1908 4019 2412
rect 4029 2328 4035 3716
rect 4045 2528 4051 3892
rect 4076 3736 4084 3744
rect 4077 3728 4083 3736
rect 4029 2108 4035 2252
rect 4045 1848 4051 2452
rect 4061 2388 4067 3432
rect 4077 3304 4083 3312
rect 4076 3296 4084 3304
rect 4093 3188 4099 4052
rect 4109 3644 4115 3672
rect 4108 3636 4116 3644
rect 4093 3124 4099 3172
rect 4092 3116 4100 3124
rect 4077 2408 4083 2752
rect 4093 2124 4099 2152
rect 4092 2116 4100 2124
rect 4077 2084 4083 2112
rect 4076 2076 4084 2084
rect 4061 1804 4067 1852
rect 4060 1796 4068 1804
rect 3996 1536 4004 1544
rect 3981 1504 3987 1512
rect 3980 1496 3988 1504
rect 4077 1464 4083 2076
rect 4125 2028 4131 4432
rect 4429 4328 4435 4592
rect 4509 4524 4515 4532
rect 4508 4516 4516 4524
rect 4508 4496 4516 4504
rect 4236 4256 4244 4264
rect 4140 4156 4148 4164
rect 4141 3708 4147 4156
rect 4172 4103 4180 4104
rect 4168 4097 4180 4103
rect 4172 4096 4180 4097
rect 4237 3808 4243 4256
rect 4141 3168 4147 3692
rect 4173 2908 4179 3232
rect 4221 2188 4227 3452
rect 4252 3363 4260 3364
rect 4252 3357 4264 3363
rect 4252 3356 4260 3357
rect 4236 3303 4244 3304
rect 4236 3297 4248 3303
rect 4236 3296 4244 3297
rect 4172 2123 4180 2124
rect 4172 2117 4184 2123
rect 4172 2116 4180 2117
rect 4237 1968 4243 2972
rect 4269 2228 4275 2672
rect 4285 2548 4291 4192
rect 4333 4184 4339 4212
rect 4509 4208 4515 4496
rect 4525 4288 4531 4532
rect 4669 4368 4675 4652
rect 4717 4468 4723 4692
rect 4684 4443 4692 4444
rect 4684 4437 4696 4443
rect 4684 4436 4692 4437
rect 4828 4423 4836 4424
rect 4824 4417 4836 4423
rect 4828 4416 4836 4417
rect 4620 4363 4628 4364
rect 4620 4357 4632 4363
rect 4620 4356 4628 4357
rect 4845 4364 4851 4492
rect 4844 4356 4852 4364
rect 4332 4176 4340 4184
rect 4316 4116 4324 4124
rect 4317 3928 4323 4116
rect 4333 3488 4339 4176
rect 4349 3828 4355 4052
rect 4365 3568 4371 4132
rect 4413 4068 4419 4092
rect 4461 4008 4467 4032
rect 4381 3888 4387 3892
rect 4301 3384 4307 3412
rect 4300 3376 4308 3384
rect 4333 3228 4339 3352
rect 4349 3288 4355 3432
rect 4365 3308 4371 3552
rect 4381 3328 4387 3872
rect 4461 3868 4467 3992
rect 4477 3908 4483 4152
rect 4541 4148 4547 4272
rect 4621 3964 4627 4052
rect 4620 3956 4628 3964
rect 4428 3863 4436 3864
rect 4428 3857 4440 3863
rect 4428 3856 4436 3857
rect 4428 3356 4436 3364
rect 4429 3348 4435 3356
rect 4477 3328 4483 3892
rect 4540 3863 4548 3864
rect 4540 3857 4552 3863
rect 4540 3856 4548 3857
rect 4620 3843 4628 3844
rect 4620 3837 4632 3843
rect 4620 3836 4628 3837
rect 4333 2848 4339 3212
rect 4349 2768 4355 3192
rect 4349 2688 4355 2752
rect 4285 2228 4291 2532
rect 4300 2316 4308 2324
rect 4237 1888 4243 1952
rect 4076 1456 4084 1464
rect 3914 1406 3920 1414
rect 3933 1368 3939 1392
rect 3948 1343 3956 1344
rect 3948 1337 3960 1343
rect 3948 1336 3956 1337
rect 3933 1324 3939 1332
rect 3932 1316 3940 1324
rect 3981 1188 3987 1412
rect 4093 1388 4099 1832
rect 3914 1006 3920 1014
rect 3869 884 3875 992
rect 4109 884 4115 1732
rect 4125 1148 4131 1872
rect 4253 1868 4259 2012
rect 4205 1388 4211 1692
rect 4253 1524 4259 1852
rect 4269 1704 4275 1912
rect 4268 1696 4276 1704
rect 4252 1516 4260 1524
rect 4173 948 4179 1372
rect 3868 876 3876 884
rect 4108 876 4116 884
rect 3788 796 3796 804
rect 3789 708 3795 796
rect 3900 696 3908 704
rect 3773 484 3779 512
rect 3772 476 3780 484
rect 3773 468 3779 476
rect 3789 424 3795 452
rect 3788 416 3796 424
rect 3820 356 3828 364
rect 3708 316 3716 324
rect 3709 308 3715 316
rect 3821 308 3827 356
rect 3869 308 3875 672
rect 3901 668 3907 696
rect 3914 606 3920 614
rect 4045 524 4051 532
rect 4253 528 4259 1492
rect 4269 1228 4275 1652
rect 4285 1484 4291 2192
rect 4301 1768 4307 2316
rect 4317 1628 4323 2092
rect 4333 1588 4339 2512
rect 4349 2368 4355 2672
rect 4365 2488 4371 3052
rect 4381 2788 4387 3312
rect 4397 3188 4403 3312
rect 4397 2944 4403 3052
rect 4396 2936 4404 2944
rect 4413 2548 4419 3292
rect 4284 1476 4292 1484
rect 4285 1228 4291 1476
rect 4349 1288 4355 2272
rect 4397 1988 4403 2312
rect 4429 2048 4435 2912
rect 4445 2284 4451 2892
rect 4477 2708 4483 3312
rect 4493 2568 4499 3452
rect 4557 3408 4563 3672
rect 4637 3644 4643 3712
rect 4636 3636 4644 3644
rect 4653 3588 4659 3712
rect 4669 3628 4675 3832
rect 4509 3188 4515 3332
rect 4588 3316 4596 3324
rect 4557 3128 4563 3312
rect 4589 3308 4595 3316
rect 4444 2276 4452 2284
rect 4381 1508 4387 1892
rect 4269 568 4275 1212
rect 4317 884 4323 912
rect 4381 904 4387 912
rect 4380 896 4388 904
rect 4316 876 4324 884
rect 4285 648 4291 712
rect 4044 516 4052 524
rect 4124 523 4132 524
rect 4120 517 4132 523
rect 4124 516 4132 517
rect 3933 368 3939 452
rect 4252 363 4260 364
rect 4248 357 4260 363
rect 4252 356 4260 357
rect 3852 283 3860 284
rect 3852 277 3864 283
rect 3852 276 3860 277
rect 3580 176 3588 184
rect 3773 128 3779 212
rect 3914 206 3920 214
rect 3933 168 3939 352
rect 3964 336 3972 344
rect 3965 288 3971 336
rect 4285 188 4291 432
rect 4301 348 4307 852
rect 4365 724 4371 732
rect 4364 716 4372 724
rect 4365 208 4371 452
rect 4381 268 4387 896
rect 4429 848 4435 1472
rect 4412 723 4420 724
rect 4408 717 4420 723
rect 4412 716 4420 717
rect 4461 588 4467 2392
rect 4493 2208 4499 2532
rect 4525 2008 4531 2692
rect 4541 2688 4547 2932
rect 4541 1748 4547 2172
rect 4557 1528 4563 2212
rect 4588 2116 4596 2124
rect 4476 1456 4484 1464
rect 4477 1148 4483 1456
rect 4541 624 4547 652
rect 4540 616 4548 624
rect 4428 316 4436 324
rect 4429 288 4435 316
rect 4380 183 4388 184
rect 4376 177 4388 183
rect 4380 176 4388 177
rect 4477 128 4483 592
rect 4557 544 4563 892
rect 4573 608 4579 1112
rect 4589 608 4595 2116
rect 4605 1908 4611 2772
rect 4637 2628 4643 2932
rect 4653 2928 4659 3572
rect 4700 3343 4708 3344
rect 4696 3337 4708 3343
rect 4700 3336 4708 3337
rect 4669 3028 4675 3132
rect 4717 3108 4723 4112
rect 4797 4108 4803 4352
rect 4812 4296 4820 4304
rect 4813 4228 4819 4296
rect 4829 3768 4835 4272
rect 4877 3928 4883 4232
rect 4893 4208 4899 4512
rect 4938 4406 4944 4414
rect 5085 4304 5091 4312
rect 5084 4296 5092 4304
rect 4988 4283 4996 4284
rect 4984 4277 4996 4283
rect 4988 4276 4996 4277
rect 4892 4136 4900 4144
rect 4893 3868 4899 4136
rect 4938 4006 4944 4014
rect 4732 3723 4740 3724
rect 4732 3717 4744 3723
rect 4732 3716 4740 3717
rect 4653 2724 4659 2872
rect 4652 2716 4660 2724
rect 4652 2563 4660 2564
rect 4652 2557 4664 2563
rect 4652 2556 4660 2557
rect 4588 576 4596 584
rect 4589 568 4595 576
rect 4556 536 4564 544
rect 4588 516 4596 524
rect 4589 508 4595 516
rect 4605 288 4611 1892
rect 4637 1704 4643 2432
rect 4717 2308 4723 3092
rect 4733 3084 4739 3092
rect 4732 3076 4740 3084
rect 4749 2668 4755 3492
rect 4781 3304 4787 3392
rect 4780 3296 4788 3304
rect 4781 2968 4787 3296
rect 4636 1696 4644 1704
rect 4637 1088 4643 1696
rect 4653 1448 4659 2272
rect 4700 2223 4708 2224
rect 4696 2217 4708 2223
rect 4700 2216 4708 2217
rect 4685 1508 4691 1532
rect 4701 1388 4707 2216
rect 4733 1488 4739 2632
rect 4749 2164 4755 2652
rect 4765 2528 4771 2792
rect 4813 2548 4819 3132
rect 4844 3036 4852 3044
rect 4845 2908 4851 3036
rect 4893 3008 4899 3772
rect 4938 3606 4944 3614
rect 4938 3206 4944 3214
rect 4957 2988 4963 4252
rect 4973 4108 4979 4272
rect 5021 4148 5027 4232
rect 5004 4096 5012 4104
rect 4973 3668 4979 4012
rect 4989 3868 4995 4072
rect 5005 3928 5011 4096
rect 5021 3688 5027 4112
rect 5036 3956 5044 3964
rect 5037 3948 5043 3956
rect 4989 3064 4995 3212
rect 4988 3056 4996 3064
rect 4938 2806 4944 2814
rect 4989 2764 4995 3056
rect 4988 2756 4996 2764
rect 4844 2596 4852 2604
rect 4812 2323 4820 2324
rect 4808 2317 4820 2323
rect 4812 2316 4820 2317
rect 4748 2156 4756 2164
rect 4749 1584 4755 1692
rect 4748 1576 4756 1584
rect 4701 1328 4707 1372
rect 4749 1328 4755 1576
rect 4829 1568 4835 2132
rect 4765 1184 4771 1472
rect 4764 1176 4772 1184
rect 4829 1068 4835 1412
rect 4652 516 4660 524
rect 4653 508 4659 516
rect 4636 503 4644 504
rect 4632 497 4644 503
rect 4636 496 4644 497
rect 4685 408 4691 792
rect 4701 748 4707 952
rect 4748 876 4756 884
rect 4749 828 4755 876
rect 4733 448 4739 652
rect 4732 296 4740 304
rect 4589 264 4595 272
rect 4733 268 4739 296
rect 4749 268 4755 812
rect 4781 548 4787 712
rect 4797 504 4803 532
rect 4796 496 4804 504
rect 4588 256 4596 264
rect 3276 103 3284 104
rect 3276 97 3288 103
rect 3276 96 3284 97
rect 4829 48 4835 1052
rect 4845 628 4851 2596
rect 4877 2508 4883 2672
rect 4938 2406 4944 2414
rect 4893 1768 4899 2392
rect 4938 2006 4944 2014
rect 4957 1848 4963 2692
rect 4938 1606 4944 1614
rect 4861 948 4867 1252
rect 4877 1108 4883 1572
rect 4989 1408 4995 2756
rect 5005 2704 5011 2752
rect 5004 2696 5012 2704
rect 5005 1788 5011 1992
rect 4938 1206 4944 1214
rect 4877 348 4883 1092
rect 4893 728 4899 1152
rect 4925 1008 4931 1032
rect 4938 806 4944 814
rect 4957 628 4963 1392
rect 5021 1328 5027 3312
rect 5053 3144 5059 3452
rect 5069 3348 5075 4192
rect 5085 3268 5091 4072
rect 5101 3468 5107 4432
rect 5116 3636 5124 3644
rect 5117 3628 5123 3636
rect 5052 3136 5060 3144
rect 5052 2696 5060 2704
rect 5053 2688 5059 2696
rect 5037 1824 5043 1872
rect 5036 1816 5044 1824
rect 4973 1148 4979 1192
rect 5053 1004 5059 1852
rect 5085 1668 5091 3212
rect 5101 2884 5107 3232
rect 5117 3028 5123 3532
rect 5100 2876 5108 2884
rect 5101 2748 5107 2876
rect 5101 1804 5107 1812
rect 5100 1796 5108 1804
rect 5117 1728 5123 3012
rect 5133 3004 5139 4692
rect 5212 4503 5220 4504
rect 5208 4497 5220 4503
rect 5212 4496 5220 4497
rect 5292 4276 5300 4284
rect 5293 4268 5299 4276
rect 5181 4008 5187 4112
rect 5197 4084 5203 4152
rect 5261 4124 5267 4132
rect 5260 4116 5268 4124
rect 5196 4076 5204 4084
rect 5165 3408 5171 3832
rect 5181 3664 5187 3992
rect 5197 3744 5203 4076
rect 5196 3736 5204 3744
rect 5180 3656 5188 3664
rect 5197 3308 5203 3736
rect 5229 3508 5235 3572
rect 5132 2996 5140 3004
rect 5133 2908 5139 2996
rect 5149 2548 5155 2672
rect 5181 2408 5187 2832
rect 5197 2048 5203 3192
rect 5213 2568 5219 2852
rect 5213 1788 5219 2552
rect 5229 1808 5235 3492
rect 5277 3428 5283 3872
rect 5293 3608 5299 3692
rect 5293 3564 5299 3592
rect 5292 3556 5300 3564
rect 5293 3368 5299 3412
rect 5309 3344 5315 3352
rect 5308 3336 5316 3344
rect 5325 3188 5331 3952
rect 5341 3108 5347 4632
rect 5421 4148 5427 4272
rect 5405 4104 5411 4112
rect 5404 4096 5412 4104
rect 5245 2708 5251 2732
rect 5261 2688 5267 3072
rect 5245 2148 5251 2672
rect 5117 1664 5123 1712
rect 5116 1656 5124 1664
rect 5261 1528 5267 2392
rect 5357 2028 5363 3212
rect 5372 3116 5380 3124
rect 5373 3108 5379 3116
rect 5373 2468 5379 3092
rect 5421 2948 5427 3372
rect 5437 3328 5443 3832
rect 5453 3748 5459 4492
rect 5517 4208 5523 4672
rect 5962 4606 5968 4614
rect 5533 4368 5539 4372
rect 5533 4188 5539 4352
rect 5645 4144 5651 4552
rect 6173 4428 6179 4452
rect 5884 4323 5892 4324
rect 5880 4317 5892 4323
rect 5884 4316 5892 4317
rect 5725 4288 5731 4312
rect 5962 4206 5968 4214
rect 5644 4136 5652 4144
rect 5421 2888 5427 2932
rect 5404 2516 5412 2524
rect 5388 2476 5396 2484
rect 5389 2208 5395 2476
rect 5405 2468 5411 2516
rect 5389 1728 5395 2052
rect 5052 996 5060 1004
rect 4957 464 4963 492
rect 4956 456 4964 464
rect 4938 406 4944 414
rect 4893 324 4899 392
rect 5005 388 5011 512
rect 5069 484 5075 1312
rect 5180 943 5188 944
rect 5176 937 5188 943
rect 5180 936 5188 937
rect 5100 776 5108 784
rect 5101 728 5107 776
rect 5164 736 5172 744
rect 5165 728 5171 736
rect 5117 704 5123 712
rect 5116 696 5124 704
rect 5165 524 5171 552
rect 5196 536 5204 544
rect 5197 528 5203 536
rect 5164 516 5172 524
rect 5068 476 5076 484
rect 4892 316 4900 324
rect 4924 303 4932 304
rect 4920 297 4932 303
rect 4924 296 4932 297
rect 4957 248 4963 292
rect 4989 168 4995 352
rect 5052 316 5060 324
rect 5053 308 5059 316
rect 5069 308 5075 476
rect 5213 428 5219 932
rect 5213 368 5219 412
rect 5229 408 5235 972
rect 5261 568 5267 612
rect 5293 408 5299 772
rect 5309 488 5315 692
rect 5341 608 5347 1552
rect 5405 1308 5411 2452
rect 5437 2388 5443 3112
rect 5453 2448 5459 3492
rect 5629 3324 5635 3332
rect 5628 3316 5636 3324
rect 5645 3308 5651 4136
rect 5693 3948 5699 4072
rect 5661 3328 5667 3752
rect 5693 3408 5699 3932
rect 5805 3588 5811 3672
rect 5485 3048 5491 3172
rect 5516 3136 5524 3144
rect 5517 3128 5523 3136
rect 5533 2768 5539 3092
rect 5468 2736 5476 2744
rect 5421 2108 5427 2292
rect 5421 1328 5427 2092
rect 5469 1908 5475 2736
rect 5500 2603 5508 2604
rect 5500 2597 5512 2603
rect 5500 2596 5508 2597
rect 5469 1208 5475 1892
rect 5485 1888 5491 2592
rect 5516 2556 5524 2564
rect 5517 2548 5523 2556
rect 5484 1816 5492 1824
rect 5485 1368 5491 1816
rect 5357 684 5363 692
rect 5356 676 5364 684
rect 5325 128 5331 252
rect 5341 168 5347 592
rect 5373 548 5379 1072
rect 5389 908 5395 1072
rect 5501 688 5507 2192
rect 5517 1908 5523 2432
rect 5533 2168 5539 2632
rect 5549 2548 5555 2852
rect 5581 2008 5587 2972
rect 5644 2883 5652 2884
rect 5640 2877 5652 2883
rect 5644 2876 5652 2877
rect 5693 2288 5699 3152
rect 5725 3088 5731 3332
rect 5772 2763 5780 2764
rect 5768 2757 5780 2763
rect 5772 2756 5780 2757
rect 5629 1248 5635 2152
rect 5693 1824 5699 2272
rect 5741 2248 5747 2392
rect 5692 1816 5700 1824
rect 5693 1308 5699 1792
rect 5757 1248 5763 2492
rect 5789 1384 5795 2712
rect 5805 1588 5811 3032
rect 5821 2708 5827 4172
rect 6044 4123 6052 4124
rect 6044 4117 6056 4123
rect 6044 4116 6052 4117
rect 5852 4076 5860 4084
rect 5853 4068 5859 4076
rect 5885 3964 5891 4112
rect 5852 3956 5860 3964
rect 5884 3956 5892 3964
rect 5837 2308 5843 3312
rect 5853 1528 5859 3956
rect 5885 3428 5891 3892
rect 5869 3324 5875 3352
rect 5868 3316 5876 3324
rect 5901 3288 5907 4032
rect 5965 4028 5971 4112
rect 6044 4096 6052 4104
rect 5962 3806 5968 3814
rect 5981 3668 5987 3872
rect 5868 2696 5876 2704
rect 5869 2688 5875 2696
rect 5869 2128 5875 2672
rect 5885 1968 5891 3192
rect 5901 2388 5907 2952
rect 5917 2744 5923 3572
rect 5962 3406 5968 3414
rect 5962 3006 5968 3014
rect 5981 2928 5987 3652
rect 6029 3548 6035 4092
rect 6045 4088 6051 4096
rect 5916 2736 5924 2744
rect 5917 2728 5923 2736
rect 5917 2628 5923 2692
rect 5962 2606 5968 2614
rect 5981 2288 5987 2892
rect 5997 2688 6003 3212
rect 6029 2983 6035 3492
rect 6045 3148 6051 4072
rect 6077 3568 6083 4112
rect 6157 3368 6163 4232
rect 6173 3508 6179 4412
rect 6269 3608 6275 3912
rect 6285 3688 6291 4132
rect 6060 3123 6068 3124
rect 6056 3117 6068 3123
rect 6060 3116 6068 3117
rect 6013 2977 6035 2983
rect 5997 2568 6003 2612
rect 5885 1748 5891 1952
rect 5901 1488 5907 2272
rect 5962 2206 5968 2214
rect 5962 1806 5968 1814
rect 5997 1728 6003 2072
rect 6013 1888 6019 2977
rect 6093 2528 6099 2772
rect 6045 2288 6051 2492
rect 6109 2248 6115 3332
rect 6205 3308 6211 3432
rect 6221 3248 6227 3492
rect 6125 2484 6131 2512
rect 6124 2476 6132 2484
rect 6189 1948 6195 2692
rect 6205 2684 6211 2692
rect 6204 2676 6212 2684
rect 5788 1376 5796 1384
rect 5901 1288 5907 1472
rect 5962 1406 5968 1414
rect 5980 1376 5988 1384
rect 5517 588 5523 1092
rect 5533 728 5539 1152
rect 5981 1028 5987 1376
rect 5962 1006 5968 1014
rect 5549 868 5555 972
rect 5629 528 5635 752
rect 5645 568 5651 912
rect 5693 508 5699 992
rect 5962 606 5968 614
rect 5773 528 5779 572
rect 5548 496 5556 504
rect 5549 468 5555 496
rect 5549 328 5555 452
rect 5468 263 5476 264
rect 5464 257 5476 263
rect 5468 256 5476 257
rect 4988 123 4996 124
rect 4988 117 5000 123
rect 4988 116 4996 117
rect 5629 48 5635 272
rect 5965 248 5971 532
rect 5917 28 5923 232
rect 5962 206 5968 214
rect 5981 104 5987 1012
rect 6013 188 6019 1872
rect 6045 1808 6051 1932
rect 6045 1648 6051 1712
rect 6125 568 6131 1012
rect 6125 548 6131 552
rect 6141 268 6147 992
rect 6189 524 6195 1852
rect 6205 1548 6211 2632
rect 6221 2528 6227 2692
rect 6237 2688 6243 3512
rect 6285 3368 6291 3672
rect 6397 3588 6403 4152
rect 6253 2648 6259 2932
rect 6413 2508 6419 2792
rect 6381 2104 6387 2112
rect 6380 2096 6388 2104
rect 6221 1548 6227 1772
rect 6205 1508 6211 1532
rect 6205 868 6211 1272
rect 6237 1168 6243 1792
rect 6221 1088 6227 1152
rect 6188 516 6196 524
rect 6333 128 6339 1372
rect 6381 988 6387 1592
rect 6397 1488 6403 2272
rect 6413 1928 6419 2292
rect 6429 2288 6435 4132
rect 6573 3728 6579 4692
rect 6445 2548 6451 3472
rect 6445 2268 6451 2532
rect 6413 1548 6419 1912
rect 6429 1408 6435 2152
rect 6445 1848 6451 2252
rect 6461 2148 6467 3612
rect 6557 2948 6563 3132
rect 6557 2148 6563 2752
rect 6445 1428 6451 1832
rect 6461 1468 6467 1892
rect 6429 1028 6435 1392
rect 6476 516 6484 524
rect 6477 508 6483 516
rect 6509 168 6515 1732
rect 6525 1328 6531 1952
rect 6525 1008 6531 1312
rect 6540 943 6548 944
rect 6536 937 6548 943
rect 6540 936 6548 937
rect 6557 868 6563 1832
rect 6573 308 6579 3712
rect 6669 3448 6675 3732
rect 6717 2928 6723 3392
rect 6589 2768 6595 2812
rect 6589 1508 6595 2752
rect 6717 2548 6723 2892
rect 6589 188 6595 1472
rect 6605 188 6611 1532
rect 6621 328 6627 2512
rect 6637 2128 6643 2192
rect 6637 1328 6643 1892
rect 6653 1728 6659 2512
rect 6701 1908 6707 2352
rect 6637 848 6643 1312
rect 6653 128 6659 1352
rect 6701 1308 6707 1492
rect 6717 1328 6723 1752
rect 6733 1508 6739 1932
rect 6733 1348 6739 1392
rect 6732 716 6740 724
rect 6733 708 6739 716
rect 6749 308 6755 3452
rect 6765 388 6771 2552
rect 6797 688 6803 3752
rect 6813 2968 6819 2992
rect 5980 103 5988 104
rect 5976 97 5988 103
rect 5980 96 5988 97
rect 826 6 832 14
rect 2890 6 2896 14
rect 4938 6 4944 14
use BUFX2  BUFX2_70
timestamp 1515852544
transform -1 0 56 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_12
timestamp 1515852544
transform -1 0 104 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_51
timestamp 1515852544
transform 1 0 104 0 1 4610
box 0 0 48 200
use INVX1  INVX1_9
timestamp 1515852544
transform -1 0 184 0 1 4610
box 0 0 32 200
use INVX1  INVX1_14
timestamp 1515852544
transform 1 0 184 0 1 4610
box 0 0 32 200
use NOR2X1  NOR2X1_55
timestamp 1515852544
transform 1 0 216 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_34
timestamp 1515852544
transform 1 0 264 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_74
timestamp 1515852544
transform 1 0 312 0 1 4610
box 0 0 48 200
use INVX1  INVX1_17
timestamp 1515852544
transform 1 0 360 0 1 4610
box 0 0 32 200
use NOR2X1  NOR2X1_59
timestamp 1515852544
transform 1 0 392 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_37
timestamp 1515852544
transform 1 0 440 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_40
timestamp 1515852544
transform 1 0 488 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_39
timestamp 1515852544
transform 1 0 536 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_36
timestamp 1515852544
transform -1 0 632 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_58
timestamp 1515852544
transform -1 0 680 0 1 4610
box 0 0 48 200
use INVX1  INVX1_16
timestamp 1515852544
transform -1 0 712 0 1 4610
box 0 0 32 200
use INVX8  INVX8_1
timestamp 1515852544
transform -1 0 792 0 1 4610
box 0 0 80 200
use BUFX2  BUFX2_67
timestamp 1515852544
transform -1 0 840 0 1 4610
box 0 0 48 200
use FILL  FILL_23_0_0
timestamp 1515852544
transform -1 0 856 0 1 4610
box 0 0 16 200
use FILL  FILL_23_0_1
timestamp 1515852544
transform -1 0 872 0 1 4610
box 0 0 16 200
use BUFX2  BUFX2_4
timestamp 1515852544
transform -1 0 920 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_62
timestamp 1515852544
transform -1 0 968 0 1 4610
box 0 0 48 200
use INVX1  INVX1_20
timestamp 1515852544
transform -1 0 1000 0 1 4610
box 0 0 32 200
use BUFX2  BUFX2_13
timestamp 1515852544
transform 1 0 1000 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_49
timestamp 1515852544
transform 1 0 1048 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_226
timestamp 1515852544
transform 1 0 1096 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_42
timestamp 1515852544
transform -1 0 1208 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_108
timestamp 1515852544
transform 1 0 1208 0 1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_80
timestamp 1515852544
transform -1 0 1592 0 1 4610
box 0 0 192 200
use BUFX2  BUFX2_11
timestamp 1515852544
transform 1 0 1592 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_48
timestamp 1515852544
transform 1 0 1640 0 1 4610
box 0 0 48 200
use INVX2  INVX2_4
timestamp 1515852544
transform -1 0 1720 0 1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_130
timestamp 1515852544
transform -1 0 1912 0 1 4610
box 0 0 192 200
use FILL  FILL_23_1_0
timestamp 1515852544
transform -1 0 1928 0 1 4610
box 0 0 16 200
use FILL  FILL_23_1_1
timestamp 1515852544
transform -1 0 1944 0 1 4610
box 0 0 16 200
use BUFX2  BUFX2_58
timestamp 1515852544
transform -1 0 1992 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_22
timestamp 1515852544
transform -1 0 2040 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_79
timestamp 1515852544
transform -1 0 2232 0 1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_153
timestamp 1515852544
transform -1 0 2424 0 1 4610
box 0 0 192 200
use BUFX2  BUFX2_47
timestamp 1515852544
transform -1 0 2472 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_10
timestamp 1515852544
transform -1 0 2520 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_183
timestamp 1515852544
transform 1 0 2520 0 1 4610
box 0 0 192 200
use NAND2X1  NAND2X1_177
timestamp 1515852544
transform 1 0 2712 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_26
timestamp 1515852544
transform -1 0 2824 0 1 4610
box 0 0 64 200
use FILL  FILL_23_2_0
timestamp 1515852544
transform 1 0 2824 0 1 4610
box 0 0 16 200
use FILL  FILL_23_2_1
timestamp 1515852544
transform 1 0 2840 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_127
timestamp 1515852544
transform 1 0 2856 0 1 4610
box 0 0 192 200
use BUFX2  BUFX2_55
timestamp 1515852544
transform 1 0 3048 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_138
timestamp 1515852544
transform -1 0 3288 0 1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_18
timestamp 1515852544
transform -1 0 3352 0 1 4610
box 0 0 64 200
use BUFX4  BUFX4_177
timestamp 1515852544
transform -1 0 3416 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_141
timestamp 1515852544
transform -1 0 3608 0 1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_21
timestamp 1515852544
transform -1 0 3672 0 1 4610
box 0 0 64 200
use BUFX4  BUFX4_167
timestamp 1515852544
transform -1 0 3736 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_174
timestamp 1515852544
transform -1 0 3928 0 1 4610
box 0 0 192 200
use FILL  FILL_23_3_0
timestamp 1515852544
transform 1 0 3928 0 1 4610
box 0 0 16 200
use FILL  FILL_23_3_1
timestamp 1515852544
transform 1 0 3944 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_235
timestamp 1515852544
transform 1 0 3960 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_51
timestamp 1515852544
transform 1 0 4008 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_185
timestamp 1515852544
transform 1 0 4072 0 1 4610
box 0 0 192 200
use AOI22X1  AOI22X1_189
timestamp 1515852544
transform 1 0 4264 0 1 4610
box 0 0 80 200
use NAND3X1  NAND3X1_100
timestamp 1515852544
transform -1 0 4408 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_19
timestamp 1515852544
transform -1 0 4456 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_119
timestamp 1515852544
transform -1 0 4648 0 1 4610
box 0 0 192 200
use INVX1  INVX1_53
timestamp 1515852544
transform 1 0 4648 0 1 4610
box 0 0 32 200
use INVX1  INVX1_52
timestamp 1515852544
transform -1 0 4712 0 1 4610
box 0 0 32 200
use NAND2X1  NAND2X1_205
timestamp 1515852544
transform 1 0 4712 0 1 4610
box 0 0 48 200
use AOI22X1  AOI22X1_73
timestamp 1515852544
transform -1 0 4840 0 1 4610
box 0 0 80 200
use NAND2X1  NAND2X1_169
timestamp 1515852544
transform 1 0 4840 0 1 4610
box 0 0 48 200
use FILL  FILL_23_4_0
timestamp 1515852544
transform 1 0 4888 0 1 4610
box 0 0 16 200
use FILL  FILL_23_4_1
timestamp 1515852544
transform 1 0 4904 0 1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_22
timestamp 1515852544
transform 1 0 4920 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_143
timestamp 1515852544
transform -1 0 5176 0 1 4610
box 0 0 192 200
use BUFX4  BUFX4_180
timestamp 1515852544
transform 1 0 5176 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_148
timestamp 1515852544
transform -1 0 5432 0 1 4610
box 0 0 192 200
use BUFX2  BUFX2_50
timestamp 1515852544
transform -1 0 5480 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_14
timestamp 1515852544
transform -1 0 5528 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_16
timestamp 1515852544
transform 1 0 5528 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_52
timestamp 1515852544
transform 1 0 5576 0 1 4610
box 0 0 48 200
use BUFX4  BUFX4_170
timestamp 1515852544
transform 1 0 5624 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1515852544
transform 1 0 5688 0 1 4610
box 0 0 192 200
use FILL  FILL_23_5_0
timestamp 1515852544
transform 1 0 5880 0 1 4610
box 0 0 16 200
use FILL  FILL_23_5_1
timestamp 1515852544
transform 1 0 5896 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1515852544
transform 1 0 5912 0 1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_99
timestamp 1515852544
transform 1 0 6104 0 1 4610
box 0 0 192 200
use BUFX2  BUFX2_63
timestamp 1515852544
transform -1 0 6344 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_28
timestamp 1515852544
transform -1 0 6392 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_26
timestamp 1515852544
transform 1 0 6392 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_61
timestamp 1515852544
transform 1 0 6440 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_30
timestamp 1515852544
transform 1 0 6488 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_65
timestamp 1515852544
transform 1 0 6536 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_42
timestamp 1515852544
transform -1 0 6632 0 1 4610
box 0 0 48 200
use BUFX2  BUFX2_3
timestamp 1515852544
transform -1 0 6680 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_61
timestamp 1515852544
transform -1 0 6728 0 1 4610
box 0 0 48 200
use INVX1  INVX1_19
timestamp 1515852544
transform -1 0 6760 0 1 4610
box 0 0 32 200
use FILL  FILL_24_1
timestamp 1515852544
transform 1 0 6760 0 1 4610
box 0 0 16 200
use FILL  FILL_24_2
timestamp 1515852544
transform 1 0 6776 0 1 4610
box 0 0 16 200
use FILL  FILL_24_3
timestamp 1515852544
transform 1 0 6792 0 1 4610
box 0 0 16 200
use BUFX2  BUFX2_60
timestamp 1515852544
transform -1 0 56 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_25
timestamp 1515852544
transform -1 0 104 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_97
timestamp 1515852544
transform -1 0 296 0 -1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_175
timestamp 1515852544
transform -1 0 488 0 -1 4610
box 0 0 192 200
use BUFX2  BUFX2_59
timestamp 1515852544
transform -1 0 536 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_24
timestamp 1515852544
transform -1 0 584 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_312
timestamp 1515852544
transform 1 0 584 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_90
timestamp 1515852544
transform -1 0 824 0 -1 4610
box 0 0 192 200
use FILL  FILL_22_0_0
timestamp 1515852544
transform -1 0 840 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_1
timestamp 1515852544
transform -1 0 856 0 -1 4610
box 0 0 16 200
use INVX8  INVX8_16
timestamp 1515852544
transform -1 0 936 0 -1 4610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_164
timestamp 1515852544
transform -1 0 1128 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_635
timestamp 1515852544
transform 1 0 1128 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_227
timestamp 1515852544
transform -1 0 1240 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_633
timestamp 1515852544
transform -1 0 1304 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_636
timestamp 1515852544
transform 1 0 1304 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_99
timestamp 1515852544
transform -1 0 1448 0 -1 4610
box 0 0 80 200
use NAND2X1  NAND2X1_311
timestamp 1515852544
transform 1 0 1448 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_92
timestamp 1515852544
transform 1 0 1496 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_180
timestamp 1515852544
transform 1 0 1560 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_63
timestamp 1515852544
transform -1 0 1704 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_310
timestamp 1515852544
transform 1 0 1704 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_61
timestamp 1515852544
transform -1 0 1816 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_1_0
timestamp 1515852544
transform 1 0 1816 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_1
timestamp 1515852544
transform 1 0 1832 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_540
timestamp 1515852544
transform 1 0 1848 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_185
timestamp 1515852544
transform -1 0 1960 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_29
timestamp 1515852544
transform 1 0 1960 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_184
timestamp 1515852544
transform 1 0 2024 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_539
timestamp 1515852544
transform 1 0 2072 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_541
timestamp 1515852544
transform 1 0 2136 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_82
timestamp 1515852544
transform -1 0 2280 0 -1 4610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_132
timestamp 1515852544
transform -1 0 2472 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_543
timestamp 1515852544
transform 1 0 2472 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_186
timestamp 1515852544
transform -1 0 2584 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_30
timestamp 1515852544
transform -1 0 2648 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_83
timestamp 1515852544
transform 1 0 2648 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_546
timestamp 1515852544
transform -1 0 2792 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_187
timestamp 1515852544
transform 1 0 2792 0 -1 4610
box 0 0 48 200
use FILL  FILL_22_2_0
timestamp 1515852544
transform -1 0 2856 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_1
timestamp 1515852544
transform -1 0 2872 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_544
timestamp 1515852544
transform -1 0 2936 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_526
timestamp 1515852544
transform -1 0 3000 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_178
timestamp 1515852544
transform 1 0 3000 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_527
timestamp 1515852544
transform -1 0 3112 0 -1 4610
box 0 0 64 200
use INVX1  INVX1_1
timestamp 1515852544
transform 1 0 3112 0 -1 4610
box 0 0 32 200
use OAI22X1  OAI22X1_1
timestamp 1515852544
transform -1 0 3224 0 -1 4610
box 0 0 80 200
use INVX1  INVX1_32
timestamp 1515852544
transform -1 0 3256 0 -1 4610
box 0 0 32 200
use AOI22X1  AOI22X1_69
timestamp 1515852544
transform 1 0 3256 0 -1 4610
box 0 0 80 200
use NAND2X1  NAND2X1_159
timestamp 1515852544
transform 1 0 3336 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_481
timestamp 1515852544
transform -1 0 3448 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_482
timestamp 1515852544
transform -1 0 3512 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_160
timestamp 1515852544
transform -1 0 3560 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_494
timestamp 1515852544
transform 1 0 3560 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_165
timestamp 1515852544
transform -1 0 3672 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_166
timestamp 1515852544
transform 1 0 3672 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_495
timestamp 1515852544
transform 1 0 3720 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_493
timestamp 1515852544
transform 1 0 3784 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_72
timestamp 1515852544
transform 1 0 3848 0 -1 4610
box 0 0 80 200
use FILL  FILL_22_3_0
timestamp 1515852544
transform -1 0 3944 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_3_1
timestamp 1515852544
transform -1 0 3960 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_496
timestamp 1515852544
transform -1 0 4024 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_101
timestamp 1515852544
transform -1 0 4088 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_112
timestamp 1515852544
transform 1 0 4088 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_113
timestamp 1515852544
transform -1 0 4232 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_90
timestamp 1515852544
transform -1 0 4296 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_224
timestamp 1515852544
transform -1 0 4344 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_18
timestamp 1515852544
transform 1 0 4344 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_116
timestamp 1515852544
transform 1 0 4392 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_117
timestamp 1515852544
transform -1 0 4520 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_115
timestamp 1515852544
transform 1 0 4520 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_118
timestamp 1515852544
transform -1 0 4648 0 -1 4610
box 0 0 64 200
use OAI22X1  OAI22X1_10
timestamp 1515852544
transform -1 0 4728 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_589
timestamp 1515852544
transform 1 0 4728 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_36
timestamp 1515852544
transform 1 0 4792 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_91
timestamp 1515852544
transform 1 0 4856 0 -1 4610
box 0 0 80 200
use FILL  FILL_22_4_0
timestamp 1515852544
transform 1 0 4936 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_4_1
timestamp 1515852544
transform 1 0 4952 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_591
timestamp 1515852544
transform 1 0 4968 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_500
timestamp 1515852544
transform 1 0 5032 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_593
timestamp 1515852544
transform -1 0 5160 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_206
timestamp 1515852544
transform -1 0 5208 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_499
timestamp 1515852544
transform 1 0 5208 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_498
timestamp 1515852544
transform 1 0 5272 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_167
timestamp 1515852544
transform -1 0 5384 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_524
timestamp 1515852544
transform -1 0 5448 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_520
timestamp 1515852544
transform 1 0 5448 0 -1 4610
box 0 0 64 200
use OR2X2  OR2X2_9
timestamp 1515852544
transform -1 0 5576 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_181
timestamp 1515852544
transform -1 0 5768 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_446
timestamp 1515852544
transform -1 0 5832 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_412
timestamp 1515852544
transform -1 0 5896 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_145
timestamp 1515852544
transform -1 0 5960 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_5_0
timestamp 1515852544
transform 1 0 5960 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_5_1
timestamp 1515852544
transform 1 0 5976 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_149
timestamp 1515852544
transform 1 0 5992 0 -1 4610
box 0 0 64 200
use AOI22X1  AOI22X1_193
timestamp 1515852544
transform -1 0 6136 0 -1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_148
timestamp 1515852544
transform -1 0 6200 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_24
timestamp 1515852544
transform 1 0 6200 0 -1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_101
timestamp 1515852544
transform -1 0 6584 0 -1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_103
timestamp 1515852544
transform -1 0 6776 0 -1 4610
box 0 0 192 200
use FILL  FILL_23_1
timestamp 1515852544
transform -1 0 6792 0 -1 4610
box 0 0 16 200
use FILL  FILL_23_2
timestamp 1515852544
transform -1 0 6808 0 -1 4610
box 0 0 16 200
use INVX1  INVX1_23
timestamp 1515852544
transform 1 0 8 0 1 4210
box 0 0 32 200
use BUFX2  BUFX2_44
timestamp 1515852544
transform -1 0 88 0 1 4210
box 0 0 48 200
use BUFX2  BUFX2_7
timestamp 1515852544
transform -1 0 136 0 1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_65
timestamp 1515852544
transform 1 0 136 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_81
timestamp 1515852544
transform 1 0 184 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_229
timestamp 1515852544
transform 1 0 376 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_639
timestamp 1515852544
transform 1 0 424 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_93
timestamp 1515852544
transform -1 0 552 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_3
timestamp 1515852544
transform 1 0 552 0 1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_181
timestamp 1515852544
transform 1 0 600 0 1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_65
timestamp 1515852544
transform 1 0 680 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_66
timestamp 1515852544
transform -1 0 808 0 1 4210
box 0 0 64 200
use FILL  FILL_21_0_0
timestamp 1515852544
transform -1 0 824 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_1
timestamp 1515852544
transform -1 0 840 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_67
timestamp 1515852544
transform -1 0 904 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_64
timestamp 1515852544
transform -1 0 968 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_62
timestamp 1515852544
transform 1 0 968 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_60
timestamp 1515852544
transform 1 0 1032 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_161
timestamp 1515852544
transform 1 0 1096 0 1 4210
box 0 0 80 200
use NAND3X1  NAND3X1_63
timestamp 1515852544
transform -1 0 1240 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_171
timestamp 1515852544
transform 1 0 1240 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_538
timestamp 1515852544
transform 1 0 1432 0 1 4210
box 0 0 64 200
use INVX2  INVX2_3
timestamp 1515852544
transform 1 0 1496 0 1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_154
timestamp 1515852544
transform -1 0 1720 0 1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_15
timestamp 1515852544
transform 1 0 1720 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_103
timestamp 1515852544
transform -1 0 1848 0 1 4210
box 0 0 64 200
use FILL  FILL_21_1_0
timestamp 1515852544
transform 1 0 1848 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_1
timestamp 1515852544
transform 1 0 1864 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_102
timestamp 1515852544
transform 1 0 1880 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_542
timestamp 1515852544
transform 1 0 1944 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_103
timestamp 1515852544
transform 1 0 2008 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_12
timestamp 1515852544
transform -1 0 2120 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_525
timestamp 1515852544
transform 1 0 2120 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_78
timestamp 1515852544
transform 1 0 2184 0 1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_528
timestamp 1515852544
transform -1 0 2328 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_88
timestamp 1515852544
transform -1 0 2392 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_187
timestamp 1515852544
transform 1 0 2392 0 1 4210
box 0 0 80 200
use NAND2X1  NAND2X1_15
timestamp 1515852544
transform 1 0 2472 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_98
timestamp 1515852544
transform 1 0 2520 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_156
timestamp 1515852544
transform -1 0 2648 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_159
timestamp 1515852544
transform 1 0 2648 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_483
timestamp 1515852544
transform 1 0 2712 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_480
timestamp 1515852544
transform 1 0 2776 0 1 4210
box 0 0 64 200
use FILL  FILL_21_2_0
timestamp 1515852544
transform 1 0 2840 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_1
timestamp 1515852544
transform 1 0 2856 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_505
timestamp 1515852544
transform 1 0 2872 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_502
timestamp 1515852544
transform 1 0 2936 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_74
timestamp 1515852544
transform -1 0 3080 0 1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_504
timestamp 1515852544
transform 1 0 3080 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_503
timestamp 1515852544
transform -1 0 3208 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_171
timestamp 1515852544
transform -1 0 3256 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_23
timestamp 1515852544
transform 1 0 3256 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_170
timestamp 1515852544
transform -1 0 3368 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_144
timestamp 1515852544
transform 1 0 3368 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1515852544
transform -1 0 3752 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_68
timestamp 1515852544
transform 1 0 3752 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_20
timestamp 1515852544
transform 1 0 3816 0 1 4210
box 0 0 48 200
use FILL  FILL_21_3_0
timestamp 1515852544
transform -1 0 3880 0 1 4210
box 0 0 16 200
use FILL  FILL_21_3_1
timestamp 1515852544
transform -1 0 3896 0 1 4210
box 0 0 16 200
use NAND3X1  NAND3X1_101
timestamp 1515852544
transform -1 0 3960 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_120
timestamp 1515852544
transform -1 0 4024 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_21
timestamp 1515852544
transform 1 0 4024 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_121
timestamp 1515852544
transform -1 0 4136 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_91
timestamp 1515852544
transform -1 0 4200 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_92
timestamp 1515852544
transform 1 0 4200 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_588
timestamp 1515852544
transform 1 0 4264 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_204
timestamp 1515852544
transform -1 0 4376 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_587
timestamp 1515852544
transform 1 0 4376 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_595
timestamp 1515852544
transform 1 0 4440 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_92
timestamp 1515852544
transform -1 0 4584 0 1 4210
box 0 0 80 200
use NAND3X1  NAND3X1_37
timestamp 1515852544
transform 1 0 4584 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_121
timestamp 1515852544
transform 1 0 4648 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_497
timestamp 1515852544
transform 1 0 4840 0 1 4210
box 0 0 64 200
use FILL  FILL_21_4_0
timestamp 1515852544
transform 1 0 4904 0 1 4210
box 0 0 16 200
use FILL  FILL_21_4_1
timestamp 1515852544
transform 1 0 4920 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_22
timestamp 1515852544
transform 1 0 4936 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_123
timestamp 1515852544
transform 1 0 4984 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_128
timestamp 1515852544
transform 1 0 5048 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1515852544
transform 1 0 5112 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_423
timestamp 1515852544
transform 1 0 5304 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_434
timestamp 1515852544
transform -1 0 5432 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_155
timestamp 1515852544
transform 1 0 5432 0 1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_144
timestamp 1515852544
transform 1 0 5512 0 1 4210
box 0 0 64 200
use INVX1  INVX1_86
timestamp 1515852544
transform -1 0 5608 0 1 4210
box 0 0 32 200
use OR2X2  OR2X2_19
timestamp 1515852544
transform 1 0 5608 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_143
timestamp 1515852544
transform 1 0 5672 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_141
timestamp 1515852544
transform 1 0 5736 0 1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_192
timestamp 1515852544
transform -1 0 5880 0 1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_142
timestamp 1515852544
transform -1 0 5944 0 1 4210
box 0 0 64 200
use FILL  FILL_21_5_0
timestamp 1515852544
transform 1 0 5944 0 1 4210
box 0 0 16 200
use FILL  FILL_21_5_1
timestamp 1515852544
transform 1 0 5960 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_147
timestamp 1515852544
transform 1 0 5976 0 1 4210
box 0 0 64 200
use INVX8  INVX8_15
timestamp 1515852544
transform -1 0 6120 0 1 4210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_136
timestamp 1515852544
transform -1 0 6312 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_147
timestamp 1515852544
transform -1 0 6504 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_46
timestamp 1515852544
transform 1 0 6504 0 1 4210
box 0 0 192 200
use BUFX2  BUFX2_29
timestamp 1515852544
transform 1 0 6696 0 1 4210
box 0 0 48 200
use BUFX2  BUFX2_64
timestamp 1515852544
transform 1 0 6744 0 1 4210
box 0 0 48 200
use FILL  FILL_22_1
timestamp 1515852544
transform 1 0 6792 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_129
timestamp 1515852544
transform -1 0 200 0 -1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_110
timestamp 1515852544
transform 1 0 200 0 -1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_43
timestamp 1515852544
transform 1 0 392 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_638
timestamp 1515852544
transform 1 0 456 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_228
timestamp 1515852544
transform -1 0 568 0 -1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_128
timestamp 1515852544
transform 1 0 568 0 -1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_180
timestamp 1515852544
transform 1 0 760 0 -1 4210
box 0 0 48 200
use FILL  FILL_20_0_0
timestamp 1515852544
transform -1 0 824 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_1
timestamp 1515852544
transform -1 0 840 0 -1 4210
box 0 0 16 200
use NAND3X1  NAND3X1_27
timestamp 1515852544
transform -1 0 904 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_80
timestamp 1515852544
transform 1 0 904 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_530
timestamp 1515852544
transform 1 0 984 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_532
timestamp 1515852544
transform -1 0 1112 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_181
timestamp 1515852544
transform 1 0 1112 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_531
timestamp 1515852544
transform -1 0 1224 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_35
timestamp 1515852544
transform 1 0 1224 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_46
timestamp 1515852544
transform 1 0 1272 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_112
timestamp 1515852544
transform 1 0 1320 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_223
timestamp 1515852544
transform -1 0 1448 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_334
timestamp 1515852544
transform -1 0 1512 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_529
timestamp 1515852544
transform -1 0 1576 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_65
timestamp 1515852544
transform 1 0 1576 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_1
timestamp 1515852544
transform -1 0 1672 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_151
timestamp 1515852544
transform 1 0 1672 0 -1 4210
box 0 0 48 200
use AOI22X1  AOI22X1_63
timestamp 1515852544
transform 1 0 1720 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_451
timestamp 1515852544
transform 1 0 1800 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_1_0
timestamp 1515852544
transform 1 0 1864 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_1
timestamp 1515852544
transform 1 0 1880 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_150
timestamp 1515852544
transform 1 0 1896 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_449
timestamp 1515852544
transform -1 0 2008 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_195
timestamp 1515852544
transform -1 0 2072 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_104
timestamp 1515852544
transform 1 0 2072 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_186
timestamp 1515852544
transform -1 0 2216 0 -1 4210
box 0 0 80 200
use NAND3X1  NAND3X1_97
timestamp 1515852544
transform 1 0 2216 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_100
timestamp 1515852544
transform -1 0 2344 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_102
timestamp 1515852544
transform -1 0 2408 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_11
timestamp 1515852544
transform -1 0 2456 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_108
timestamp 1515852544
transform 1 0 2456 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_107
timestamp 1515852544
transform -1 0 2584 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_105
timestamp 1515852544
transform 1 0 2584 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_106
timestamp 1515852544
transform -1 0 2712 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_14
timestamp 1515852544
transform -1 0 2760 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_688
timestamp 1515852544
transform 1 0 2760 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_57
timestamp 1515852544
transform -1 0 2904 0 -1 4210
box 0 0 80 200
use FILL  FILL_20_2_0
timestamp 1515852544
transform 1 0 2904 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_1
timestamp 1515852544
transform 1 0 2920 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_666
timestamp 1515852544
transform 1 0 2936 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_113
timestamp 1515852544
transform -1 0 3048 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_74
timestamp 1515852544
transform -1 0 3112 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_135
timestamp 1515852544
transform 1 0 3112 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_677
timestamp 1515852544
transform -1 0 3224 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_445
timestamp 1515852544
transform -1 0 3288 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_57
timestamp 1515852544
transform -1 0 3352 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_51
timestamp 1515852544
transform -1 0 3384 0 -1 4210
box 0 0 32 200
use NOR2X1  NOR2X1_27
timestamp 1515852544
transform -1 0 3432 0 -1 4210
box 0 0 48 200
use BUFX4  BUFX4_131
timestamp 1515852544
transform -1 0 3496 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_184
timestamp 1515852544
transform 1 0 3496 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_217
timestamp 1515852544
transform 1 0 3560 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_50
timestamp 1515852544
transform -1 0 3656 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_224
timestamp 1515852544
transform 1 0 3656 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_130
timestamp 1515852544
transform -1 0 3800 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_212
timestamp 1515852544
transform 1 0 3800 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_3_0
timestamp 1515852544
transform 1 0 3864 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_3_1
timestamp 1515852544
transform 1 0 3880 0 -1 4210
box 0 0 16 200
use AOI22X1  AOI22X1_190
timestamp 1515852544
transform 1 0 3896 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_122
timestamp 1515852544
transform -1 0 4040 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_119
timestamp 1515852544
transform -1 0 4104 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_130
timestamp 1515852544
transform 1 0 4104 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_158
timestamp 1515852544
transform 1 0 4168 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_87
timestamp 1515852544
transform 1 0 4232 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_548
timestamp 1515852544
transform 1 0 4296 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_592
timestamp 1515852544
transform 1 0 4360 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_594
timestamp 1515852544
transform 1 0 4424 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_207
timestamp 1515852544
transform -1 0 4536 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_29
timestamp 1515852544
transform 1 0 4536 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_126
timestamp 1515852544
transform 1 0 4584 0 -1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_9
timestamp 1515852544
transform 1 0 4648 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_26
timestamp 1515852544
transform -1 0 4760 0 -1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_23
timestamp 1515852544
transform -1 0 4808 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_125
timestamp 1515852544
transform -1 0 4872 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_521
timestamp 1515852544
transform 1 0 4872 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_4_0
timestamp 1515852544
transform -1 0 4952 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_4_1
timestamp 1515852544
transform -1 0 4968 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_522
timestamp 1515852544
transform -1 0 5032 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_152
timestamp 1515852544
transform 1 0 5032 0 -1 4210
box 0 0 80 200
use AOI22X1  AOI22X1_77
timestamp 1515852544
transform 1 0 5112 0 -1 4210
box 0 0 80 200
use AOI21X1  AOI21X1_49
timestamp 1515852544
transform 1 0 5192 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_368
timestamp 1515852544
transform 1 0 5256 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_146
timestamp 1515852544
transform -1 0 5400 0 -1 4210
box 0 0 80 200
use OAI21X1  OAI21X1_346
timestamp 1515852544
transform 1 0 5400 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1515852544
transform 1 0 5464 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_140
timestamp 1515852544
transform 1 0 5656 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_139
timestamp 1515852544
transform 1 0 5720 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_81
timestamp 1515852544
transform -1 0 5816 0 -1 4210
box 0 0 32 200
use AOI21X1  AOI21X1_11
timestamp 1515852544
transform -1 0 5880 0 -1 4210
box 0 0 64 200
use OAI22X1  OAI22X1_21
timestamp 1515852544
transform -1 0 5960 0 -1 4210
box 0 0 80 200
use FILL  FILL_20_5_0
timestamp 1515852544
transform 1 0 5960 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_5_1
timestamp 1515852544
transform 1 0 5976 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_567
timestamp 1515852544
transform 1 0 5992 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_566
timestamp 1515852544
transform 1 0 6056 0 -1 4210
box 0 0 64 200
use AOI22X1  AOI22X1_85
timestamp 1515852544
transform -1 0 6200 0 -1 4210
box 0 0 80 200
use INVX1  INVX1_80
timestamp 1515852544
transform 1 0 6200 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_569
timestamp 1515852544
transform -1 0 6296 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_565
timestamp 1515852544
transform 1 0 6296 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_35
timestamp 1515852544
transform 1 0 6360 0 -1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_102
timestamp 1515852544
transform 1 0 6552 0 -1 4210
box 0 0 192 200
use BUFX2  BUFX2_18
timestamp 1515852544
transform 1 0 6744 0 -1 4210
box 0 0 48 200
use FILL  FILL_21_1
timestamp 1515852544
transform -1 0 6808 0 -1 4210
box 0 0 16 200
use BUFX2  BUFX2_57
timestamp 1515852544
transform -1 0 56 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_21
timestamp 1515852544
transform -1 0 104 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_68
timestamp 1515852544
transform -1 0 296 0 1 3810
box 0 0 192 200
use NAND3X1  NAND3X1_28
timestamp 1515852544
transform 1 0 296 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_81
timestamp 1515852544
transform 1 0 360 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_533
timestamp 1515852544
transform -1 0 504 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_640
timestamp 1515852544
transform 1 0 504 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_100
timestamp 1515852544
transform -1 0 648 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_637
timestamp 1515852544
transform -1 0 712 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_231
timestamp 1515852544
transform 1 0 712 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_643
timestamp 1515852544
transform 1 0 760 0 1 3810
box 0 0 64 200
use FILL  FILL_19_0_0
timestamp 1515852544
transform 1 0 824 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_1
timestamp 1515852544
transform 1 0 840 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_642
timestamp 1515852544
transform 1 0 856 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_230
timestamp 1515852544
transform -1 0 968 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_644
timestamp 1515852544
transform 1 0 968 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_102
timestamp 1515852544
transform -1 0 1112 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_641
timestamp 1515852544
transform -1 0 1176 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_127
timestamp 1515852544
transform -1 0 1256 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_632
timestamp 1515852544
transform 1 0 1256 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_220
timestamp 1515852544
transform -1 0 1384 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_221
timestamp 1515852544
transform 1 0 1384 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_133
timestamp 1515852544
transform -1 0 1512 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_114
timestamp 1515852544
transform -1 0 1592 0 1 3810
box 0 0 80 200
use BUFX4  BUFX4_9
timestamp 1515852544
transform -1 0 1656 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_8
timestamp 1515852544
transform -1 0 1704 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_89
timestamp 1515852544
transform -1 0 1768 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_7
timestamp 1515852544
transform -1 0 1832 0 1 3810
box 0 0 64 200
use FILL  FILL_19_1_0
timestamp 1515852544
transform 1 0 1832 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_1
timestamp 1515852544
transform 1 0 1848 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_450
timestamp 1515852544
transform 1 0 1864 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_448
timestamp 1515852544
transform -1 0 1992 0 1 3810
box 0 0 64 200
use INVX1  INVX1_49
timestamp 1515852544
transform 1 0 1992 0 1 3810
box 0 0 32 200
use NAND2X1  NAND2X1_145
timestamp 1515852544
transform 1 0 2024 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_439
timestamp 1515852544
transform -1 0 2136 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_24
timestamp 1515852544
transform -1 0 2200 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_113
timestamp 1515852544
transform 1 0 2200 0 1 3810
box 0 0 80 200
use AND2X2  AND2X2_23
timestamp 1515852544
transform 1 0 2280 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_182
timestamp 1515852544
transform 1 0 2344 0 1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_139
timestamp 1515852544
transform -1 0 2728 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_484
timestamp 1515852544
transform 1 0 2728 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_485
timestamp 1515852544
transform 1 0 2792 0 1 3810
box 0 0 64 200
use FILL  FILL_19_2_0
timestamp 1515852544
transform -1 0 2872 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_1
timestamp 1515852544
transform -1 0 2888 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_161
timestamp 1515852544
transform -1 0 2936 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_19
timestamp 1515852544
transform -1 0 3000 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_70
timestamp 1515852544
transform 1 0 3000 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_487
timestamp 1515852544
transform -1 0 3144 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_486
timestamp 1515852544
transform -1 0 3208 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_162
timestamp 1515852544
transform -1 0 3256 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_172
timestamp 1515852544
transform -1 0 3448 0 1 3810
box 0 0 192 200
use BUFX4  BUFX4_143
timestamp 1515852544
transform -1 0 3512 0 1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_12
timestamp 1515852544
transform 1 0 3512 0 1 3810
box 0 0 128 200
use BUFX4  BUFX4_219
timestamp 1515852544
transform -1 0 3704 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_240
timestamp 1515852544
transform 1 0 3704 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_146
timestamp 1515852544
transform -1 0 3816 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_179
timestamp 1515852544
transform -1 0 3880 0 1 3810
box 0 0 64 200
use FILL  FILL_19_3_0
timestamp 1515852544
transform 1 0 3880 0 1 3810
box 0 0 16 200
use FILL  FILL_19_3_1
timestamp 1515852544
transform 1 0 3896 0 1 3810
box 0 0 16 200
use AOI22X1  AOI22X1_120
timestamp 1515852544
transform 1 0 3912 0 1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_168
timestamp 1515852544
transform -1 0 4056 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_124
timestamp 1515852544
transform -1 0 4120 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_61
timestamp 1515852544
transform -1 0 4184 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_244
timestamp 1515852544
transform -1 0 4232 0 1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_243
timestamp 1515852544
transform 1 0 4232 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_201
timestamp 1515852544
transform -1 0 4344 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_550
timestamp 1515852544
transform 1 0 4344 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_549
timestamp 1515852544
transform -1 0 4472 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_191
timestamp 1515852544
transform -1 0 4520 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_36
timestamp 1515852544
transform 1 0 4520 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_192
timestamp 1515852544
transform -1 0 4632 0 1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_125
timestamp 1515852544
transform 1 0 4632 0 1 3810
box 0 0 80 200
use NAND2X1  NAND2X1_189
timestamp 1515852544
transform 1 0 4712 0 1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_210
timestamp 1515852544
transform 1 0 4760 0 1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_211
timestamp 1515852544
transform 1 0 4808 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_599
timestamp 1515852544
transform 1 0 4856 0 1 3810
box 0 0 64 200
use FILL  FILL_19_4_0
timestamp 1515852544
transform 1 0 4920 0 1 3810
box 0 0 16 200
use FILL  FILL_19_4_1
timestamp 1515852544
transform 1 0 4936 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_598
timestamp 1515852544
transform 1 0 4952 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_39
timestamp 1515852544
transform 1 0 5016 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_127
timestamp 1515852544
transform -1 0 5144 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_25
timestamp 1515852544
transform -1 0 5192 0 1 3810
box 0 0 48 200
use BUFX4  BUFX4_2
timestamp 1515852544
transform 1 0 5192 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_571
timestamp 1515852544
transform 1 0 5256 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_572
timestamp 1515852544
transform -1 0 5384 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_125
timestamp 1515852544
transform -1 0 5448 0 1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_86
timestamp 1515852544
transform 1 0 5448 0 1 3810
box 0 0 80 200
use INVX1  INVX1_84
timestamp 1515852544
transform 1 0 5528 0 1 3810
box 0 0 32 200
use AOI21X1  AOI21X1_48
timestamp 1515852544
transform -1 0 5624 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_379
timestamp 1515852544
transform 1 0 5624 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_180
timestamp 1515852544
transform -1 0 5880 0 1 3810
box 0 0 192 200
use BUFX4  BUFX4_140
timestamp 1515852544
transform 1 0 5880 0 1 3810
box 0 0 64 200
use FILL  FILL_19_5_0
timestamp 1515852544
transform -1 0 5960 0 1 3810
box 0 0 16 200
use FILL  FILL_19_5_1
timestamp 1515852544
transform -1 0 5976 0 1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_38
timestamp 1515852544
transform -1 0 6040 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_34
timestamp 1515852544
transform -1 0 6104 0 1 3810
box 0 0 64 200
use AOI21X1  AOI21X1_42
timestamp 1515852544
transform -1 0 6168 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_126
timestamp 1515852544
transform 1 0 6168 0 1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_125
timestamp 1515852544
transform -1 0 6552 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_614
timestamp 1515852544
transform -1 0 6616 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_564
timestamp 1515852544
transform -1 0 6680 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_17
timestamp 1515852544
transform 1 0 6680 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_53
timestamp 1515852544
transform 1 0 6728 0 1 3810
box 0 0 48 200
use FILL  FILL_20_1
timestamp 1515852544
transform 1 0 6776 0 1 3810
box 0 0 16 200
use FILL  FILL_20_2
timestamp 1515852544
transform 1 0 6792 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_142
timestamp 1515852544
transform 1 0 8 0 -1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_183
timestamp 1515852544
transform 1 0 200 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_536
timestamp 1515852544
transform 1 0 248 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_182
timestamp 1515852544
transform 1 0 312 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_535
timestamp 1515852544
transform -1 0 424 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_537
timestamp 1515852544
transform -1 0 488 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_619
timestamp 1515852544
transform -1 0 552 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_76
timestamp 1515852544
transform -1 0 616 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_73
timestamp 1515852544
transform 1 0 616 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_111
timestamp 1515852544
transform 1 0 680 0 -1 3810
box 0 0 192 200
use FILL  FILL_18_0_0
timestamp 1515852544
transform 1 0 872 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_1
timestamp 1515852544
transform 1 0 888 0 -1 3810
box 0 0 16 200
use NAND3X1  NAND3X1_44
timestamp 1515852544
transform 1 0 904 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_197
timestamp 1515852544
transform -1 0 1032 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_75
timestamp 1515852544
transform 1 0 1032 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_65
timestamp 1515852544
transform -1 0 1160 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_98
timestamp 1515852544
transform 1 0 1160 0 -1 3810
box 0 0 192 200
use XNOR2X1  XNOR2X1_1
timestamp 1515852544
transform -1 0 1464 0 -1 3810
box 0 0 112 200
use NAND2X1  NAND2X1_9
timestamp 1515852544
transform 1 0 1464 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_92
timestamp 1515852544
transform 1 0 1512 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_44
timestamp 1515852544
transform -1 0 1624 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_91
timestamp 1515852544
transform -1 0 1688 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_43
timestamp 1515852544
transform -1 0 1736 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_147
timestamp 1515852544
transform 1 0 1736 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_440
timestamp 1515852544
transform 1 0 1784 0 -1 3810
box 0 0 64 200
use FILL  FILL_18_1_0
timestamp 1515852544
transform 1 0 1848 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_1
timestamp 1515852544
transform 1 0 1864 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_441
timestamp 1515852544
transform 1 0 1880 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_61
timestamp 1515852544
transform -1 0 2024 0 -1 3810
box 0 0 80 200
use NAND3X1  NAND3X1_12
timestamp 1515852544
transform 1 0 2024 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_438
timestamp 1515852544
transform -1 0 2152 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_151
timestamp 1515852544
transform 1 0 2152 0 -1 3810
box 0 0 192 200
use AOI22X1  AOI22X1_107
timestamp 1515852544
transform 1 0 2344 0 -1 3810
box 0 0 80 200
use INVX1  INVX1_43
timestamp 1515852544
transform 1 0 2424 0 -1 3810
box 0 0 32 200
use NOR2X1  NOR2X1_25
timestamp 1515852544
transform 1 0 2456 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_54
timestamp 1515852544
transform 1 0 2504 0 -1 3810
box 0 0 32 200
use INVX1  INVX1_76
timestamp 1515852544
transform -1 0 2568 0 -1 3810
box 0 0 32 200
use OAI22X1  OAI22X1_12
timestamp 1515852544
transform 1 0 2568 0 -1 3810
box 0 0 80 200
use AOI22X1  AOI22X1_108
timestamp 1515852544
transform -1 0 2728 0 -1 3810
box 0 0 80 200
use INVX1  INVX1_98
timestamp 1515852544
transform 1 0 2728 0 -1 3810
box 0 0 32 200
use OAI22X1  OAI22X1_25
timestamp 1515852544
transform 1 0 2760 0 -1 3810
box 0 0 80 200
use INVX1  INVX1_87
timestamp 1515852544
transform -1 0 2872 0 -1 3810
box 0 0 32 200
use FILL  FILL_18_2_0
timestamp 1515852544
transform 1 0 2872 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_1
timestamp 1515852544
transform 1 0 2888 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_17
timestamp 1515852544
transform 1 0 2904 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_111
timestamp 1515852544
transform -1 0 3016 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_191
timestamp 1515852544
transform -1 0 3080 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_53
timestamp 1515852544
transform 1 0 3080 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_21
timestamp 1515852544
transform 1 0 3144 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_206
timestamp 1515852544
transform 1 0 3208 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_58
timestamp 1515852544
transform 1 0 3272 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_22
timestamp 1515852544
transform -1 0 3400 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_212
timestamp 1515852544
transform -1 0 3448 0 -1 3810
box 0 0 48 200
use NOR3X1  NOR3X1_13
timestamp 1515852544
transform 1 0 3448 0 -1 3810
box 0 0 128 200
use OAI21X1  OAI21X1_157
timestamp 1515852544
transform 1 0 3576 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_241
timestamp 1515852544
transform -1 0 3688 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_56
timestamp 1515852544
transform 1 0 3688 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_177
timestamp 1515852544
transform -1 0 3944 0 -1 3810
box 0 0 192 200
use FILL  FILL_18_3_0
timestamp 1515852544
transform 1 0 3944 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_1
timestamp 1515852544
transform 1 0 3960 0 -1 3810
box 0 0 16 200
use AOI22X1  AOI22X1_115
timestamp 1515852544
transform 1 0 3976 0 -1 3810
box 0 0 80 200
use NAND3X1  NAND3X1_53
timestamp 1515852544
transform 1 0 4056 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_43
timestamp 1515852544
transform 1 0 4120 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_89
timestamp 1515852544
transform 1 0 4184 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_62
timestamp 1515852544
transform 1 0 4248 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_133
timestamp 1515852544
transform -1 0 4504 0 -1 3810
box 0 0 192 200
use BUFX4  BUFX4_112
timestamp 1515852544
transform -1 0 4568 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_551
timestamp 1515852544
transform -1 0 4632 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_547
timestamp 1515852544
transform 1 0 4632 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_188
timestamp 1515852544
transform -1 0 4744 0 -1 3810
box 0 0 48 200
use BUFX4  BUFX4_190
timestamp 1515852544
transform 1 0 4744 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_209
timestamp 1515852544
transform -1 0 4856 0 -1 3810
box 0 0 48 200
use AOI22X1  AOI22X1_116
timestamp 1515852544
transform -1 0 4936 0 -1 3810
box 0 0 80 200
use FILL  FILL_18_4_0
timestamp 1515852544
transform -1 0 4952 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_4_1
timestamp 1515852544
transform -1 0 4968 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_597
timestamp 1515852544
transform -1 0 5032 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_157
timestamp 1515852544
transform 1 0 5032 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_17
timestamp 1515852544
transform -1 0 5160 0 -1 3810
box 0 0 64 200
use INVX8  INVX8_18
timestamp 1515852544
transform -1 0 5240 0 -1 3810
box 0 0 80 200
use BUFX4  BUFX4_104
timestamp 1515852544
transform -1 0 5304 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_10
timestamp 1515852544
transform 1 0 5304 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_570
timestamp 1515852544
transform -1 0 5432 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_573
timestamp 1515852544
transform 1 0 5432 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_105
timestamp 1515852544
transform 1 0 5496 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_137
timestamp 1515852544
transform -1 0 5752 0 -1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_178
timestamp 1515852544
transform -1 0 5944 0 -1 3810
box 0 0 192 200
use FILL  FILL_18_5_0
timestamp 1515852544
transform 1 0 5944 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_5_1
timestamp 1515852544
transform 1 0 5960 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_18
timestamp 1515852544
transform 1 0 5976 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_615
timestamp 1515852544
transform 1 0 6040 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_11
timestamp 1515852544
transform -1 0 6168 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_618
timestamp 1515852544
transform 1 0 6168 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_95
timestamp 1515852544
transform 1 0 6232 0 -1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_611
timestamp 1515852544
transform 1 0 6312 0 -1 3810
box 0 0 64 200
use AOI22X1  AOI22X1_94
timestamp 1515852544
transform -1 0 6456 0 -1 3810
box 0 0 80 200
use OAI21X1  OAI21X1_613
timestamp 1515852544
transform 1 0 6456 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_4
timestamp 1515852544
transform 1 0 6520 0 -1 3810
box 0 0 32 200
use AOI21X1  AOI21X1_41
timestamp 1515852544
transform -1 0 6616 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_57
timestamp 1515852544
transform -1 0 6664 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_15
timestamp 1515852544
transform -1 0 6696 0 -1 3810
box 0 0 32 200
use BUFX2  BUFX2_35
timestamp 1515852544
transform 1 0 6696 0 -1 3810
box 0 0 48 200
use BUFX2  BUFX2_38
timestamp 1515852544
transform 1 0 6744 0 -1 3810
box 0 0 48 200
use FILL  FILL_19_1
timestamp 1515852544
transform -1 0 6808 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_105
timestamp 1515852544
transform 1 0 8 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_218
timestamp 1515852544
transform 1 0 200 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_39
timestamp 1515852544
transform -1 0 312 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_219
timestamp 1515852544
transform 1 0 312 0 1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_96
timestamp 1515852544
transform 1 0 360 0 1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_622
timestamp 1515852544
transform 1 0 440 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_621
timestamp 1515852544
transform -1 0 568 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_620
timestamp 1515852544
transform -1 0 632 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_220
timestamp 1515852544
transform 1 0 632 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_625
timestamp 1515852544
transform -1 0 744 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_221
timestamp 1515852544
transform 1 0 744 0 1 3410
box 0 0 48 200
use FILL  FILL_17_0_0
timestamp 1515852544
transform -1 0 808 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_1
timestamp 1515852544
transform -1 0 824 0 1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_626
timestamp 1515852544
transform -1 0 888 0 1 3410
box 0 0 64 200
use INVX1  INVX1_27
timestamp 1515852544
transform -1 0 920 0 1 3410
box 0 0 32 200
use AOI22X1  AOI22X1_98
timestamp 1515852544
transform -1 0 1000 0 1 3410
box 0 0 80 200
use NAND3X1  NAND3X1_41
timestamp 1515852544
transform -1 0 1064 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_225
timestamp 1515852544
transform -1 0 1112 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_107
timestamp 1515852544
transform -1 0 1304 0 1 3410
box 0 0 192 200
use BUFX4  BUFX4_175
timestamp 1515852544
transform -1 0 1368 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_131
timestamp 1515852544
transform 1 0 1368 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_93
timestamp 1515852544
transform -1 0 1624 0 1 3410
box 0 0 64 200
use INVX2  INVX2_5
timestamp 1515852544
transform 1 0 1624 0 1 3410
box 0 0 32 200
use AND2X2  AND2X2_15
timestamp 1515852544
transform 1 0 1656 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_99
timestamp 1515852544
transform -1 0 1784 0 1 3410
box 0 0 64 200
use FILL  FILL_17_1_0
timestamp 1515852544
transform -1 0 1800 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_1
timestamp 1515852544
transform -1 0 1816 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_120
timestamp 1515852544
transform -1 0 2008 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_96
timestamp 1515852544
transform 1 0 2008 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_13
timestamp 1515852544
transform -1 0 2136 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_95
timestamp 1515852544
transform -1 0 2200 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_10
timestamp 1515852544
transform 1 0 2200 0 1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_4
timestamp 1515852544
transform 1 0 2248 0 1 3410
box 0 0 48 200
use BUFX4  BUFX4_224
timestamp 1515852544
transform -1 0 2360 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_98
timestamp 1515852544
transform -1 0 2424 0 1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_8
timestamp 1515852544
transform -1 0 2488 0 1 3410
box 0 0 64 200
use OAI22X1  OAI22X1_23
timestamp 1515852544
transform -1 0 2568 0 1 3410
box 0 0 80 200
use NOR2X1  NOR2X1_3
timestamp 1515852544
transform -1 0 2616 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_246
timestamp 1515852544
transform 1 0 2616 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_2
timestamp 1515852544
transform -1 0 2712 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_52
timestamp 1515852544
transform -1 0 2776 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_106
timestamp 1515852544
transform -1 0 2840 0 1 3410
box 0 0 64 200
use FILL  FILL_17_2_0
timestamp 1515852544
transform -1 0 2856 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_1
timestamp 1515852544
transform -1 0 2872 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_160
timestamp 1515852544
transform -1 0 2936 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_1
timestamp 1515852544
transform -1 0 2984 0 1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_26
timestamp 1515852544
transform 1 0 2984 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_50
timestamp 1515852544
transform -1 0 3096 0 1 3410
box 0 0 64 200
use BUFX2  BUFX2_19
timestamp 1515852544
transform -1 0 3144 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_99
timestamp 1515852544
transform 1 0 3144 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_16
timestamp 1515852544
transform 1 0 3208 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_110
timestamp 1515852544
transform -1 0 3320 0 1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_188
timestamp 1515852544
transform 1 0 3320 0 1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_114
timestamp 1515852544
transform -1 0 3464 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_116
timestamp 1515852544
transform -1 0 3656 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_576
timestamp 1515852544
transform 1 0 3656 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_198
timestamp 1515852544
transform 1 0 3720 0 1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_32
timestamp 1515852544
transform 1 0 3768 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_197
timestamp 1515852544
transform 1 0 3832 0 1 3410
box 0 0 48 200
use FILL  FILL_17_3_0
timestamp 1515852544
transform -1 0 3896 0 1 3410
box 0 0 16 200
use FILL  FILL_17_3_1
timestamp 1515852544
transform -1 0 3912 0 1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_575
timestamp 1515852544
transform -1 0 3976 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_176
timestamp 1515852544
transform 1 0 3976 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_199
timestamp 1515852544
transform 1 0 4168 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_580
timestamp 1515852544
transform -1 0 4280 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_390
timestamp 1515852544
transform 1 0 4280 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_117
timestamp 1515852544
transform 1 0 4344 0 1 3410
box 0 0 192 200
use BUFX4  BUFX4_173
timestamp 1515852544
transform -1 0 4600 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_42
timestamp 1515852544
transform -1 0 4664 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_162
timestamp 1515852544
transform 1 0 4664 0 1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_126
timestamp 1515852544
transform 1 0 4728 0 1 3410
box 0 0 80 200
use BUFX4  BUFX4_214
timestamp 1515852544
transform 1 0 4808 0 1 3410
box 0 0 64 200
use FILL  FILL_17_4_0
timestamp 1515852544
transform -1 0 4888 0 1 3410
box 0 0 16 200
use FILL  FILL_17_4_1
timestamp 1515852544
transform -1 0 4904 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_122
timestamp 1515852544
transform -1 0 5096 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_600
timestamp 1515852544
transform -1 0 5160 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_596
timestamp 1515852544
transform 1 0 5160 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_208
timestamp 1515852544
transform -1 0 5272 0 1 3410
box 0 0 48 200
use BUFX4  BUFX4_185
timestamp 1515852544
transform -1 0 5336 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_61
timestamp 1515852544
transform 1 0 5336 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_158
timestamp 1515852544
transform -1 0 5592 0 1 3410
box 0 0 192 200
use BUFX4  BUFX4_155
timestamp 1515852544
transform -1 0 5656 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_149
timestamp 1515852544
transform 1 0 5656 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_248
timestamp 1515852544
transform -1 0 5768 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_257
timestamp 1515852544
transform 1 0 5768 0 1 3410
box 0 0 64 200
use INVX1  INVX1_69
timestamp 1515852544
transform -1 0 5864 0 1 3410
box 0 0 32 200
use NAND3X1  NAND3X1_65
timestamp 1515852544
transform 1 0 5864 0 1 3410
box 0 0 64 200
use FILL  FILL_17_5_0
timestamp 1515852544
transform 1 0 5928 0 1 3410
box 0 0 16 200
use FILL  FILL_17_5_1
timestamp 1515852544
transform 1 0 5944 0 1 3410
box 0 0 16 200
use AOI22X1  AOI22X1_135
timestamp 1515852544
transform 1 0 5960 0 1 3410
box 0 0 80 200
use AOI22X1  AOI22X1_76
timestamp 1515852544
transform -1 0 6120 0 1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_517
timestamp 1515852544
transform -1 0 6184 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_617
timestamp 1515852544
transform 1 0 6184 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_616
timestamp 1515852544
transform -1 0 6312 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_181
timestamp 1515852544
transform 1 0 6312 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_519
timestamp 1515852544
transform 1 0 6376 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_134
timestamp 1515852544
transform 1 0 6440 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_217
timestamp 1515852544
transform -1 0 6680 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_196
timestamp 1515852544
transform 1 0 6680 0 1 3410
box 0 0 48 200
use AND2X2  AND2X2_37
timestamp 1515852544
transform 1 0 6728 0 1 3410
box 0 0 64 200
use FILL  FILL_18_1
timestamp 1515852544
transform 1 0 6792 0 1 3410
box 0 0 16 200
use NAND3X1  NAND3X1_20
timestamp 1515852544
transform -1 0 72 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_71
timestamp 1515852544
transform 1 0 72 0 -1 3410
box 0 0 80 200
use INVX1  INVX1_28
timestamp 1515852544
transform 1 0 152 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_488
timestamp 1515852544
transform -1 0 248 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_492
timestamp 1515852544
transform -1 0 312 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_97
timestamp 1515852544
transform 1 0 312 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_627
timestamp 1515852544
transform 1 0 392 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_40
timestamp 1515852544
transform -1 0 520 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_624
timestamp 1515852544
transform -1 0 584 0 -1 3410
box 0 0 64 200
use OAI22X1  OAI22X1_28
timestamp 1515852544
transform -1 0 664 0 -1 3410
box 0 0 80 200
use BUFX4  BUFX4_74
timestamp 1515852544
transform 1 0 664 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_629
timestamp 1515852544
transform 1 0 728 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_0_0
timestamp 1515852544
transform 1 0 792 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_1
timestamp 1515852544
transform 1 0 808 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_628
timestamp 1515852544
transform 1 0 824 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_631
timestamp 1515852544
transform 1 0 888 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_222
timestamp 1515852544
transform -1 0 1000 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_630
timestamp 1515852544
transform -1 0 1064 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_59
timestamp 1515852544
transform -1 0 1128 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_48
timestamp 1515852544
transform -1 0 1192 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_20
timestamp 1515852544
transform -1 0 1256 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_109
timestamp 1515852544
transform 1 0 1256 0 -1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_280
timestamp 1515852544
transform 1 0 1448 0 -1 3410
box 0 0 48 200
use OR2X2  OR2X2_12
timestamp 1515852544
transform -1 0 1560 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_14
timestamp 1515852544
transform -1 0 1624 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_97
timestamp 1515852544
transform -1 0 1688 0 -1 3410
box 0 0 64 200
use INVX4  INVX4_2
timestamp 1515852544
transform -1 0 1736 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_95
timestamp 1515852544
transform -1 0 1800 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_47
timestamp 1515852544
transform 1 0 1800 0 -1 3410
box 0 0 48 200
use FILL  FILL_16_1_0
timestamp 1515852544
transform 1 0 1848 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_1
timestamp 1515852544
transform 1 0 1864 0 -1 3410
box 0 0 16 200
use NOR2X1  NOR2X1_46
timestamp 1515852544
transform 1 0 1880 0 -1 3410
box 0 0 48 200
use INVX4  INVX4_1
timestamp 1515852544
transform -1 0 1976 0 -1 3410
box 0 0 48 200
use INVX4  INVX4_4
timestamp 1515852544
transform -1 0 2024 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_1
timestamp 1515852544
transform 1 0 2024 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_157
timestamp 1515852544
transform -1 0 2136 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_94
timestamp 1515852544
transform 1 0 2136 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_2
timestamp 1515852544
transform 1 0 2200 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_72
timestamp 1515852544
transform 1 0 2248 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_24
timestamp 1515852544
transform -1 0 2376 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_302
timestamp 1515852544
transform 1 0 2376 0 -1 3410
box 0 0 48 200
use NOR3X1  NOR3X1_7
timestamp 1515852544
transform -1 0 2552 0 -1 3410
box 0 0 128 200
use DFFPOSX1  DFFPOSX1_184
timestamp 1515852544
transform -1 0 2744 0 -1 3410
box 0 0 192 200
use BUFX4  BUFX4_138
timestamp 1515852544
transform -1 0 2808 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_2_0
timestamp 1515852544
transform 1 0 2808 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_1
timestamp 1515852544
transform 1 0 2824 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_118
timestamp 1515852544
transform 1 0 2840 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_109
timestamp 1515852544
transform 1 0 3032 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_583
timestamp 1515852544
transform -1 0 3160 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_1
timestamp 1515852544
transform -1 0 3224 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_574
timestamp 1515852544
transform 1 0 3224 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_87
timestamp 1515852544
transform 1 0 3288 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_577
timestamp 1515852544
transform -1 0 3432 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_151
timestamp 1515852544
transform 1 0 3432 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_239
timestamp 1515852544
transform 1 0 3496 0 -1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_88
timestamp 1515852544
transform 1 0 3544 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_582
timestamp 1515852544
transform 1 0 3624 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_581
timestamp 1515852544
transform 1 0 3688 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_200
timestamp 1515852544
transform -1 0 3800 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_33
timestamp 1515852544
transform 1 0 3800 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_3_0
timestamp 1515852544
transform -1 0 3880 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_3_1
timestamp 1515852544
transform -1 0 3896 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_578
timestamp 1515852544
transform -1 0 3960 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_152
timestamp 1515852544
transform 1 0 3960 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_155
timestamp 1515852544
transform 1 0 4008 0 -1 3410
box 0 0 192 200
use NAND3X1  NAND3X1_16
timestamp 1515852544
transform -1 0 4264 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_64
timestamp 1515852544
transform 1 0 4264 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_455
timestamp 1515852544
transform -1 0 4408 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_153
timestamp 1515852544
transform 1 0 4408 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_454
timestamp 1515852544
transform -1 0 4520 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_452
timestamp 1515852544
transform -1 0 4584 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_58
timestamp 1515852544
transform 1 0 4584 0 -1 3410
box 0 0 64 200
use OAI22X1  OAI22X1_22
timestamp 1515852544
transform 1 0 4648 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_467
timestamp 1515852544
transform 1 0 4728 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_82
timestamp 1515852544
transform -1 0 4824 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_470
timestamp 1515852544
transform 1 0 4824 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_4_0
timestamp 1515852544
transform -1 0 4904 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_4_1
timestamp 1515852544
transform -1 0 4920 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_469
timestamp 1515852544
transform -1 0 4984 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_471
timestamp 1515852544
transform 1 0 4984 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_66
timestamp 1515852544
transform -1 0 5128 0 -1 3410
box 0 0 80 200
use OAI21X1  OAI21X1_473
timestamp 1515852544
transform 1 0 5128 0 -1 3410
box 0 0 64 200
use AOI22X1  AOI22X1_129
timestamp 1515852544
transform 1 0 5192 0 -1 3410
box 0 0 80 200
use BUFX4  BUFX4_121
timestamp 1515852544
transform -1 0 5336 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_19
timestamp 1515852544
transform -1 0 5400 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_142
timestamp 1515852544
transform -1 0 5464 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_123
timestamp 1515852544
transform 1 0 5464 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_45
timestamp 1515852544
transform -1 0 5592 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_70
timestamp 1515852544
transform -1 0 5656 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_235
timestamp 1515852544
transform 1 0 5656 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_43
timestamp 1515852544
transform 1 0 5720 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_252
timestamp 1515852544
transform -1 0 5832 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_250
timestamp 1515852544
transform 1 0 5832 0 -1 3410
box 0 0 48 200
use AOI22X1  AOI22X1_145
timestamp 1515852544
transform -1 0 5960 0 -1 3410
box 0 0 80 200
use FILL  FILL_16_5_0
timestamp 1515852544
transform -1 0 5976 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_5_1
timestamp 1515852544
transform -1 0 5992 0 -1 3410
box 0 0 16 200
use NOR2X1  NOR2X1_23
timestamp 1515852544
transform -1 0 6040 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_516
timestamp 1515852544
transform 1 0 6040 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_117
timestamp 1515852544
transform 1 0 6104 0 -1 3410
box 0 0 32 200
use AOI21X1  AOI21X1_35
timestamp 1515852544
transform -1 0 6200 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_608
timestamp 1515852544
transform 1 0 6200 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_40
timestamp 1515852544
transform 1 0 6264 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_607
timestamp 1515852544
transform 1 0 6328 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_609
timestamp 1515852544
transform -1 0 6456 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_39
timestamp 1515852544
transform -1 0 6520 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_561
timestamp 1515852544
transform 1 0 6520 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_37
timestamp 1515852544
transform 1 0 6584 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_560
timestamp 1515852544
transform 1 0 6648 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_562
timestamp 1515852544
transform 1 0 6712 0 -1 3410
box 0 0 64 200
use FILL  FILL_17_1
timestamp 1515852544
transform -1 0 6792 0 -1 3410
box 0 0 16 200
use FILL  FILL_17_2
timestamp 1515852544
transform -1 0 6808 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_140
timestamp 1515852544
transform 1 0 8 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_163
timestamp 1515852544
transform 1 0 200 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_489
timestamp 1515852544
transform -1 0 312 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_164
timestamp 1515852544
transform 1 0 312 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_491
timestamp 1515852544
transform -1 0 424 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_106
timestamp 1515852544
transform 1 0 424 0 1 3010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1515852544
transform 1 0 616 0 1 3010
box 0 0 192 200
use FILL  FILL_15_0_0
timestamp 1515852544
transform 1 0 808 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_1
timestamp 1515852544
transform 1 0 824 0 1 3010
box 0 0 16 200
use AOI22X1  AOI22X1_33
timestamp 1515852544
transform 1 0 840 0 1 3010
box 0 0 80 200
use NAND3X1  NAND3X1_128
timestamp 1515852544
transform -1 0 984 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_89
timestamp 1515852544
transform 1 0 984 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_91
timestamp 1515852544
transform 1 0 1032 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_300
timestamp 1515852544
transform -1 0 1144 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_299
timestamp 1515852544
transform -1 0 1208 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_302
timestamp 1515852544
transform -1 0 1272 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_298
timestamp 1515852544
transform -1 0 1336 0 1 3010
box 0 0 64 200
use INVX1  INVX1_26
timestamp 1515852544
transform 1 0 1336 0 1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_14
timestamp 1515852544
transform 1 0 1368 0 1 3010
box 0 0 48 200
use OR2X2  OR2X2_1
timestamp 1515852544
transform 1 0 1416 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_41
timestamp 1515852544
transform -1 0 1544 0 1 3010
box 0 0 64 200
use NOR3X1  NOR3X1_11
timestamp 1515852544
transform -1 0 1672 0 1 3010
box 0 0 128 200
use BUFX4  BUFX4_136
timestamp 1515852544
transform 1 0 1672 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_1
timestamp 1515852544
transform 1 0 1736 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_13
timestamp 1515852544
transform 1 0 1800 0 1 3010
box 0 0 48 200
use FILL  FILL_15_1_0
timestamp 1515852544
transform -1 0 1864 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_1
timestamp 1515852544
transform -1 0 1880 0 1 3010
box 0 0 16 200
use NAND3X1  NAND3X1_2
timestamp 1515852544
transform -1 0 1944 0 1 3010
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1515852544
transform -1 0 2072 0 1 3010
box 0 0 128 200
use NAND2X1  NAND2X1_269
timestamp 1515852544
transform 1 0 2072 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_556
timestamp 1515852544
transform -1 0 2184 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_101
timestamp 1515852544
transform 1 0 2184 0 1 3010
box 0 0 48 200
use NOR3X1  NOR3X1_9
timestamp 1515852544
transform -1 0 2360 0 1 3010
box 0 0 128 200
use NOR3X1  NOR3X1_8
timestamp 1515852544
transform -1 0 2488 0 1 3010
box 0 0 128 200
use OAI22X1  OAI22X1_30
timestamp 1515852544
transform 1 0 2488 0 1 3010
box 0 0 80 200
use INVX1  INVX1_33
timestamp 1515852544
transform -1 0 2600 0 1 3010
box 0 0 32 200
use INVX1  INVX1_31
timestamp 1515852544
transform -1 0 2632 0 1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_101
timestamp 1515852544
transform -1 0 2712 0 1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_586
timestamp 1515852544
transform 1 0 2712 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_89
timestamp 1515852544
transform -1 0 2856 0 1 3010
box 0 0 80 200
use FILL  FILL_15_2_0
timestamp 1515852544
transform -1 0 2872 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_1
timestamp 1515852544
transform -1 0 2888 0 1 3010
box 0 0 16 200
use NAND3X1  NAND3X1_34
timestamp 1515852544
transform -1 0 2952 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_203
timestamp 1515852544
transform 1 0 2952 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_585
timestamp 1515852544
transform -1 0 3064 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_202
timestamp 1515852544
transform 1 0 3064 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_584
timestamp 1515852544
transform -1 0 3176 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_657
timestamp 1515852544
transform 1 0 3176 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_655
timestamp 1515852544
transform 1 0 3240 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_663
timestamp 1515852544
transform 1 0 3304 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_664
timestamp 1515852544
transform 1 0 3368 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_105
timestamp 1515852544
transform 1 0 3432 0 1 3010
box 0 0 80 200
use INVX1  INVX1_83
timestamp 1515852544
transform -1 0 3544 0 1 3010
box 0 0 32 200
use BUFX4  BUFX4_134
timestamp 1515852544
transform -1 0 3608 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_44
timestamp 1515852544
transform -1 0 3672 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_218
timestamp 1515852544
transform -1 0 3736 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_225
timestamp 1515852544
transform 1 0 3736 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_168
timestamp 1515852544
transform 1 0 3800 0 1 3010
box 0 0 64 200
use FILL  FILL_15_3_0
timestamp 1515852544
transform 1 0 3864 0 1 3010
box 0 0 16 200
use FILL  FILL_15_3_1
timestamp 1515852544
transform 1 0 3880 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_44
timestamp 1515852544
transform 1 0 3896 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_453
timestamp 1515852544
transform 1 0 3960 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_37
timestamp 1515852544
transform 1 0 4024 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_132
timestamp 1515852544
transform 1 0 4088 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_159
timestamp 1515852544
transform 1 0 4152 0 1 3010
box 0 0 192 200
use BUFX4  BUFX4_223
timestamp 1515852544
transform 1 0 4344 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_32
timestamp 1515852544
transform 1 0 4408 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_476
timestamp 1515852544
transform -1 0 4520 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_477
timestamp 1515852544
transform -1 0 4584 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_4
timestamp 1515852544
transform -1 0 4648 0 1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_67
timestamp 1515852544
transform 1 0 4648 0 1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_478
timestamp 1515852544
transform -1 0 4792 0 1 3010
box 0 0 64 200
use NOR3X1  NOR3X1_3
timestamp 1515852544
transform -1 0 4920 0 1 3010
box 0 0 128 200
use FILL  FILL_15_4_0
timestamp 1515852544
transform 1 0 4920 0 1 3010
box 0 0 16 200
use FILL  FILL_15_4_1
timestamp 1515852544
transform 1 0 4936 0 1 3010
box 0 0 16 200
use INVX1  INVX1_115
timestamp 1515852544
transform 1 0 4952 0 1 3010
box 0 0 32 200
use AOI21X1  AOI21X1_12
timestamp 1515852544
transform 1 0 4984 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_246
timestamp 1515852544
transform -1 0 5112 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_183
timestamp 1515852544
transform -1 0 5176 0 1 3010
box 0 0 64 200
use INVX2  INVX2_1
timestamp 1515852544
transform -1 0 5208 0 1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_68
timestamp 1515852544
transform -1 0 5272 0 1 3010
box 0 0 64 200
use INVX1  INVX1_73
timestamp 1515852544
transform 1 0 5272 0 1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_15
timestamp 1515852544
transform 1 0 5304 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_275
timestamp 1515852544
transform 1 0 5352 0 1 3010
box 0 0 48 200
use AND2X2  AND2X2_6
timestamp 1515852544
transform 1 0 5400 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_673
timestamp 1515852544
transform 1 0 5464 0 1 3010
box 0 0 64 200
use INVX1  INVX1_91
timestamp 1515852544
transform -1 0 5560 0 1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_132
timestamp 1515852544
transform 1 0 5560 0 1 3010
box 0 0 80 200
use AND2X2  AND2X2_36
timestamp 1515852544
transform 1 0 5640 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_251
timestamp 1515852544
transform 1 0 5704 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_249
timestamp 1515852544
transform -1 0 5800 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_553
timestamp 1515852544
transform -1 0 5864 0 1 3010
box 0 0 64 200
use INVX1  INVX1_119
timestamp 1515852544
transform -1 0 5896 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_552
timestamp 1515852544
transform 1 0 5896 0 1 3010
box 0 0 64 200
use FILL  FILL_15_5_0
timestamp 1515852544
transform -1 0 5976 0 1 3010
box 0 0 16 200
use FILL  FILL_15_5_1
timestamp 1515852544
transform -1 0 5992 0 1 3010
box 0 0 16 200
use NAND3X1  NAND3X1_31
timestamp 1515852544
transform -1 0 6056 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_193
timestamp 1515852544
transform -1 0 6104 0 1 3010
box 0 0 48 200
use BUFX4  BUFX4_182
timestamp 1515852544
transform 1 0 6104 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_122
timestamp 1515852544
transform 1 0 6168 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_610
timestamp 1515852544
transform 1 0 6232 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_124
timestamp 1515852544
transform 1 0 6296 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_563
timestamp 1515852544
transform 1 0 6488 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_135
timestamp 1515852544
transform 1 0 6552 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_195
timestamp 1515852544
transform -1 0 6792 0 1 3010
box 0 0 48 200
use FILL  FILL_16_1
timestamp 1515852544
transform 1 0 6792 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_43
timestamp 1515852544
transform 1 0 8 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_2
timestamp 1515852544
transform -1 0 232 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_57
timestamp 1515852544
transform 1 0 232 0 -1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_41
timestamp 1515852544
transform 1 0 280 0 -1 3010
box 0 0 80 200
use NAND3X1  NAND3X1_134
timestamp 1515852544
transform -1 0 424 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_344
timestamp 1515852544
transform 1 0 424 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_341
timestamp 1515852544
transform -1 0 552 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_342
timestamp 1515852544
transform -1 0 616 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_107
timestamp 1515852544
transform -1 0 664 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_120
timestamp 1515852544
transform -1 0 728 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_0_0
timestamp 1515852544
transform 1 0 728 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_1
timestamp 1515852544
transform 1 0 744 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_92
timestamp 1515852544
transform 1 0 760 0 -1 3010
box 0 0 192 200
use BUFX4  BUFX4_192
timestamp 1515852544
transform -1 0 1016 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_150
timestamp 1515852544
transform 1 0 1016 0 -1 3010
box 0 0 80 200
use AOI22X1  AOI22X1_35
timestamp 1515852544
transform 1 0 1096 0 -1 3010
box 0 0 80 200
use BUFX4  BUFX4_47
timestamp 1515852544
transform -1 0 1240 0 -1 3010
box 0 0 64 200
use NOR3X1  NOR3X1_6
timestamp 1515852544
transform -1 0 1368 0 -1 3010
box 0 0 128 200
use BUFX4  BUFX4_213
timestamp 1515852544
transform 1 0 1368 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_85
timestamp 1515852544
transform 1 0 1432 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_12
timestamp 1515852544
transform -1 0 1560 0 -1 3010
box 0 0 64 200
use INVX4  INVX4_3
timestamp 1515852544
transform -1 0 1608 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_96
timestamp 1515852544
transform 1 0 1608 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_112
timestamp 1515852544
transform -1 0 1720 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_44
timestamp 1515852544
transform 1 0 1720 0 -1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_129
timestamp 1515852544
transform -1 0 1816 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_17
timestamp 1515852544
transform -1 0 1864 0 -1 3010
box 0 0 48 200
use FILL  FILL_14_1_0
timestamp 1515852544
transform -1 0 1880 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_1
timestamp 1515852544
transform -1 0 1896 0 -1 3010
box 0 0 16 200
use NAND3X1  NAND3X1_35
timestamp 1515852544
transform -1 0 1960 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_19
timestamp 1515852544
transform -1 0 2008 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_47
timestamp 1515852544
transform -1 0 2072 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_14
timestamp 1515852544
transform -1 0 2136 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_13
timestamp 1515852544
transform -1 0 2184 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_90
timestamp 1515852544
transform -1 0 2232 0 -1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_46
timestamp 1515852544
transform -1 0 2312 0 -1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_24
timestamp 1515852544
transform 1 0 2312 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_55
timestamp 1515852544
transform -1 0 2424 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_468
timestamp 1515852544
transform 1 0 2424 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_262
timestamp 1515852544
transform -1 0 2536 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_479
timestamp 1515852544
transform 1 0 2536 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_263
timestamp 1515852544
transform -1 0 2648 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_72
timestamp 1515852544
transform 1 0 2648 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_53
timestamp 1515852544
transform 1 0 2712 0 -1 3010
box 0 0 192 200
use FILL  FILL_14_2_0
timestamp 1515852544
transform 1 0 2904 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_1
timestamp 1515852544
transform 1 0 2920 0 -1 3010
box 0 0 16 200
use OAI22X1  OAI22X1_4
timestamp 1515852544
transform 1 0 2936 0 -1 3010
box 0 0 80 200
use INVX1  INVX1_39
timestamp 1515852544
transform -1 0 3048 0 -1 3010
box 0 0 32 200
use INVX1  INVX1_38
timestamp 1515852544
transform -1 0 3080 0 -1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_183
timestamp 1515852544
transform -1 0 3160 0 -1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_659
timestamp 1515852544
transform 1 0 3160 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_658
timestamp 1515852544
transform 1 0 3224 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_661
timestamp 1515852544
transform 1 0 3288 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_85
timestamp 1515852544
transform 1 0 3352 0 -1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_104
timestamp 1515852544
transform 1 0 3384 0 -1 3010
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_115
timestamp 1515852544
transform -1 0 3656 0 -1 3010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_54
timestamp 1515852544
transform -1 0 3848 0 -1 3010
box 0 0 192 200
use FILL  FILL_14_3_0
timestamp 1515852544
transform -1 0 3864 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_3_1
timestamp 1515852544
transform -1 0 3880 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_59
timestamp 1515852544
transform -1 0 4072 0 -1 3010
box 0 0 192 200
use NOR2X1  NOR2X1_31
timestamp 1515852544
transform -1 0 4120 0 -1 3010
box 0 0 48 200
use OR2X2  OR2X2_18
timestamp 1515852544
transform 1 0 4120 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_58
timestamp 1515852544
transform -1 0 4376 0 -1 3010
box 0 0 192 200
use BUFX4  BUFX4_31
timestamp 1515852544
transform -1 0 4440 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_89
timestamp 1515852544
transform 1 0 4440 0 -1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_5
timestamp 1515852544
transform 1 0 4472 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_474
timestamp 1515852544
transform -1 0 4584 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_153
timestamp 1515852544
transform 1 0 4584 0 -1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_475
timestamp 1515852544
transform -1 0 4728 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_190
timestamp 1515852544
transform 1 0 4728 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_60
timestamp 1515852544
transform -1 0 4856 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_135
timestamp 1515852544
transform 1 0 4856 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_4_0
timestamp 1515852544
transform 1 0 4920 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_4_1
timestamp 1515852544
transform 1 0 4936 0 -1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_1
timestamp 1515852544
transform 1 0 4952 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_59
timestamp 1515852544
transform 1 0 5016 0 -1 3010
box 0 0 32 200
use NAND3X1  NAND3X1_59
timestamp 1515852544
transform -1 0 5112 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_35
timestamp 1515852544
transform 1 0 5112 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_279
timestamp 1515852544
transform 1 0 5176 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_254
timestamp 1515852544
transform 1 0 5240 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_60
timestamp 1515852544
transform -1 0 5480 0 -1 3010
box 0 0 192 200
use NAND3X1  NAND3X1_79
timestamp 1515852544
transform 1 0 5480 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_278
timestamp 1515852544
transform 1 0 5544 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_279
timestamp 1515852544
transform -1 0 5640 0 -1 3010
box 0 0 48 200
use AOI22X1  AOI22X1_163
timestamp 1515852544
transform -1 0 5720 0 -1 3010
box 0 0 80 200
use NAND2X1  NAND2X1_277
timestamp 1515852544
transform 1 0 5720 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_276
timestamp 1515852544
transform -1 0 5816 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_118
timestamp 1515852544
transform -1 0 5848 0 -1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_194
timestamp 1515852544
transform 1 0 5848 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_555
timestamp 1515852544
transform -1 0 5960 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_5_0
timestamp 1515852544
transform -1 0 5976 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_5_1
timestamp 1515852544
transform -1 0 5992 0 -1 3010
box 0 0 16 200
use INVX1  INVX1_60
timestamp 1515852544
transform -1 0 6024 0 -1 3010
box 0 0 32 200
use AOI22X1  AOI22X1_84
timestamp 1515852544
transform -1 0 6104 0 -1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_554
timestamp 1515852544
transform -1 0 6168 0 -1 3010
box 0 0 64 200
use INVX8  INVX8_7
timestamp 1515852544
transform 1 0 6168 0 -1 3010
box 0 0 80 200
use OAI21X1  OAI21X1_606
timestamp 1515852544
transform 1 0 6248 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_605
timestamp 1515852544
transform -1 0 6376 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_216
timestamp 1515852544
transform 1 0 6376 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_558
timestamp 1515852544
transform 1 0 6424 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_559
timestamp 1515852544
transform -1 0 6552 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_312
timestamp 1515852544
transform 1 0 6552 0 -1 3010
box 0 0 64 200
use AOI22X1  AOI22X1_140
timestamp 1515852544
transform -1 0 6696 0 -1 3010
box 0 0 80 200
use BUFX2  BUFX2_15
timestamp 1515852544
transform 1 0 6696 0 -1 3010
box 0 0 48 200
use BUFX2  BUFX2_51
timestamp 1515852544
transform 1 0 6744 0 -1 3010
box 0 0 48 200
use FILL  FILL_15_1
timestamp 1515852544
transform -1 0 6808 0 -1 3010
box 0 0 16 200
use BUFX2  BUFX2_46
timestamp 1515852544
transform -1 0 56 0 1 2610
box 0 0 48 200
use BUFX2  BUFX2_9
timestamp 1515852544
transform -1 0 104 0 1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_105
timestamp 1515852544
transform 1 0 104 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_88
timestamp 1515852544
transform 1 0 168 0 1 2610
box 0 0 192 200
use AOI22X1  AOI22X1_5
timestamp 1515852544
transform 1 0 360 0 1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_162
timestamp 1515852544
transform -1 0 504 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_45
timestamp 1515852544
transform 1 0 504 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_352
timestamp 1515852544
transform 1 0 696 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_114
timestamp 1515852544
transform -1 0 808 0 1 2610
box 0 0 48 200
use FILL  FILL_13_0_0
timestamp 1515852544
transform 1 0 808 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_1
timestamp 1515852544
transform 1 0 824 0 1 2610
box 0 0 16 200
use NAND3X1  NAND3X1_136
timestamp 1515852544
transform 1 0 840 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_43
timestamp 1515852544
transform 1 0 904 0 1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_353
timestamp 1515852544
transform -1 0 1048 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_111
timestamp 1515852544
transform 1 0 1048 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_351
timestamp 1515852544
transform -1 0 1160 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_44
timestamp 1515852544
transform 1 0 1160 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_174
timestamp 1515852544
transform -1 0 1272 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_109
timestamp 1515852544
transform 1 0 1272 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_43
timestamp 1515852544
transform -1 0 1384 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_173
timestamp 1515852544
transform -1 0 1448 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_175
timestamp 1515852544
transform 1 0 1448 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_8
timestamp 1515852544
transform -1 0 1592 0 1 2610
box 0 0 80 200
use BUFX4  BUFX4_171
timestamp 1515852544
transform 1 0 1592 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_292
timestamp 1515852544
transform 1 0 1656 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_86
timestamp 1515852544
transform -1 0 1768 0 1 2610
box 0 0 48 200
use BUFX4  BUFX4_90
timestamp 1515852544
transform -1 0 1832 0 1 2610
box 0 0 64 200
use FILL  FILL_13_1_0
timestamp 1515852544
transform 1 0 1832 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_1
timestamp 1515852544
transform 1 0 1848 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_179
timestamp 1515852544
transform 1 0 1864 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_24
timestamp 1515852544
transform -1 0 1976 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_63
timestamp 1515852544
transform 1 0 1976 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_223
timestamp 1515852544
transform -1 0 2088 0 1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_118
timestamp 1515852544
transform -1 0 2152 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_146
timestamp 1515852544
transform 1 0 2152 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_258
timestamp 1515852544
transform 1 0 2200 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_168
timestamp 1515852544
transform -1 0 2296 0 1 2610
box 0 0 48 200
use OR2X2  OR2X2_15
timestamp 1515852544
transform -1 0 2360 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_20
timestamp 1515852544
transform -1 0 2408 0 1 2610
box 0 0 48 200
use OR2X2  OR2X2_16
timestamp 1515852544
transform -1 0 2472 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_28
timestamp 1515852544
transform 1 0 2472 0 1 2610
box 0 0 48 200
use NOR3X1  NOR3X1_2
timestamp 1515852544
transform -1 0 2648 0 1 2610
box 0 0 128 200
use NOR2X1  NOR2X1_21
timestamp 1515852544
transform -1 0 2696 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_13
timestamp 1515852544
transform -1 0 2760 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_22
timestamp 1515852544
transform 1 0 2760 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_79
timestamp 1515852544
transform 1 0 2808 0 1 2610
box 0 0 64 200
use FILL  FILL_13_2_0
timestamp 1515852544
transform 1 0 2872 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_1
timestamp 1515852544
transform 1 0 2888 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_457
timestamp 1515852544
transform 1 0 2904 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_17
timestamp 1515852544
transform 1 0 2968 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_68
timestamp 1515852544
transform -1 0 3080 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_490
timestamp 1515852544
transform -1 0 3144 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_156
timestamp 1515852544
transform -1 0 3224 0 1 2610
box 0 0 80 200
use AOI22X1  AOI22X1_106
timestamp 1515852544
transform 1 0 3224 0 1 2610
box 0 0 80 200
use BUFX4  BUFX4_84
timestamp 1515852544
transform -1 0 3368 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_660
timestamp 1515852544
transform 1 0 3368 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_114
timestamp 1515852544
transform 1 0 3432 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_665
timestamp 1515852544
transform -1 0 3688 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_662
timestamp 1515852544
transform -1 0 3752 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_73
timestamp 1515852544
transform -1 0 3816 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_122
timestamp 1515852544
transform -1 0 3896 0 1 2610
box 0 0 80 200
use FILL  FILL_13_3_0
timestamp 1515852544
transform 1 0 3896 0 1 2610
box 0 0 16 200
use FILL  FILL_13_3_1
timestamp 1515852544
transform 1 0 3912 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_85
timestamp 1515852544
transform 1 0 3928 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_78
timestamp 1515852544
transform -1 0 4056 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_671
timestamp 1515852544
transform 1 0 4056 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_162
timestamp 1515852544
transform -1 0 4200 0 1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_668
timestamp 1515852544
transform -1 0 4264 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_154
timestamp 1515852544
transform 1 0 4264 0 1 2610
box 0 0 80 200
use AOI22X1  AOI22X1_160
timestamp 1515852544
transform -1 0 4424 0 1 2610
box 0 0 80 200
use NAND3X1  NAND3X1_77
timestamp 1515852544
transform 1 0 4424 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_5
timestamp 1515852544
transform -1 0 4552 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_3
timestamp 1515852544
transform -1 0 4616 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_15
timestamp 1515852544
transform -1 0 4680 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_63
timestamp 1515852544
transform 1 0 4680 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_472
timestamp 1515852544
transform 1 0 4872 0 1 2610
box 0 0 64 200
use FILL  FILL_13_4_0
timestamp 1515852544
transform 1 0 4936 0 1 2610
box 0 0 16 200
use FILL  FILL_13_4_1
timestamp 1515852544
transform 1 0 4952 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_604
timestamp 1515852544
transform 1 0 4968 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_93
timestamp 1515852544
transform 1 0 5032 0 1 2610
box 0 0 80 200
use NAND2X1  NAND2X1_215
timestamp 1515852544
transform 1 0 5112 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_214
timestamp 1515852544
transform -1 0 5208 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_38
timestamp 1515852544
transform -1 0 5272 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_401
timestamp 1515852544
transform 1 0 5272 0 1 2610
box 0 0 64 200
use INVX1  INVX1_90
timestamp 1515852544
transform 1 0 5336 0 1 2610
box 0 0 32 200
use NAND3X1  NAND3X1_71
timestamp 1515852544
transform -1 0 5432 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_50
timestamp 1515852544
transform 1 0 5432 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_41
timestamp 1515852544
transform 1 0 5496 0 1 2610
box 0 0 48 200
use INVX2  INVX2_2
timestamp 1515852544
transform 1 0 5544 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_672
timestamp 1515852544
transform -1 0 5640 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_16
timestamp 1515852544
transform 1 0 5640 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_357
timestamp 1515852544
transform 1 0 5704 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_47
timestamp 1515852544
transform -1 0 5832 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_518
timestamp 1515852544
transform -1 0 5896 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_141
timestamp 1515852544
transform 1 0 5896 0 1 2610
box 0 0 64 200
use FILL  FILL_13_5_0
timestamp 1515852544
transform 1 0 5960 0 1 2610
box 0 0 16 200
use FILL  FILL_13_5_1
timestamp 1515852544
transform 1 0 5976 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_462
timestamp 1515852544
transform 1 0 5992 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_676
timestamp 1515852544
transform 1 0 6056 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_461
timestamp 1515852544
transform -1 0 6184 0 1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_149
timestamp 1515852544
transform -1 0 6264 0 1 2610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_61
timestamp 1515852544
transform -1 0 6456 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_679
timestamp 1515852544
transform 1 0 6456 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_7
timestamp 1515852544
transform 1 0 6520 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_678
timestamp 1515852544
transform 1 0 6584 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_42
timestamp 1515852544
transform -1 0 6696 0 1 2610
box 0 0 48 200
use AOI21X1  AOI21X1_2
timestamp 1515852544
transform 1 0 6696 0 1 2610
box 0 0 64 200
use FILL  FILL_14_1
timestamp 1515852544
transform 1 0 6760 0 1 2610
box 0 0 16 200
use FILL  FILL_14_2
timestamp 1515852544
transform 1 0 6776 0 1 2610
box 0 0 16 200
use FILL  FILL_14_3
timestamp 1515852544
transform 1 0 6792 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_37
timestamp 1515852544
transform 1 0 8 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_38
timestamp 1515852544
transform 1 0 56 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_161
timestamp 1515852544
transform -1 0 168 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_160
timestamp 1515852544
transform -1 0 232 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_42
timestamp 1515852544
transform 1 0 232 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_159
timestamp 1515852544
transform -1 0 488 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_108
timestamp 1515852544
transform 1 0 488 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_343
timestamp 1515852544
transform -1 0 600 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_119
timestamp 1515852544
transform -1 0 664 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_350
timestamp 1515852544
transform 1 0 664 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_154
timestamp 1515852544
transform 1 0 728 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_0_0
timestamp 1515852544
transform -1 0 808 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_1
timestamp 1515852544
transform -1 0 824 0 -1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_156
timestamp 1515852544
transform -1 0 888 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_26
timestamp 1515852544
transform -1 0 952 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_36
timestamp 1515852544
transform -1 0 1000 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_193
timestamp 1515852544
transform 1 0 1000 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_146
timestamp 1515852544
transform -1 0 1128 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_172
timestamp 1515852544
transform 1 0 1128 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_85
timestamp 1515852544
transform 1 0 1192 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_126
timestamp 1515852544
transform -1 0 1304 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_173
timestamp 1515852544
transform 1 0 1304 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_35
timestamp 1515852544
transform 1 0 1496 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_201
timestamp 1515852544
transform -1 0 1608 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_48
timestamp 1515852544
transform 1 0 1608 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_109
timestamp 1515852544
transform 1 0 1672 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_46
timestamp 1515852544
transform -1 0 1816 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_1_0
timestamp 1515852544
transform 1 0 1816 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_1
timestamp 1515852544
transform 1 0 1832 0 -1 2610
box 0 0 16 200
use AOI22X1  AOI22X1_90
timestamp 1515852544
transform 1 0 1848 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_2
timestamp 1515852544
transform -1 0 1992 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_38
timestamp 1515852544
transform -1 0 2056 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_114
timestamp 1515852544
transform 1 0 2056 0 -1 2610
box 0 0 64 200
use OAI22X1  OAI22X1_6
timestamp 1515852544
transform 1 0 2120 0 -1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_10
timestamp 1515852544
transform -1 0 2248 0 -1 2610
box 0 0 48 200
use NOR3X1  NOR3X1_10
timestamp 1515852544
transform -1 0 2376 0 -1 2610
box 0 0 128 200
use OR2X2  OR2X2_13
timestamp 1515852544
transform 1 0 2376 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_270
timestamp 1515852544
transform 1 0 2440 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_76
timestamp 1515852544
transform 1 0 2488 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_268
timestamp 1515852544
transform 1 0 2552 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_612
timestamp 1515852544
transform 1 0 2600 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_601
timestamp 1515852544
transform -1 0 2728 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_590
timestamp 1515852544
transform -1 0 2792 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_623
timestamp 1515852544
transform -1 0 2856 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_2_0
timestamp 1515852544
transform -1 0 2872 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_1
timestamp 1515852544
transform -1 0 2888 0 -1 2610
box 0 0 16 200
use AOI22X1  AOI22X1_159
timestamp 1515852544
transform -1 0 2968 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_429
timestamp 1515852544
transform 1 0 2968 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_59
timestamp 1515852544
transform 1 0 3032 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_432
timestamp 1515852544
transform -1 0 3176 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_10
timestamp 1515852544
transform -1 0 3240 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_141
timestamp 1515852544
transform 1 0 3240 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_430
timestamp 1515852544
transform -1 0 3352 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_431
timestamp 1515852544
transform -1 0 3416 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_142
timestamp 1515852544
transform -1 0 3464 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_534
timestamp 1515852544
transform -1 0 3528 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_157
timestamp 1515852544
transform -1 0 3608 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_512
timestamp 1515852544
transform 1 0 3608 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_523
timestamp 1515852544
transform -1 0 3736 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_264
timestamp 1515852544
transform -1 0 3784 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_265
timestamp 1515852544
transform -1 0 3832 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_273
timestamp 1515852544
transform 1 0 3832 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_3_0
timestamp 1515852544
transform 1 0 3880 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_3_1
timestamp 1515852544
transform 1 0 3896 0 -1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_669
timestamp 1515852544
transform 1 0 3912 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_83
timestamp 1515852544
transform 1 0 3976 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_274
timestamp 1515852544
transform 1 0 4040 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_670
timestamp 1515852544
transform -1 0 4152 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_667
timestamp 1515852544
transform 1 0 4152 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_634
timestamp 1515852544
transform 1 0 4216 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_656
timestamp 1515852544
transform 1 0 4280 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_272
timestamp 1515852544
transform 1 0 4344 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_645
timestamp 1515852544
transform -1 0 4456 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_271
timestamp 1515852544
transform -1 0 4504 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_686
timestamp 1515852544
transform 1 0 4504 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_42
timestamp 1515852544
transform 1 0 4568 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_34
timestamp 1515852544
transform -1 0 4680 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_690
timestamp 1515852544
transform 1 0 4680 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_153
timestamp 1515852544
transform -1 0 4808 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_602
timestamp 1515852544
transform 1 0 4808 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_213
timestamp 1515852544
transform 1 0 4872 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_4_0
timestamp 1515852544
transform 1 0 4920 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_4_1
timestamp 1515852544
transform 1 0 4936 0 -1 2610
box 0 0 16 200
use NAND3X1  NAND3X1_38
timestamp 1515852544
transform 1 0 4952 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_603
timestamp 1515852544
transform -1 0 5080 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_3
timestamp 1515852544
transform -1 0 5112 0 -1 2610
box 0 0 32 200
use NOR3X1  NOR3X1_4
timestamp 1515852544
transform -1 0 5240 0 -1 2610
box 0 0 128 200
use NAND2X1  NAND2X1_155
timestamp 1515852544
transform 1 0 5240 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_187
timestamp 1515852544
transform -1 0 5352 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_649
timestamp 1515852544
transform 1 0 5352 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_12
timestamp 1515852544
transform 1 0 5416 0 -1 2610
box 0 0 64 200
use OAI22X1  OAI22X1_14
timestamp 1515852544
transform -1 0 5560 0 -1 2610
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_157
timestamp 1515852544
transform 1 0 5560 0 -1 2610
box 0 0 192 200
use NOR2X1  NOR2X1_38
timestamp 1515852544
transform -1 0 5800 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_466
timestamp 1515852544
transform -1 0 5864 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_12
timestamp 1515852544
transform 1 0 5864 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_1
timestamp 1515852544
transform -1 0 5960 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_5_0
timestamp 1515852544
transform -1 0 5976 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_5_1
timestamp 1515852544
transform -1 0 5992 0 -1 2610
box 0 0 16 200
use AOI22X1  AOI22X1_138
timestamp 1515852544
transform -1 0 6072 0 -1 2610
box 0 0 80 200
use NAND3X1  NAND3X1_67
timestamp 1515852544
transform 1 0 6072 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_45
timestamp 1515852544
transform -1 0 6200 0 -1 2610
box 0 0 64 200
use AOI22X1  AOI22X1_142
timestamp 1515852544
transform 1 0 6200 0 -1 2610
box 0 0 80 200
use OAI21X1  OAI21X1_674
timestamp 1515852544
transform 1 0 6280 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_675
timestamp 1515852544
transform -1 0 6408 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_282
timestamp 1515852544
transform 1 0 6408 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_283
timestamp 1515852544
transform 1 0 6456 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_257
timestamp 1515852544
transform 1 0 6504 0 -1 2610
box 0 0 48 200
use AND2X2  AND2X2_2
timestamp 1515852544
transform 1 0 6552 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_323
timestamp 1515852544
transform 1 0 6616 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_256
timestamp 1515852544
transform -1 0 6728 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_39
timestamp 1515852544
transform -1 0 6776 0 -1 2610
box 0 0 48 200
use FILL  FILL_13_1
timestamp 1515852544
transform -1 0 6792 0 -1 2610
box 0 0 16 200
use FILL  FILL_13_2
timestamp 1515852544
transform -1 0 6808 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_41
timestamp 1515852544
transform 1 0 8 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_108
timestamp 1515852544
transform -1 0 120 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_42
timestamp 1515852544
transform 1 0 120 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_170
timestamp 1515852544
transform 1 0 168 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_7
timestamp 1515852544
transform 1 0 232 0 1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_171
timestamp 1515852544
transform -1 0 376 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_167
timestamp 1515852544
transform -1 0 440 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_169
timestamp 1515852544
transform -1 0 504 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_133
timestamp 1515852544
transform 1 0 504 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_340
timestamp 1515852544
transform 1 0 568 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_40
timestamp 1515852544
transform -1 0 712 0 1 2210
box 0 0 80 200
use BUFX4  BUFX4_117
timestamp 1515852544
transform -1 0 776 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_337
timestamp 1515852544
transform -1 0 840 0 1 2210
box 0 0 64 200
use FILL  FILL_11_0_0
timestamp 1515852544
transform -1 0 856 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1515852544
transform -1 0 872 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_27
timestamp 1515852544
transform -1 0 936 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_158
timestamp 1515852544
transform 1 0 936 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_4
timestamp 1515852544
transform -1 0 1080 0 1 2210
box 0 0 80 200
use NAND3X1  NAND3X1_104
timestamp 1515852544
transform 1 0 1080 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_155
timestamp 1515852544
transform -1 0 1208 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_34
timestamp 1515852544
transform -1 0 1256 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_87
timestamp 1515852544
transform 1 0 1256 0 1 2210
box 0 0 192 200
use AOI22X1  AOI22X1_31
timestamp 1515852544
transform 1 0 1448 0 1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_289
timestamp 1515852544
transform 1 0 1528 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_293
timestamp 1515852544
transform -1 0 1656 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_291
timestamp 1515852544
transform -1 0 1720 0 1 2210
box 0 0 64 200
use INVX1  INVX1_35
timestamp 1515852544
transform 1 0 1720 0 1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_2
timestamp 1515852544
transform 1 0 1752 0 1 2210
box 0 0 80 200
use FILL  FILL_11_1_0
timestamp 1515852544
transform -1 0 1848 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1515852544
transform -1 0 1864 0 1 2210
box 0 0 16 200
use INVX1  INVX1_34
timestamp 1515852544
transform -1 0 1896 0 1 2210
box 0 0 32 200
use INVX1  INVX1_41
timestamp 1515852544
transform 1 0 1896 0 1 2210
box 0 0 32 200
use INVX1  INVX1_40
timestamp 1515852544
transform 1 0 1928 0 1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_5
timestamp 1515852544
transform -1 0 2040 0 1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_291
timestamp 1515852544
transform 1 0 2040 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_79
timestamp 1515852544
transform 1 0 2088 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_57
timestamp 1515852544
transform 1 0 2136 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_46
timestamp 1515852544
transform -1 0 2264 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_226
timestamp 1515852544
transform -1 0 2328 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_18
timestamp 1515852544
transform 1 0 2328 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_13
timestamp 1515852544
transform -1 0 2440 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_16
timestamp 1515852544
transform -1 0 2488 0 1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_68
timestamp 1515852544
transform -1 0 2536 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_247
timestamp 1515852544
transform -1 0 2584 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_56
timestamp 1515852544
transform 1 0 2584 0 1 2210
box 0 0 192 200
use BUFX4  BUFX4_86
timestamp 1515852544
transform 1 0 2776 0 1 2210
box 0 0 64 200
use FILL  FILL_11_2_0
timestamp 1515852544
transform 1 0 2840 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1515852544
transform 1 0 2856 0 1 2210
box 0 0 16 200
use AOI22X1  AOI22X1_1
timestamp 1515852544
transform 1 0 2872 0 1 2210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_149
timestamp 1515852544
transform -1 0 3144 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_266
timestamp 1515852544
transform 1 0 3144 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_557
timestamp 1515852544
transform 1 0 3192 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_568
timestamp 1515852544
transform 1 0 3256 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_267
timestamp 1515852544
transform -1 0 3368 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_501
timestamp 1515852544
transform -1 0 3432 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_150
timestamp 1515852544
transform 1 0 3432 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_436
timestamp 1515852544
transform 1 0 3624 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_144
timestamp 1515852544
transform -1 0 3736 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_11
timestamp 1515852544
transform 1 0 3736 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_143
timestamp 1515852544
transform 1 0 3800 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_435
timestamp 1515852544
transform -1 0 3912 0 1 2210
box 0 0 64 200
use FILL  FILL_11_3_0
timestamp 1515852544
transform 1 0 3912 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_1
timestamp 1515852544
transform 1 0 3928 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_82
timestamp 1515852544
transform 1 0 3944 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_196
timestamp 1515852544
transform 1 0 4008 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_137
timestamp 1515852544
transform 1 0 4072 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_186
timestamp 1515852544
transform -1 0 4200 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_107
timestamp 1515852544
transform 1 0 4200 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_216
timestamp 1515852544
transform -1 0 4328 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_45
timestamp 1515852544
transform 1 0 4328 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_227
timestamp 1515852544
transform 1 0 4392 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_14
timestamp 1515852544
transform -1 0 4520 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_2
timestamp 1515852544
transform 1 0 4520 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_687
timestamp 1515852544
transform 1 0 4584 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_689
timestamp 1515852544
transform -1 0 4712 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_165
timestamp 1515852544
transform 1 0 4712 0 1 2210
box 0 0 80 200
use BUFX4  BUFX4_139
timestamp 1515852544
transform -1 0 4856 0 1 2210
box 0 0 64 200
use FILL  FILL_11_4_0
timestamp 1515852544
transform 1 0 4856 0 1 2210
box 0 0 16 200
use FILL  FILL_11_4_1
timestamp 1515852544
transform 1 0 4872 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_123
timestamp 1515852544
transform 1 0 4888 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_456
timestamp 1515852544
transform 1 0 5080 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_459
timestamp 1515852544
transform -1 0 5208 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_65
timestamp 1515852544
transform 1 0 5208 0 1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_460
timestamp 1515852544
transform -1 0 5352 0 1 2210
box 0 0 64 200
use INVX1  INVX1_61
timestamp 1515852544
transform -1 0 5384 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_650
timestamp 1515852544
transform -1 0 5448 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_654
timestamp 1515852544
transform 1 0 5448 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_652
timestamp 1515852544
transform 1 0 5512 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_43
timestamp 1515852544
transform 1 0 5576 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_651
timestamp 1515852544
transform -1 0 5704 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_464
timestamp 1515852544
transform 1 0 5704 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_32
timestamp 1515852544
transform 1 0 5768 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_41
timestamp 1515852544
transform -1 0 5896 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_32
timestamp 1515852544
transform -1 0 5960 0 1 2210
box 0 0 64 200
use FILL  FILL_11_5_0
timestamp 1515852544
transform -1 0 5976 0 1 2210
box 0 0 16 200
use FILL  FILL_11_5_1
timestamp 1515852544
transform -1 0 5992 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_463
timestamp 1515852544
transform -1 0 6056 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_158
timestamp 1515852544
transform -1 0 6104 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_4
timestamp 1515852544
transform -1 0 6168 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_3
timestamp 1515852544
transform 1 0 6168 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_169
timestamp 1515852544
transform -1 0 6424 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_290
timestamp 1515852544
transform 1 0 6424 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_301
timestamp 1515852544
transform -1 0 6552 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_335
timestamp 1515852544
transform 1 0 6552 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_179
timestamp 1515852544
transform 1 0 6616 0 1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_91
timestamp 1515852544
transform 1 0 8 0 -1 2210
box 0 0 192 200
use OAI22X1  OAI22X1_26
timestamp 1515852544
transform 1 0 200 0 -1 2210
box 0 0 80 200
use NOR2X1  NOR2X1_11
timestamp 1515852544
transform -1 0 328 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_24
timestamp 1515852544
transform 1 0 328 0 -1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_27
timestamp 1515852544
transform 1 0 360 0 -1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_106
timestamp 1515852544
transform 1 0 440 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_339
timestamp 1515852544
transform -1 0 552 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_105
timestamp 1515852544
transform -1 0 600 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_338
timestamp 1515852544
transform -1 0 664 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_361
timestamp 1515852544
transform 1 0 664 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_118
timestamp 1515852544
transform -1 0 776 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_0_0
timestamp 1515852544
transform 1 0 776 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1515852544
transform 1 0 792 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_48
timestamp 1515852544
transform 1 0 808 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_65
timestamp 1515852544
transform 1 0 1000 0 -1 2210
box 0 0 192 200
use BUFX4  BUFX4_111
timestamp 1515852544
transform -1 0 1256 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1515852544
transform 1 0 1256 0 -1 2210
box 0 0 192 200
use AOI22X1  AOI22X1_123
timestamp 1515852544
transform 1 0 1448 0 -1 2210
box 0 0 80 200
use AND2X2  AND2X2_34
timestamp 1515852544
transform 1 0 1528 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_124
timestamp 1515852544
transform -1 0 1672 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_101
timestamp 1515852544
transform 1 0 1672 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_128
timestamp 1515852544
transform 1 0 1736 0 -1 2210
box 0 0 80 200
use FILL  FILL_10_1_0
timestamp 1515852544
transform 1 0 1816 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1515852544
transform 1 0 1832 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_209
timestamp 1515852544
transform 1 0 1848 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_13
timestamp 1515852544
transform 1 0 1912 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_442
timestamp 1515852544
transform 1 0 1992 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_444
timestamp 1515852544
transform -1 0 2120 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_447
timestamp 1515852544
transform 1 0 2120 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_443
timestamp 1515852544
transform -1 0 2248 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_24
timestamp 1515852544
transform 1 0 2248 0 -1 2210
box 0 0 80 200
use INVX1  INVX1_37
timestamp 1515852544
transform 1 0 2328 0 -1 2210
box 0 0 32 200
use OAI22X1  OAI22X1_3
timestamp 1515852544
transform 1 0 2360 0 -1 2210
box 0 0 80 200
use INVX1  INVX1_36
timestamp 1515852544
transform -1 0 2472 0 -1 2210
box 0 0 32 200
use BUFX4  BUFX4_8
timestamp 1515852544
transform -1 0 2536 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_76
timestamp 1515852544
transform -1 0 2728 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_47
timestamp 1515852544
transform 1 0 2728 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_50
timestamp 1515852544
transform 1 0 2792 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_2_0
timestamp 1515852544
transform -1 0 2872 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1515852544
transform -1 0 2888 0 -1 2210
box 0 0 16 200
use AOI22X1  AOI22X1_177
timestamp 1515852544
transform -1 0 2968 0 -1 2210
box 0 0 80 200
use NAND3X1  NAND3X1_89
timestamp 1515852544
transform -1 0 3032 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_304
timestamp 1515852544
transform 1 0 3032 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_48
timestamp 1515852544
transform -1 0 3144 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_49
timestamp 1515852544
transform -1 0 3208 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_305
timestamp 1515852544
transform -1 0 3256 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_75
timestamp 1515852544
transform -1 0 3320 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_158
timestamp 1515852544
transform 1 0 3320 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_545
timestamp 1515852544
transform 1 0 3400 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_579
timestamp 1515852544
transform -1 0 3528 0 -1 2210
box 0 0 64 200
use OAI22X1  OAI22X1_24
timestamp 1515852544
transform 1 0 3528 0 -1 2210
box 0 0 80 200
use AOI22X1  AOI22X1_172
timestamp 1515852544
transform 1 0 3608 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_437
timestamp 1515852544
transform 1 0 3688 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_60
timestamp 1515852544
transform -1 0 3832 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_433
timestamp 1515852544
transform -1 0 3896 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_3_0
timestamp 1515852544
transform -1 0 3912 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_3_1
timestamp 1515852544
transform -1 0 3928 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_10
timestamp 1515852544
transform -1 0 3992 0 -1 2210
box 0 0 64 200
use OAI22X1  OAI22X1_9
timestamp 1515852544
transform -1 0 4072 0 -1 2210
box 0 0 80 200
use INVX1  INVX1_48
timestamp 1515852544
transform -1 0 4104 0 -1 2210
box 0 0 32 200
use NOR3X1  NOR3X1_5
timestamp 1515852544
transform -1 0 4232 0 -1 2210
box 0 0 128 200
use OAI21X1  OAI21X1_59
timestamp 1515852544
transform 1 0 4232 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_179
timestamp 1515852544
transform -1 0 4376 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_56
timestamp 1515852544
transform 1 0 4376 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_58
timestamp 1515852544
transform 1 0 4440 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_309
timestamp 1515852544
transform -1 0 4552 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_91
timestamp 1515852544
transform 1 0 4552 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_308
timestamp 1515852544
transform -1 0 4664 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_78
timestamp 1515852544
transform -1 0 4856 0 -1 2210
box 0 0 192 200
use FILL  FILL_10_4_0
timestamp 1515852544
transform 1 0 4856 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_4_1
timestamp 1515852544
transform 1 0 4872 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_166
timestamp 1515852544
transform 1 0 4888 0 -1 2210
box 0 0 192 200
use AND2X2  AND2X2_31
timestamp 1515852544
transform 1 0 5080 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_114
timestamp 1515852544
transform 1 0 5144 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_458
timestamp 1515852544
transform 1 0 5176 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_17
timestamp 1515852544
transform -1 0 5304 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_154
timestamp 1515852544
transform -1 0 5352 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_156
timestamp 1515852544
transform -1 0 5544 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_113
timestamp 1515852544
transform 1 0 5544 0 -1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_236
timestamp 1515852544
transform 1 0 5736 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_653
timestamp 1515852544
transform -1 0 5848 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_237
timestamp 1515852544
transform 1 0 5848 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_465
timestamp 1515852544
transform 1 0 5896 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_5_0
timestamp 1515852544
transform -1 0 5976 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_5_1
timestamp 1515852544
transform -1 0 5992 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_156
timestamp 1515852544
transform -1 0 6040 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_421
timestamp 1515852544
transform -1 0 6104 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_112
timestamp 1515852544
transform 1 0 6104 0 -1 2210
box 0 0 32 200
use AOI22X1  AOI22X1_141
timestamp 1515852544
transform -1 0 6216 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_5
timestamp 1515852544
transform -1 0 6280 0 -1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_56
timestamp 1515852544
transform -1 0 6360 0 -1 2210
box 0 0 80 200
use OAI21X1  OAI21X1_419
timestamp 1515852544
transform 1 0 6360 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_420
timestamp 1515852544
transform -1 0 6488 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_6
timestamp 1515852544
transform -1 0 6552 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_422
timestamp 1515852544
transform -1 0 6616 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_111
timestamp 1515852544
transform 1 0 6616 0 -1 2210
box 0 0 32 200
use AOI21X1  AOI21X1_31
timestamp 1515852544
transform -1 0 6712 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_189
timestamp 1515852544
transform 1 0 6712 0 -1 2210
box 0 0 64 200
use FILL  FILL_11_1
timestamp 1515852544
transform -1 0 6792 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_2
timestamp 1515852544
transform -1 0 6808 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_44
timestamp 1515852544
transform 1 0 8 0 1 1810
box 0 0 192 200
use NAND2X1  NAND2X1_110
timestamp 1515852544
transform 1 0 200 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_135
timestamp 1515852544
transform 1 0 248 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_42
timestamp 1515852544
transform 1 0 312 0 1 1810
box 0 0 80 200
use INVX1  INVX1_13
timestamp 1515852544
transform 1 0 392 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_349
timestamp 1515852544
transform 1 0 424 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_347
timestamp 1515852544
transform -1 0 552 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_348
timestamp 1515852544
transform -1 0 616 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_345
timestamp 1515852544
transform -1 0 680 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_360
timestamp 1515852544
transform 1 0 680 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_117
timestamp 1515852544
transform 1 0 744 0 1 1810
box 0 0 48 200
use FILL  FILL_9_0_0
timestamp 1515852544
transform 1 0 792 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1515852544
transform 1 0 808 0 1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_138
timestamp 1515852544
transform 1 0 824 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_362
timestamp 1515852544
transform 1 0 888 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_45
timestamp 1515852544
transform -1 0 1032 0 1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_81
timestamp 1515852544
transform 1 0 1032 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_359
timestamp 1515852544
transform -1 0 1160 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1515852544
transform 1 0 1160 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_313
timestamp 1515852544
transform 1 0 1352 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_98
timestamp 1515852544
transform -1 0 1464 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_315
timestamp 1515852544
transform -1 0 1528 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_314
timestamp 1515852544
transform -1 0 1592 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_21
timestamp 1515852544
transform 1 0 1592 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_316
timestamp 1515852544
transform -1 0 1720 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_40
timestamp 1515852544
transform -1 0 1784 0 1 1810
box 0 0 64 200
use OAI22X1  OAI22X1_7
timestamp 1515852544
transform 1 0 1784 0 1 1810
box 0 0 80 200
use FILL  FILL_9_1_0
timestamp 1515852544
transform 1 0 1864 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1515852544
transform 1 0 1880 0 1 1810
box 0 0 16 200
use INVX1  INVX1_42
timestamp 1515852544
transform 1 0 1896 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_24
timestamp 1515852544
transform 1 0 1928 0 1 1810
box 0 0 48 200
use BUFX4  BUFX4_52
timestamp 1515852544
transform -1 0 2040 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_49
timestamp 1515852544
transform -1 0 2104 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_62
timestamp 1515852544
transform 1 0 2104 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_148
timestamp 1515852544
transform -1 0 2232 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_149
timestamp 1515852544
transform -1 0 2280 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_107
timestamp 1515852544
transform 1 0 2280 0 1 1810
box 0 0 64 200
use INVX1  INVX1_30
timestamp 1515852544
transform 1 0 2344 0 1 1810
box 0 0 32 200
use OAI22X1  OAI22X1_29
timestamp 1515852544
transform 1 0 2376 0 1 1810
box 0 0 80 200
use INVX1  INVX1_29
timestamp 1515852544
transform -1 0 2488 0 1 1810
box 0 0 32 200
use AOI22X1  AOI22X1_139
timestamp 1515852544
transform -1 0 2568 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_303
timestamp 1515852544
transform 1 0 2568 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_44
timestamp 1515852544
transform 1 0 2616 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_301
timestamp 1515852544
transform 1 0 2680 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_43
timestamp 1515852544
transform -1 0 2792 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_45
timestamp 1515852544
transform 1 0 2792 0 1 1810
box 0 0 64 200
use FILL  FILL_9_2_0
timestamp 1515852544
transform 1 0 2856 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1515852544
transform 1 0 2872 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_42
timestamp 1515852544
transform 1 0 2888 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_125
timestamp 1515852544
transform 1 0 2952 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_385
timestamp 1515852544
transform -1 0 3064 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_383
timestamp 1515852544
transform -1 0 3128 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_39
timestamp 1515852544
transform 1 0 3128 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_111
timestamp 1515852544
transform 1 0 3192 0 1 1810
box 0 0 80 200
use AOI22X1  AOI22X1_79
timestamp 1515852544
transform -1 0 3352 0 1 1810
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_55
timestamp 1515852544
transform 1 0 3352 0 1 1810
box 0 0 192 200
use INVX1  INVX1_25
timestamp 1515852544
transform -1 0 3576 0 1 1810
box 0 0 32 200
use BUFX4  BUFX4_55
timestamp 1515852544
transform -1 0 3640 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_32
timestamp 1515852544
transform 1 0 3640 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_161
timestamp 1515852544
transform -1 0 3896 0 1 1810
box 0 0 192 200
use FILL  FILL_9_3_0
timestamp 1515852544
transform -1 0 3912 0 1 1810
box 0 0 16 200
use FILL  FILL_9_3_1
timestamp 1515852544
transform -1 0 3928 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_176
timestamp 1515852544
transform -1 0 3992 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_36
timestamp 1515852544
transform -1 0 4056 0 1 1810
box 0 0 64 200
use INVX1  INVX1_47
timestamp 1515852544
transform -1 0 4088 0 1 1810
box 0 0 32 200
use AOI22X1  AOI22X1_119
timestamp 1515852544
transform -1 0 4168 0 1 1810
box 0 0 80 200
use BUFX4  BUFX4_154
timestamp 1515852544
transform -1 0 4232 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_163
timestamp 1515852544
transform 1 0 4232 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_165
timestamp 1515852544
transform 1 0 4296 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_9
timestamp 1515852544
transform 1 0 4360 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_40
timestamp 1515852544
transform -1 0 4456 0 1 1810
box 0 0 48 200
use BUFX4  BUFX4_33
timestamp 1515852544
transform 1 0 4456 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_55
timestamp 1515852544
transform -1 0 4584 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_408
timestamp 1515852544
transform 1 0 4584 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_55
timestamp 1515852544
transform -1 0 4728 0 1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_405
timestamp 1515852544
transform 1 0 4728 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_407
timestamp 1515852544
transform -1 0 4856 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1515852544
transform -1 0 4920 0 1 1810
box 0 0 64 200
use FILL  FILL_9_4_0
timestamp 1515852544
transform -1 0 4936 0 1 1810
box 0 0 16 200
use FILL  FILL_9_4_1
timestamp 1515852544
transform -1 0 4952 0 1 1810
box 0 0 16 200
use INVX1  INVX1_92
timestamp 1515852544
transform -1 0 4984 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_136
timestamp 1515852544
transform -1 0 5032 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_506
timestamp 1515852544
transform 1 0 5032 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_133
timestamp 1515852544
transform 1 0 5096 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_172
timestamp 1515852544
transform 1 0 5176 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_508
timestamp 1515852544
transform 1 0 5224 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_75
timestamp 1515852544
transform 1 0 5288 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_174
timestamp 1515852544
transform 1 0 5368 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_173
timestamp 1515852544
transform -1 0 5464 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_33
timestamp 1515852544
transform 1 0 5464 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_62
timestamp 1515852544
transform -1 0 5576 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_188
timestamp 1515852544
transform 1 0 5576 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_16
timestamp 1515852544
transform 1 0 5640 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_424
timestamp 1515852544
transform 1 0 5704 0 1 1810
box 0 0 64 200
use INVX1  INVX1_113
timestamp 1515852544
transform -1 0 5800 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_425
timestamp 1515852544
transform -1 0 5864 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_426
timestamp 1515852544
transform 1 0 5864 0 1 1810
box 0 0 64 200
use FILL  FILL_9_5_0
timestamp 1515852544
transform -1 0 5944 0 1 1810
box 0 0 16 200
use FILL  FILL_9_5_1
timestamp 1515852544
transform -1 0 5960 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_427
timestamp 1515852544
transform -1 0 6024 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_58
timestamp 1515852544
transform 1 0 6024 0 1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_428
timestamp 1515852544
transform 1 0 6104 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_170
timestamp 1515852544
transform -1 0 6360 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_415
timestamp 1515852544
transform 1 0 6360 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_139
timestamp 1515852544
transform 1 0 6424 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_140
timestamp 1515852544
transform 1 0 6472 0 1 1810
box 0 0 48 200
use AND2X2  AND2X2_30
timestamp 1515852544
transform 1 0 6520 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_418
timestamp 1515852544
transform 1 0 6584 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_23
timestamp 1515852544
transform -1 0 6712 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_255
timestamp 1515852544
transform -1 0 6760 0 1 1810
box 0 0 48 200
use FILL  FILL_10_1
timestamp 1515852544
transform 1 0 6760 0 1 1810
box 0 0 16 200
use FILL  FILL_10_2
timestamp 1515852544
transform 1 0 6776 0 1 1810
box 0 0 16 200
use FILL  FILL_10_3
timestamp 1515852544
transform 1 0 6792 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_66
timestamp 1515852544
transform 1 0 8 0 -1 1810
box 0 0 192 200
use INVX1  INVX1_109
timestamp 1515852544
transform 1 0 200 0 -1 1810
box 0 0 32 200
use AOI22X1  AOI22X1_168
timestamp 1515852544
transform 1 0 232 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_6
timestamp 1515852544
transform -1 0 376 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_3
timestamp 1515852544
transform -1 0 440 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_109
timestamp 1515852544
transform 1 0 440 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_151
timestamp 1515852544
transform 1 0 488 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_32
timestamp 1515852544
transform -1 0 600 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_150
timestamp 1515852544
transform -1 0 664 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_696
timestamp 1515852544
transform 1 0 664 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_286
timestamp 1515852544
transform -1 0 776 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_697
timestamp 1515852544
transform 1 0 776 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_0_0
timestamp 1515852544
transform -1 0 856 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1515852544
transform -1 0 872 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_287
timestamp 1515852544
transform -1 0 920 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_45
timestamp 1515852544
transform 1 0 920 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_695
timestamp 1515852544
transform 1 0 952 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_698
timestamp 1515852544
transform -1 0 1080 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_167
timestamp 1515852544
transform -1 0 1160 0 -1 1810
box 0 0 80 200
use BUFX4  BUFX4_124
timestamp 1515852544
transform -1 0 1224 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_210
timestamp 1515852544
transform -1 0 1288 0 -1 1810
box 0 0 64 200
use OAI22X1  OAI22X1_8
timestamp 1515852544
transform -1 0 1368 0 -1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_97
timestamp 1515852544
transform 1 0 1368 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_99
timestamp 1515852544
transform -1 0 1464 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_290
timestamp 1515852544
transform 1 0 1464 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_8
timestamp 1515852544
transform 1 0 1512 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1515852544
transform 1 0 1576 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_292
timestamp 1515852544
transform -1 0 1688 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_311
timestamp 1515852544
transform 1 0 1688 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_83
timestamp 1515852544
transform 1 0 1752 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_1_0
timestamp 1515852544
transform 1 0 1816 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1515852544
transform 1 0 1832 0 -1 1810
box 0 0 16 200
use AOI22X1  AOI22X1_169
timestamp 1515852544
transform 1 0 1848 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_10
timestamp 1515852544
transform -1 0 1992 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_29
timestamp 1515852544
transform -1 0 2056 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_110
timestamp 1515852544
transform -1 0 2136 0 -1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_14
timestamp 1515852544
transform -1 0 2200 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_68
timestamp 1515852544
transform 1 0 2200 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_694
timestamp 1515852544
transform -1 0 2344 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_166
timestamp 1515852544
transform -1 0 2424 0 -1 1810
box 0 0 80 200
use BUFX4  BUFX4_194
timestamp 1515852544
transform -1 0 2488 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_75
timestamp 1515852544
transform -1 0 2680 0 -1 1810
box 0 0 192 200
use NAND3X1  NAND3X1_88
timestamp 1515852544
transform 1 0 2680 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_176
timestamp 1515852544
transform 1 0 2744 0 -1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_66
timestamp 1515852544
transform 1 0 2824 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_2_0
timestamp 1515852544
transform -1 0 2888 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1515852544
transform -1 0 2904 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_3
timestamp 1515852544
transform -1 0 2968 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_50
timestamp 1515852544
transform 1 0 2968 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_386
timestamp 1515852544
transform -1 0 3112 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_395
timestamp 1515852544
transform 1 0 3112 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_52
timestamp 1515852544
transform -1 0 3256 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_392
timestamp 1515852544
transform 1 0 3256 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_394
timestamp 1515852544
transform -1 0 3384 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1515852544
transform -1 0 3448 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_129
timestamp 1515852544
transform -1 0 3496 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_162
timestamp 1515852544
transform -1 0 3688 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_391
timestamp 1515852544
transform 1 0 3688 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_51
timestamp 1515852544
transform -1 0 3832 0 -1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_4
timestamp 1515852544
transform -1 0 3896 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_3_0
timestamp 1515852544
transform -1 0 3912 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_3_1
timestamp 1515852544
transform -1 0 3928 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_387
timestamp 1515852544
transform -1 0 3992 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_389
timestamp 1515852544
transform -1 0 4056 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_127
timestamp 1515852544
transform -1 0 4104 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_396
timestamp 1515852544
transform 1 0 4104 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_397
timestamp 1515852544
transform -1 0 4232 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_164
timestamp 1515852544
transform 1 0 4232 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_166
timestamp 1515852544
transform 1 0 4296 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_6
timestamp 1515852544
transform -1 0 4440 0 -1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_106
timestamp 1515852544
transform 1 0 4440 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_39
timestamp 1515852544
transform -1 0 4552 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_400
timestamp 1515852544
transform -1 0 4616 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_89
timestamp 1515852544
transform -1 0 4808 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_406
timestamp 1515852544
transform -1 0 4872 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_134
timestamp 1515852544
transform -1 0 4920 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_4_0
timestamp 1515852544
transform -1 0 4936 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_4_1
timestamp 1515852544
transform -1 0 4952 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_684
timestamp 1515852544
transform -1 0 5016 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_57
timestamp 1515852544
transform -1 0 5080 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_7
timestamp 1515852544
transform -1 0 5128 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_174
timestamp 1515852544
transform -1 0 5192 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_145
timestamp 1515852544
transform -1 0 5384 0 -1 1810
box 0 0 192 200
use NAND3X1  NAND3X1_25
timestamp 1515852544
transform 1 0 5384 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_36
timestamp 1515852544
transform -1 0 5496 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_116
timestamp 1515852544
transform 1 0 5496 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_507
timestamp 1515852544
transform -1 0 5592 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_33
timestamp 1515852544
transform -1 0 5656 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_178
timestamp 1515852544
transform 1 0 5656 0 -1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_131
timestamp 1515852544
transform -1 0 5800 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_130
timestamp 1515852544
transform 1 0 5800 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_95
timestamp 1515852544
transform -1 0 5896 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_27
timestamp 1515852544
transform 1 0 5896 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_5_0
timestamp 1515852544
transform 1 0 5944 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_5_1
timestamp 1515852544
transform 1 0 5960 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_102
timestamp 1515852544
transform 1 0 5976 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_129
timestamp 1515852544
transform -1 0 6104 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_409
timestamp 1515852544
transform 1 0 6104 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1515852544
transform -1 0 6360 0 -1 1810
box 0 0 192 200
use BUFX4  BUFX4_78
timestamp 1515852544
transform 1 0 6360 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_167
timestamp 1515852544
transform 1 0 6424 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_417
timestamp 1515852544
transform 1 0 6616 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_30
timestamp 1515852544
transform -1 0 6744 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_416
timestamp 1515852544
transform -1 0 6808 0 -1 1810
box 0 0 64 200
use INVX8  INVX8_14
timestamp 1515852544
transform 1 0 8 0 1 1410
box 0 0 80 200
use INVX1  INVX1_8
timestamp 1515852544
transform 1 0 88 0 1 1410
box 0 0 32 200
use INVX8  INVX8_17
timestamp 1515852544
transform 1 0 120 0 1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_82
timestamp 1515852544
transform -1 0 264 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_289
timestamp 1515852544
transform 1 0 264 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_5
timestamp 1515852544
transform -1 0 376 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_288
timestamp 1515852544
transform 1 0 376 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_4
timestamp 1515852544
transform -1 0 488 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_153
timestamp 1515852544
transform 1 0 488 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_103
timestamp 1515852544
transform -1 0 616 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_3
timestamp 1515852544
transform -1 0 696 0 1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_152
timestamp 1515852544
transform -1 0 760 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_33
timestamp 1515852544
transform -1 0 808 0 1 1410
box 0 0 48 200
use FILL  FILL_7_0_0
timestamp 1515852544
transform 1 0 808 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1515852544
transform 1 0 824 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_211
timestamp 1515852544
transform 1 0 840 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_215
timestamp 1515852544
transform -1 0 968 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_56
timestamp 1515852544
transform 1 0 968 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_213
timestamp 1515852544
transform -1 0 1080 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_214
timestamp 1515852544
transform 1 0 1080 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_58
timestamp 1515852544
transform -1 0 1192 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_66
timestamp 1515852544
transform 1 0 1192 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_93
timestamp 1515852544
transform 1 0 1256 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_305
timestamp 1515852544
transform 1 0 1304 0 1 1410
box 0 0 64 200
use INVX1  INVX1_46
timestamp 1515852544
transform -1 0 1400 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_303
timestamp 1515852544
transform 1 0 1400 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_306
timestamp 1515852544
transform 1 0 1464 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_34
timestamp 1515852544
transform -1 0 1608 0 1 1410
box 0 0 80 200
use NAND2X1  NAND2X1_92
timestamp 1515852544
transform 1 0 1608 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_304
timestamp 1515852544
transform -1 0 1720 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_67
timestamp 1515852544
transform 1 0 1720 0 1 1410
box 0 0 192 200
use FILL  FILL_7_1_0
timestamp 1515852544
transform -1 0 1928 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1515852544
transform -1 0 1944 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_7
timestamp 1515852544
transform -1 0 2008 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_152
timestamp 1515852544
transform -1 0 2200 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_692
timestamp 1515852544
transform 1 0 2200 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_693
timestamp 1515852544
transform 1 0 2264 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_285
timestamp 1515852544
transform -1 0 2376 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_691
timestamp 1515852544
transform -1 0 2440 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_46
timestamp 1515852544
transform -1 0 2504 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_54
timestamp 1515852544
transform 1 0 2504 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_13
timestamp 1515852544
transform -1 0 2632 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_108
timestamp 1515852544
transform -1 0 2696 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_30
timestamp 1515852544
transform 1 0 2696 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_160
timestamp 1515852544
transform 1 0 2760 0 1 1410
box 0 0 192 200
use FILL  FILL_7_2_0
timestamp 1515852544
transform 1 0 2952 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1515852544
transform 1 0 2968 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_123
timestamp 1515852544
transform 1 0 2984 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_384
timestamp 1515852544
transform -1 0 3096 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_393
timestamp 1515852544
transform 1 0 3096 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_128
timestamp 1515852544
transform -1 0 3208 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_37
timestamp 1515852544
transform 1 0 3208 0 1 1410
box 0 0 64 200
use INVX1  INVX1_88
timestamp 1515852544
transform 1 0 3272 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_38
timestamp 1515852544
transform -1 0 3368 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_129
timestamp 1515852544
transform -1 0 3432 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_39
timestamp 1515852544
transform -1 0 3496 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_34
timestamp 1515852544
transform -1 0 3560 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_126
timestamp 1515852544
transform 1 0 3560 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_126
timestamp 1515852544
transform 1 0 3624 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_388
timestamp 1515852544
transform 1 0 3672 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_4
timestamp 1515852544
transform -1 0 3800 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_398
timestamp 1515852544
transform 1 0 3800 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_8
timestamp 1515852544
transform -1 0 3912 0 1 1410
box 0 0 48 200
use FILL  FILL_7_3_0
timestamp 1515852544
transform 1 0 3912 0 1 1410
box 0 0 16 200
use FILL  FILL_7_3_1
timestamp 1515852544
transform 1 0 3928 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_399
timestamp 1515852544
transform 1 0 3944 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_131
timestamp 1515852544
transform -1 0 4056 0 1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_53
timestamp 1515852544
transform -1 0 4136 0 1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_6
timestamp 1515852544
transform 1 0 4136 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_130
timestamp 1515852544
transform -1 0 4248 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_201
timestamp 1515852544
transform -1 0 4312 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_132
timestamp 1515852544
transform 1 0 4312 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_7
timestamp 1515852544
transform -1 0 4424 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_133
timestamp 1515852544
transform 1 0 4424 0 1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_54
timestamp 1515852544
transform 1 0 4472 0 1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_404
timestamp 1515852544
transform -1 0 4616 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_403
timestamp 1515852544
transform -1 0 4680 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_402
timestamp 1515852544
transform -1 0 4744 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_127
timestamp 1515852544
transform 1 0 4744 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_62
timestamp 1515852544
transform 1 0 4808 0 1 1410
box 0 0 192 200
use FILL  FILL_7_4_0
timestamp 1515852544
transform -1 0 5016 0 1 1410
box 0 0 16 200
use FILL  FILL_7_4_1
timestamp 1515852544
transform -1 0 5032 0 1 1410
box 0 0 16 200
use AOI22X1  AOI22X1_164
timestamp 1515852544
transform -1 0 5112 0 1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_685
timestamp 1515852544
transform -1 0 5176 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_64
timestamp 1515852544
transform 1 0 5176 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_648
timestamp 1515852544
transform 1 0 5240 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_103
timestamp 1515852544
transform 1 0 5304 0 1 1410
box 0 0 80 200
use NAND2X1  NAND2X1_232
timestamp 1515852544
transform -1 0 5432 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_45
timestamp 1515852544
transform 1 0 5432 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_647
timestamp 1515852544
transform -1 0 5560 0 1 1410
box 0 0 64 200
use INVX1  INVX1_5
timestamp 1515852544
transform -1 0 5592 0 1 1410
box 0 0 32 200
use INVX8  INVX8_10
timestamp 1515852544
transform -1 0 5672 0 1 1410
box 0 0 80 200
use BUFX4  BUFX4_128
timestamp 1515852544
transform 1 0 5672 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_29
timestamp 1515852544
transform 1 0 5736 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_138
timestamp 1515852544
transform -1 0 5848 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_131
timestamp 1515852544
transform 1 0 5848 0 1 1410
box 0 0 64 200
use FILL  FILL_7_5_0
timestamp 1515852544
transform 1 0 5912 0 1 1410
box 0 0 16 200
use FILL  FILL_7_5_1
timestamp 1515852544
transform 1 0 5928 0 1 1410
box 0 0 16 200
use AOI22X1  AOI22X1_191
timestamp 1515852544
transform 1 0 5944 0 1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_410
timestamp 1515852544
transform -1 0 6088 0 1 1410
box 0 0 64 200
use INVX1  INVX1_110
timestamp 1515852544
transform -1 0 6120 0 1 1410
box 0 0 32 200
use AOI21X1  AOI21X1_28
timestamp 1515852544
transform 1 0 6120 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_411
timestamp 1515852544
transform -1 0 6248 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_29
timestamp 1515852544
transform -1 0 6312 0 1 1410
box 0 0 64 200
use INVX8  INVX8_6
timestamp 1515852544
transform 1 0 6312 0 1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_9
timestamp 1515852544
transform -1 0 6456 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_137
timestamp 1515852544
transform -1 0 6504 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1515852544
transform 1 0 6504 0 1 1410
box 0 0 192 200
use BUFX2  BUFX2_27
timestamp 1515852544
transform 1 0 6696 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_414
timestamp 1515852544
transform 1 0 6744 0 1 1410
box 0 0 64 200
use BUFX2  BUFX2_69
timestamp 1515852544
transform -1 0 56 0 -1 1410
box 0 0 48 200
use BUFX2  BUFX2_1
timestamp 1515852544
transform -1 0 104 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_50
timestamp 1515852544
transform 1 0 104 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_124
timestamp 1515852544
transform 1 0 152 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_21
timestamp 1515852544
transform 1 0 200 0 -1 1410
box 0 0 192 200
use INVX1  INVX1_56
timestamp 1515852544
transform 1 0 392 0 -1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_86
timestamp 1515852544
transform 1 0 424 0 -1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_23
timestamp 1515852544
transform -1 0 808 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_0_0
timestamp 1515852544
transform 1 0 808 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1515852544
transform 1 0 824 0 -1 1410
box 0 0 16 200
use AOI22X1  AOI22X1_16
timestamp 1515852544
transform 1 0 840 0 -1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_114
timestamp 1515852544
transform -1 0 984 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_50
timestamp 1515852544
transform 1 0 984 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_199
timestamp 1515852544
transform -1 0 1096 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_10
timestamp 1515852544
transform 1 0 1096 0 -1 1410
box 0 0 192 200
use AOI22X1  AOI22X1_32
timestamp 1515852544
transform 1 0 1288 0 -1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_127
timestamp 1515852544
transform -1 0 1432 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_87
timestamp 1515852544
transform 1 0 1432 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_295
timestamp 1515852544
transform 1 0 1480 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_294
timestamp 1515852544
transform 1 0 1544 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_130
timestamp 1515852544
transform 1 0 1608 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_113
timestamp 1515852544
transform -1 0 1736 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_28
timestamp 1515852544
transform -1 0 1800 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_1_0
timestamp 1515852544
transform -1 0 1816 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1515852544
transform -1 0 1832 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1515852544
transform -1 0 2024 0 -1 1410
box 0 0 192 200
use AOI22X1  AOI22X1_2
timestamp 1515852544
transform -1 0 2104 0 -1 1410
box 0 0 80 200
use NAND2X1  NAND2X1_96
timestamp 1515852544
transform -1 0 2152 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_172
timestamp 1515852544
transform 1 0 2152 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_284
timestamp 1515852544
transform 1 0 2216 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_179
timestamp 1515852544
transform 1 0 2264 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_80
timestamp 1515852544
transform -1 0 2392 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_205
timestamp 1515852544
transform -1 0 2456 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_204
timestamp 1515852544
transform -1 0 2520 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_64
timestamp 1515852544
transform -1 0 2712 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_261
timestamp 1515852544
transform 1 0 2712 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_75
timestamp 1515852544
transform -1 0 2824 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_262
timestamp 1515852544
transform 1 0 2824 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_2_0
timestamp 1515852544
transform -1 0 2904 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1515852544
transform -1 0 2920 0 -1 1410
box 0 0 16 200
use AOI22X1  AOI22X1_26
timestamp 1515852544
transform -1 0 3000 0 -1 1410
box 0 0 80 200
use NAND3X1  NAND3X1_122
timestamp 1515852544
transform 1 0 3000 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_74
timestamp 1515852544
transform 1 0 3064 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_260
timestamp 1515852544
transform -1 0 3176 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_74
timestamp 1515852544
transform -1 0 3368 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_41
timestamp 1515852544
transform 1 0 3368 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_40
timestamp 1515852544
transform -1 0 3496 0 -1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_175
timestamp 1515852544
transform -1 0 3576 0 -1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_33
timestamp 1515852544
transform 1 0 3576 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_34
timestamp 1515852544
transform -1 0 3704 0 -1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_174
timestamp 1515852544
transform -1 0 3784 0 -1 1410
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_73
timestamp 1515852544
transform -1 0 3976 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_3_0
timestamp 1515852544
transform -1 0 3992 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_3_1
timestamp 1515852544
transform -1 0 4008 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_36
timestamp 1515852544
transform -1 0 4072 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_75
timestamp 1515852544
transform 1 0 4072 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_32
timestamp 1515852544
transform 1 0 4104 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_31
timestamp 1515852544
transform -1 0 4232 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_163
timestamp 1515852544
transform -1 0 4424 0 -1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_165
timestamp 1515852544
transform 1 0 4424 0 -1 1410
box 0 0 192 200
use OAI22X1  OAI22X1_19
timestamp 1515852544
transform -1 0 4696 0 -1 1410
box 0 0 80 200
use BUFX4  BUFX4_169
timestamp 1515852544
transform -1 0 4760 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_38
timestamp 1515852544
transform 1 0 4760 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_4_0
timestamp 1515852544
transform -1 0 4968 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_4_1
timestamp 1515852544
transform -1 0 4984 0 -1 1410
box 0 0 16 200
use INVX1  INVX1_77
timestamp 1515852544
transform -1 0 5016 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_683
timestamp 1515852544
transform 1 0 5016 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_682
timestamp 1515852544
transform -1 0 5144 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_681
timestamp 1515852544
transform 1 0 5144 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_680
timestamp 1515852544
transform -1 0 5272 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_56
timestamp 1515852544
transform 1 0 5272 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_64
timestamp 1515852544
transform 1 0 5336 0 -1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_134
timestamp 1515852544
transform -1 0 5480 0 -1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_646
timestamp 1515852544
transform 1 0 5480 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_40
timestamp 1515852544
transform -1 0 5608 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_234
timestamp 1515852544
transform 1 0 5608 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_233
timestamp 1515852544
transform -1 0 5704 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_112
timestamp 1515852544
transform -1 0 5896 0 -1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_28
timestamp 1515852544
transform 1 0 5896 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_5_0
timestamp 1515852544
transform -1 0 5960 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_5_1
timestamp 1515852544
transform -1 0 5976 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_29
timestamp 1515852544
transform -1 0 6024 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_511
timestamp 1515852544
transform 1 0 6024 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_80
timestamp 1515852544
transform -1 0 6152 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_513
timestamp 1515852544
transform -1 0 6216 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_176
timestamp 1515852544
transform 1 0 6216 0 -1 1410
box 0 0 48 200
use AND2X2  AND2X2_35
timestamp 1515852544
transform 1 0 6264 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_514
timestamp 1515852544
transform 1 0 6328 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_175
timestamp 1515852544
transform -1 0 6440 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_33
timestamp 1515852544
transform -1 0 6504 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_509
timestamp 1515852544
transform 1 0 6504 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_510
timestamp 1515852544
transform -1 0 6632 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_515
timestamp 1515852544
transform 1 0 6632 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_74
timestamp 1515852544
transform 1 0 6696 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_413
timestamp 1515852544
transform 1 0 6728 0 -1 1410
box 0 0 64 200
use FILL  FILL_7_1
timestamp 1515852544
transform -1 0 6808 0 -1 1410
box 0 0 16 200
use NAND3X1  NAND3X1_112
timestamp 1515852544
transform -1 0 72 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_14
timestamp 1515852544
transform -1 0 152 0 1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_206
timestamp 1515852544
transform -1 0 216 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_52
timestamp 1515852544
transform -1 0 264 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_204
timestamp 1515852544
transform -1 0 328 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_203
timestamp 1515852544
transform -1 0 392 0 1 1010
box 0 0 64 200
use INVX1  INVX1_55
timestamp 1515852544
transform 1 0 392 0 1 1010
box 0 0 32 200
use OAI22X1  OAI22X1_11
timestamp 1515852544
transform 1 0 424 0 1 1010
box 0 0 80 200
use BUFX4  BUFX4_166
timestamp 1515852544
transform -1 0 568 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_163
timestamp 1515852544
transform -1 0 632 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_69
timestamp 1515852544
transform 1 0 632 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_248
timestamp 1515852544
transform -1 0 744 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_165
timestamp 1515852544
transform 1 0 744 0 1 1010
box 0 0 64 200
use FILL  FILL_5_0_0
timestamp 1515852544
transform 1 0 808 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1515852544
transform 1 0 824 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_202
timestamp 1515852544
transform 1 0 840 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_12
timestamp 1515852544
transform -1 0 984 0 1 1010
box 0 0 80 200
use NAND3X1  NAND3X1_111
timestamp 1515852544
transform -1 0 1048 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_20
timestamp 1515852544
transform 1 0 1048 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_198
timestamp 1515852544
transform -1 0 1304 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_200
timestamp 1515852544
transform -1 0 1368 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_30
timestamp 1515852544
transform -1 0 1416 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_88
timestamp 1515852544
transform 1 0 1416 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_296
timestamp 1515852544
transform 1 0 1464 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_297
timestamp 1515852544
transform -1 0 1592 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_79
timestamp 1515852544
transform -1 0 1656 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_121
timestamp 1515852544
transform 1 0 1656 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_33
timestamp 1515852544
transform 1 0 1720 0 1 1010
box 0 0 192 200
use FILL  FILL_5_1_0
timestamp 1515852544
transform -1 0 1928 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1515852544
transform -1 0 1944 0 1 1010
box 0 0 16 200
use AOI22X1  AOI22X1_117
timestamp 1515852544
transform -1 0 2024 0 1 1010
box 0 0 80 200
use BUFX4  BUFX4_70
timestamp 1515852544
transform -1 0 2088 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_49
timestamp 1515852544
transform 1 0 2088 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_109
timestamp 1515852544
transform -1 0 2216 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_68
timestamp 1515852544
transform 1 0 2216 0 1 1010
box 0 0 64 200
use INVX8  INVX8_2
timestamp 1515852544
transform 1 0 2280 0 1 1010
box 0 0 80 200
use BUFX4  BUFX4_60
timestamp 1515852544
transform 1 0 2360 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_95
timestamp 1515852544
transform 1 0 2424 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_19
timestamp 1515852544
transform -1 0 2568 0 1 1010
box 0 0 80 200
use BUFX4  BUFX4_164
timestamp 1515852544
transform -1 0 2632 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_64
timestamp 1515852544
transform 1 0 2632 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_229
timestamp 1515852544
transform -1 0 2744 0 1 1010
box 0 0 64 200
use INVX1  INVX1_64
timestamp 1515852544
transform 1 0 2744 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_226
timestamp 1515852544
transform -1 0 2840 0 1 1010
box 0 0 64 200
use FILL  FILL_5_2_0
timestamp 1515852544
transform -1 0 2856 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1515852544
transform -1 0 2872 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_228
timestamp 1515852544
transform -1 0 2936 0 1 1010
box 0 0 64 200
use OAI22X1  OAI22X1_16
timestamp 1515852544
transform 1 0 2936 0 1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_259
timestamp 1515852544
transform -1 0 3080 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_161
timestamp 1515852544
transform 1 0 3080 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_113
timestamp 1515852544
transform -1 0 3208 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_22
timestamp 1515852544
transform -1 0 3400 0 1 1010
box 0 0 192 200
use NOR2X1  NOR2X1_35
timestamp 1515852544
transform 1 0 3400 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_34
timestamp 1515852544
transform 1 0 3448 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_53
timestamp 1515852544
transform 1 0 3640 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_307
timestamp 1515852544
transform -1 0 3752 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_135
timestamp 1515852544
transform 1 0 3752 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_54
timestamp 1515852544
transform -1 0 3880 0 1 1010
box 0 0 64 200
use FILL  FILL_5_3_0
timestamp 1515852544
transform 1 0 3880 0 1 1010
box 0 0 16 200
use FILL  FILL_5_3_1
timestamp 1515852544
transform 1 0 3896 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_50
timestamp 1515852544
transform 1 0 3912 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_23
timestamp 1515852544
transform -1 0 4040 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_51
timestamp 1515852544
transform -1 0 4104 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_69
timestamp 1515852544
transform 1 0 4104 0 1 1010
box 0 0 64 200
use INVX1  INVX1_94
timestamp 1515852544
transform 1 0 4168 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_70
timestamp 1515852544
transform 1 0 4200 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_4
timestamp 1515852544
transform 1 0 4264 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_94
timestamp 1515852544
transform 1 0 4312 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_82
timestamp 1515852544
transform 1 0 4376 0 1 1010
box 0 0 192 200
use BUFX4  BUFX4_51
timestamp 1515852544
transform 1 0 4568 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_25
timestamp 1515852544
transform 1 0 4632 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_7
timestamp 1515852544
transform -1 0 4760 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_110
timestamp 1515852544
transform -1 0 4824 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_6
timestamp 1515852544
transform 1 0 4824 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_212
timestamp 1515852544
transform 1 0 4872 0 1 1010
box 0 0 64 200
use FILL  FILL_5_4_0
timestamp 1515852544
transform -1 0 4952 0 1 1010
box 0 0 16 200
use FILL  FILL_5_4_1
timestamp 1515852544
transform -1 0 4968 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_273
timestamp 1515852544
transform -1 0 5032 0 1 1010
box 0 0 64 200
use INVX1  INVX1_102
timestamp 1515852544
transform -1 0 5064 0 1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_125
timestamp 1515852544
transform -1 0 5128 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_81
timestamp 1515852544
transform -1 0 5176 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_115
timestamp 1515852544
transform 1 0 5176 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_11
timestamp 1515852544
transform 1 0 5240 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_272
timestamp 1515852544
transform -1 0 5368 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_84
timestamp 1515852544
transform 1 0 5368 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_67
timestamp 1515852544
transform 1 0 5416 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_83
timestamp 1515852544
transform -1 0 5528 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_276
timestamp 1515852544
transform 1 0 5528 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_275
timestamp 1515852544
transform -1 0 5656 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_136
timestamp 1515852544
transform -1 0 5736 0 1 1010
box 0 0 80 200
use NAND3X1  NAND3X1_66
timestamp 1515852544
transform 1 0 5736 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_37
timestamp 1515852544
transform -1 0 5848 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_121
timestamp 1515852544
transform -1 0 5896 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_148
timestamp 1515852544
transform 1 0 5896 0 1 1010
box 0 0 64 200
use FILL  FILL_5_5_0
timestamp 1515852544
transform -1 0 5976 0 1 1010
box 0 0 16 200
use FILL  FILL_5_5_1
timestamp 1515852544
transform -1 0 5992 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_7
timestamp 1515852544
transform -1 0 6040 0 1 1010
box 0 0 48 200
use INVX8  INVX8_13
timestamp 1515852544
transform 1 0 6040 0 1 1010
box 0 0 80 200
use INVX1  INVX1_71
timestamp 1515852544
transform 1 0 6120 0 1 1010
box 0 0 32 200
use OAI22X1  OAI22X1_18
timestamp 1515852544
transform 1 0 6152 0 1 1010
box 0 0 80 200
use INVX1  INVX1_72
timestamp 1515852544
transform -1 0 6264 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_134
timestamp 1515852544
transform 1 0 6264 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_31
timestamp 1515852544
transform 1 0 6328 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_17
timestamp 1515852544
transform 1 0 6376 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_136
timestamp 1515852544
transform -1 0 6504 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_10
timestamp 1515852544
transform -1 0 6568 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_146
timestamp 1515852544
transform -1 0 6760 0 1 1010
box 0 0 192 200
use FILL  FILL_6_1
timestamp 1515852544
transform 1 0 6760 0 1 1010
box 0 0 16 200
use FILL  FILL_6_2
timestamp 1515852544
transform 1 0 6776 0 1 1010
box 0 0 16 200
use FILL  FILL_6_3
timestamp 1515852544
transform 1 0 6792 0 1 1010
box 0 0 16 200
use INVX1  INVX1_21
timestamp 1515852544
transform 1 0 8 0 -1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_53
timestamp 1515852544
transform -1 0 88 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_60
timestamp 1515852544
transform 1 0 88 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_205
timestamp 1515852544
transform -1 0 200 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_218
timestamp 1515852544
transform 1 0 200 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_17
timestamp 1515852544
transform 1 0 264 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_219
timestamp 1515852544
transform -1 0 408 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_31
timestamp 1515852544
transform 1 0 408 0 -1 1010
box 0 0 192 200
use NAND3X1  NAND3X1_119
timestamp 1515852544
transform -1 0 664 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_67
timestamp 1515852544
transform 1 0 664 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_247
timestamp 1515852544
transform -1 0 776 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_22
timestamp 1515852544
transform 1 0 776 0 -1 1010
box 0 0 80 200
use FILL  FILL_4_0_0
timestamp 1515852544
transform -1 0 872 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1515852544
transform -1 0 888 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_249
timestamp 1515852544
transform -1 0 952 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_251
timestamp 1515852544
transform 1 0 952 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_252
timestamp 1515852544
transform -1 0 1080 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_245
timestamp 1515852544
transform -1 0 1144 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_118
timestamp 1515852544
transform -1 0 1208 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_51
timestamp 1515852544
transform 1 0 1208 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_198
timestamp 1515852544
transform -1 0 1320 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_215
timestamp 1515852544
transform -1 0 1384 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_254
timestamp 1515852544
transform 1 0 1384 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_256
timestamp 1515852544
transform 1 0 1448 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_73
timestamp 1515852544
transform -1 0 1560 0 -1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_25
timestamp 1515852544
transform 1 0 1560 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_258
timestamp 1515852544
transform -1 0 1704 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_255
timestamp 1515852544
transform -1 0 1768 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_72
timestamp 1515852544
transform -1 0 1816 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_1_0
timestamp 1515852544
transform 1 0 1816 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1515852544
transform 1 0 1832 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_222
timestamp 1515852544
transform 1 0 1848 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_70
timestamp 1515852544
transform 1 0 1912 0 -1 1010
box 0 0 192 200
use AOI22X1  AOI22X1_121
timestamp 1515852544
transform -1 0 2184 0 -1 1010
box 0 0 80 200
use BUFX4  BUFX4_116
timestamp 1515852544
transform 1 0 2184 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_94
timestamp 1515852544
transform -1 0 2312 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_45
timestamp 1515852544
transform 1 0 2312 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_227
timestamp 1515852544
transform -1 0 2424 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_99
timestamp 1515852544
transform -1 0 2456 0 -1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_117
timestamp 1515852544
transform -1 0 2520 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_63
timestamp 1515852544
transform -1 0 2568 0 -1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_27
timestamp 1515852544
transform 1 0 2568 0 -1 1010
box 0 0 192 200
use BUFX4  BUFX4_207
timestamp 1515852544
transform 1 0 2760 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_207
timestamp 1515852544
transform 1 0 2824 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_2_0
timestamp 1515852544
transform 1 0 2888 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1515852544
transform 1 0 2904 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_208
timestamp 1515852544
transform 1 0 2920 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_54
timestamp 1515852544
transform -1 0 3032 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_210
timestamp 1515852544
transform 1 0 3032 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_15
timestamp 1515852544
transform -1 0 3176 0 -1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_55
timestamp 1515852544
transform 1 0 3176 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_209
timestamp 1515852544
transform -1 0 3288 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_68
timestamp 1515852544
transform 1 0 3288 0 -1 1010
box 0 0 32 200
use OAI22X1  OAI22X1_17
timestamp 1515852544
transform -1 0 3400 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_23
timestamp 1515852544
transform 1 0 3400 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_298
timestamp 1515852544
transform 1 0 3464 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_199
timestamp 1515852544
transform 1 0 3512 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_306
timestamp 1515852544
transform 1 0 3576 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_52
timestamp 1515852544
transform 1 0 3624 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_90
timestamp 1515852544
transform -1 0 3752 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_77
timestamp 1515852544
transform 1 0 3752 0 -1 1010
box 0 0 192 200
use FILL  FILL_4_3_0
timestamp 1515852544
transform 1 0 3944 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_1
timestamp 1515852544
transform 1 0 3960 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_54
timestamp 1515852544
transform 1 0 3976 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_178
timestamp 1515852544
transform 1 0 4040 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_71
timestamp 1515852544
transform 1 0 4120 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_10
timestamp 1515852544
transform -1 0 4248 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_182
timestamp 1515852544
transform 1 0 4248 0 -1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_5
timestamp 1515852544
transform 1 0 4328 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_72
timestamp 1515852544
transform -1 0 4440 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_63
timestamp 1515852544
transform -1 0 4472 0 -1 1010
box 0 0 32 200
use OAI22X1  OAI22X1_15
timestamp 1515852544
transform -1 0 4552 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_232
timestamp 1515852544
transform -1 0 4616 0 -1 1010
box 0 0 64 200
use INVX8  INVX8_5
timestamp 1515852544
transform -1 0 4696 0 -1 1010
box 0 0 80 200
use BUFX4  BUFX4_200
timestamp 1515852544
transform 1 0 4696 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_268
timestamp 1515852544
transform -1 0 4824 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_70
timestamp 1515852544
transform -1 0 4856 0 -1 1010
box 0 0 32 200
use AND2X2  AND2X2_22
timestamp 1515852544
transform 1 0 4856 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_4_0
timestamp 1515852544
transform 1 0 4920 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_4_1
timestamp 1515852544
transform 1 0 4936 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_82
timestamp 1515852544
transform 1 0 4952 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_16
timestamp 1515852544
transform -1 0 5064 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_17
timestamp 1515852544
transform -1 0 5128 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_274
timestamp 1515852544
transform -1 0 5192 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_278
timestamp 1515852544
transform 1 0 5192 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_18
timestamp 1515852544
transform 1 0 5256 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_277
timestamp 1515852544
transform 1 0 5320 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_24
timestamp 1515852544
transform 1 0 5384 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_280
timestamp 1515852544
transform 1 0 5448 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_324
timestamp 1515852544
transform 1 0 5512 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_370
timestamp 1515852544
transform 1 0 5576 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_321
timestamp 1515852544
transform 1 0 5640 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_322
timestamp 1515852544
transform -1 0 5768 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_137
timestamp 1515852544
transform -1 0 5848 0 -1 1010
box 0 0 80 200
use OAI21X1  OAI21X1_75
timestamp 1515852544
transform 1 0 5848 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_5_0
timestamp 1515852544
transform -1 0 5928 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_5_1
timestamp 1515852544
transform -1 0 5944 0 -1 1010
box 0 0 16 200
use AND2X2  AND2X2_11
timestamp 1515852544
transform -1 0 6008 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_77
timestamp 1515852544
transform 1 0 6008 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_6
timestamp 1515852544
transform -1 0 6120 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_77
timestamp 1515852544
transform -1 0 6184 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_81
timestamp 1515852544
transform -1 0 6248 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_132
timestamp 1515852544
transform 1 0 6248 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_133
timestamp 1515852544
transform -1 0 6376 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_30
timestamp 1515852544
transform 1 0 6376 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_48
timestamp 1515852544
transform 1 0 6424 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_137
timestamp 1515852544
transform 1 0 6472 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_138
timestamp 1515852544
transform 1 0 6536 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1515852544
transform -1 0 6792 0 -1 1010
box 0 0 192 200
use FILL  FILL_5_1
timestamp 1515852544
transform -1 0 6808 0 -1 1010
box 0 0 16 200
use BUFX2  BUFX2_68
timestamp 1515852544
transform -1 0 56 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_5
timestamp 1515852544
transform -1 0 104 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_63
timestamp 1515852544
transform 1 0 104 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_115
timestamp 1515852544
transform 1 0 152 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_25
timestamp 1515852544
transform 1 0 216 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_216
timestamp 1515852544
transform -1 0 472 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_59
timestamp 1515852544
transform 1 0 472 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_217
timestamp 1515852544
transform -1 0 584 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_61
timestamp 1515852544
transform 1 0 584 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_221
timestamp 1515852544
transform -1 0 696 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_32
timestamp 1515852544
transform 1 0 696 0 1 610
box 0 0 192 200
use FILL  FILL_3_0_0
timestamp 1515852544
transform 1 0 888 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1515852544
transform 1 0 904 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_70
timestamp 1515852544
transform 1 0 920 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_120
timestamp 1515852544
transform -1 0 1032 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_71
timestamp 1515852544
transform -1 0 1080 0 1 610
box 0 0 48 200
use AOI22X1  AOI22X1_23
timestamp 1515852544
transform 1 0 1080 0 1 610
box 0 0 80 200
use INVX1  INVX1_57
timestamp 1515852544
transform 1 0 1160 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_253
timestamp 1515852544
transform -1 0 1256 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_250
timestamp 1515852544
transform -1 0 1320 0 1 610
box 0 0 64 200
use OAI22X1  OAI22X1_13
timestamp 1515852544
transform 1 0 1320 0 1 610
box 0 0 80 200
use INVX1  INVX1_58
timestamp 1515852544
transform -1 0 1432 0 1 610
box 0 0 32 200
use BUFX4  BUFX4_144
timestamp 1515852544
transform -1 0 1496 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_11
timestamp 1515852544
transform -1 0 1560 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_208
timestamp 1515852544
transform -1 0 1624 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_211
timestamp 1515852544
transform 1 0 1624 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_295
timestamp 1515852544
transform 1 0 1688 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_17
timestamp 1515852544
transform 1 0 1736 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_18
timestamp 1515852544
transform 1 0 1800 0 1 610
box 0 0 64 200
use FILL  FILL_3_1_0
timestamp 1515852544
transform -1 0 1880 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1515852544
transform -1 0 1896 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_296
timestamp 1515852544
transform -1 0 1944 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_86
timestamp 1515852544
transform 1 0 1944 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_16
timestamp 1515852544
transform 1 0 2008 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_19
timestamp 1515852544
transform -1 0 2136 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_171
timestamp 1515852544
transform -1 0 2216 0 1 610
box 0 0 80 200
use NAND2X1  NAND2X1_100
timestamp 1515852544
transform -1 0 2264 0 1 610
box 0 0 48 200
use AND2X2  AND2X2_25
timestamp 1515852544
transform -1 0 2328 0 1 610
box 0 0 64 200
use INVX1  INVX1_66
timestamp 1515852544
transform 1 0 2328 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_320
timestamp 1515852544
transform 1 0 2360 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_102
timestamp 1515852544
transform -1 0 2472 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_93
timestamp 1515852544
transform 1 0 2472 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_147
timestamp 1515852544
transform -1 0 2600 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_178
timestamp 1515852544
transform 1 0 2600 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_9
timestamp 1515852544
transform 1 0 2664 0 1 610
box 0 0 80 200
use NAND2X1  NAND2X1_45
timestamp 1515852544
transform -1 0 2792 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_176
timestamp 1515852544
transform -1 0 2856 0 1 610
box 0 0 64 200
use FILL  FILL_3_2_0
timestamp 1515852544
transform 1 0 2856 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1515852544
transform 1 0 2872 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_47
timestamp 1515852544
transform 1 0 2888 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_180
timestamp 1515852544
transform -1 0 3000 0 1 610
box 0 0 64 200
use INVX1  INVX1_67
timestamp 1515852544
transform 1 0 3000 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_297
timestamp 1515852544
transform 1 0 3032 0 1 610
box 0 0 48 200
use AOI22X1  AOI22X1_173
timestamp 1515852544
transform -1 0 3160 0 1 610
box 0 0 80 200
use OAI21X1  OAI21X1_22
timestamp 1515852544
transform 1 0 3160 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_20
timestamp 1515852544
transform 1 0 3224 0 1 610
box 0 0 64 200
use INVX1  INVX1_93
timestamp 1515852544
transform 1 0 3288 0 1 610
box 0 0 32 200
use BUFX4  BUFX4_145
timestamp 1515852544
transform 1 0 3320 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_67
timestamp 1515852544
transform -1 0 3432 0 1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_19
timestamp 1515852544
transform 1 0 3432 0 1 610
box 0 0 192 200
use BUFX4  BUFX4_202
timestamp 1515852544
transform 1 0 3624 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_336
timestamp 1515852544
transform -1 0 3752 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_331
timestamp 1515852544
transform 1 0 3752 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_7
timestamp 1515852544
transform -1 0 3880 0 1 610
box 0 0 64 200
use FILL  FILL_3_3_0
timestamp 1515852544
transform 1 0 3880 0 1 610
box 0 0 16 200
use FILL  FILL_3_3_1
timestamp 1515852544
transform 1 0 3896 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_28
timestamp 1515852544
transform 1 0 3912 0 1 610
box 0 0 192 200
use NAND2X1  NAND2X1_65
timestamp 1515852544
transform -1 0 4152 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_236
timestamp 1515852544
transform -1 0 4216 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_231
timestamp 1515852544
transform -1 0 4280 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_14
timestamp 1515852544
transform 1 0 4280 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_230
timestamp 1515852544
transform -1 0 4408 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_234
timestamp 1515852544
transform -1 0 4472 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_233
timestamp 1515852544
transform 1 0 4472 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_21
timestamp 1515852544
transform -1 0 4600 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_253
timestamp 1515852544
transform 1 0 4600 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_66
timestamp 1515852544
transform -1 0 4696 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_27
timestamp 1515852544
transform 1 0 4696 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_28
timestamp 1515852544
transform 1 0 4760 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1515852544
transform 1 0 4824 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_299
timestamp 1515852544
transform 1 0 4888 0 1 610
box 0 0 48 200
use FILL  FILL_3_4_0
timestamp 1515852544
transform -1 0 4952 0 1 610
box 0 0 16 200
use FILL  FILL_3_4_1
timestamp 1515852544
transform -1 0 4968 0 1 610
box 0 0 16 200
use OAI21X1  OAI21X1_29
timestamp 1515852544
transform -1 0 5032 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_9
timestamp 1515852544
transform -1 0 5096 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_25
timestamp 1515852544
transform -1 0 5160 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_203
timestamp 1515852544
transform 1 0 5160 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_104
timestamp 1515852544
transform 1 0 5224 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_281
timestamp 1515852544
transform -1 0 5336 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_325
timestamp 1515852544
transform 1 0 5336 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_26
timestamp 1515852544
transform 1 0 5400 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_326
timestamp 1515852544
transform 1 0 5464 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_103
timestamp 1515852544
transform -1 0 5576 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_22
timestamp 1515852544
transform -1 0 5640 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_371
timestamp 1515852544
transform 1 0 5640 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_327
timestamp 1515852544
transform 1 0 5704 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_28
timestamp 1515852544
transform 1 0 5768 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_372
timestamp 1515852544
transform 1 0 5832 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_76
timestamp 1515852544
transform 1 0 5896 0 1 610
box 0 0 64 200
use FILL  FILL_3_5_0
timestamp 1515852544
transform 1 0 5960 0 1 610
box 0 0 16 200
use FILL  FILL_3_5_1
timestamp 1515852544
transform 1 0 5976 0 1 610
box 0 0 16 200
use AOI21X1  AOI21X1_5
timestamp 1515852544
transform 1 0 5992 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_17
timestamp 1515852544
transform -1 0 6248 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_78
timestamp 1515852544
transform 1 0 6248 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_83
timestamp 1515852544
transform -1 0 6504 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_185
timestamp 1515852544
transform -1 0 6568 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_186
timestamp 1515852544
transform -1 0 6632 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_182
timestamp 1515852544
transform 1 0 6632 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_181
timestamp 1515852544
transform -1 0 6760 0 1 610
box 0 0 64 200
use FILL  FILL_4_1
timestamp 1515852544
transform 1 0 6760 0 1 610
box 0 0 16 200
use FILL  FILL_4_2
timestamp 1515852544
transform 1 0 6776 0 1 610
box 0 0 16 200
use FILL  FILL_4_3
timestamp 1515852544
transform 1 0 6792 0 1 610
box 0 0 16 200
use BUFX2  BUFX2_43
timestamp 1515852544
transform -1 0 56 0 -1 610
box 0 0 48 200
use INVX1  INVX1_22
timestamp 1515852544
transform 1 0 56 0 -1 610
box 0 0 32 200
use BUFX2  BUFX2_6
timestamp 1515852544
transform -1 0 136 0 -1 610
box 0 0 48 200
use NOR2X1  NOR2X1_64
timestamp 1515852544
transform 1 0 136 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_222
timestamp 1515852544
transform 1 0 184 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_62
timestamp 1515852544
transform -1 0 296 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_116
timestamp 1515852544
transform 1 0 296 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_18
timestamp 1515852544
transform 1 0 360 0 -1 610
box 0 0 80 200
use OAI21X1  OAI21X1_225
timestamp 1515852544
transform -1 0 504 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_220
timestamp 1515852544
transform -1 0 568 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_37
timestamp 1515852544
transform 1 0 568 0 -1 610
box 0 0 192 200
use AOI22X1  AOI22X1_28
timestamp 1515852544
transform 1 0 760 0 -1 610
box 0 0 80 200
use FILL  FILL_2_0_0
timestamp 1515852544
transform -1 0 856 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1515852544
transform -1 0 872 0 -1 610
box 0 0 16 200
use NAND3X1  NAND3X1_124
timestamp 1515852544
transform -1 0 936 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_78
timestamp 1515852544
transform 1 0 936 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_80
timestamp 1515852544
transform -1 0 1032 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_269
timestamp 1515852544
transform 1 0 1032 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_270
timestamp 1515852544
transform -1 0 1160 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_271
timestamp 1515852544
transform -1 0 1224 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_267
timestamp 1515852544
transform -1 0 1288 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_98
timestamp 1515852544
transform -1 0 1352 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_100
timestamp 1515852544
transform 1 0 1352 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_294
timestamp 1515852544
transform 1 0 1416 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_14
timestamp 1515852544
transform -1 0 1528 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_69
timestamp 1515852544
transform -1 0 1720 0 -1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1515852544
transform 1 0 1720 0 -1 610
box 0 0 192 200
use FILL  FILL_2_1_0
timestamp 1515852544
transform -1 0 1928 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1515852544
transform -1 0 1944 0 -1 610
box 0 0 16 200
use NAND3X1  NAND3X1_132
timestamp 1515852544
transform -1 0 2008 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_318
timestamp 1515852544
transform -1 0 2072 0 -1 610
box 0 0 64 200
use INVX1  INVX1_104
timestamp 1515852544
transform -1 0 2104 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_317
timestamp 1515852544
transform -1 0 2168 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_37
timestamp 1515852544
transform -1 0 2248 0 -1 610
box 0 0 80 200
use OAI21X1  OAI21X1_319
timestamp 1515852544
transform -1 0 2312 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_56
timestamp 1515852544
transform 1 0 2312 0 -1 610
box 0 0 48 200
use AND2X2  AND2X2_20
timestamp 1515852544
transform -1 0 2424 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_96
timestamp 1515852544
transform 1 0 2424 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_18
timestamp 1515852544
transform 1 0 2488 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_177
timestamp 1515852544
transform 1 0 2552 0 -1 610
box 0 0 64 200
use INVX1  INVX1_96
timestamp 1515852544
transform -1 0 2648 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_110
timestamp 1515852544
transform -1 0 2712 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_93
timestamp 1515852544
transform 1 0 2712 0 -1 610
box 0 0 192 200
use FILL  FILL_2_2_0
timestamp 1515852544
transform -1 0 2920 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1515852544
transform -1 0 2936 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_71
timestamp 1515852544
transform -1 0 3128 0 -1 610
box 0 0 192 200
use NAND3X1  NAND3X1_87
timestamp 1515852544
transform 1 0 3128 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_8
timestamp 1515852544
transform 1 0 3192 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_21
timestamp 1515852544
transform 1 0 3256 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_18
timestamp 1515852544
transform 1 0 3320 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_328
timestamp 1515852544
transform 1 0 3512 0 -1 610
box 0 0 64 200
use INVX1  INVX1_105
timestamp 1515852544
transform 1 0 3576 0 -1 610
box 0 0 32 200
use AOI21X1  AOI21X1_24
timestamp 1515852544
transform -1 0 3672 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_330
timestamp 1515852544
transform 1 0 3672 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_329
timestamp 1515852544
transform -1 0 3800 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_242
timestamp 1515852544
transform -1 0 3864 0 -1 610
box 0 0 64 200
use FILL  FILL_2_3_0
timestamp 1515852544
transform 1 0 3864 0 -1 610
box 0 0 16 200
use FILL  FILL_2_3_1
timestamp 1515852544
transform 1 0 3880 0 -1 610
box 0 0 16 200
use AOI22X1  AOI22X1_38
timestamp 1515852544
transform 1 0 3896 0 -1 610
box 0 0 80 200
use OAI21X1  OAI21X1_332
timestamp 1515852544
transform 1 0 3976 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_39
timestamp 1515852544
transform 1 0 4040 0 -1 610
box 0 0 80 200
use OAI21X1  OAI21X1_333
timestamp 1515852544
transform -1 0 4184 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_143
timestamp 1515852544
transform -1 0 4264 0 -1 610
box 0 0 80 200
use AOI21X1  AOI21X1_25
timestamp 1515852544
transform -1 0 4328 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_152
timestamp 1515852544
transform 1 0 4328 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_151
timestamp 1515852544
transform 1 0 4392 0 -1 610
box 0 0 80 200
use AOI21X1  AOI21X1_20
timestamp 1515852544
transform -1 0 4536 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_148
timestamp 1515852544
transform -1 0 4616 0 -1 610
box 0 0 80 200
use NAND3X1  NAND3X1_69
timestamp 1515852544
transform 1 0 4616 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_40
timestamp 1515852544
transform -1 0 4728 0 -1 610
box 0 0 48 200
use OAI22X1  OAI22X1_20
timestamp 1515852544
transform -1 0 4808 0 -1 610
box 0 0 80 200
use NAND2X1  NAND2X1_260
timestamp 1515852544
transform -1 0 4856 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_30
timestamp 1515852544
transform -1 0 4920 0 -1 610
box 0 0 64 200
use FILL  FILL_2_4_0
timestamp 1515852544
transform -1 0 4936 0 -1 610
box 0 0 16 200
use FILL  FILL_2_4_1
timestamp 1515852544
transform -1 0 4952 0 -1 610
box 0 0 16 200
use OR2X2  OR2X2_4
timestamp 1515852544
transform -1 0 5016 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1515852544
transform 1 0 5016 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_300
timestamp 1515852544
transform -1 0 5128 0 -1 610
box 0 0 48 200
use AOI22X1  AOI22X1_147
timestamp 1515852544
transform -1 0 5208 0 -1 610
box 0 0 80 200
use BUFX4  BUFX4_71
timestamp 1515852544
transform -1 0 5272 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_39
timestamp 1515852544
transform 1 0 5272 0 -1 610
box 0 0 192 200
use BUFX4  BUFX4_150
timestamp 1515852544
transform -1 0 5528 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_367
timestamp 1515852544
transform 1 0 5528 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_369
timestamp 1515852544
transform -1 0 5656 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_122
timestamp 1515852544
transform 1 0 5656 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_373
timestamp 1515852544
transform 1 0 5704 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_26
timestamp 1515852544
transform 1 0 5768 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_189
timestamp 1515852544
transform -1 0 5896 0 -1 610
box 0 0 64 200
use FILL  FILL_2_5_0
timestamp 1515852544
transform -1 0 5912 0 -1 610
box 0 0 16 200
use FILL  FILL_2_5_1
timestamp 1515852544
transform -1 0 5928 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_50
timestamp 1515852544
transform -1 0 6120 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_73
timestamp 1515852544
transform 1 0 6120 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_74
timestamp 1515852544
transform -1 0 6248 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_183
timestamp 1515852544
transform 1 0 6248 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_184
timestamp 1515852544
transform 1 0 6312 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_13
timestamp 1515852544
transform 1 0 6376 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_49
timestamp 1515852544
transform 1 0 6440 0 -1 610
box 0 0 48 200
use AND2X2  AND2X2_19
timestamp 1515852544
transform 1 0 6488 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_94
timestamp 1515852544
transform 1 0 6552 0 -1 610
box 0 0 192 200
use INVX1  INVX1_10
timestamp 1515852544
transform -1 0 6776 0 -1 610
box 0 0 32 200
use FILL  FILL_3_1
timestamp 1515852544
transform -1 0 6792 0 -1 610
box 0 0 16 200
use FILL  FILL_3_2
timestamp 1515852544
transform -1 0 6808 0 -1 610
box 0 0 16 200
use INVX8  INVX8_4
timestamp 1515852544
transform 1 0 8 0 1 210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_26
timestamp 1515852544
transform -1 0 280 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_310
timestamp 1515852544
transform -1 0 344 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_36
timestamp 1515852544
transform -1 0 424 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_308
timestamp 1515852544
transform -1 0 488 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_94
timestamp 1515852544
transform -1 0 536 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_309
timestamp 1515852544
transform -1 0 600 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_307
timestamp 1515852544
transform -1 0 664 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_115
timestamp 1515852544
transform 1 0 664 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_355
timestamp 1515852544
transform 1 0 712 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_354
timestamp 1515852544
transform -1 0 840 0 1 210
box 0 0 64 200
use FILL  FILL_1_0_0
timestamp 1515852544
transform 1 0 840 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1515852544
transform 1 0 856 0 1 210
box 0 0 16 200
use OAI21X1  OAI21X1_264
timestamp 1515852544
transform 1 0 872 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_76
timestamp 1515852544
transform -1 0 984 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_266
timestamp 1515852544
transform 1 0 984 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_27
timestamp 1515852544
transform -1 0 1128 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_263
timestamp 1515852544
transform -1 0 1192 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_15
timestamp 1515852544
transform 1 0 1192 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_170
timestamp 1515852544
transform -1 0 1336 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_12
timestamp 1515852544
transform 1 0 1336 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_293
timestamp 1515852544
transform -1 0 1448 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_84
timestamp 1515852544
transform 1 0 1448 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_104
timestamp 1515852544
transform 1 0 1512 0 1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_57
timestamp 1515852544
transform -1 0 1896 0 1 210
box 0 0 192 200
use FILL  FILL_1_1_0
timestamp 1515852544
transform -1 0 1912 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1515852544
transform -1 0 1928 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_69
timestamp 1515852544
transform -1 0 1992 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_364
timestamp 1515852544
transform -1 0 2056 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_27
timestamp 1515852544
transform -1 0 2120 0 1 210
box 0 0 64 200
use INVX1  INVX1_106
timestamp 1515852544
transform -1 0 2152 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_363
timestamp 1515852544
transform -1 0 2216 0 1 210
box 0 0 64 200
use INVX1  INVX1_62
timestamp 1515852544
transform 1 0 2216 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_374
timestamp 1515852544
transform 1 0 2248 0 1 210
box 0 0 64 200
use INVX1  INVX1_107
timestamp 1515852544
transform 1 0 2312 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_375
timestamp 1515852544
transform -1 0 2408 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_283
timestamp 1515852544
transform 1 0 2408 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_282
timestamp 1515852544
transform 1 0 2472 0 1 210
box 0 0 64 200
use INVX1  INVX1_103
timestamp 1515852544
transform 1 0 2536 0 1 210
box 0 0 32 200
use AOI22X1  AOI22X1_29
timestamp 1515852544
transform -1 0 2648 0 1 210
box 0 0 80 200
use AOI22X1  AOI22X1_144
timestamp 1515852544
transform -1 0 2728 0 1 210
box 0 0 80 200
use AOI22X1  AOI22X1_48
timestamp 1515852544
transform 1 0 2728 0 1 210
box 0 0 80 200
use AOI21X1  AOI21X1_27
timestamp 1515852544
transform -1 0 2872 0 1 210
box 0 0 64 200
use FILL  FILL_1_2_0
timestamp 1515852544
transform 1 0 2872 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1515852544
transform 1 0 2888 0 1 210
box 0 0 16 200
use OAI21X1  OAI21X1_286
timestamp 1515852544
transform 1 0 2904 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_287
timestamp 1515852544
transform -1 0 3032 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_30
timestamp 1515852544
transform -1 0 3112 0 1 210
box 0 0 80 200
use AOI21X1  AOI21X1_15
timestamp 1515852544
transform 1 0 3112 0 1 210
box 0 0 64 200
use INVX1  INVX1_100
timestamp 1515852544
transform -1 0 3208 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_240
timestamp 1515852544
transform 1 0 3208 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_238
timestamp 1515852544
transform 1 0 3272 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_20
timestamp 1515852544
transform 1 0 3336 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_237
timestamp 1515852544
transform -1 0 3480 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_243
timestamp 1515852544
transform 1 0 3480 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_21
timestamp 1515852544
transform 1 0 3544 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_381
timestamp 1515852544
transform 1 0 3624 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_380
timestamp 1515852544
transform 1 0 3688 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_49
timestamp 1515852544
transform 1 0 3752 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_382
timestamp 1515852544
transform -1 0 3896 0 1 210
box 0 0 64 200
use FILL  FILL_1_3_0
timestamp 1515852544
transform -1 0 3912 0 1 210
box 0 0 16 200
use FILL  FILL_1_3_1
timestamp 1515852544
transform -1 0 3928 0 1 210
box 0 0 16 200
use OAI21X1  OAI21X1_378
timestamp 1515852544
transform -1 0 3992 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_8
timestamp 1515852544
transform -1 0 4056 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_52
timestamp 1515852544
transform 1 0 4056 0 1 210
box 0 0 192 200
use INVX1  INVX1_108
timestamp 1515852544
transform -1 0 4280 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_376
timestamp 1515852544
transform 1 0 4280 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_72
timestamp 1515852544
transform 1 0 4344 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_195
timestamp 1515852544
transform 1 0 4536 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_196
timestamp 1515852544
transform -1 0 4664 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_80
timestamp 1515852544
transform 1 0 4664 0 1 210
box 0 0 64 200
use INVX1  INVX1_79
timestamp 1515852544
transform -1 0 4760 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_82
timestamp 1515852544
transform 1 0 4760 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_194
timestamp 1515852544
transform 1 0 4824 0 1 210
box 0 0 64 200
use FILL  FILL_1_4_0
timestamp 1515852544
transform -1 0 4904 0 1 210
box 0 0 16 200
use FILL  FILL_1_4_1
timestamp 1515852544
transform -1 0 4920 0 1 210
box 0 0 16 200
use OAI21X1  OAI21X1_81
timestamp 1515852544
transform -1 0 4984 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_84
timestamp 1515852544
transform 1 0 4984 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_83
timestamp 1515852544
transform -1 0 5112 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_184
timestamp 1515852544
transform -1 0 5192 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_86
timestamp 1515852544
transform 1 0 5192 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_87
timestamp 1515852544
transform -1 0 5320 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_185
timestamp 1515852544
transform -1 0 5400 0 1 210
box 0 0 80 200
use AOI21X1  AOI21X1_6
timestamp 1515852544
transform -1 0 5464 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_187
timestamp 1515852544
transform 1 0 5464 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_188
timestamp 1515852544
transform -1 0 5592 0 1 210
box 0 0 64 200
use INVX1  INVX1_78
timestamp 1515852544
transform -1 0 5624 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_191
timestamp 1515852544
transform 1 0 5624 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_192
timestamp 1515852544
transform 1 0 5688 0 1 210
box 0 0 64 200
use INVX8  INVX8_11
timestamp 1515852544
transform 1 0 5752 0 1 210
box 0 0 80 200
use INVX8  INVX8_12
timestamp 1515852544
transform 1 0 5832 0 1 210
box 0 0 80 200
use NAND2X1  NAND2X1_259
timestamp 1515852544
transform -1 0 5960 0 1 210
box 0 0 48 200
use FILL  FILL_1_5_0
timestamp 1515852544
transform 1 0 5960 0 1 210
box 0 0 16 200
use FILL  FILL_1_5_1
timestamp 1515852544
transform 1 0 5976 0 1 210
box 0 0 16 200
use NOR2X1  NOR2X1_48
timestamp 1515852544
transform 1 0 5992 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_238
timestamp 1515852544
transform -1 0 6088 0 1 210
box 0 0 48 200
use AOI21X1  AOI21X1_46
timestamp 1515852544
transform 1 0 6088 0 1 210
box 0 0 64 200
use INVX1  INVX1_7
timestamp 1515852544
transform -1 0 6184 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1515852544
transform -1 0 6376 0 1 210
box 0 0 192 200
use INVX1  INVX1_6
timestamp 1515852544
transform 1 0 6376 0 1 210
box 0 0 32 200
use NOR2X1  NOR2X1_49
timestamp 1515852544
transform 1 0 6408 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_20
timestamp 1515852544
transform 1 0 6456 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_56
timestamp 1515852544
transform 1 0 6504 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_52
timestamp 1515852544
transform -1 0 6600 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_23
timestamp 1515852544
transform 1 0 6600 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_71
timestamp 1515852544
transform 1 0 6648 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_54
timestamp 1515852544
transform -1 0 6744 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_281
timestamp 1515852544
transform -1 0 6792 0 1 210
box 0 0 48 200
use FILL  FILL_2_1
timestamp 1515852544
transform 1 0 6792 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_72
timestamp 1515852544
transform -1 0 56 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_32
timestamp 1515852544
transform -1 0 104 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_53
timestamp 1515852544
transform 1 0 104 0 -1 210
box 0 0 48 200
use INVX1  INVX1_11
timestamp 1515852544
transform -1 0 184 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_60
timestamp 1515852544
transform -1 0 232 0 -1 210
box 0 0 48 200
use INVX1  INVX1_18
timestamp 1515852544
transform -1 0 264 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_2
timestamp 1515852544
transform 1 0 264 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_41
timestamp 1515852544
transform 1 0 312 0 -1 210
box 0 0 48 200
use INVX8  INVX8_3
timestamp 1515852544
transform -1 0 440 0 -1 210
box 0 0 80 200
use NAND3X1  NAND3X1_131
timestamp 1515852544
transform -1 0 504 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_95
timestamp 1515852544
transform 1 0 504 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_14
timestamp 1515852544
transform 1 0 552 0 -1 210
box 0 0 192 200
use FILL  FILL_0_0_0
timestamp 1515852544
transform -1 0 760 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1515852544
transform -1 0 776 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_47
timestamp 1515852544
transform -1 0 968 0 -1 210
box 0 0 192 200
use NAND3X1  NAND3X1_137
timestamp 1515852544
transform -1 0 1032 0 -1 210
box 0 0 64 200
use AOI22X1  AOI22X1_44
timestamp 1515852544
transform 1 0 1032 0 -1 210
box 0 0 80 200
use OAI21X1  OAI21X1_358
timestamp 1515852544
transform -1 0 1176 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_116
timestamp 1515852544
transform 1 0 1176 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_356
timestamp 1515852544
transform -1 0 1288 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_265
timestamp 1515852544
transform -1 0 1352 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_77
timestamp 1515852544
transform -1 0 1400 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_123
timestamp 1515852544
transform 1 0 1400 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_36
timestamp 1515852544
transform 1 0 1464 0 -1 210
box 0 0 192 200
use AOI22X1  AOI22X1_118
timestamp 1515852544
transform 1 0 1656 0 -1 210
box 0 0 80 200
use BUFX4  BUFX4_99
timestamp 1515852544
transform -1 0 1800 0 -1 210
box 0 0 64 200
use INVX8  INVX8_9
timestamp 1515852544
transform 1 0 1800 0 -1 210
box 0 0 80 200
use FILL  FILL_0_1_0
timestamp 1515852544
transform -1 0 1896 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1515852544
transform -1 0 1912 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_66
timestamp 1515852544
transform -1 0 1960 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_31
timestamp 1515852544
transform -1 0 2008 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_49
timestamp 1515852544
transform 1 0 2008 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_119
timestamp 1515852544
transform 1 0 2200 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_139
timestamp 1515852544
transform 1 0 2248 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_365
timestamp 1515852544
transform -1 0 2376 0 -1 210
box 0 0 64 200
use AOI22X1  AOI22X1_47
timestamp 1515852544
transform 1 0 2376 0 -1 210
box 0 0 80 200
use NAND2X1  NAND2X1_120
timestamp 1515852544
transform 1 0 2456 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_366
timestamp 1515852544
transform -1 0 2568 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_97
timestamp 1515852544
transform 1 0 2568 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_40
timestamp 1515852544
transform -1 0 2824 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_284
timestamp 1515852544
transform -1 0 2888 0 -1 210
box 0 0 64 200
use FILL  FILL_0_2_0
timestamp 1515852544
transform -1 0 2904 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1515852544
transform -1 0 2920 0 -1 210
box 0 0 16 200
use AOI21X1  AOI21X1_19
timestamp 1515852544
transform -1 0 2984 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_377
timestamp 1515852544
transform 1 0 2984 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_51
timestamp 1515852544
transform -1 0 3240 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_190
timestamp 1515852544
transform 1 0 3240 0 -1 210
box 0 0 48 200
use OR2X2  OR2X2_6
timestamp 1515852544
transform 1 0 3288 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_285
timestamp 1515852544
transform -1 0 3416 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_288
timestamp 1515852544
transform 1 0 3416 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_29
timestamp 1515852544
transform 1 0 3480 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_41
timestamp 1515852544
transform 1 0 3672 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_8
timestamp 1515852544
transform 1 0 3864 0 -1 210
box 0 0 48 200
use FILL  FILL_0_3_0
timestamp 1515852544
transform 1 0 3912 0 -1 210
box 0 0 16 200
use FILL  FILL_0_3_1
timestamp 1515852544
transform 1 0 3928 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_45
timestamp 1515852544
transform 1 0 3944 0 -1 210
box 0 0 48 200
use OR2X2  OR2X2_5
timestamp 1515852544
transform 1 0 3992 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_241
timestamp 1515852544
transform -1 0 4120 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_244
timestamp 1515852544
transform 1 0 4120 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_30
timestamp 1515852544
transform 1 0 4184 0 -1 210
box 0 0 192 200
use INVX1  INVX1_101
timestamp 1515852544
transform -1 0 4408 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_239
timestamp 1515852544
transform -1 0 4472 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_242
timestamp 1515852544
transform -1 0 4520 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_44
timestamp 1515852544
transform -1 0 4584 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_245
timestamp 1515852544
transform -1 0 4632 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_96
timestamp 1515852544
transform -1 0 4824 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_197
timestamp 1515852544
transform -1 0 4888 0 -1 210
box 0 0 64 200
use FILL  FILL_0_4_0
timestamp 1515852544
transform 1 0 4888 0 -1 210
box 0 0 16 200
use FILL  FILL_0_4_1
timestamp 1515852544
transform 1 0 4904 0 -1 210
box 0 0 16 200
use AOI22X1  AOI22X1_11
timestamp 1515852544
transform 1 0 4920 0 -1 210
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_84
timestamp 1515852544
transform 1 0 5000 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_85
timestamp 1515852544
transform -1 0 5384 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_88
timestamp 1515852544
transform -1 0 5448 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_3
timestamp 1515852544
transform 1 0 5448 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_85
timestamp 1515852544
transform -1 0 5576 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_193
timestamp 1515852544
transform 1 0 5576 0 -1 210
box 0 0 64 200
use AOI22X1  AOI22X1_10
timestamp 1515852544
transform 1 0 5640 0 -1 210
box 0 0 80 200
use INVX1  INVX1_97
timestamp 1515852544
transform 1 0 5720 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_95
timestamp 1515852544
transform 1 0 5752 0 -1 210
box 0 0 192 200
use FILL  FILL_0_5_0
timestamp 1515852544
transform -1 0 5960 0 -1 210
box 0 0 16 200
use FILL  FILL_0_5_1
timestamp 1515852544
transform -1 0 5976 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_261
timestamp 1515852544
transform -1 0 6024 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_46
timestamp 1515852544
transform -1 0 6088 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_73
timestamp 1515852544
transform -1 0 6136 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_33
timestamp 1515852544
transform -1 0 6184 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_54
timestamp 1515852544
transform -1 0 6232 0 -1 210
box 0 0 48 200
use INVX1  INVX1_12
timestamp 1515852544
transform -1 0 6264 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_100
timestamp 1515852544
transform 1 0 6264 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_168
timestamp 1515852544
transform 1 0 6456 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_62
timestamp 1515852544
transform 1 0 6648 0 -1 210
box 0 0 48 200
use INVX8  INVX8_8
timestamp 1515852544
transform 1 0 6696 0 -1 210
box 0 0 80 200
use FILL  FILL_1_1
timestamp 1515852544
transform -1 0 6792 0 -1 210
box 0 0 16 200
use FILL  FILL_1_2
timestamp 1515852544
transform -1 0 6808 0 -1 210
box 0 0 16 200
<< labels >>
flabel space 1028 42 1036 136 6 FreeSans 48 0 0 0 vdd
port 0 nsew
flabel space 2068 42 2076 136 6 FreeSans 48 0 0 0 gnd
port 1 nsew
flabel metal3 -48 1460 -48 1460 7 FreeSans 48 0 0 0 IDATA_CORE_out<0>
port 2 nsew
flabel metal2 176 4860 176 4860 3 FreeSans 48 90 0 0 IDATA_CORE_out<1>
port 3 nsew
flabel metal3 6864 560 6864 560 3 FreeSans 48 0 0 0 IDATA_CORE_out<2>
port 4 nsew
flabel metal2 176 -40 176 -40 7 FreeSans 48 270 0 0 IDATA_CORE_out<3>
port 5 nsew
flabel metal2 6256 -40 6256 -40 7 FreeSans 48 270 0 0 IDATA_CORE_out<4>
port 6 nsew
flabel metal2 224 4860 224 4860 3 FreeSans 48 90 0 0 IDATA_CORE_out<5>
port 7 nsew
flabel metal3 6864 3800 6864 3800 3 FreeSans 48 0 0 0 IDATA_CORE_out<6>
port 8 nsew
flabel metal2 704 4860 704 4860 3 FreeSans 48 90 0 0 IDATA_CORE_out<7>
port 9 nsew
flabel metal2 400 4860 400 4860 3 FreeSans 48 90 0 0 IDATA_CORE_out<8>
port 10 nsew
flabel metal2 256 -40 256 -40 7 FreeSans 48 270 0 0 IDATA_CORE_out<9>
port 11 nsew
flabel metal2 6752 4860 6752 4860 3 FreeSans 48 90 0 0 IDATA_CORE_out<10>
port 12 nsew
flabel metal2 960 4860 960 4860 3 FreeSans 48 90 0 0 IDATA_CORE_out<11>
port 13 nsew
flabel metal3 -48 960 -48 960 7 FreeSans 48 0 0 0 IDATA_CORE_out<12>
port 14 nsew
flabel metal3 -48 560 -48 560 7 FreeSans 48 0 0 0 IDATA_CORE_out<13>
port 15 nsew
flabel metal3 -48 4260 -48 4260 7 FreeSans 48 0 0 0 IDATA_CORE_out<14>
port 16 nsew
flabel metal2 3872 -40 3872 -40 7 FreeSans 48 270 0 0 IDATA_CORE_out<15>
port 17 nsew
flabel metal2 4464 -40 4464 -40 7 FreeSans 48 270 0 0 CORE_PC_ctrl<0>
port 18 nsew
flabel metal2 6176 -40 6176 -40 7 FreeSans 48 270 0 0 CORE_PC_ctrl<1>
port 19 nsew
flabel metal2 1504 4860 1504 4860 3 FreeSans 48 90 0 0 CORE_STACK_ctrl<0>
port 20 nsew
flabel metal2 1728 4860 1728 4860 3 FreeSans 48 90 0 0 CORE_STACK_ctrl<1>
port 21 nsew
flabel metal3 -48 2940 -48 2940 7 FreeSans 48 0 0 0 ULA_OUT<0>
port 22 nsew
flabel metal3 -48 1360 -48 1360 7 FreeSans 48 0 0 0 ULA_OUT<1>
port 23 nsew
flabel metal2 3248 -40 3248 -40 7 FreeSans 48 270 0 0 ULA_OUT<2>
port 24 nsew
flabel metal2 3504 4860 3504 4860 3 FreeSans 48 90 0 0 ULA_OUT<3>
port 25 nsew
flabel metal2 4512 -40 4512 -40 7 FreeSans 48 270 0 0 ULA_OUT<4>
port 26 nsew
flabel metal2 4624 -40 4624 -40 7 FreeSans 48 270 0 0 ULA_OUT<5>
port 27 nsew
flabel metal2 4560 -40 4560 -40 7 FreeSans 48 270 0 0 ULA_OUT<6>
port 28 nsew
flabel metal2 6032 -40 6032 -40 7 FreeSans 48 270 0 0 ULA_OUT<7>
port 29 nsew
flabel metal2 5952 -40 5952 -40 7 FreeSans 48 270 0 0 ULA_OUT<8>
port 30 nsew
flabel metal2 6000 -40 6000 -40 7 FreeSans 48 270 0 0 ULA_OUT<9>
port 31 nsew
flabel metal2 784 4860 784 4860 3 FreeSans 48 90 0 0 INTERRUPT_ch<0>
port 32 nsew
flabel metal3 -48 1500 -48 1500 7 FreeSans 48 0 0 0 INTERRUPT_ch<1>
port 33 nsew
flabel metal2 896 4860 896 4860 3 FreeSans 48 90 0 0 INTERRUPT_ch<2>
port 34 nsew
flabel metal3 -48 1540 -48 1540 7 FreeSans 48 0 0 0 INTERRUPT_ch<3>
port 35 nsew
flabel metal2 432 -40 432 -40 7 FreeSans 48 270 0 0 INTERRUPT_ch<4>
port 36 nsew
flabel metal3 -48 320 -48 320 7 FreeSans 48 0 0 0 INTERRUPT_ch<5>
port 37 nsew
flabel metal3 6864 2960 6864 2960 3 FreeSans 48 0 0 0 INTERRUPT_ch<6>
port 38 nsew
flabel metal3 6864 280 6864 280 3 FreeSans 48 0 0 0 INTERRUPT_ch<7>
port 39 nsew
flabel metal2 4432 -40 4432 -40 7 FreeSans 48 270 0 0 INTERRUPT_flag
port 40 nsew
flabel metal2 5232 4860 5232 4860 3 FreeSans 48 90 0 0 clk
port 41 nsew
flabel metal3 6864 2120 6864 2120 3 FreeSans 48 0 0 0 rst
port 42 nsew
flabel metal3 -48 2720 -48 2720 7 FreeSans 48 0 0 0 IDATA_CORE_addr<0>
port 43 nsew
flabel metal2 2432 4860 2432 4860 3 FreeSans 48 90 0 0 IDATA_CORE_addr<1>
port 44 nsew
flabel metal2 1680 4860 1680 4860 3 FreeSans 48 90 0 0 IDATA_CORE_addr<2>
port 45 nsew
flabel metal2 1088 4860 1088 4860 3 FreeSans 48 90 0 0 IDATA_CORE_addr<3>
port 46 nsew
flabel metal2 5440 4860 5440 4860 3 FreeSans 48 90 0 0 IDATA_CORE_addr<4>
port 47 nsew
flabel metal3 6864 2920 6864 2920 3 FreeSans 48 0 0 0 IDATA_CORE_addr<5>
port 48 nsew
flabel metal2 5616 4860 5616 4860 3 FreeSans 48 90 0 0 IDATA_CORE_addr<6>
port 49 nsew
flabel metal3 6864 3920 6864 3920 3 FreeSans 48 0 0 0 IDATA_CORE_addr<7>
port 50 nsew
flabel metal3 6864 3760 6864 3760 3 FreeSans 48 0 0 0 IDATA_CORE_addr<8>
port 51 nsew
flabel metal2 3088 4860 3088 4860 3 FreeSans 48 90 0 0 IDATA_CORE_addr<9>
port 52 nsew
flabel metal2 6544 -40 6544 -40 7 FreeSans 48 270 0 0 IDATA_clk
port 53 nsew
flabel metal3 -48 1320 -48 1320 7 FreeSans 48 0 0 0 CORE_InstructionIN<0>
port 54 nsew
flabel metal3 -48 4720 -48 4720 7 FreeSans 48 0 0 0 CORE_InstructionIN<1>
port 55 nsew
flabel metal3 6864 320 6864 320 3 FreeSans 48 0 0 0 CORE_InstructionIN<2>
port 56 nsew
flabel metal3 -48 120 -48 120 7 FreeSans 48 0 0 0 CORE_InstructionIN<3>
port 57 nsew
flabel metal2 6080 -40 6080 -40 7 FreeSans 48 270 0 0 CORE_InstructionIN<4>
port 58 nsew
flabel metal2 352 4860 352 4860 3 FreeSans 48 90 0 0 CORE_InstructionIN<5>
port 59 nsew
flabel metal3 6864 3720 6864 3720 3 FreeSans 48 0 0 0 CORE_InstructionIN<6>
port 60 nsew
flabel metal2 576 4860 576 4860 3 FreeSans 48 90 0 0 CORE_InstructionIN<7>
port 61 nsew
flabel metal2 544 4860 544 4860 3 FreeSans 48 90 0 0 CORE_InstructionIN<8>
port 62 nsew
flabel metal2 352 -40 352 -40 7 FreeSans 48 270 0 0 CORE_InstructionIN<9>
port 63 nsew
flabel metal2 6624 4860 6624 4860 3 FreeSans 48 90 0 0 CORE_InstructionIN<10>
port 64 nsew
flabel metal2 832 4860 832 4860 3 FreeSans 48 90 0 0 CORE_InstructionIN<11>
port 65 nsew
flabel metal3 -48 720 -48 720 7 FreeSans 48 0 0 0 CORE_InstructionIN<12>
port 66 nsew
flabel metal3 -48 520 -48 520 7 FreeSans 48 0 0 0 CORE_InstructionIN<13>
port 67 nsew
flabel metal3 -48 4320 -48 4320 7 FreeSans 48 0 0 0 CORE_InstructionIN<14>
port 68 nsew
flabel metal2 3952 -40 3952 -40 7 FreeSans 48 270 0 0 CORE_InstructionIN<15>
port 69 nsew
flabel metal3 -48 3920 -48 3920 7 FreeSans 48 0 0 0 REG_R0<0>
port 70 nsew
flabel metal2 1920 4860 1920 4860 3 FreeSans 48 90 0 0 REG_R0<1>
port 71 nsew
flabel metal2 496 4860 496 4860 3 FreeSans 48 90 0 0 REG_R0<2>
port 72 nsew
flabel metal3 -48 4520 -48 4520 7 FreeSans 48 0 0 0 REG_R0<3>
port 73 nsew
flabel metal2 6480 4860 6480 4860 3 FreeSans 48 90 0 0 REG_R0<4>
port 74 nsew
flabel metal3 6864 120 6864 120 3 FreeSans 48 0 0 0 REG_R0<5>
port 75 nsew
flabel metal2 6304 4860 6304 4860 3 FreeSans 48 90 0 0 REG_R0<6>
port 76 nsew
flabel metal3 6864 4320 6864 4320 3 FreeSans 48 0 0 0 REG_R0<7>
port 77 nsew
flabel metal2 6576 4860 6576 4860 3 FreeSans 48 90 0 0 REG_R0<8>
port 78 nsew
flabel metal2 1888 -40 1888 -40 7 FreeSans 48 270 0 0 REG_R0<9>
port 79 nsew
<< end >>
