magic
tech scmos
timestamp 1514851247
<< metal1 >>
rect 206 1166 210 1168
rect 558 1166 562 1168
rect 774 1158 785 1161
rect 1102 1158 1113 1161
rect 1298 1158 1305 1161
rect 418 1148 425 1151
rect 622 1148 630 1151
rect 818 1148 822 1151
rect 918 1148 926 1151
rect 1026 1148 1033 1151
rect 1262 1146 1266 1148
rect 1406 1146 1410 1148
rect 1630 1146 1634 1148
rect 198 1138 214 1141
rect 598 1138 614 1141
rect 634 1138 649 1141
rect 966 1138 974 1141
rect 1198 1138 1209 1141
rect 1478 1138 1497 1141
rect 1686 1138 1697 1141
rect 1750 1138 1761 1141
rect 1005 1128 1006 1132
rect 1170 1128 1177 1131
rect 1326 1128 1337 1131
rect 1862 1118 1886 1121
rect 694 1078 705 1081
rect 166 1068 174 1071
rect 190 1068 198 1071
rect 502 1068 510 1071
rect 594 1068 601 1071
rect 798 1068 806 1071
rect 1574 1068 1593 1071
rect 1646 1068 1654 1071
rect 758 1062 762 1064
rect 186 1058 201 1061
rect 438 1058 446 1061
rect 586 1058 601 1061
rect 910 1061 914 1064
rect 1550 1062 1554 1064
rect 1774 1062 1778 1064
rect 910 1058 921 1061
rect 982 1058 990 1061
rect 662 1056 666 1058
rect 1022 1048 1033 1051
rect 1490 958 1497 961
rect 1682 958 1689 961
rect 502 952 506 954
rect 46 948 57 951
rect 194 948 202 951
rect 282 948 290 951
rect 818 948 825 951
rect 1394 948 1402 951
rect 1598 948 1606 951
rect 198 946 202 948
rect 286 946 290 948
rect 438 946 442 948
rect 982 946 986 948
rect 1230 946 1234 948
rect 1398 946 1402 948
rect 1838 946 1842 948
rect 66 938 81 941
rect 438 938 449 941
rect 570 938 585 941
rect 654 938 670 941
rect 1126 938 1137 941
rect 1518 938 1529 941
rect 1542 938 1558 941
rect 1766 938 1785 941
rect 1798 938 1806 941
rect 1322 928 1323 932
rect 1374 928 1385 931
rect 486 918 494 921
rect 1581 918 1582 922
rect 1858 888 1859 892
rect 1242 878 1243 882
rect 1418 878 1425 881
rect 1666 878 1667 882
rect 426 868 433 871
rect 474 868 478 871
rect 494 868 513 871
rect 798 868 809 871
rect 1170 868 1177 871
rect 1426 868 1433 871
rect 1534 868 1542 871
rect 46 858 57 861
rect 142 858 153 861
rect 318 861 322 864
rect 350 862 354 864
rect 414 862 418 864
rect 1022 862 1026 864
rect 318 858 329 861
rect 1582 856 1586 858
rect 962 848 969 851
rect 1578 848 1585 851
rect 1722 848 1729 851
rect 1534 768 1542 771
rect 1786 768 1793 771
rect 490 758 497 761
rect 554 758 561 761
rect 46 748 57 751
rect 138 748 158 751
rect 678 748 686 751
rect 422 746 426 748
rect 454 746 458 748
rect 678 746 682 748
rect 742 746 746 748
rect 830 746 834 748
rect 1326 748 1334 751
rect 1374 748 1382 751
rect 902 746 906 748
rect 150 738 166 741
rect 294 738 305 741
rect 510 738 518 741
rect 610 738 625 741
rect 714 738 721 741
rect 986 738 993 741
rect 1006 738 1025 741
rect 1038 738 1046 741
rect 1090 738 1097 741
rect 1110 738 1118 741
rect 1150 738 1158 741
rect 1278 738 1286 741
rect 1470 738 1478 741
rect 1782 738 1793 741
rect 698 718 699 722
rect 1234 678 1238 681
rect 386 668 401 671
rect 446 668 454 671
rect 734 668 745 671
rect 834 668 841 671
rect 1118 668 1137 671
rect 1146 668 1161 671
rect 1234 668 1249 671
rect 1278 668 1297 671
rect 1310 668 1318 671
rect 1854 668 1870 671
rect 1566 662 1570 664
rect 46 658 57 661
rect 870 658 878 661
rect 934 658 953 661
rect 1054 658 1065 661
rect 706 648 713 651
rect 1354 648 1361 651
rect 1821 578 1822 582
rect 218 558 225 561
rect 282 558 289 561
rect 738 558 745 561
rect 802 558 809 561
rect 46 548 57 551
rect 510 546 514 548
rect 582 546 586 548
rect 830 546 834 548
rect 1486 548 1494 551
rect 1742 548 1750 551
rect 838 546 842 548
rect 926 546 930 548
rect 1742 546 1746 548
rect 1870 546 1874 548
rect 310 538 321 541
rect 334 538 342 541
rect 758 538 766 541
rect 1086 538 1105 541
rect 1158 538 1177 541
rect 1354 538 1369 541
rect 1558 538 1569 541
rect 1189 528 1190 532
rect 986 488 987 492
rect 454 468 462 471
rect 626 468 633 471
rect 182 462 186 464
rect 134 458 145 461
rect 430 458 449 461
rect 662 461 665 471
rect 774 468 785 471
rect 818 468 825 471
rect 838 468 849 471
rect 1046 468 1065 471
rect 1090 468 1097 471
rect 1114 468 1121 471
rect 1366 468 1382 471
rect 1534 468 1542 471
rect 1590 468 1598 471
rect 1730 468 1734 471
rect 1782 468 1793 471
rect 1022 462 1026 464
rect 654 458 665 461
rect 1174 462 1178 464
rect 1238 462 1242 464
rect 1302 462 1306 464
rect 1694 461 1698 464
rect 1670 458 1698 461
rect 430 448 433 458
rect 622 448 630 451
rect 686 448 705 451
rect 46 442 50 444
rect 990 442 994 444
rect 446 438 454 441
rect 1110 442 1114 444
rect 1242 438 1249 441
rect 386 368 401 371
rect 1342 368 1358 371
rect 58 348 62 351
rect 206 351 209 361
rect 374 358 385 361
rect 458 358 465 361
rect 554 358 561 361
rect 1562 358 1569 361
rect 190 348 209 351
rect 214 348 233 351
rect 382 351 386 354
rect 378 348 386 351
rect 782 348 793 351
rect 1110 348 1118 351
rect 1166 348 1177 351
rect 54 338 62 341
rect 70 338 89 341
rect 110 338 121 341
rect 234 338 241 341
rect 614 338 633 341
rect 782 338 785 348
rect 814 346 818 348
rect 1110 346 1114 348
rect 990 338 1001 341
rect 1166 338 1169 348
rect 1198 346 1202 348
rect 1466 348 1473 351
rect 1770 348 1777 351
rect 1854 348 1878 351
rect 1238 346 1242 348
rect 1198 338 1209 341
rect 1294 338 1313 341
rect 1438 338 1457 341
rect 1518 338 1526 341
rect 1614 338 1633 341
rect 1650 338 1657 341
rect 86 328 89 338
rect 286 328 297 331
rect 318 328 329 331
rect 614 328 617 338
rect 170 278 177 281
rect 126 268 137 271
rect 606 268 617 271
rect 630 268 638 271
rect 742 268 753 271
rect 926 268 934 271
rect 1026 268 1041 271
rect 1046 268 1054 271
rect 1366 268 1377 271
rect 1762 268 1777 271
rect 1822 268 1830 271
rect 1862 268 1886 271
rect 510 262 514 264
rect 518 262 522 264
rect 686 262 690 264
rect 966 261 970 264
rect 1454 262 1458 264
rect 966 258 977 261
rect 1054 258 1073 261
rect 1734 261 1738 264
rect 1734 258 1745 261
rect 54 256 58 258
rect 422 241 425 251
rect 1338 248 1345 251
rect 462 246 466 248
rect 422 238 433 241
rect 1194 168 1202 171
rect 1198 166 1202 168
rect 574 158 585 161
rect 942 158 950 161
rect 1098 158 1105 161
rect 1310 158 1318 161
rect 1778 158 1785 161
rect 198 152 202 154
rect 518 148 526 151
rect 758 146 762 148
rect 910 146 914 148
rect 1278 148 1289 151
rect 1518 148 1526 151
rect 918 146 922 148
rect 126 138 134 141
rect 310 138 318 141
rect 342 138 361 141
rect 1286 138 1289 148
rect 1414 146 1418 148
rect 1630 146 1634 148
rect 1630 138 1641 141
rect 1702 138 1710 141
rect 110 71 113 81
rect 538 78 553 81
rect 94 68 113 71
rect 134 68 145 71
rect 414 68 425 71
rect 758 68 766 71
rect 990 68 998 71
rect 1134 68 1145 71
rect 166 58 174 61
rect 190 58 209 61
rect 454 61 458 64
rect 450 58 458 61
rect 490 58 513 61
rect 558 58 569 61
rect 734 58 745 61
rect 1006 58 1017 61
rect 1170 58 1177 61
rect 1270 61 1273 71
rect 1318 68 1334 71
rect 1446 71 1449 81
rect 1418 68 1425 71
rect 1430 68 1449 71
rect 1494 68 1510 71
rect 1614 68 1633 71
rect 1262 58 1273 61
rect 1398 58 1417 61
rect 1542 58 1553 61
rect 54 56 58 58
rect 190 48 193 58
rect 402 48 417 51
rect 1294 48 1305 51
rect 702 42 706 44
rect 878 42 882 44
rect 1510 42 1514 44
<< m2contact >>
rect 54 1188 58 1192
rect 102 1188 106 1192
rect 342 1188 346 1192
rect 742 1188 746 1192
rect 1118 1178 1122 1182
rect 6 1168 10 1172
rect 206 1168 210 1172
rect 558 1168 562 1172
rect 1126 1168 1130 1172
rect 1142 1168 1146 1172
rect 414 1158 418 1162
rect 1294 1158 1298 1162
rect 1438 1158 1442 1162
rect 22 1148 26 1152
rect 70 1148 74 1152
rect 94 1148 98 1152
rect 118 1148 122 1152
rect 142 1148 146 1152
rect 230 1148 234 1152
rect 278 1148 282 1152
rect 358 1148 362 1152
rect 382 1148 386 1152
rect 398 1148 402 1152
rect 414 1148 418 1152
rect 438 1148 442 1152
rect 550 1148 554 1152
rect 582 1148 586 1152
rect 614 1148 618 1152
rect 630 1148 634 1152
rect 678 1148 682 1152
rect 694 1148 698 1152
rect 702 1148 706 1152
rect 726 1148 730 1152
rect 758 1148 762 1152
rect 814 1148 818 1152
rect 822 1148 826 1152
rect 846 1148 850 1152
rect 854 1148 858 1152
rect 862 1148 866 1152
rect 886 1148 890 1152
rect 894 1148 898 1152
rect 926 1148 930 1152
rect 934 1148 938 1152
rect 942 1148 946 1152
rect 966 1148 970 1152
rect 990 1148 994 1152
rect 1014 1148 1018 1152
rect 1022 1148 1026 1152
rect 1038 1148 1042 1152
rect 1062 1148 1066 1152
rect 1118 1148 1122 1152
rect 1214 1148 1218 1152
rect 1230 1148 1234 1152
rect 1254 1148 1258 1152
rect 1262 1148 1266 1152
rect 1286 1148 1290 1152
rect 1350 1148 1354 1152
rect 1366 1148 1370 1152
rect 1374 1148 1378 1152
rect 1390 1148 1394 1152
rect 1398 1148 1402 1152
rect 1406 1148 1410 1152
rect 1526 1148 1530 1152
rect 1558 1148 1562 1152
rect 1566 1148 1570 1152
rect 1582 1148 1586 1152
rect 1590 1148 1594 1152
rect 1630 1148 1634 1152
rect 1638 1148 1642 1152
rect 1742 1148 1746 1152
rect 30 1138 34 1142
rect 78 1138 82 1142
rect 126 1138 130 1142
rect 150 1138 154 1142
rect 214 1138 218 1142
rect 222 1138 226 1142
rect 270 1138 274 1142
rect 286 1138 290 1142
rect 334 1138 338 1142
rect 366 1138 370 1142
rect 390 1138 394 1142
rect 430 1138 434 1142
rect 470 1140 474 1144
rect 478 1138 482 1142
rect 486 1138 490 1142
rect 534 1138 538 1142
rect 574 1138 578 1142
rect 590 1138 594 1142
rect 614 1138 618 1142
rect 630 1138 634 1142
rect 670 1138 674 1142
rect 718 1138 722 1142
rect 750 1138 754 1142
rect 766 1138 770 1142
rect 798 1138 802 1142
rect 822 1138 826 1142
rect 878 1138 882 1142
rect 974 1138 978 1142
rect 1086 1138 1090 1142
rect 1158 1138 1162 1142
rect 1182 1138 1186 1142
rect 1294 1138 1298 1142
rect 1318 1138 1322 1142
rect 1414 1140 1418 1144
rect 1446 1138 1450 1142
rect 1462 1138 1466 1142
rect 1518 1138 1522 1142
rect 1614 1140 1618 1144
rect 1622 1138 1626 1142
rect 1670 1138 1674 1142
rect 1702 1140 1706 1144
rect 1774 1138 1778 1142
rect 1798 1138 1802 1142
rect 1814 1138 1818 1142
rect 1830 1138 1834 1142
rect 86 1127 90 1131
rect 246 1128 250 1132
rect 254 1128 258 1132
rect 446 1128 450 1132
rect 542 1128 546 1132
rect 566 1128 570 1132
rect 606 1128 610 1132
rect 630 1128 634 1132
rect 638 1128 642 1132
rect 806 1128 810 1132
rect 1006 1128 1010 1132
rect 1078 1128 1082 1132
rect 1166 1128 1170 1132
rect 1454 1128 1458 1132
rect 1486 1128 1490 1132
rect 1662 1128 1666 1132
rect 1782 1128 1786 1132
rect 1790 1128 1794 1132
rect 1822 1128 1826 1132
rect 1854 1128 1858 1132
rect 174 1118 178 1122
rect 238 1118 242 1122
rect 262 1118 266 1122
rect 310 1118 314 1122
rect 414 1118 418 1122
rect 454 1118 458 1122
rect 510 1118 514 1122
rect 662 1118 666 1122
rect 910 1118 914 1122
rect 1054 1118 1058 1122
rect 1238 1118 1242 1122
rect 1270 1118 1274 1122
rect 1334 1118 1338 1122
rect 1430 1118 1434 1122
rect 1510 1118 1514 1122
rect 1542 1118 1546 1122
rect 1598 1118 1602 1122
rect 1654 1118 1658 1122
rect 1718 1118 1722 1122
rect 1726 1118 1730 1122
rect 1846 1118 1850 1122
rect 1886 1118 1890 1122
rect 142 1088 146 1092
rect 294 1088 298 1092
rect 398 1088 402 1092
rect 582 1088 586 1092
rect 734 1088 738 1092
rect 1238 1088 1242 1092
rect 1414 1088 1418 1092
rect 1622 1088 1626 1092
rect 1678 1088 1682 1092
rect 1686 1088 1690 1092
rect 1766 1088 1770 1092
rect 1798 1088 1802 1092
rect 86 1078 90 1082
rect 238 1078 242 1082
rect 350 1078 354 1082
rect 510 1078 514 1082
rect 726 1078 730 1082
rect 998 1078 1002 1082
rect 1086 1078 1090 1082
rect 1230 1078 1234 1082
rect 1582 1078 1586 1082
rect 1614 1078 1618 1082
rect 1710 1078 1714 1082
rect 6 1068 10 1072
rect 78 1068 82 1072
rect 94 1068 98 1072
rect 134 1068 138 1072
rect 174 1068 178 1072
rect 198 1068 202 1072
rect 206 1068 210 1072
rect 222 1068 226 1072
rect 246 1068 250 1072
rect 270 1068 274 1072
rect 278 1066 282 1070
rect 358 1068 362 1072
rect 382 1068 386 1072
rect 438 1068 442 1072
rect 478 1068 482 1072
rect 510 1068 514 1072
rect 566 1068 570 1072
rect 590 1068 594 1072
rect 686 1068 690 1072
rect 718 1068 722 1072
rect 806 1068 810 1072
rect 814 1068 818 1072
rect 942 1068 946 1072
rect 982 1068 986 1072
rect 1006 1068 1010 1072
rect 1078 1068 1082 1072
rect 1142 1068 1146 1072
rect 1174 1068 1178 1072
rect 1222 1068 1226 1072
rect 1262 1068 1266 1072
rect 1302 1068 1306 1072
rect 1438 1068 1442 1072
rect 1518 1068 1522 1072
rect 1606 1068 1610 1072
rect 1654 1068 1658 1072
rect 1718 1068 1722 1072
rect 1742 1068 1746 1072
rect 1838 1068 1842 1072
rect 46 1058 50 1062
rect 158 1058 162 1062
rect 182 1058 186 1062
rect 214 1058 218 1062
rect 230 1058 234 1062
rect 310 1058 314 1062
rect 334 1058 338 1062
rect 342 1058 346 1062
rect 406 1058 410 1062
rect 414 1058 418 1062
rect 446 1058 450 1062
rect 462 1058 466 1062
rect 470 1058 474 1062
rect 526 1058 530 1062
rect 550 1058 554 1062
rect 558 1058 562 1062
rect 582 1058 586 1062
rect 622 1058 626 1062
rect 630 1058 634 1062
rect 654 1058 658 1062
rect 662 1058 666 1062
rect 670 1058 674 1062
rect 750 1058 754 1062
rect 758 1058 762 1062
rect 766 1058 770 1062
rect 774 1058 778 1062
rect 798 1058 802 1062
rect 830 1058 834 1062
rect 838 1058 842 1062
rect 846 1058 850 1062
rect 870 1058 874 1062
rect 902 1058 906 1062
rect 934 1058 938 1062
rect 950 1058 954 1062
rect 958 1058 962 1062
rect 990 1058 994 1062
rect 1038 1058 1042 1062
rect 1102 1058 1106 1062
rect 1126 1058 1130 1062
rect 1134 1058 1138 1062
rect 1150 1058 1154 1062
rect 1182 1058 1186 1062
rect 1198 1058 1202 1062
rect 1254 1058 1258 1062
rect 1270 1058 1274 1062
rect 1278 1058 1282 1062
rect 1302 1058 1306 1062
rect 1326 1058 1330 1062
rect 1334 1058 1338 1062
rect 1350 1058 1354 1062
rect 1358 1058 1362 1062
rect 1366 1058 1370 1062
rect 1374 1058 1378 1062
rect 1398 1058 1402 1062
rect 1430 1058 1434 1062
rect 1454 1058 1458 1062
rect 1462 1058 1466 1062
rect 1478 1058 1482 1062
rect 1486 1058 1490 1062
rect 1510 1058 1514 1062
rect 1526 1058 1530 1062
rect 1542 1058 1546 1062
rect 1550 1058 1554 1062
rect 1638 1058 1642 1062
rect 1662 1058 1666 1062
rect 1702 1058 1706 1062
rect 1750 1058 1754 1062
rect 1774 1058 1778 1062
rect 1782 1058 1786 1062
rect 1814 1058 1818 1062
rect 1830 1058 1834 1062
rect 1846 1058 1850 1062
rect 22 1048 26 1052
rect 54 1048 58 1052
rect 62 1048 66 1052
rect 118 1048 122 1052
rect 174 1048 178 1052
rect 398 1048 402 1052
rect 486 1048 490 1052
rect 582 1048 586 1052
rect 1494 1048 1498 1052
rect 1806 1048 1810 1052
rect 38 1038 42 1042
rect 374 1038 378 1042
rect 454 1038 458 1042
rect 646 1038 650 1042
rect 886 1038 890 1042
rect 1046 1038 1050 1042
rect 1062 1038 1066 1042
rect 1110 1038 1114 1042
rect 1822 1038 1826 1042
rect 14 1028 18 1032
rect 654 1028 658 1032
rect 46 1018 50 1022
rect 70 1018 74 1022
rect 110 1018 114 1022
rect 126 1018 130 1022
rect 262 1018 266 1022
rect 318 1018 322 1022
rect 534 1018 538 1022
rect 862 1018 866 1022
rect 1038 1018 1042 1022
rect 1166 1018 1170 1022
rect 1206 1018 1210 1022
rect 1390 1018 1394 1022
rect 1558 1018 1562 1022
rect 1734 1018 1738 1022
rect 1862 1018 1866 1022
rect 510 988 514 992
rect 598 988 602 992
rect 798 988 802 992
rect 910 988 914 992
rect 1054 988 1058 992
rect 1430 988 1434 992
rect 1574 988 1578 992
rect 1630 988 1634 992
rect 1750 988 1754 992
rect 1102 978 1106 982
rect 6 968 10 972
rect 166 968 170 972
rect 486 968 490 972
rect 750 968 754 972
rect 1654 968 1658 972
rect 262 958 266 962
rect 734 958 738 962
rect 1022 958 1026 962
rect 1070 958 1074 962
rect 1198 958 1202 962
rect 1486 958 1490 962
rect 1678 958 1682 962
rect 22 948 26 952
rect 70 948 74 952
rect 118 948 122 952
rect 142 948 146 952
rect 174 948 178 952
rect 182 948 186 952
rect 190 948 194 952
rect 206 948 210 952
rect 246 948 250 952
rect 270 948 274 952
rect 278 948 282 952
rect 294 948 298 952
rect 318 948 322 952
rect 390 948 394 952
rect 438 948 442 952
rect 454 948 458 952
rect 494 948 498 952
rect 502 948 506 952
rect 542 948 546 952
rect 638 948 642 952
rect 678 948 682 952
rect 702 948 706 952
rect 742 948 746 952
rect 814 948 818 952
rect 854 948 858 952
rect 894 948 898 952
rect 926 948 930 952
rect 950 948 954 952
rect 958 948 962 952
rect 974 948 978 952
rect 982 948 986 952
rect 998 948 1002 952
rect 1086 948 1090 952
rect 1118 948 1122 952
rect 1230 948 1234 952
rect 1238 948 1242 952
rect 1262 948 1266 952
rect 1302 948 1306 952
rect 1310 948 1314 952
rect 1334 948 1338 952
rect 1390 948 1394 952
rect 1406 948 1410 952
rect 1478 948 1482 952
rect 1510 948 1514 952
rect 1566 948 1570 952
rect 1590 948 1594 952
rect 1606 948 1610 952
rect 1614 948 1618 952
rect 1638 948 1642 952
rect 1670 948 1674 952
rect 1814 948 1818 952
rect 1830 948 1834 952
rect 1838 948 1842 952
rect 1862 948 1866 952
rect 30 938 34 942
rect 62 938 66 942
rect 126 938 130 942
rect 134 938 138 942
rect 190 938 194 942
rect 254 938 258 942
rect 278 938 282 942
rect 334 938 338 942
rect 350 938 354 942
rect 358 940 362 944
rect 382 938 386 942
rect 430 940 434 944
rect 526 938 530 942
rect 558 938 562 942
rect 566 938 570 942
rect 614 938 618 942
rect 670 938 674 942
rect 718 940 722 944
rect 726 938 730 942
rect 766 938 770 942
rect 782 938 786 942
rect 846 938 850 942
rect 902 938 906 942
rect 990 938 994 942
rect 1038 938 1042 942
rect 1094 938 1098 942
rect 1150 938 1154 942
rect 1174 938 1178 942
rect 1214 938 1218 942
rect 1366 938 1370 942
rect 1446 938 1450 942
rect 1486 938 1490 942
rect 1558 938 1562 942
rect 1678 938 1682 942
rect 1702 938 1706 942
rect 1718 938 1722 942
rect 1734 938 1738 942
rect 1806 938 1810 942
rect 1870 938 1874 942
rect 62 928 66 932
rect 94 928 98 932
rect 342 928 346 932
rect 534 928 538 932
rect 566 928 570 932
rect 574 928 578 932
rect 606 928 610 932
rect 662 928 666 932
rect 750 928 754 932
rect 790 928 794 932
rect 1046 928 1050 932
rect 1062 928 1066 932
rect 1158 928 1162 932
rect 1166 928 1170 932
rect 1190 928 1194 932
rect 1222 928 1226 932
rect 1294 928 1298 932
rect 1318 928 1322 932
rect 1390 928 1394 932
rect 1454 928 1458 932
rect 1550 928 1554 932
rect 1710 928 1714 932
rect 1742 928 1746 932
rect 1774 928 1778 932
rect 1806 928 1810 932
rect 86 918 90 922
rect 102 918 106 922
rect 158 918 162 922
rect 222 918 226 922
rect 230 918 234 922
rect 310 918 314 922
rect 374 918 378 922
rect 406 918 410 922
rect 414 918 418 922
rect 470 918 474 922
rect 494 918 498 922
rect 630 918 634 922
rect 694 918 698 922
rect 838 918 842 922
rect 870 918 874 922
rect 878 918 882 922
rect 934 918 938 922
rect 1014 918 1018 922
rect 1070 918 1074 922
rect 1254 918 1258 922
rect 1278 918 1282 922
rect 1286 918 1290 922
rect 1350 918 1354 922
rect 1382 918 1386 922
rect 1422 918 1426 922
rect 1462 918 1466 922
rect 1582 918 1586 922
rect 1846 918 1850 922
rect 294 888 298 892
rect 390 888 394 892
rect 526 888 530 892
rect 774 888 778 892
rect 998 888 1002 892
rect 1190 888 1194 892
rect 1302 888 1306 892
rect 1334 888 1338 892
rect 1358 888 1362 892
rect 1390 888 1394 892
rect 1518 888 1522 892
rect 1694 888 1698 892
rect 1758 888 1762 892
rect 1790 888 1794 892
rect 1854 888 1858 892
rect 6 878 10 882
rect 62 878 66 882
rect 158 878 162 882
rect 166 878 170 882
rect 382 878 386 882
rect 422 878 426 882
rect 462 878 466 882
rect 470 878 474 882
rect 502 878 506 882
rect 534 878 538 882
rect 646 878 650 882
rect 734 878 738 882
rect 830 878 834 882
rect 870 878 874 882
rect 1102 878 1106 882
rect 1166 878 1170 882
rect 1214 878 1218 882
rect 1238 878 1242 882
rect 1294 878 1298 882
rect 1414 878 1418 882
rect 1454 878 1458 882
rect 1542 878 1546 882
rect 1598 878 1602 882
rect 1638 878 1642 882
rect 1662 878 1666 882
rect 1750 878 1754 882
rect 1798 878 1802 882
rect 1830 878 1834 882
rect 30 868 34 872
rect 70 868 74 872
rect 102 868 106 872
rect 126 868 130 872
rect 174 868 178 872
rect 190 868 194 872
rect 222 868 226 872
rect 254 868 258 872
rect 262 868 266 872
rect 342 866 346 870
rect 374 868 378 872
rect 422 868 426 872
rect 470 868 474 872
rect 478 868 482 872
rect 542 868 546 872
rect 582 866 586 870
rect 590 868 594 872
rect 606 868 610 872
rect 614 868 618 872
rect 654 868 658 872
rect 678 868 682 872
rect 710 868 714 872
rect 726 868 730 872
rect 822 868 826 872
rect 862 868 866 872
rect 878 868 882 872
rect 926 868 930 872
rect 958 868 962 872
rect 982 866 986 870
rect 990 868 994 872
rect 1078 868 1082 872
rect 1094 868 1098 872
rect 1158 868 1162 872
rect 1166 868 1170 872
rect 1206 868 1210 872
rect 1286 868 1290 872
rect 1326 868 1330 872
rect 1374 866 1378 870
rect 1382 868 1386 872
rect 1406 868 1410 872
rect 1422 868 1426 872
rect 1462 868 1466 872
rect 1542 868 1546 872
rect 1566 866 1570 870
rect 1574 868 1578 872
rect 1614 868 1618 872
rect 1630 868 1634 872
rect 1718 868 1722 872
rect 1742 868 1746 872
rect 1782 868 1786 872
rect 1806 868 1810 872
rect 1822 868 1826 872
rect 22 858 26 862
rect 78 858 82 862
rect 118 858 122 862
rect 214 858 218 862
rect 230 858 234 862
rect 246 858 250 862
rect 270 858 274 862
rect 310 858 314 862
rect 350 858 354 862
rect 406 858 410 862
rect 414 858 418 862
rect 566 858 570 862
rect 622 858 626 862
rect 670 858 674 862
rect 686 858 690 862
rect 750 858 754 862
rect 790 858 794 862
rect 838 858 842 862
rect 854 858 858 862
rect 902 858 906 862
rect 918 858 922 862
rect 934 858 938 862
rect 950 858 954 862
rect 1014 858 1018 862
rect 1022 858 1026 862
rect 1030 858 1034 862
rect 1038 858 1042 862
rect 1062 858 1066 862
rect 1126 858 1130 862
rect 1142 858 1146 862
rect 1222 858 1226 862
rect 1230 858 1234 862
rect 1254 858 1258 862
rect 1318 858 1322 862
rect 1350 858 1354 862
rect 1494 858 1498 862
rect 1550 858 1554 862
rect 1582 858 1586 862
rect 1590 858 1594 862
rect 1646 858 1650 862
rect 1654 858 1658 862
rect 1678 858 1682 862
rect 1710 858 1714 862
rect 1774 858 1778 862
rect 1838 858 1842 862
rect 1846 858 1850 862
rect 1870 858 1874 862
rect 702 848 706 852
rect 742 848 746 852
rect 958 848 962 852
rect 1110 848 1114 852
rect 1182 848 1186 852
rect 1486 848 1490 852
rect 1574 848 1578 852
rect 1718 848 1722 852
rect 758 838 762 842
rect 1126 838 1130 842
rect 1502 838 1506 842
rect 1598 838 1602 842
rect 454 828 458 832
rect 598 828 602 832
rect 94 818 98 822
rect 198 818 202 822
rect 286 818 290 822
rect 358 818 362 822
rect 446 818 450 822
rect 494 818 498 822
rect 526 818 530 822
rect 558 818 562 822
rect 638 818 642 822
rect 710 818 714 822
rect 750 818 754 822
rect 894 818 898 822
rect 1054 818 1058 822
rect 1118 818 1122 822
rect 1270 818 1274 822
rect 1334 818 1338 822
rect 1446 818 1450 822
rect 1478 818 1482 822
rect 1494 818 1498 822
rect 238 788 242 792
rect 334 788 338 792
rect 366 788 370 792
rect 1254 788 1258 792
rect 1702 788 1706 792
rect 6 778 10 782
rect 1126 778 1130 782
rect 1542 768 1546 772
rect 1734 768 1738 772
rect 1782 768 1786 772
rect 214 758 218 762
rect 486 758 490 762
rect 550 758 554 762
rect 702 758 706 762
rect 1094 758 1098 762
rect 1406 758 1410 762
rect 22 748 26 752
rect 134 748 138 752
rect 158 748 162 752
rect 190 748 194 752
rect 254 748 258 752
rect 270 748 274 752
rect 286 748 290 752
rect 414 748 418 752
rect 422 748 426 752
rect 430 748 434 752
rect 446 748 450 752
rect 454 748 458 752
rect 478 748 482 752
rect 526 748 530 752
rect 542 748 546 752
rect 670 748 674 752
rect 686 748 690 752
rect 742 748 746 752
rect 750 748 754 752
rect 830 748 834 752
rect 902 748 906 752
rect 910 748 914 752
rect 966 748 970 752
rect 1054 748 1058 752
rect 1070 748 1074 752
rect 1086 748 1090 752
rect 1118 748 1122 752
rect 1166 748 1170 752
rect 1222 748 1226 752
rect 1238 748 1242 752
rect 1270 748 1274 752
rect 1294 748 1298 752
rect 1318 748 1322 752
rect 1334 748 1338 752
rect 1342 748 1346 752
rect 1366 748 1370 752
rect 1382 748 1386 752
rect 1390 748 1394 752
rect 1414 748 1418 752
rect 1446 748 1450 752
rect 1502 748 1506 752
rect 1518 748 1522 752
rect 1550 748 1554 752
rect 1574 748 1578 752
rect 1606 748 1610 752
rect 1654 748 1658 752
rect 1670 748 1674 752
rect 1686 748 1690 752
rect 1750 748 1754 752
rect 1830 748 1834 752
rect 30 738 34 742
rect 86 740 90 744
rect 94 738 98 742
rect 102 738 106 742
rect 166 738 170 742
rect 222 738 226 742
rect 230 738 234 742
rect 262 738 266 742
rect 318 738 322 742
rect 350 738 354 742
rect 366 738 370 742
rect 382 738 386 742
rect 486 738 490 742
rect 518 738 522 742
rect 550 738 554 742
rect 574 738 578 742
rect 590 738 594 742
rect 606 738 610 742
rect 638 738 642 742
rect 686 738 690 742
rect 710 738 714 742
rect 782 738 786 742
rect 822 740 826 744
rect 846 738 850 742
rect 862 738 866 742
rect 886 740 890 744
rect 894 738 898 742
rect 942 738 946 742
rect 982 738 986 742
rect 1046 738 1050 742
rect 1078 738 1082 742
rect 1086 738 1090 742
rect 1118 738 1122 742
rect 1142 740 1146 744
rect 1158 738 1162 742
rect 1198 738 1202 742
rect 1246 738 1250 742
rect 1286 738 1290 742
rect 1342 738 1346 742
rect 1454 738 1458 742
rect 1478 738 1482 742
rect 1510 738 1514 742
rect 1542 738 1546 742
rect 1582 738 1586 742
rect 1622 738 1626 742
rect 1662 738 1666 742
rect 1694 738 1698 742
rect 1718 738 1722 742
rect 1774 740 1778 744
rect 1806 738 1810 742
rect 1822 738 1826 742
rect 1854 738 1858 742
rect 1862 740 1866 744
rect 62 728 66 732
rect 182 728 186 732
rect 206 728 210 732
rect 326 728 330 732
rect 358 728 362 732
rect 390 728 394 732
rect 518 728 522 732
rect 582 728 586 732
rect 614 728 618 732
rect 646 728 650 732
rect 710 728 714 732
rect 774 728 778 732
rect 838 728 842 732
rect 934 728 938 732
rect 982 728 986 732
rect 1014 728 1018 732
rect 1046 728 1050 732
rect 1190 728 1194 732
rect 1478 728 1482 732
rect 1598 728 1602 732
rect 1630 728 1634 732
rect 1726 728 1730 732
rect 1814 728 1818 732
rect 70 718 74 722
rect 126 718 130 722
rect 174 718 178 722
rect 198 718 202 722
rect 398 718 402 722
rect 462 718 466 722
rect 654 718 658 722
rect 694 718 698 722
rect 734 718 738 722
rect 766 718 770 722
rect 798 718 802 722
rect 806 718 810 722
rect 870 718 874 722
rect 926 718 930 722
rect 958 718 962 722
rect 974 718 978 722
rect 1182 718 1186 722
rect 1214 718 1218 722
rect 1302 718 1306 722
rect 1430 718 1434 722
rect 1486 718 1490 722
rect 1566 718 1570 722
rect 1590 718 1594 722
rect 1638 718 1642 722
rect 1758 718 1762 722
rect 1846 718 1850 722
rect 1878 718 1882 722
rect 86 688 90 692
rect 206 688 210 692
rect 270 688 274 692
rect 326 688 330 692
rect 366 688 370 692
rect 422 688 426 692
rect 526 688 530 692
rect 622 688 626 692
rect 678 688 682 692
rect 774 688 778 692
rect 918 688 922 692
rect 1078 688 1082 692
rect 1102 688 1106 692
rect 1182 688 1186 692
rect 1406 688 1410 692
rect 1462 688 1466 692
rect 1606 688 1610 692
rect 1678 688 1682 692
rect 1790 688 1794 692
rect 1798 688 1802 692
rect 1830 688 1834 692
rect 174 678 178 682
rect 358 678 362 682
rect 390 678 394 682
rect 454 678 458 682
rect 462 678 466 682
rect 582 678 586 682
rect 614 678 618 682
rect 766 678 770 682
rect 822 678 826 682
rect 830 678 834 682
rect 878 678 882 682
rect 974 678 978 682
rect 1006 678 1010 682
rect 1046 678 1050 682
rect 1166 678 1170 682
rect 1174 678 1178 682
rect 1230 678 1234 682
rect 1238 678 1242 682
rect 1254 678 1258 682
rect 1286 678 1290 682
rect 1318 678 1322 682
rect 1510 678 1514 682
rect 1598 678 1602 682
rect 1670 678 1674 682
rect 1726 678 1730 682
rect 1758 678 1762 682
rect 6 668 10 672
rect 30 668 34 672
rect 78 668 82 672
rect 110 668 114 672
rect 134 668 138 672
rect 166 668 170 672
rect 182 668 186 672
rect 198 668 202 672
rect 230 668 234 672
rect 238 668 242 672
rect 294 668 298 672
rect 302 668 306 672
rect 350 668 354 672
rect 382 668 386 672
rect 406 666 410 670
rect 454 668 458 672
rect 470 668 474 672
rect 518 668 522 672
rect 550 668 554 672
rect 574 668 578 672
rect 606 668 610 672
rect 702 668 706 672
rect 726 666 730 670
rect 758 668 762 672
rect 814 668 818 672
rect 830 668 834 672
rect 910 668 914 672
rect 942 668 946 672
rect 966 668 970 672
rect 982 668 986 672
rect 998 668 1002 672
rect 1014 668 1018 672
rect 1070 668 1074 672
rect 1086 668 1090 672
rect 1142 668 1146 672
rect 1190 668 1194 672
rect 1222 668 1226 672
rect 1230 668 1234 672
rect 1262 668 1266 672
rect 1318 668 1322 672
rect 1350 668 1354 672
rect 1382 668 1386 672
rect 1502 668 1506 672
rect 1590 668 1594 672
rect 1630 668 1634 672
rect 1662 668 1666 672
rect 1686 668 1690 672
rect 1718 668 1722 672
rect 1750 668 1754 672
rect 1766 668 1770 672
rect 1774 666 1778 670
rect 1822 668 1826 672
rect 1846 666 1850 670
rect 1870 668 1874 672
rect 22 658 26 662
rect 70 658 74 662
rect 102 658 106 662
rect 126 658 130 662
rect 142 658 146 662
rect 158 658 162 662
rect 222 658 226 662
rect 246 658 250 662
rect 286 658 290 662
rect 310 658 314 662
rect 430 658 434 662
rect 494 658 498 662
rect 510 658 514 662
rect 542 658 546 662
rect 638 658 642 662
rect 662 658 666 662
rect 694 658 698 662
rect 790 658 794 662
rect 862 658 866 662
rect 878 658 882 662
rect 902 658 906 662
rect 1022 658 1026 662
rect 1030 658 1034 662
rect 1094 658 1098 662
rect 1150 658 1154 662
rect 1198 658 1202 662
rect 1238 658 1242 662
rect 1326 658 1330 662
rect 1342 658 1346 662
rect 1374 658 1378 662
rect 1398 658 1402 662
rect 1422 658 1426 662
rect 1430 658 1434 662
rect 1438 658 1442 662
rect 1446 658 1450 662
rect 1470 658 1474 662
rect 1518 658 1522 662
rect 1542 658 1546 662
rect 1558 658 1562 662
rect 1566 658 1570 662
rect 1574 658 1578 662
rect 1622 658 1626 662
rect 1654 658 1658 662
rect 1694 658 1698 662
rect 1702 658 1706 662
rect 1814 658 1818 662
rect 118 648 122 652
rect 262 648 266 652
rect 334 648 338 652
rect 670 648 674 652
rect 702 648 706 652
rect 854 648 858 652
rect 918 648 922 652
rect 1038 648 1042 652
rect 1102 648 1106 652
rect 1126 648 1130 652
rect 1350 648 1354 652
rect 1638 648 1642 652
rect 654 638 658 642
rect 1734 638 1738 642
rect 366 618 370 622
rect 486 618 490 622
rect 558 618 562 622
rect 590 618 594 622
rect 662 618 666 622
rect 798 618 802 622
rect 886 618 890 622
rect 1206 618 1210 622
rect 1486 618 1490 622
rect 1534 618 1538 622
rect 190 588 194 592
rect 430 588 434 592
rect 710 588 714 592
rect 1062 588 1066 592
rect 1422 588 1426 592
rect 1614 588 1618 592
rect 1670 588 1674 592
rect 1686 588 1690 592
rect 1766 588 1770 592
rect 894 578 898 582
rect 1326 578 1330 582
rect 1822 578 1826 582
rect 6 568 10 572
rect 422 568 426 572
rect 478 568 482 572
rect 1030 568 1034 572
rect 70 558 74 562
rect 214 558 218 562
rect 278 558 282 562
rect 438 558 442 562
rect 590 558 594 562
rect 638 558 642 562
rect 734 558 738 562
rect 798 558 802 562
rect 22 548 26 552
rect 118 548 122 552
rect 134 548 138 552
rect 150 548 154 552
rect 166 548 170 552
rect 182 548 186 552
rect 206 548 210 552
rect 238 548 242 552
rect 302 548 306 552
rect 350 548 354 552
rect 366 548 370 552
rect 382 548 386 552
rect 430 548 434 552
rect 494 548 498 552
rect 510 548 514 552
rect 518 548 522 552
rect 558 548 562 552
rect 574 548 578 552
rect 582 548 586 552
rect 606 548 610 552
rect 670 548 674 552
rect 702 548 706 552
rect 726 548 730 552
rect 774 548 778 552
rect 790 548 794 552
rect 822 548 826 552
rect 830 548 834 552
rect 838 548 842 552
rect 902 548 906 552
rect 926 548 930 552
rect 934 548 938 552
rect 1046 548 1050 552
rect 1070 548 1074 552
rect 1150 548 1154 552
rect 1174 548 1178 552
rect 1198 548 1202 552
rect 1206 548 1210 552
rect 1222 548 1226 552
rect 1246 548 1250 552
rect 1254 548 1258 552
rect 1278 548 1282 552
rect 1310 548 1314 552
rect 1342 548 1346 552
rect 1366 548 1370 552
rect 1390 548 1394 552
rect 1398 548 1402 552
rect 1414 548 1418 552
rect 1438 548 1442 552
rect 1446 548 1450 552
rect 1454 548 1458 552
rect 1462 548 1466 552
rect 1494 548 1498 552
rect 1518 548 1522 552
rect 1598 548 1602 552
rect 1622 548 1626 552
rect 1630 548 1634 552
rect 1654 548 1658 552
rect 1734 548 1738 552
rect 1750 548 1754 552
rect 1758 548 1762 552
rect 1782 548 1786 552
rect 1790 548 1794 552
rect 1806 548 1810 552
rect 1830 548 1834 552
rect 1838 548 1842 552
rect 1862 548 1866 552
rect 1870 548 1874 552
rect 30 538 34 542
rect 86 538 90 542
rect 102 538 106 542
rect 126 538 130 542
rect 158 538 162 542
rect 214 538 218 542
rect 246 538 250 542
rect 270 540 274 544
rect 278 538 282 542
rect 342 538 346 542
rect 374 538 378 542
rect 398 538 402 542
rect 454 538 458 542
rect 502 538 506 542
rect 542 538 546 542
rect 614 538 618 542
rect 622 538 626 542
rect 662 538 666 542
rect 686 538 690 542
rect 734 538 738 542
rect 766 538 770 542
rect 798 538 802 542
rect 846 540 850 544
rect 878 538 882 542
rect 918 540 922 544
rect 950 538 954 542
rect 982 538 986 542
rect 998 538 1002 542
rect 1014 538 1018 542
rect 1118 538 1122 542
rect 1286 538 1290 542
rect 1318 538 1322 542
rect 1350 538 1354 542
rect 1486 538 1490 542
rect 1526 538 1530 542
rect 1542 538 1546 542
rect 1574 540 1578 544
rect 1702 538 1706 542
rect 62 528 66 532
rect 78 528 82 532
rect 94 528 98 532
rect 342 528 346 532
rect 406 528 410 532
rect 446 528 450 532
rect 550 528 554 532
rect 646 528 650 532
rect 654 528 658 532
rect 678 528 682 532
rect 766 528 770 532
rect 870 528 874 532
rect 958 528 962 532
rect 966 528 970 532
rect 990 528 994 532
rect 1022 528 1026 532
rect 1054 528 1058 532
rect 1094 528 1098 532
rect 1126 528 1130 532
rect 1190 528 1194 532
rect 1534 528 1538 532
rect 1678 528 1682 532
rect 1710 528 1714 532
rect 254 518 258 522
rect 470 518 474 522
rect 534 518 538 522
rect 638 518 642 522
rect 862 518 866 522
rect 1062 518 1066 522
rect 1134 518 1138 522
rect 1230 518 1234 522
rect 1262 518 1266 522
rect 1294 518 1298 522
rect 1502 518 1506 522
rect 1590 518 1594 522
rect 1646 518 1650 522
rect 1718 518 1722 522
rect 1846 518 1850 522
rect 46 488 50 492
rect 102 488 106 492
rect 158 488 162 492
rect 214 488 218 492
rect 278 488 282 492
rect 374 488 378 492
rect 430 488 434 492
rect 582 488 586 492
rect 622 488 626 492
rect 870 488 874 492
rect 910 488 914 492
rect 942 488 946 492
rect 982 488 986 492
rect 998 488 1002 492
rect 1110 488 1114 492
rect 1150 488 1154 492
rect 1214 488 1218 492
rect 1278 488 1282 492
rect 1326 488 1330 492
rect 1510 488 1514 492
rect 1566 488 1570 492
rect 1574 488 1578 492
rect 1814 488 1818 492
rect 1878 488 1882 492
rect 62 478 66 482
rect 110 478 114 482
rect 150 478 154 482
rect 222 478 226 482
rect 246 478 250 482
rect 310 478 314 482
rect 342 478 346 482
rect 382 478 386 482
rect 462 478 466 482
rect 502 478 506 482
rect 526 478 530 482
rect 590 478 594 482
rect 750 478 754 482
rect 814 478 818 482
rect 878 478 882 482
rect 934 478 938 482
rect 1054 478 1058 482
rect 1086 478 1090 482
rect 1142 478 1146 482
rect 1206 478 1210 482
rect 1270 478 1274 482
rect 1438 478 1442 482
rect 1470 478 1474 482
rect 1598 478 1602 482
rect 1726 478 1730 482
rect 1758 478 1762 482
rect 1854 478 1858 482
rect 6 468 10 472
rect 30 468 34 472
rect 94 468 98 472
rect 118 468 122 472
rect 174 466 178 470
rect 190 468 194 472
rect 238 468 242 472
rect 254 468 258 472
rect 286 468 290 472
rect 302 468 306 472
rect 334 468 338 472
rect 350 468 354 472
rect 390 468 394 472
rect 414 468 418 472
rect 462 468 466 472
rect 470 468 474 472
rect 534 468 538 472
rect 558 468 562 472
rect 598 468 602 472
rect 606 468 610 472
rect 622 468 626 472
rect 638 466 642 470
rect 22 458 26 462
rect 70 458 74 462
rect 86 458 90 462
rect 182 458 186 462
rect 198 458 202 462
rect 262 458 266 462
rect 318 458 322 462
rect 358 458 362 462
rect 486 458 490 462
rect 502 458 506 462
rect 566 458 570 462
rect 694 468 698 472
rect 718 468 722 472
rect 758 468 762 472
rect 814 468 818 472
rect 886 468 890 472
rect 926 468 930 472
rect 966 468 970 472
rect 974 468 978 472
rect 1078 468 1082 472
rect 1086 468 1090 472
rect 1110 468 1114 472
rect 1134 468 1138 472
rect 1166 466 1170 470
rect 1198 468 1202 472
rect 1262 468 1266 472
rect 1382 468 1386 472
rect 1430 468 1434 472
rect 1462 468 1466 472
rect 1494 466 1498 470
rect 1502 468 1506 472
rect 1526 466 1530 470
rect 1542 468 1546 472
rect 1598 468 1602 472
rect 1630 468 1634 472
rect 1638 468 1642 472
rect 1686 468 1690 472
rect 1726 468 1730 472
rect 1734 468 1738 472
rect 1766 468 1770 472
rect 1846 468 1850 472
rect 1862 468 1866 472
rect 670 458 674 462
rect 678 458 682 462
rect 726 458 730 462
rect 790 458 794 462
rect 806 458 810 462
rect 854 458 858 462
rect 958 458 962 462
rect 1014 458 1018 462
rect 1022 458 1026 462
rect 1174 458 1178 462
rect 1230 458 1234 462
rect 1238 458 1242 462
rect 1294 458 1298 462
rect 1302 458 1306 462
rect 1310 458 1314 462
rect 1334 458 1338 462
rect 1342 458 1346 462
rect 1366 458 1370 462
rect 1390 458 1394 462
rect 1406 458 1410 462
rect 1478 458 1482 462
rect 1550 458 1554 462
rect 1606 458 1610 462
rect 1622 458 1626 462
rect 1702 458 1706 462
rect 1718 458 1722 462
rect 1750 458 1754 462
rect 1798 458 1802 462
rect 1838 458 1842 462
rect 78 448 82 452
rect 438 448 442 452
rect 518 448 522 452
rect 630 448 634 452
rect 710 448 714 452
rect 742 448 746 452
rect 1030 448 1034 452
rect 46 438 50 442
rect 62 438 66 442
rect 454 438 458 442
rect 502 438 506 442
rect 990 438 994 442
rect 1110 438 1114 442
rect 1238 438 1242 442
rect 406 428 410 432
rect 1414 428 1418 432
rect 550 418 554 422
rect 902 418 906 422
rect 1182 418 1186 422
rect 1446 418 1450 422
rect 1574 418 1578 422
rect 1822 418 1826 422
rect 1878 418 1882 422
rect 174 388 178 392
rect 366 388 370 392
rect 390 388 394 392
rect 502 388 506 392
rect 590 388 594 392
rect 646 388 650 392
rect 670 388 674 392
rect 702 388 706 392
rect 1142 388 1146 392
rect 1414 388 1418 392
rect 1502 388 1506 392
rect 1830 388 1834 392
rect 414 378 418 382
rect 958 378 962 382
rect 1838 378 1842 382
rect 382 368 386 372
rect 510 368 514 372
rect 1358 368 1362 372
rect 1614 368 1618 372
rect 198 358 202 362
rect 54 348 58 352
rect 62 348 66 352
rect 126 348 130 352
rect 142 348 146 352
rect 158 348 162 352
rect 454 358 458 362
rect 494 358 498 362
rect 550 358 554 362
rect 758 358 762 362
rect 768 358 772 362
rect 1038 358 1042 362
rect 1334 358 1338 362
rect 1358 358 1362 362
rect 1558 358 1562 362
rect 1686 358 1690 362
rect 246 348 250 352
rect 374 348 378 352
rect 390 348 394 352
rect 446 348 450 352
rect 478 348 482 352
rect 502 348 506 352
rect 574 348 578 352
rect 638 348 642 352
rect 662 348 666 352
rect 718 348 722 352
rect 726 348 730 352
rect 774 348 778 352
rect 806 348 810 352
rect 814 348 818 352
rect 854 348 858 352
rect 942 348 946 352
rect 966 348 970 352
rect 982 348 986 352
rect 1046 348 1050 352
rect 1102 348 1106 352
rect 1118 348 1122 352
rect 1190 348 1194 352
rect 1198 348 1202 352
rect 6 338 10 342
rect 62 338 66 342
rect 94 338 98 342
rect 150 338 154 342
rect 182 338 186 342
rect 222 338 226 342
rect 230 338 234 342
rect 278 338 282 342
rect 310 338 314 342
rect 342 338 346 342
rect 358 338 362 342
rect 454 338 458 342
rect 486 338 490 342
rect 542 340 546 344
rect 550 338 554 342
rect 582 338 586 342
rect 606 338 610 342
rect 686 338 690 342
rect 742 338 746 342
rect 830 338 834 342
rect 846 338 850 342
rect 870 338 874 342
rect 886 338 890 342
rect 934 338 938 342
rect 1014 338 1018 342
rect 1070 338 1074 342
rect 1118 338 1122 342
rect 1238 348 1242 352
rect 1246 348 1250 352
rect 1350 348 1354 352
rect 1382 348 1386 352
rect 1462 348 1466 352
rect 1550 348 1554 352
rect 1582 348 1586 352
rect 1598 348 1602 352
rect 1662 348 1666 352
rect 1726 348 1730 352
rect 1766 348 1770 352
rect 1878 348 1882 352
rect 1222 338 1226 342
rect 1278 338 1282 342
rect 1366 338 1370 342
rect 1398 338 1402 342
rect 1526 338 1530 342
rect 1558 338 1562 342
rect 1590 338 1594 342
rect 1646 338 1650 342
rect 1702 338 1706 342
rect 1718 338 1722 342
rect 1750 338 1754 342
rect 1798 338 1802 342
rect 1814 338 1818 342
rect 78 328 82 332
rect 254 328 258 332
rect 350 328 354 332
rect 422 328 426 332
rect 622 328 626 332
rect 694 328 698 332
rect 750 328 754 332
rect 822 328 826 332
rect 878 328 882 332
rect 1022 328 1026 332
rect 1030 328 1034 332
rect 1078 328 1082 332
rect 1230 328 1234 332
rect 1270 328 1274 332
rect 1302 328 1306 332
rect 1390 328 1394 332
rect 1446 328 1450 332
rect 1462 328 1466 332
rect 1526 328 1530 332
rect 1622 328 1626 332
rect 1710 328 1714 332
rect 1806 328 1810 332
rect 30 318 34 322
rect 262 318 266 322
rect 430 318 434 322
rect 526 318 530 322
rect 670 318 674 322
rect 790 318 794 322
rect 910 318 914 322
rect 1054 318 1058 322
rect 1086 318 1090 322
rect 1262 318 1266 322
rect 1326 318 1330 322
rect 1422 318 1426 322
rect 1486 318 1490 322
rect 1534 318 1538 322
rect 1614 318 1618 322
rect 1678 318 1682 322
rect 1742 318 1746 322
rect 70 288 74 292
rect 214 288 218 292
rect 222 288 226 292
rect 294 288 298 292
rect 326 288 330 292
rect 366 288 370 292
rect 486 288 490 292
rect 542 288 546 292
rect 582 288 586 292
rect 710 288 714 292
rect 1118 288 1122 292
rect 1150 288 1154 292
rect 1278 288 1282 292
rect 1430 288 1434 292
rect 1526 288 1530 292
rect 1646 288 1650 292
rect 1710 288 1714 292
rect 1798 288 1802 292
rect 1838 288 1842 292
rect 94 278 98 282
rect 102 278 106 282
rect 166 278 170 282
rect 182 278 186 282
rect 302 278 306 282
rect 358 278 362 282
rect 406 278 410 282
rect 446 278 450 282
rect 574 278 578 282
rect 638 278 642 282
rect 654 278 658 282
rect 718 278 722 282
rect 806 278 810 282
rect 838 278 842 282
rect 846 278 850 282
rect 878 278 882 282
rect 910 278 914 282
rect 934 278 938 282
rect 1014 278 1018 282
rect 1030 278 1034 282
rect 1110 278 1114 282
rect 1174 278 1178 282
rect 1182 278 1186 282
rect 1270 278 1274 282
rect 1302 278 1306 282
rect 1398 278 1402 282
rect 1486 278 1490 282
rect 1494 278 1498 282
rect 1574 278 1578 282
rect 1614 278 1618 282
rect 1702 278 1706 282
rect 1742 278 1746 282
rect 1830 278 1834 282
rect 6 268 10 272
rect 30 268 34 272
rect 110 268 114 272
rect 190 268 194 272
rect 270 268 274 272
rect 310 268 314 272
rect 334 268 338 272
rect 390 268 394 272
rect 462 268 466 272
rect 566 268 570 272
rect 638 268 642 272
rect 678 268 682 272
rect 726 268 730 272
rect 798 268 802 272
rect 830 268 834 272
rect 854 268 858 272
rect 886 268 890 272
rect 934 268 938 272
rect 958 266 962 270
rect 998 268 1002 272
rect 1006 268 1010 272
rect 1022 268 1026 272
rect 1054 268 1058 272
rect 1062 268 1066 272
rect 1102 268 1106 272
rect 1142 268 1146 272
rect 1166 268 1170 272
rect 1190 268 1194 272
rect 1238 268 1242 272
rect 1262 268 1266 272
rect 1294 268 1298 272
rect 1334 268 1338 272
rect 1390 268 1394 272
rect 1406 268 1410 272
rect 1446 266 1450 270
rect 1478 268 1482 272
rect 1510 268 1514 272
rect 1550 268 1554 272
rect 1606 268 1610 272
rect 1622 268 1626 272
rect 1670 268 1674 272
rect 1694 268 1698 272
rect 1726 266 1730 270
rect 1758 268 1762 272
rect 1782 266 1786 270
rect 1830 268 1834 272
rect 1886 268 1890 272
rect 22 258 26 262
rect 46 258 50 262
rect 54 258 58 262
rect 62 258 66 262
rect 86 258 90 262
rect 142 258 146 262
rect 166 258 170 262
rect 198 258 202 262
rect 238 258 242 262
rect 262 258 266 262
rect 278 258 282 262
rect 342 258 346 262
rect 382 258 386 262
rect 414 258 418 262
rect 430 258 434 262
rect 470 258 474 262
rect 502 258 506 262
rect 510 258 514 262
rect 518 258 522 262
rect 526 258 530 262
rect 598 258 602 262
rect 646 258 650 262
rect 662 258 666 262
rect 686 258 690 262
rect 694 258 698 262
rect 758 258 762 262
rect 942 258 946 262
rect 990 258 994 262
rect 1134 258 1138 262
rect 1214 258 1218 262
rect 1230 258 1234 262
rect 1246 258 1250 262
rect 1310 258 1314 262
rect 1326 258 1330 262
rect 1358 258 1362 262
rect 1422 258 1426 262
rect 1454 258 1458 262
rect 1518 258 1522 262
rect 1542 258 1546 262
rect 1566 258 1570 262
rect 1766 258 1770 262
rect 1806 258 1810 262
rect 1846 258 1850 262
rect 158 248 162 252
rect 358 248 362 252
rect 70 238 74 242
rect 406 238 410 242
rect 438 248 442 252
rect 462 248 466 252
rect 478 248 482 252
rect 550 248 554 252
rect 774 248 778 252
rect 1022 248 1026 252
rect 1078 248 1082 252
rect 1086 248 1090 252
rect 1334 248 1338 252
rect 1558 248 1562 252
rect 1590 248 1594 252
rect 1494 238 1498 242
rect 1574 238 1578 242
rect 1678 238 1682 242
rect 246 218 250 222
rect 782 218 786 222
rect 814 218 818 222
rect 870 218 874 222
rect 902 218 906 222
rect 1206 218 1210 222
rect 1278 218 1282 222
rect 1462 218 1466 222
rect 1742 218 1746 222
rect 110 188 114 192
rect 174 188 178 192
rect 222 188 226 192
rect 238 188 242 192
rect 286 188 290 192
rect 374 188 378 192
rect 390 188 394 192
rect 398 188 402 192
rect 446 188 450 192
rect 534 188 538 192
rect 886 188 890 192
rect 1070 188 1074 192
rect 1142 188 1146 192
rect 1350 188 1354 192
rect 1494 188 1498 192
rect 1742 188 1746 192
rect 1750 188 1754 192
rect 1838 188 1842 192
rect 694 178 698 182
rect 798 178 802 182
rect 86 168 90 172
rect 182 168 186 172
rect 214 168 218 172
rect 438 168 442 172
rect 806 168 810 172
rect 1150 168 1154 172
rect 1190 168 1194 172
rect 1550 168 1554 172
rect 102 158 106 162
rect 230 158 234 162
rect 454 158 458 162
rect 638 158 642 162
rect 790 158 794 162
rect 950 158 954 162
rect 1094 158 1098 162
rect 1134 158 1138 162
rect 1318 158 1322 162
rect 1574 158 1578 162
rect 1774 158 1778 162
rect 78 148 82 152
rect 94 148 98 152
rect 142 148 146 152
rect 190 148 194 152
rect 198 148 202 152
rect 222 148 226 152
rect 302 148 306 152
rect 414 148 418 152
rect 446 148 450 152
rect 486 148 490 152
rect 502 148 506 152
rect 526 148 530 152
rect 558 148 562 152
rect 566 148 570 152
rect 670 148 674 152
rect 686 148 690 152
rect 710 148 714 152
rect 758 148 762 152
rect 766 148 770 152
rect 798 148 802 152
rect 830 148 834 152
rect 910 148 914 152
rect 918 148 922 152
rect 926 148 930 152
rect 958 148 962 152
rect 982 148 986 152
rect 1086 148 1090 152
rect 1142 148 1146 152
rect 1182 148 1186 152
rect 1206 148 1210 152
rect 1294 148 1298 152
rect 1326 148 1330 152
rect 1342 148 1346 152
rect 1366 148 1370 152
rect 1390 148 1394 152
rect 1406 148 1410 152
rect 1414 148 1418 152
rect 1446 148 1450 152
rect 1462 148 1466 152
rect 1486 148 1490 152
rect 1510 148 1514 152
rect 1526 148 1530 152
rect 1534 148 1538 152
rect 1558 148 1562 152
rect 1606 148 1610 152
rect 1622 148 1626 152
rect 1630 148 1634 152
rect 1646 148 1650 152
rect 1670 148 1674 152
rect 1678 148 1682 152
rect 1702 148 1706 152
rect 1766 148 1770 152
rect 1814 148 1818 152
rect 1822 148 1826 152
rect 1846 148 1850 152
rect 6 138 10 142
rect 54 138 58 142
rect 134 138 138 142
rect 150 138 154 142
rect 254 138 258 142
rect 318 138 322 142
rect 326 138 330 142
rect 422 138 426 142
rect 470 138 474 142
rect 494 138 498 142
rect 542 138 546 142
rect 550 138 554 142
rect 598 138 602 142
rect 622 138 626 142
rect 662 138 666 142
rect 718 138 722 142
rect 742 138 746 142
rect 822 138 826 142
rect 854 138 858 142
rect 870 138 874 142
rect 902 140 906 144
rect 950 138 954 142
rect 998 138 1002 142
rect 1014 138 1018 142
rect 1062 138 1066 142
rect 1094 138 1098 142
rect 1118 138 1122 142
rect 1190 138 1194 142
rect 1214 138 1218 142
rect 1230 138 1234 142
rect 1254 138 1258 142
rect 1262 140 1266 144
rect 1310 138 1314 142
rect 1318 138 1322 142
rect 1374 138 1378 142
rect 1382 138 1386 142
rect 1422 140 1426 144
rect 1470 138 1474 142
rect 1590 138 1594 142
rect 1710 138 1714 142
rect 1726 138 1730 142
rect 1774 138 1778 142
rect 1798 138 1802 142
rect 70 128 74 132
rect 110 128 114 132
rect 134 128 138 132
rect 158 128 162 132
rect 166 128 170 132
rect 262 128 266 132
rect 278 128 282 132
rect 318 128 322 132
rect 350 128 354 132
rect 382 128 386 132
rect 462 128 466 132
rect 606 128 610 132
rect 614 128 618 132
rect 646 128 650 132
rect 654 128 658 132
rect 726 128 730 132
rect 750 128 754 132
rect 878 128 882 132
rect 1006 128 1010 132
rect 1126 128 1130 132
rect 1222 128 1226 132
rect 1246 128 1250 132
rect 1598 128 1602 132
rect 1718 128 1722 132
rect 1806 128 1810 132
rect 30 118 34 122
rect 62 118 66 122
rect 270 118 274 122
rect 286 118 290 122
rect 390 118 394 122
rect 534 118 538 122
rect 782 118 786 122
rect 846 118 850 122
rect 974 118 978 122
rect 1038 118 1042 122
rect 1166 118 1170 122
rect 1438 118 1442 122
rect 1662 118 1666 122
rect 1750 118 1754 122
rect 246 88 250 92
rect 302 88 306 92
rect 334 88 338 92
rect 374 88 378 92
rect 478 88 482 92
rect 518 88 522 92
rect 638 88 642 92
rect 670 88 674 92
rect 774 88 778 92
rect 934 88 938 92
rect 966 88 970 92
rect 1038 88 1042 92
rect 1102 88 1106 92
rect 1110 88 1114 92
rect 1382 88 1386 92
rect 1478 88 1482 92
rect 1510 88 1514 92
rect 1670 88 1674 92
rect 1718 88 1722 92
rect 1742 88 1746 92
rect 1798 88 1802 92
rect 1806 88 1810 92
rect 1830 88 1834 92
rect 102 78 106 82
rect 6 68 10 72
rect 30 68 34 72
rect 182 78 186 82
rect 406 78 410 82
rect 494 78 498 82
rect 534 78 538 82
rect 726 78 730 82
rect 766 78 770 82
rect 998 78 1002 82
rect 1198 78 1202 82
rect 1294 78 1298 82
rect 1326 78 1330 82
rect 1438 78 1442 82
rect 118 68 122 72
rect 174 68 178 72
rect 214 68 218 72
rect 222 68 226 72
rect 270 68 274 72
rect 278 68 282 72
rect 310 68 314 72
rect 390 66 394 70
rect 398 68 402 72
rect 502 68 506 72
rect 582 68 586 72
rect 614 68 618 72
rect 662 68 666 72
rect 694 68 698 72
rect 718 68 722 72
rect 766 68 770 72
rect 782 68 786 72
rect 830 68 834 72
rect 838 68 842 72
rect 894 68 898 72
rect 902 68 906 72
rect 958 68 962 72
rect 982 66 986 70
rect 998 68 1002 72
rect 1030 68 1034 72
rect 1126 66 1130 70
rect 1166 68 1170 72
rect 1190 68 1194 72
rect 1238 68 1242 72
rect 1246 66 1250 70
rect 22 58 26 62
rect 46 58 50 62
rect 54 58 58 62
rect 62 58 66 62
rect 78 58 82 62
rect 86 58 90 62
rect 150 58 154 62
rect 174 58 178 62
rect 286 58 290 62
rect 318 58 322 62
rect 358 58 362 62
rect 430 58 434 62
rect 446 58 450 62
rect 462 58 466 62
rect 486 58 490 62
rect 590 58 594 62
rect 686 58 690 62
rect 710 58 714 62
rect 790 58 794 62
rect 798 58 802 62
rect 854 58 858 62
rect 910 58 914 62
rect 926 58 930 62
rect 950 58 954 62
rect 1054 58 1058 62
rect 1062 58 1066 62
rect 1086 58 1090 62
rect 1158 58 1162 62
rect 1166 58 1170 62
rect 1214 58 1218 62
rect 1230 58 1234 62
rect 1334 68 1338 72
rect 1342 68 1346 72
rect 1350 68 1354 72
rect 1358 68 1362 72
rect 1406 68 1410 72
rect 1414 68 1418 72
rect 1502 78 1506 82
rect 1534 78 1538 82
rect 1622 78 1626 82
rect 1638 78 1642 82
rect 1854 78 1858 82
rect 1454 68 1458 72
rect 1470 68 1474 72
rect 1510 68 1514 72
rect 1526 68 1530 72
rect 1566 68 1570 72
rect 1694 68 1698 72
rect 1774 68 1778 72
rect 1782 66 1786 70
rect 1846 68 1850 72
rect 1278 58 1282 62
rect 1366 58 1370 62
rect 1574 58 1578 62
rect 1646 58 1650 62
rect 1654 58 1658 62
rect 1678 58 1682 62
rect 1702 58 1706 62
rect 1734 58 1738 62
rect 1758 58 1762 62
rect 1766 58 1770 62
rect 1822 58 1826 62
rect 198 48 202 52
rect 342 48 346 52
rect 366 48 370 52
rect 398 48 402 52
rect 822 48 826 52
rect 846 48 850 52
rect 886 48 890 52
rect 1142 48 1146 52
rect 1206 48 1210 52
rect 1334 48 1338 52
rect 1390 48 1394 52
rect 1598 48 1602 52
rect 70 38 74 42
rect 350 38 354 42
rect 702 38 706 42
rect 862 38 866 42
rect 878 38 882 42
rect 1222 38 1226 42
rect 1510 38 1514 42
rect 870 28 874 32
rect 606 18 610 22
rect 814 18 818 22
rect 1078 18 1082 22
rect 1590 18 1594 22
<< metal2 >>
rect 54 1192 57 1231
rect 102 1192 105 1231
rect 206 1172 209 1231
rect 342 1192 345 1231
rect 558 1182 561 1231
rect 574 1228 585 1231
rect 558 1172 561 1178
rect 6 1162 9 1168
rect 206 1152 209 1168
rect 26 1148 33 1151
rect 74 1148 81 1151
rect 30 1142 33 1148
rect 78 1142 81 1148
rect 122 1148 129 1151
rect 94 1131 97 1148
rect 126 1142 129 1148
rect 274 1148 278 1151
rect 46 1082 49 1088
rect 6 1072 9 1078
rect 46 1062 49 1078
rect 78 1072 81 1128
rect 90 1128 97 1131
rect 86 1082 89 1088
rect 134 1072 137 1118
rect 142 1092 145 1148
rect 286 1142 289 1148
rect 334 1142 337 1158
rect 150 1132 153 1138
rect 222 1122 225 1138
rect 246 1122 249 1128
rect 198 1072 201 1108
rect 22 1052 25 1058
rect 38 1042 41 1058
rect 54 1042 57 1048
rect 6 962 9 968
rect 26 948 33 951
rect 30 942 33 948
rect 30 861 33 868
rect 26 858 33 861
rect 26 748 33 751
rect 30 742 33 748
rect 6 662 9 668
rect 30 661 33 668
rect 26 658 33 661
rect 38 622 41 1038
rect 62 1032 65 1048
rect 62 942 65 1018
rect 70 952 73 1018
rect 62 922 65 928
rect 62 882 65 888
rect 70 872 73 918
rect 78 912 81 1068
rect 94 1062 97 1068
rect 118 1018 126 1021
rect 118 952 121 1018
rect 134 942 137 998
rect 142 952 145 1028
rect 166 972 169 1018
rect 174 1012 177 1048
rect 182 952 185 958
rect 102 932 105 938
rect 98 928 102 931
rect 126 922 129 938
rect 78 862 81 888
rect 86 882 89 918
rect 94 851 97 908
rect 102 862 105 868
rect 126 861 129 868
rect 122 858 129 861
rect 94 848 105 851
rect 94 742 97 818
rect 102 742 105 848
rect 134 752 137 938
rect 158 922 161 928
rect 158 872 161 878
rect 174 792 177 868
rect 86 732 89 740
rect 102 731 105 738
rect 94 728 105 731
rect 70 662 73 718
rect 86 692 89 728
rect 6 562 9 568
rect 26 548 33 551
rect 30 542 33 548
rect 46 492 49 558
rect 62 532 65 548
rect 78 541 81 598
rect 94 542 97 728
rect 130 718 137 721
rect 110 672 113 678
rect 134 672 137 718
rect 158 712 161 748
rect 182 732 185 948
rect 206 942 209 948
rect 190 932 193 938
rect 214 871 217 1058
rect 222 1052 225 1068
rect 230 1062 233 1098
rect 238 1082 241 1118
rect 246 1072 249 1078
rect 254 1062 257 1128
rect 262 1082 265 1118
rect 270 1072 273 1098
rect 222 882 225 918
rect 230 892 233 918
rect 214 868 222 871
rect 190 752 193 758
rect 198 732 201 818
rect 238 801 241 968
rect 254 962 257 1058
rect 286 1042 289 1138
rect 294 1092 297 1118
rect 310 1112 313 1118
rect 350 1112 353 1168
rect 418 1158 425 1161
rect 422 1152 425 1158
rect 362 1148 369 1151
rect 366 1142 369 1148
rect 554 1148 558 1151
rect 382 1122 385 1148
rect 390 1142 393 1148
rect 398 1112 401 1148
rect 574 1142 577 1228
rect 622 1212 625 1231
rect 742 1192 745 1231
rect 614 1152 617 1178
rect 822 1152 825 1231
rect 878 1212 881 1231
rect 846 1152 849 1168
rect 862 1152 865 1208
rect 886 1152 889 1158
rect 934 1152 937 1158
rect 634 1148 641 1151
rect 718 1148 726 1151
rect 882 1148 886 1151
rect 582 1142 585 1148
rect 334 1082 337 1088
rect 310 1062 313 1068
rect 334 1062 337 1078
rect 342 1062 345 1088
rect 350 1082 353 1108
rect 350 1072 353 1078
rect 382 1072 385 1108
rect 398 1092 401 1108
rect 414 1102 417 1118
rect 430 1112 433 1138
rect 446 1122 449 1128
rect 454 1102 457 1118
rect 470 1112 473 1140
rect 618 1138 630 1141
rect 486 1132 489 1138
rect 534 1132 537 1138
rect 542 1122 545 1128
rect 574 1122 577 1138
rect 590 1132 593 1138
rect 638 1132 641 1148
rect 694 1142 697 1148
rect 718 1142 721 1148
rect 758 1132 761 1148
rect 790 1138 798 1141
rect 502 1118 510 1121
rect 398 1052 401 1068
rect 406 1062 409 1088
rect 478 1072 481 1098
rect 262 962 265 1008
rect 254 932 257 938
rect 262 892 265 958
rect 278 952 281 1018
rect 286 941 289 1028
rect 318 962 321 1018
rect 350 942 353 958
rect 282 938 289 941
rect 294 892 297 918
rect 262 872 265 878
rect 310 872 313 918
rect 334 912 337 938
rect 346 928 350 931
rect 358 922 361 940
rect 230 798 241 801
rect 214 752 217 758
rect 230 742 233 798
rect 230 732 233 738
rect 246 732 249 858
rect 270 792 273 858
rect 350 822 353 858
rect 286 752 289 818
rect 318 742 321 748
rect 350 742 353 778
rect 358 772 361 818
rect 366 792 369 908
rect 374 872 377 918
rect 390 881 393 888
rect 386 878 393 881
rect 398 842 401 1048
rect 414 1022 417 1058
rect 438 952 441 1068
rect 446 1012 449 1058
rect 462 1042 465 1058
rect 450 948 454 951
rect 430 922 433 940
rect 406 902 409 918
rect 406 862 409 878
rect 414 871 417 918
rect 430 902 433 918
rect 422 882 425 898
rect 414 868 422 871
rect 166 701 169 728
rect 158 698 169 701
rect 142 662 145 668
rect 158 662 161 698
rect 174 691 177 718
rect 198 692 201 718
rect 326 692 329 728
rect 350 721 353 738
rect 374 731 377 768
rect 414 752 417 838
rect 438 832 441 888
rect 446 882 449 948
rect 462 882 465 958
rect 470 892 473 918
rect 478 872 481 978
rect 486 972 489 1038
rect 494 962 497 1118
rect 502 1032 505 1118
rect 510 1082 513 1098
rect 510 992 513 1068
rect 550 1062 553 1098
rect 558 1062 561 1088
rect 566 1072 569 1098
rect 574 1081 577 1118
rect 582 1092 585 1108
rect 574 1078 585 1081
rect 582 1062 585 1078
rect 526 1052 529 1058
rect 534 982 537 1018
rect 582 1002 585 1048
rect 494 952 497 958
rect 558 942 561 948
rect 530 938 534 941
rect 566 932 569 938
rect 518 928 534 931
rect 518 922 521 928
rect 574 922 577 928
rect 526 892 529 918
rect 582 892 585 898
rect 534 882 537 888
rect 470 862 473 868
rect 502 842 505 878
rect 582 870 585 888
rect 590 872 593 1068
rect 606 1062 609 1128
rect 630 1122 633 1128
rect 622 1062 625 1108
rect 662 1102 665 1118
rect 766 1102 769 1138
rect 670 1091 673 1098
rect 662 1088 673 1091
rect 630 1062 633 1088
rect 662 1062 665 1088
rect 734 1081 737 1088
rect 730 1078 737 1081
rect 686 1062 689 1068
rect 650 1058 654 1061
rect 674 1058 678 1061
rect 622 972 625 1058
rect 718 1042 721 1068
rect 766 1062 769 1088
rect 774 1062 777 1118
rect 646 992 649 1038
rect 654 1032 657 1038
rect 606 932 609 938
rect 606 872 609 928
rect 614 922 617 938
rect 566 862 569 868
rect 622 862 625 878
rect 422 752 425 808
rect 382 742 385 748
rect 362 728 369 731
rect 374 728 385 731
rect 394 728 401 731
rect 350 718 361 721
rect 174 688 185 691
rect 166 681 169 688
rect 166 678 174 681
rect 182 672 185 688
rect 206 682 209 688
rect 270 682 273 688
rect 230 672 233 678
rect 294 672 297 688
rect 358 682 361 718
rect 366 692 369 728
rect 358 672 361 678
rect 382 672 385 728
rect 398 722 401 728
rect 406 671 409 678
rect 414 671 417 748
rect 422 682 425 688
rect 406 670 417 671
rect 118 632 121 648
rect 190 592 193 668
rect 302 662 305 668
rect 350 662 353 668
rect 410 668 417 670
rect 286 652 289 658
rect 310 622 313 658
rect 102 542 105 558
rect 70 538 81 541
rect 90 538 94 541
rect 30 472 33 478
rect 70 472 73 538
rect 82 528 89 531
rect 98 528 105 531
rect 6 462 9 468
rect 70 462 73 468
rect 86 462 89 528
rect 102 492 105 528
rect 110 482 113 578
rect 218 538 222 541
rect 94 472 97 478
rect 62 352 65 438
rect 54 342 57 348
rect 70 341 73 458
rect 78 362 81 448
rect 110 412 113 478
rect 118 462 121 468
rect 66 338 73 341
rect 70 331 73 338
rect 70 328 78 331
rect 6 262 9 268
rect 30 261 33 268
rect 54 262 57 318
rect 102 291 105 368
rect 126 362 129 538
rect 158 492 161 538
rect 238 532 241 548
rect 246 542 249 608
rect 366 562 369 618
rect 278 542 281 558
rect 302 532 305 548
rect 350 541 353 548
rect 346 538 353 541
rect 374 542 377 568
rect 214 492 217 528
rect 254 482 257 518
rect 278 492 281 528
rect 366 522 369 528
rect 174 470 177 478
rect 238 472 241 478
rect 94 288 105 291
rect 94 282 97 288
rect 110 272 113 338
rect 126 292 129 348
rect 150 342 153 408
rect 174 392 177 448
rect 182 372 185 458
rect 190 452 193 468
rect 114 268 121 271
rect 26 258 33 261
rect 62 162 65 258
rect 70 232 73 238
rect 110 192 113 258
rect 54 142 57 158
rect 6 92 9 138
rect 30 112 33 118
rect 6 62 9 68
rect 30 61 33 68
rect 26 58 33 61
rect 46 62 49 118
rect 54 62 57 108
rect 62 62 65 68
rect 70 42 73 108
rect 86 92 89 168
rect 102 162 105 168
rect 94 142 97 148
rect 86 62 89 88
rect 94 82 97 138
rect 118 72 121 268
rect 134 142 137 318
rect 150 292 153 338
rect 182 302 185 338
rect 182 282 185 298
rect 198 282 201 358
rect 214 292 217 468
rect 222 342 225 418
rect 246 352 249 478
rect 306 468 310 471
rect 262 462 265 468
rect 334 462 337 468
rect 342 412 345 478
rect 342 342 345 388
rect 214 262 217 278
rect 142 192 145 258
rect 198 252 201 258
rect 182 172 185 228
rect 214 172 217 258
rect 230 251 233 338
rect 246 251 249 338
rect 222 248 233 251
rect 238 248 249 251
rect 254 272 257 328
rect 262 292 265 318
rect 326 292 329 338
rect 222 192 225 248
rect 230 172 233 238
rect 238 192 241 248
rect 254 241 257 268
rect 262 262 265 288
rect 294 281 297 288
rect 342 282 345 338
rect 350 332 353 468
rect 358 372 361 458
rect 366 392 369 518
rect 374 492 377 508
rect 390 481 393 658
rect 430 592 433 648
rect 438 632 441 828
rect 450 818 457 821
rect 454 762 457 818
rect 494 812 497 818
rect 478 758 486 761
rect 454 752 457 758
rect 478 752 481 758
rect 510 752 513 828
rect 526 761 529 818
rect 518 758 529 761
rect 542 758 550 761
rect 462 712 465 718
rect 454 662 457 668
rect 398 542 401 558
rect 386 478 393 481
rect 390 392 393 468
rect 414 422 417 468
rect 422 412 425 568
rect 438 562 441 628
rect 430 492 433 548
rect 454 542 457 548
rect 462 532 465 678
rect 470 672 473 738
rect 510 662 513 748
rect 518 742 521 758
rect 542 752 545 758
rect 526 742 529 748
rect 518 682 521 728
rect 526 692 529 728
rect 550 672 553 688
rect 558 672 561 818
rect 574 742 577 758
rect 582 682 585 728
rect 606 672 609 738
rect 622 692 625 838
rect 630 732 633 918
rect 638 902 641 948
rect 670 942 673 948
rect 678 942 681 948
rect 662 932 665 938
rect 726 932 729 938
rect 646 882 649 928
rect 638 751 641 818
rect 646 782 649 878
rect 638 748 649 751
rect 638 732 641 738
rect 646 732 649 748
rect 662 742 665 928
rect 678 872 681 928
rect 694 882 697 918
rect 734 911 737 958
rect 742 952 745 1048
rect 750 1042 753 1058
rect 750 972 753 988
rect 742 921 745 948
rect 742 918 753 921
rect 734 908 745 911
rect 726 872 729 878
rect 742 862 745 908
rect 750 862 753 918
rect 758 912 761 1058
rect 790 1002 793 1138
rect 806 1112 809 1128
rect 814 1112 817 1148
rect 846 1142 849 1148
rect 814 1072 817 1088
rect 798 1062 801 1068
rect 798 992 801 998
rect 790 912 793 928
rect 742 852 745 858
rect 750 842 753 858
rect 758 842 761 888
rect 774 882 777 888
rect 790 832 793 858
rect 806 832 809 1068
rect 814 1062 817 1068
rect 814 952 817 998
rect 822 942 825 1138
rect 846 1062 849 1068
rect 830 1032 833 1058
rect 846 1012 849 1058
rect 862 1032 865 1148
rect 878 1142 881 1148
rect 894 1142 897 1148
rect 910 1092 913 1118
rect 870 1062 873 1078
rect 926 1062 929 1148
rect 934 1082 937 1148
rect 950 1141 953 1178
rect 942 1138 953 1141
rect 942 1072 945 1138
rect 950 1062 953 1078
rect 958 1062 961 1231
rect 982 1152 985 1231
rect 966 1072 969 1148
rect 990 1142 993 1148
rect 998 1142 1001 1231
rect 1022 1152 1025 1158
rect 1062 1152 1065 1231
rect 1286 1158 1294 1161
rect 1286 1152 1289 1158
rect 1350 1152 1353 1231
rect 1342 1148 1350 1151
rect 974 1132 977 1138
rect 1006 1132 1009 1138
rect 1014 1112 1017 1148
rect 978 1068 982 1071
rect 990 1062 993 1108
rect 998 1082 1001 1098
rect 902 1032 905 1058
rect 862 962 865 1018
rect 894 952 897 1008
rect 910 992 913 1008
rect 838 912 841 918
rect 854 912 857 948
rect 902 942 905 958
rect 934 952 937 1058
rect 958 1052 961 1058
rect 982 952 985 1018
rect 998 992 1001 1078
rect 1006 1072 1009 1088
rect 1054 1082 1057 1118
rect 1062 1072 1065 1148
rect 1078 1102 1081 1128
rect 1078 1072 1081 1078
rect 1054 992 1057 1058
rect 1086 1052 1089 1078
rect 1102 1062 1105 1118
rect 1118 1062 1121 1148
rect 1186 1138 1193 1141
rect 1158 1132 1161 1138
rect 1166 1072 1169 1128
rect 1174 1072 1177 1078
rect 1126 1062 1129 1068
rect 1150 1062 1153 1068
rect 1150 1052 1153 1058
rect 1086 1012 1089 1048
rect 998 952 1001 958
rect 1070 952 1073 958
rect 1118 952 1121 958
rect 1166 951 1169 1018
rect 1182 982 1185 1058
rect 1190 1042 1193 1138
rect 1198 1062 1201 1068
rect 1206 962 1209 1018
rect 1214 992 1217 1148
rect 1230 1142 1233 1148
rect 1238 1112 1241 1118
rect 1254 1112 1257 1148
rect 1254 1102 1257 1108
rect 1238 1081 1241 1088
rect 1234 1078 1241 1081
rect 1254 1062 1257 1098
rect 1262 1092 1265 1148
rect 1318 1132 1321 1138
rect 1270 1102 1273 1118
rect 1278 1062 1281 1118
rect 1334 1112 1337 1118
rect 1262 1002 1265 1028
rect 1206 952 1209 958
rect 1230 952 1233 958
rect 1238 952 1241 988
rect 1262 952 1265 998
rect 1166 948 1177 951
rect 830 872 833 878
rect 822 862 825 868
rect 742 818 750 821
rect 686 752 689 808
rect 670 741 673 748
rect 670 738 681 741
rect 542 652 545 658
rect 582 618 590 621
rect 486 582 489 618
rect 494 552 497 588
rect 510 552 513 578
rect 542 542 545 618
rect 558 592 561 618
rect 582 552 585 618
rect 606 552 609 578
rect 622 542 625 658
rect 638 652 641 658
rect 446 522 449 528
rect 474 518 481 521
rect 462 482 465 488
rect 462 472 465 478
rect 438 452 441 468
rect 382 372 385 378
rect 358 342 361 368
rect 390 352 393 368
rect 374 342 377 348
rect 366 292 369 328
rect 390 312 393 348
rect 406 282 409 408
rect 438 372 441 448
rect 438 352 441 368
rect 446 352 449 358
rect 422 332 425 348
rect 454 342 457 358
rect 462 352 465 468
rect 478 352 481 518
rect 526 492 529 518
rect 526 482 529 488
rect 502 472 505 478
rect 534 472 537 518
rect 502 392 505 408
rect 518 392 521 448
rect 534 422 537 458
rect 510 372 513 378
rect 294 278 302 281
rect 302 272 305 278
rect 406 272 409 278
rect 246 238 257 241
rect 246 222 249 238
rect 142 102 145 148
rect 150 142 153 148
rect 182 122 185 168
rect 190 142 193 148
rect 174 72 177 118
rect 182 82 185 98
rect 190 72 193 138
rect 198 102 201 148
rect 214 91 217 168
rect 230 162 233 168
rect 222 152 225 158
rect 246 132 249 218
rect 278 162 281 258
rect 286 192 289 268
rect 310 222 313 268
rect 390 262 393 268
rect 422 261 425 328
rect 446 282 449 308
rect 486 292 489 338
rect 462 262 465 268
rect 422 258 430 261
rect 342 222 345 258
rect 382 232 385 258
rect 254 132 257 138
rect 278 132 281 158
rect 306 148 313 151
rect 246 112 249 128
rect 262 102 265 128
rect 286 122 289 138
rect 274 118 278 121
rect 246 92 249 98
rect 214 88 225 91
rect 118 52 121 68
rect 198 52 201 88
rect 214 72 217 78
rect 222 72 225 88
rect 278 72 281 118
rect 222 -22 225 68
rect 270 -22 273 68
rect 286 62 289 118
rect 302 92 305 138
rect 310 131 313 148
rect 318 142 321 148
rect 310 128 318 131
rect 310 72 313 108
rect 318 82 321 128
rect 326 122 329 138
rect 334 92 337 208
rect 390 192 393 258
rect 398 238 406 241
rect 398 232 401 238
rect 398 192 401 228
rect 342 52 345 168
rect 414 152 417 158
rect 350 132 353 148
rect 350 42 353 118
rect 358 62 361 148
rect 382 142 385 148
rect 382 132 385 138
rect 414 122 417 148
rect 422 142 425 148
rect 374 92 377 98
rect 390 72 393 118
rect 422 82 425 138
rect 430 131 433 258
rect 470 241 473 258
rect 482 248 486 251
rect 494 242 497 358
rect 526 312 529 318
rect 470 238 481 241
rect 478 222 481 238
rect 446 192 449 198
rect 438 162 441 168
rect 454 142 457 158
rect 430 128 441 131
rect 398 62 401 68
rect 430 62 433 118
rect 358 -19 361 58
rect 438 -19 441 128
rect 454 61 457 138
rect 462 102 465 128
rect 470 112 473 138
rect 478 92 481 218
rect 502 212 505 258
rect 510 252 513 258
rect 518 232 521 258
rect 518 192 521 228
rect 526 202 529 258
rect 534 192 537 418
rect 542 372 545 538
rect 582 492 585 518
rect 590 482 593 508
rect 606 462 609 468
rect 566 392 569 458
rect 550 342 553 358
rect 574 352 577 428
rect 542 292 545 308
rect 582 292 585 338
rect 606 322 609 338
rect 574 272 577 278
rect 566 222 569 268
rect 598 182 601 258
rect 614 222 617 538
rect 622 512 625 538
rect 646 532 649 708
rect 654 692 657 718
rect 670 652 673 698
rect 678 692 681 738
rect 702 731 705 758
rect 710 742 713 818
rect 742 752 745 818
rect 750 742 753 748
rect 702 728 710 731
rect 694 702 697 718
rect 694 682 697 698
rect 710 682 713 728
rect 750 692 753 738
rect 758 681 761 778
rect 790 742 793 828
rect 782 732 785 738
rect 766 728 774 731
rect 766 722 769 728
rect 806 722 809 728
rect 758 678 766 681
rect 698 658 705 661
rect 702 652 705 658
rect 654 562 657 638
rect 662 542 665 618
rect 670 572 673 648
rect 710 632 713 678
rect 798 672 801 718
rect 814 672 817 748
rect 846 742 849 898
rect 854 862 857 888
rect 870 882 873 918
rect 878 872 881 918
rect 902 882 905 938
rect 926 912 929 948
rect 862 832 865 868
rect 902 862 905 868
rect 910 861 913 908
rect 926 882 929 898
rect 934 892 937 918
rect 950 912 953 948
rect 958 942 961 948
rect 966 882 969 918
rect 998 892 1001 928
rect 1038 922 1041 938
rect 1062 932 1065 938
rect 926 872 929 878
rect 910 858 918 861
rect 954 858 961 861
rect 894 752 897 818
rect 902 752 905 828
rect 910 752 913 858
rect 958 852 961 858
rect 942 742 945 778
rect 966 752 969 878
rect 974 870 985 871
rect 974 868 982 870
rect 974 852 977 868
rect 1014 862 1017 918
rect 1030 862 1033 888
rect 1038 862 1041 898
rect 1062 882 1065 928
rect 1086 922 1089 948
rect 1150 942 1153 948
rect 1174 942 1177 948
rect 1166 932 1169 938
rect 1214 932 1217 938
rect 1226 928 1230 931
rect 1070 882 1073 918
rect 1158 882 1161 928
rect 1166 882 1169 928
rect 822 732 825 740
rect 830 728 838 731
rect 926 728 934 731
rect 822 702 825 708
rect 822 682 825 698
rect 830 682 833 728
rect 926 722 929 728
rect 718 670 729 671
rect 718 668 726 670
rect 622 492 625 498
rect 638 470 641 518
rect 622 452 625 468
rect 638 451 641 466
rect 634 448 641 451
rect 646 392 649 528
rect 670 502 673 548
rect 678 542 681 628
rect 710 592 713 608
rect 678 532 681 538
rect 678 482 681 528
rect 686 402 689 538
rect 694 481 697 568
rect 718 522 721 668
rect 790 652 793 658
rect 790 618 798 621
rect 726 558 734 561
rect 726 552 729 558
rect 790 552 793 618
rect 774 541 777 548
rect 770 538 777 541
rect 798 542 801 558
rect 838 552 841 718
rect 862 662 865 678
rect 870 572 873 718
rect 914 688 918 691
rect 942 682 945 698
rect 958 692 961 718
rect 966 681 969 748
rect 986 738 990 741
rect 1014 732 1017 798
rect 958 678 969 681
rect 974 682 977 718
rect 878 672 881 678
rect 910 672 913 678
rect 938 668 942 671
rect 902 652 905 658
rect 918 642 921 648
rect 766 492 769 528
rect 766 482 769 488
rect 814 482 817 498
rect 846 492 849 540
rect 866 528 870 531
rect 694 478 705 481
rect 670 392 673 398
rect 702 392 705 478
rect 762 468 766 471
rect 806 468 814 471
rect 710 452 713 468
rect 718 441 721 468
rect 806 462 809 468
rect 794 458 798 461
rect 854 452 857 458
rect 710 438 721 441
rect 638 352 641 378
rect 622 332 625 348
rect 498 138 502 141
rect 518 132 521 158
rect 558 152 561 158
rect 566 152 569 178
rect 486 62 489 118
rect 518 92 521 128
rect 526 81 529 148
rect 542 92 545 138
rect 550 82 553 138
rect 526 78 534 81
rect 494 72 497 78
rect 502 72 505 78
rect 454 58 462 61
rect 486 12 489 58
rect 350 -22 361 -19
rect 430 -22 441 -19
rect 502 -22 505 68
rect 582 61 585 68
rect 582 58 590 61
rect 598 52 601 138
rect 606 132 609 178
rect 622 172 625 318
rect 654 282 657 318
rect 662 292 665 348
rect 690 338 694 341
rect 698 328 702 331
rect 710 292 713 438
rect 758 372 761 428
rect 758 362 761 368
rect 766 362 769 368
rect 766 358 768 362
rect 806 352 809 368
rect 814 352 817 418
rect 718 322 721 348
rect 642 268 657 271
rect 654 262 657 268
rect 662 262 665 288
rect 678 262 681 268
rect 686 252 689 258
rect 686 181 689 218
rect 694 192 697 258
rect 718 232 721 278
rect 726 272 729 338
rect 742 252 745 338
rect 754 328 758 331
rect 758 262 761 268
rect 774 262 777 348
rect 834 338 838 341
rect 790 282 793 318
rect 822 312 825 328
rect 838 282 841 328
rect 846 282 849 288
rect 862 271 865 518
rect 870 492 873 518
rect 886 482 889 618
rect 894 582 897 628
rect 926 552 929 608
rect 902 542 905 548
rect 950 542 953 678
rect 918 522 921 540
rect 958 532 961 678
rect 978 668 982 671
rect 994 668 998 671
rect 966 662 969 668
rect 910 492 913 508
rect 958 482 961 528
rect 974 521 977 588
rect 982 542 985 568
rect 994 538 998 541
rect 1006 531 1009 678
rect 1022 672 1025 858
rect 1062 832 1065 858
rect 1058 818 1065 821
rect 1054 741 1057 748
rect 1050 738 1057 741
rect 1062 742 1065 818
rect 1070 752 1073 758
rect 1046 722 1049 728
rect 1014 662 1017 668
rect 1034 658 1038 661
rect 1022 652 1025 658
rect 1042 648 1046 651
rect 1030 562 1033 568
rect 1018 538 1022 541
rect 998 528 1009 531
rect 966 518 977 521
rect 966 472 969 518
rect 982 492 985 518
rect 870 342 873 348
rect 878 342 881 458
rect 902 402 905 418
rect 926 412 929 468
rect 958 452 961 458
rect 974 432 977 468
rect 990 462 993 528
rect 998 492 1001 528
rect 886 342 889 378
rect 982 352 985 378
rect 990 362 993 438
rect 1014 432 1017 458
rect 878 332 881 338
rect 906 278 910 281
rect 858 268 865 271
rect 886 272 889 278
rect 938 268 945 271
rect 798 262 801 268
rect 830 262 833 268
rect 942 262 945 268
rect 958 270 961 348
rect 966 342 969 348
rect 990 332 993 358
rect 998 272 1001 398
rect 1006 272 1009 428
rect 1022 402 1025 458
rect 1038 362 1041 648
rect 1062 642 1065 718
rect 1070 672 1073 748
rect 1078 742 1081 768
rect 1098 758 1102 761
rect 1086 752 1089 758
rect 1078 732 1081 738
rect 1078 692 1081 698
rect 1102 692 1105 738
rect 1046 552 1049 618
rect 1046 452 1049 548
rect 1054 532 1057 638
rect 1062 592 1065 638
rect 1066 548 1070 551
rect 1086 522 1089 668
rect 1102 532 1105 648
rect 1062 502 1065 518
rect 1054 482 1057 488
rect 1078 472 1081 508
rect 1086 482 1089 498
rect 1094 482 1097 528
rect 1110 492 1113 848
rect 1130 838 1137 841
rect 1118 752 1121 758
rect 1118 722 1121 738
rect 1134 702 1137 838
rect 1166 752 1169 868
rect 1182 852 1185 908
rect 1190 892 1193 898
rect 1254 882 1257 918
rect 1218 878 1222 881
rect 1242 878 1246 881
rect 1210 868 1214 871
rect 1222 862 1225 868
rect 1234 858 1238 861
rect 1198 742 1201 748
rect 1238 742 1241 748
rect 1262 741 1265 948
rect 1270 932 1273 1058
rect 1302 972 1305 1058
rect 1310 1052 1313 1068
rect 1322 1058 1326 1061
rect 1310 952 1313 1048
rect 1342 1032 1345 1148
rect 1366 1102 1369 1148
rect 1350 1062 1353 1098
rect 1358 1062 1361 1088
rect 1390 1082 1393 1148
rect 1398 1092 1401 1148
rect 1422 1141 1425 1158
rect 1558 1152 1561 1168
rect 1638 1152 1641 1158
rect 1418 1140 1425 1141
rect 1414 1138 1425 1140
rect 1430 1122 1433 1128
rect 1414 1092 1417 1098
rect 1446 1072 1449 1138
rect 1462 1132 1465 1138
rect 1518 1132 1521 1138
rect 1486 1112 1489 1128
rect 1366 1062 1369 1068
rect 1438 1062 1441 1068
rect 1454 1062 1457 1078
rect 1486 1062 1489 1088
rect 1510 1081 1513 1118
rect 1518 1092 1521 1128
rect 1526 1082 1529 1148
rect 1582 1142 1585 1148
rect 1590 1132 1593 1148
rect 1638 1142 1641 1148
rect 1674 1138 1681 1141
rect 1622 1132 1625 1138
rect 1590 1102 1593 1128
rect 1582 1082 1585 1088
rect 1510 1078 1521 1081
rect 1518 1072 1521 1078
rect 1598 1071 1601 1118
rect 1678 1092 1681 1138
rect 1702 1102 1705 1138
rect 1710 1112 1713 1128
rect 1686 1092 1689 1098
rect 1710 1082 1713 1108
rect 1614 1072 1617 1078
rect 1718 1072 1721 1118
rect 1598 1068 1606 1071
rect 1726 1071 1729 1118
rect 1742 1082 1745 1148
rect 1834 1138 1838 1141
rect 1790 1122 1793 1128
rect 1798 1092 1801 1138
rect 1818 1128 1822 1131
rect 1766 1082 1769 1088
rect 1726 1068 1742 1071
rect 1542 1062 1545 1068
rect 1654 1062 1657 1068
rect 1782 1062 1785 1068
rect 1814 1062 1817 1128
rect 1838 1118 1846 1121
rect 1402 1058 1406 1061
rect 1278 912 1281 918
rect 1302 912 1305 948
rect 1318 932 1321 938
rect 1278 872 1281 908
rect 1326 891 1329 978
rect 1326 888 1334 891
rect 1302 881 1305 888
rect 1298 878 1305 881
rect 1326 881 1329 888
rect 1318 878 1329 881
rect 1270 772 1273 818
rect 1262 738 1273 741
rect 1158 732 1161 738
rect 1182 728 1190 731
rect 1182 722 1185 728
rect 1182 692 1185 698
rect 1142 672 1145 678
rect 1118 542 1121 568
rect 1126 542 1129 648
rect 1086 432 1089 468
rect 1014 342 1017 348
rect 1046 342 1049 348
rect 1030 312 1033 328
rect 1046 322 1049 338
rect 1078 332 1081 388
rect 1086 342 1089 428
rect 1102 352 1105 368
rect 1110 362 1113 438
rect 1118 432 1121 528
rect 1126 502 1129 528
rect 1134 512 1137 518
rect 1142 501 1145 648
rect 1150 582 1153 658
rect 1166 622 1169 678
rect 1174 642 1177 678
rect 1190 662 1193 668
rect 1198 662 1201 678
rect 1214 671 1217 718
rect 1230 682 1233 708
rect 1214 668 1222 671
rect 1238 662 1241 678
rect 1206 592 1209 618
rect 1246 592 1249 738
rect 1254 612 1257 678
rect 1270 632 1273 738
rect 1206 562 1209 568
rect 1206 552 1209 558
rect 1246 552 1249 588
rect 1254 552 1257 558
rect 1278 552 1281 868
rect 1294 742 1297 748
rect 1286 702 1289 738
rect 1286 642 1289 678
rect 1294 551 1297 698
rect 1310 681 1313 878
rect 1318 862 1321 878
rect 1326 862 1329 868
rect 1334 752 1337 818
rect 1342 762 1345 968
rect 1366 942 1369 968
rect 1390 952 1393 1018
rect 1430 992 1433 1058
rect 1478 1052 1481 1058
rect 1494 1052 1497 1058
rect 1406 932 1409 948
rect 1350 922 1353 928
rect 1390 922 1393 928
rect 1358 872 1361 888
rect 1374 870 1377 908
rect 1382 882 1385 918
rect 1390 892 1393 898
rect 1414 891 1417 978
rect 1478 962 1481 1048
rect 1510 1032 1513 1058
rect 1406 888 1417 891
rect 1406 872 1409 888
rect 1422 872 1425 918
rect 1446 892 1449 938
rect 1478 932 1481 948
rect 1486 942 1489 958
rect 1462 872 1465 918
rect 1350 852 1353 858
rect 1406 762 1409 858
rect 1486 852 1489 888
rect 1494 862 1497 928
rect 1502 922 1505 1028
rect 1510 952 1513 1018
rect 1550 992 1553 1058
rect 1638 1042 1641 1058
rect 1566 952 1569 958
rect 1638 952 1641 1038
rect 1662 962 1665 1058
rect 1670 958 1678 961
rect 1670 952 1673 958
rect 1702 952 1705 1058
rect 1602 948 1606 951
rect 1618 948 1625 951
rect 1590 942 1593 948
rect 1502 842 1505 918
rect 1550 912 1553 928
rect 1518 892 1521 898
rect 1546 868 1553 871
rect 1446 772 1449 818
rect 1342 752 1345 758
rect 1390 752 1393 758
rect 1318 732 1321 748
rect 1382 742 1385 748
rect 1342 732 1345 738
rect 1406 692 1409 698
rect 1310 678 1318 681
rect 1322 668 1329 671
rect 1326 662 1329 668
rect 1342 662 1345 678
rect 1374 622 1377 658
rect 1398 652 1401 658
rect 1414 652 1417 748
rect 1478 742 1481 818
rect 1430 722 1433 738
rect 1482 728 1489 731
rect 1486 722 1489 728
rect 1430 662 1433 718
rect 1462 692 1465 708
rect 1494 682 1497 818
rect 1518 752 1521 848
rect 1502 732 1505 748
rect 1510 692 1513 738
rect 1510 672 1513 678
rect 1498 668 1502 671
rect 1518 662 1521 748
rect 1526 722 1529 868
rect 1550 862 1553 868
rect 1546 768 1553 771
rect 1550 752 1553 768
rect 1558 752 1561 938
rect 1566 870 1569 878
rect 1582 862 1585 908
rect 1574 752 1577 848
rect 1286 548 1297 551
rect 1310 552 1313 558
rect 1150 542 1153 548
rect 1174 512 1177 548
rect 1222 532 1225 548
rect 1134 498 1145 501
rect 1134 472 1137 498
rect 1214 492 1217 498
rect 1150 481 1153 488
rect 1146 478 1153 481
rect 1206 472 1209 478
rect 1198 462 1201 468
rect 1118 352 1121 428
rect 1182 402 1185 418
rect 1198 402 1201 458
rect 1054 292 1057 318
rect 686 178 694 181
rect 622 142 625 168
rect 690 148 710 151
rect 742 142 745 208
rect 758 152 761 168
rect 790 162 793 198
rect 798 172 801 178
rect 766 152 769 158
rect 654 132 657 138
rect 662 132 665 138
rect 718 122 721 138
rect 638 92 641 98
rect 614 72 617 88
rect 670 82 673 88
rect 726 82 729 128
rect 766 82 769 108
rect 774 92 777 128
rect 782 122 785 128
rect 790 122 793 158
rect 798 112 801 148
rect 806 142 809 168
rect 830 152 833 218
rect 822 132 825 138
rect 718 72 721 78
rect 662 62 665 68
rect 766 62 769 68
rect 702 42 705 48
rect 526 -22 529 8
rect 606 -22 609 18
rect 702 -22 705 38
rect 782 32 785 68
rect 790 62 793 68
rect 822 52 825 108
rect 838 102 841 228
rect 990 222 993 258
rect 902 212 905 218
rect 886 192 889 208
rect 910 152 913 218
rect 1030 192 1033 278
rect 1086 272 1089 318
rect 1150 292 1153 318
rect 1182 291 1185 398
rect 1190 382 1193 388
rect 1190 352 1193 378
rect 1206 342 1209 468
rect 1254 462 1257 548
rect 1278 542 1281 548
rect 1286 542 1289 548
rect 1366 542 1369 548
rect 1318 532 1321 538
rect 1262 481 1265 518
rect 1278 482 1281 488
rect 1262 478 1270 481
rect 1294 472 1297 518
rect 1326 492 1329 498
rect 1334 462 1337 498
rect 1342 462 1345 538
rect 1350 532 1353 538
rect 1366 512 1369 528
rect 1366 462 1369 508
rect 1238 451 1241 458
rect 1238 448 1249 451
rect 1238 412 1241 438
rect 1246 412 1249 448
rect 1238 352 1241 408
rect 1222 342 1225 348
rect 1246 342 1249 348
rect 1302 341 1305 458
rect 1310 452 1313 458
rect 1302 338 1313 341
rect 1222 332 1225 338
rect 1230 332 1233 338
rect 1182 288 1193 291
rect 1118 281 1121 288
rect 1114 278 1121 281
rect 1054 202 1057 268
rect 1062 232 1065 268
rect 1134 262 1137 278
rect 1070 192 1073 218
rect 926 152 929 168
rect 950 142 953 158
rect 998 142 1001 188
rect 1014 142 1017 158
rect 1078 152 1081 248
rect 1086 158 1094 161
rect 1086 152 1089 158
rect 1118 142 1121 248
rect 846 112 849 118
rect 838 72 841 98
rect 846 52 849 88
rect 854 62 857 98
rect 814 -22 817 18
rect 854 -22 857 58
rect 870 42 873 138
rect 878 102 881 128
rect 894 72 897 98
rect 902 72 905 108
rect 934 92 937 138
rect 1006 122 1009 128
rect 966 82 969 88
rect 974 71 977 118
rect 1014 92 1017 138
rect 1062 122 1065 138
rect 1110 92 1113 138
rect 1126 132 1129 258
rect 1166 252 1169 268
rect 1182 262 1185 278
rect 1190 272 1193 288
rect 1262 281 1265 318
rect 1278 312 1281 338
rect 1278 292 1281 298
rect 1302 292 1305 328
rect 1310 282 1313 338
rect 1326 292 1329 318
rect 1262 278 1270 281
rect 1230 262 1233 278
rect 1302 272 1305 278
rect 1290 268 1294 271
rect 1262 262 1265 268
rect 1326 242 1329 258
rect 1334 252 1337 268
rect 1142 192 1145 198
rect 1142 152 1145 158
rect 982 71 985 78
rect 974 70 985 71
rect 974 68 982 70
rect 910 62 913 68
rect 926 62 929 68
rect 1046 68 1065 71
rect 1030 62 1033 68
rect 1046 62 1049 68
rect 1062 62 1065 68
rect 1126 70 1129 78
rect 1150 72 1153 168
rect 1198 162 1201 168
rect 1206 162 1209 218
rect 1166 72 1169 118
rect 1190 112 1193 138
rect 1198 82 1201 158
rect 1214 142 1217 168
rect 1278 142 1281 218
rect 1342 172 1345 458
rect 1350 352 1353 378
rect 1374 372 1377 618
rect 1398 602 1401 648
rect 1382 472 1385 578
rect 1438 572 1441 658
rect 1446 652 1449 658
rect 1398 552 1401 568
rect 1454 552 1457 568
rect 1462 552 1465 658
rect 1482 618 1486 621
rect 1518 552 1521 558
rect 1390 532 1393 548
rect 1438 542 1441 548
rect 1446 532 1449 548
rect 1494 542 1497 548
rect 1526 542 1529 718
rect 1542 712 1545 738
rect 1542 662 1545 668
rect 1538 618 1542 621
rect 1542 542 1545 608
rect 1550 552 1553 748
rect 1574 742 1577 748
rect 1582 742 1585 748
rect 1590 732 1593 858
rect 1606 772 1609 948
rect 1622 762 1625 948
rect 1734 942 1737 1018
rect 1750 992 1753 1058
rect 1774 992 1777 1058
rect 1782 1042 1785 1058
rect 1814 972 1817 1058
rect 1822 1042 1825 1098
rect 1838 1072 1841 1118
rect 1638 862 1641 878
rect 1654 862 1657 918
rect 1662 872 1665 878
rect 1678 852 1681 858
rect 1702 792 1705 938
rect 1746 928 1761 931
rect 1742 872 1745 918
rect 1758 892 1761 928
rect 1790 892 1793 928
rect 1798 882 1801 968
rect 1814 941 1817 948
rect 1810 938 1817 941
rect 1822 922 1825 1038
rect 1830 952 1833 1038
rect 1838 952 1841 1048
rect 1854 1012 1857 1128
rect 1830 882 1833 948
rect 1710 851 1713 858
rect 1710 848 1718 851
rect 1654 752 1657 758
rect 1622 742 1625 748
rect 1662 742 1665 768
rect 1634 728 1641 731
rect 1558 662 1561 728
rect 1638 722 1641 728
rect 1686 722 1689 748
rect 1742 742 1745 868
rect 1750 842 1753 878
rect 1818 868 1822 871
rect 1774 831 1777 858
rect 1766 828 1777 831
rect 1694 732 1697 738
rect 1566 672 1569 718
rect 1590 682 1593 718
rect 1718 702 1721 738
rect 1726 722 1729 728
rect 1606 681 1609 688
rect 1742 682 1745 738
rect 1766 722 1769 828
rect 1782 772 1785 868
rect 1830 862 1833 878
rect 1838 872 1841 948
rect 1846 922 1849 928
rect 1854 892 1857 998
rect 1862 982 1865 1018
rect 1862 922 1865 948
rect 1846 862 1849 878
rect 1870 862 1873 938
rect 1798 738 1806 741
rect 1758 691 1761 718
rect 1750 688 1761 691
rect 1602 678 1609 681
rect 1662 672 1665 678
rect 1486 532 1489 538
rect 1526 532 1529 538
rect 1390 522 1393 528
rect 1502 512 1505 518
rect 1406 462 1409 468
rect 1438 462 1441 478
rect 1462 472 1465 508
rect 1510 482 1513 488
rect 1382 352 1385 438
rect 1390 382 1393 458
rect 1502 452 1505 468
rect 1414 392 1417 408
rect 1350 312 1353 348
rect 1358 262 1361 318
rect 1382 222 1385 348
rect 1390 332 1393 368
rect 1398 322 1401 338
rect 1398 282 1401 308
rect 1430 292 1433 358
rect 1462 352 1465 448
rect 1502 392 1505 398
rect 1446 332 1449 348
rect 1526 342 1529 358
rect 1534 342 1537 528
rect 1542 472 1545 508
rect 1550 462 1553 548
rect 1558 492 1561 658
rect 1566 642 1569 658
rect 1598 552 1601 628
rect 1622 591 1625 658
rect 1618 588 1625 591
rect 1622 562 1625 588
rect 1630 632 1633 668
rect 1630 582 1633 628
rect 1670 592 1673 678
rect 1694 662 1697 678
rect 1750 672 1753 688
rect 1766 672 1769 698
rect 1774 670 1777 718
rect 1798 692 1801 738
rect 1822 732 1825 738
rect 1854 732 1857 738
rect 1814 722 1817 728
rect 1790 682 1793 688
rect 1822 672 1825 728
rect 1850 718 1854 721
rect 1830 692 1833 718
rect 1686 592 1689 608
rect 1718 592 1721 668
rect 1846 670 1849 708
rect 1870 682 1873 858
rect 1814 632 1817 658
rect 1814 601 1817 628
rect 1806 598 1817 601
rect 1574 532 1577 540
rect 1590 502 1593 518
rect 1598 491 1601 548
rect 1622 542 1625 548
rect 1654 542 1657 548
rect 1590 488 1601 491
rect 1566 482 1569 488
rect 1462 322 1465 328
rect 1390 272 1393 278
rect 1446 270 1449 318
rect 1486 312 1489 318
rect 1478 272 1481 288
rect 1486 282 1489 298
rect 1494 282 1497 338
rect 1530 328 1537 331
rect 1534 322 1537 328
rect 1510 282 1513 288
rect 1526 282 1529 288
rect 1510 272 1513 278
rect 1390 192 1393 268
rect 1318 152 1321 158
rect 1390 152 1393 158
rect 1254 112 1257 138
rect 1262 122 1265 140
rect 1294 112 1297 148
rect 1326 142 1329 148
rect 1342 142 1345 148
rect 1318 132 1321 138
rect 1154 58 1158 61
rect 950 52 953 58
rect 878 -22 881 38
rect 1054 12 1057 58
rect 1166 51 1169 58
rect 1146 48 1169 51
rect 966 -22 969 8
rect 1078 -22 1081 18
rect 1190 -22 1193 68
rect 1198 12 1201 78
rect 1206 52 1209 88
rect 1238 72 1241 108
rect 1230 62 1233 68
rect 1278 62 1281 108
rect 1382 92 1385 138
rect 1326 62 1329 78
rect 1358 72 1361 78
rect 1398 71 1401 228
rect 1422 222 1425 258
rect 1446 222 1449 266
rect 1414 152 1417 208
rect 1446 182 1449 218
rect 1462 152 1465 218
rect 1478 202 1481 268
rect 1406 142 1409 148
rect 1430 141 1433 148
rect 1426 140 1433 141
rect 1422 138 1433 140
rect 1438 112 1441 118
rect 1438 82 1441 88
rect 1454 72 1457 108
rect 1478 92 1481 128
rect 1486 72 1489 148
rect 1518 142 1521 258
rect 1534 182 1537 308
rect 1550 292 1553 348
rect 1558 342 1561 348
rect 1550 272 1553 278
rect 1566 262 1569 368
rect 1574 302 1577 418
rect 1582 352 1585 368
rect 1590 351 1593 488
rect 1606 481 1609 518
rect 1646 512 1649 518
rect 1602 478 1609 481
rect 1630 472 1633 488
rect 1686 472 1689 558
rect 1734 552 1737 558
rect 1806 552 1809 598
rect 1822 591 1825 668
rect 1814 588 1825 591
rect 1602 468 1609 471
rect 1606 462 1609 468
rect 1638 462 1641 468
rect 1622 352 1625 458
rect 1662 352 1665 388
rect 1590 348 1598 351
rect 1590 322 1593 338
rect 1606 322 1609 348
rect 1622 322 1625 328
rect 1606 272 1609 318
rect 1614 282 1617 318
rect 1622 312 1625 318
rect 1646 292 1649 328
rect 1678 271 1681 318
rect 1674 268 1681 271
rect 1694 272 1697 548
rect 1714 528 1721 531
rect 1718 522 1721 528
rect 1702 462 1705 478
rect 1734 472 1737 548
rect 1758 512 1761 548
rect 1814 492 1817 588
rect 1822 572 1825 578
rect 1830 552 1833 558
rect 1862 552 1865 558
rect 1870 552 1873 668
rect 1754 478 1758 481
rect 1718 462 1721 468
rect 1702 392 1705 458
rect 1726 352 1729 468
rect 1766 352 1769 468
rect 1830 452 1833 548
rect 1878 542 1881 718
rect 1838 462 1841 498
rect 1878 492 1881 528
rect 1846 451 1849 468
rect 1838 448 1849 451
rect 1714 338 1718 341
rect 1702 321 1705 338
rect 1742 322 1745 328
rect 1702 318 1713 321
rect 1710 292 1713 318
rect 1726 272 1729 288
rect 1742 282 1745 318
rect 1750 282 1753 338
rect 1798 322 1801 338
rect 1758 272 1761 298
rect 1798 292 1801 308
rect 1542 242 1545 258
rect 1558 252 1561 258
rect 1574 222 1577 238
rect 1534 161 1537 178
rect 1526 158 1537 161
rect 1526 152 1529 158
rect 1534 132 1537 148
rect 1510 92 1513 118
rect 1534 102 1537 128
rect 1398 68 1406 71
rect 1466 68 1470 71
rect 1214 32 1217 58
rect 1214 -22 1217 8
rect 1230 -22 1233 38
rect 1254 12 1257 28
rect 1326 12 1329 58
rect 1334 52 1337 68
rect 1342 52 1345 68
rect 1350 62 1353 68
rect 1366 62 1369 68
rect 1334 42 1337 48
rect 1254 -22 1257 8
rect 1430 -22 1433 68
rect 1486 62 1489 68
rect 1502 62 1505 78
rect 1510 42 1513 68
rect 1526 62 1529 68
rect 1558 62 1561 148
rect 1590 142 1593 198
rect 1590 82 1593 138
rect 1598 132 1601 198
rect 1606 162 1609 268
rect 1630 152 1633 208
rect 1646 152 1649 218
rect 1670 152 1673 178
rect 1606 142 1609 148
rect 1622 132 1625 148
rect 1646 132 1649 148
rect 1670 102 1673 148
rect 1566 61 1569 68
rect 1646 62 1649 98
rect 1654 62 1657 68
rect 1678 62 1681 148
rect 1694 72 1697 258
rect 1710 142 1713 268
rect 1742 202 1745 218
rect 1750 192 1753 268
rect 1718 132 1721 138
rect 1726 121 1729 138
rect 1718 118 1729 121
rect 1718 92 1721 118
rect 1734 62 1737 128
rect 1742 92 1745 158
rect 1758 142 1761 268
rect 1766 262 1769 268
rect 1806 262 1809 318
rect 1814 312 1817 338
rect 1766 192 1769 258
rect 1822 162 1825 418
rect 1830 392 1833 398
rect 1838 382 1841 448
rect 1830 378 1838 381
rect 1830 302 1833 378
rect 1854 372 1857 478
rect 1838 292 1841 368
rect 1878 352 1881 418
rect 1830 262 1833 268
rect 1766 158 1774 161
rect 1766 152 1769 158
rect 1814 152 1817 158
rect 1846 152 1849 168
rect 1750 82 1753 118
rect 1758 62 1761 78
rect 1766 62 1769 98
rect 1782 82 1785 148
rect 1798 92 1801 138
rect 1806 122 1809 128
rect 1854 82 1857 158
rect 1782 70 1785 78
rect 1846 72 1849 78
rect 1878 62 1881 348
rect 1886 322 1889 1118
rect 1886 262 1889 268
rect 1566 58 1574 61
rect 1594 48 1598 51
rect 1510 -22 1513 38
rect 1590 -22 1593 18
rect 1678 -22 1681 58
rect 1734 -22 1737 58
<< m3contact >>
rect 558 1178 562 1182
rect 350 1168 354 1172
rect 6 1158 10 1162
rect 334 1158 338 1162
rect 78 1128 82 1132
rect 206 1148 210 1152
rect 230 1148 234 1152
rect 270 1148 274 1152
rect 286 1148 290 1152
rect 46 1088 50 1092
rect 6 1078 10 1082
rect 46 1078 50 1082
rect 134 1118 138 1122
rect 86 1088 90 1092
rect 214 1138 218 1142
rect 270 1138 274 1142
rect 150 1128 154 1132
rect 174 1118 178 1122
rect 222 1118 226 1122
rect 246 1118 250 1122
rect 198 1108 202 1112
rect 230 1098 234 1102
rect 174 1068 178 1072
rect 206 1068 210 1072
rect 22 1058 26 1062
rect 38 1058 42 1062
rect 54 1038 58 1042
rect 14 1028 18 1032
rect 6 958 10 962
rect 6 878 10 882
rect 6 778 10 782
rect 6 658 10 662
rect 62 1028 66 1032
rect 46 1018 50 1022
rect 62 1018 66 1022
rect 62 918 66 922
rect 70 918 74 922
rect 62 888 66 892
rect 94 1058 98 1062
rect 158 1058 162 1062
rect 182 1058 186 1062
rect 118 1048 122 1052
rect 174 1048 178 1052
rect 142 1028 146 1032
rect 110 1018 114 1022
rect 134 998 138 1002
rect 166 1018 170 1022
rect 174 1008 178 1012
rect 182 958 186 962
rect 174 948 178 952
rect 190 948 194 952
rect 102 938 106 942
rect 102 928 106 932
rect 102 918 106 922
rect 126 918 130 922
rect 78 908 82 912
rect 78 888 82 892
rect 94 908 98 912
rect 86 878 90 882
rect 102 858 106 862
rect 158 928 162 932
rect 166 878 170 882
rect 158 868 162 872
rect 174 788 178 792
rect 62 728 66 732
rect 86 728 90 732
rect 78 668 82 672
rect 38 618 42 622
rect 78 598 82 602
rect 6 558 10 562
rect 46 558 50 562
rect 70 558 74 562
rect 62 548 66 552
rect 110 678 114 682
rect 166 738 170 742
rect 206 938 210 942
rect 190 928 194 932
rect 190 868 194 872
rect 246 1078 250 1082
rect 270 1098 274 1102
rect 262 1078 266 1082
rect 278 1070 282 1072
rect 278 1068 282 1070
rect 254 1058 258 1062
rect 222 1048 226 1052
rect 238 968 242 972
rect 230 888 234 892
rect 222 878 226 882
rect 214 858 218 862
rect 230 858 234 862
rect 190 758 194 762
rect 190 748 194 752
rect 294 1118 298 1122
rect 390 1148 394 1152
rect 414 1148 418 1152
rect 422 1148 426 1152
rect 438 1148 442 1152
rect 558 1148 562 1152
rect 382 1118 386 1122
rect 622 1208 626 1212
rect 614 1178 618 1182
rect 862 1208 866 1212
rect 878 1208 882 1212
rect 846 1168 850 1172
rect 950 1178 954 1182
rect 886 1158 890 1162
rect 934 1158 938 1162
rect 678 1148 682 1152
rect 702 1148 706 1152
rect 854 1148 858 1152
rect 878 1148 882 1152
rect 926 1148 930 1152
rect 942 1148 946 1152
rect 310 1108 314 1112
rect 350 1108 354 1112
rect 382 1108 386 1112
rect 398 1108 402 1112
rect 334 1088 338 1092
rect 342 1088 346 1092
rect 334 1078 338 1082
rect 310 1068 314 1072
rect 446 1118 450 1122
rect 430 1108 434 1112
rect 478 1138 482 1142
rect 582 1138 586 1142
rect 486 1128 490 1132
rect 534 1128 538 1132
rect 566 1128 570 1132
rect 670 1138 674 1142
rect 694 1138 698 1142
rect 750 1138 754 1142
rect 590 1128 594 1132
rect 606 1128 610 1132
rect 758 1128 762 1132
rect 494 1118 498 1122
rect 542 1118 546 1122
rect 574 1118 578 1122
rect 470 1108 474 1112
rect 414 1098 418 1102
rect 454 1098 458 1102
rect 478 1098 482 1102
rect 406 1088 410 1092
rect 350 1068 354 1072
rect 358 1068 362 1072
rect 398 1068 402 1072
rect 286 1038 290 1042
rect 374 1038 378 1042
rect 286 1028 290 1032
rect 262 1018 266 1022
rect 278 1018 282 1022
rect 262 1008 266 1012
rect 254 958 258 962
rect 246 948 250 952
rect 254 928 258 932
rect 270 948 274 952
rect 318 958 322 962
rect 350 958 354 962
rect 294 948 298 952
rect 318 948 322 952
rect 390 948 394 952
rect 350 938 354 942
rect 294 918 298 922
rect 262 888 266 892
rect 262 878 266 882
rect 350 928 354 932
rect 382 938 386 942
rect 358 918 362 922
rect 334 908 338 912
rect 366 908 370 912
rect 254 868 258 872
rect 310 868 314 872
rect 342 870 346 872
rect 342 868 346 870
rect 310 858 314 862
rect 214 748 218 752
rect 238 788 242 792
rect 222 738 226 742
rect 350 818 354 822
rect 270 788 274 792
rect 334 788 338 792
rect 350 778 354 782
rect 254 748 258 752
rect 270 748 274 752
rect 318 748 322 752
rect 414 1018 418 1022
rect 470 1058 474 1062
rect 486 1048 490 1052
rect 454 1038 458 1042
rect 462 1038 466 1042
rect 486 1038 490 1042
rect 446 1008 450 1012
rect 478 978 482 982
rect 462 958 466 962
rect 446 948 450 952
rect 430 918 434 922
rect 406 898 410 902
rect 406 878 410 882
rect 422 898 426 902
rect 430 898 434 902
rect 438 888 442 892
rect 414 858 418 862
rect 398 838 402 842
rect 414 838 418 842
rect 358 768 362 772
rect 374 768 378 772
rect 262 738 266 742
rect 366 738 370 742
rect 166 728 170 732
rect 198 728 202 732
rect 206 728 210 732
rect 230 728 234 732
rect 246 728 250 732
rect 158 708 162 712
rect 142 668 146 672
rect 166 688 170 692
rect 470 888 474 892
rect 446 878 450 882
rect 470 878 474 882
rect 510 1098 514 1102
rect 550 1098 554 1102
rect 566 1098 570 1102
rect 502 1028 506 1032
rect 558 1088 562 1092
rect 582 1108 586 1112
rect 526 1048 530 1052
rect 582 998 586 1002
rect 534 978 538 982
rect 494 958 498 962
rect 502 948 506 952
rect 542 948 546 952
rect 558 948 562 952
rect 534 938 538 942
rect 566 928 570 932
rect 494 918 498 922
rect 518 918 522 922
rect 526 918 530 922
rect 574 918 578 922
rect 582 898 586 902
rect 534 888 538 892
rect 582 888 586 892
rect 470 858 474 862
rect 542 868 546 872
rect 566 868 570 872
rect 630 1118 634 1122
rect 622 1108 626 1112
rect 774 1118 778 1122
rect 662 1098 666 1102
rect 670 1098 674 1102
rect 766 1098 770 1102
rect 630 1088 634 1092
rect 766 1088 770 1092
rect 606 1058 610 1062
rect 646 1058 650 1062
rect 678 1058 682 1062
rect 686 1058 690 1062
rect 598 988 602 992
rect 742 1048 746 1052
rect 654 1038 658 1042
rect 718 1038 722 1042
rect 646 988 650 992
rect 622 968 626 972
rect 638 948 642 952
rect 670 948 674 952
rect 702 948 706 952
rect 606 938 610 942
rect 614 918 618 922
rect 630 918 634 922
rect 622 878 626 882
rect 590 868 594 872
rect 614 868 618 872
rect 502 838 506 842
rect 622 838 626 842
rect 438 828 442 832
rect 454 828 458 832
rect 510 828 514 832
rect 598 828 602 832
rect 422 808 426 812
rect 382 748 386 752
rect 430 748 434 752
rect 198 688 202 692
rect 294 688 298 692
rect 206 678 210 682
rect 230 678 234 682
rect 270 678 274 682
rect 390 678 394 682
rect 406 678 410 682
rect 166 668 170 672
rect 190 668 194 672
rect 198 668 202 672
rect 238 668 242 672
rect 358 668 362 672
rect 422 678 426 682
rect 102 658 106 662
rect 126 658 130 662
rect 118 628 122 632
rect 222 658 226 662
rect 246 658 250 662
rect 302 658 306 662
rect 350 658 354 662
rect 390 658 394 662
rect 430 658 434 662
rect 262 648 266 652
rect 286 648 290 652
rect 334 648 338 652
rect 310 618 314 622
rect 246 608 250 612
rect 110 578 114 582
rect 102 558 106 562
rect 94 538 98 542
rect 30 478 34 482
rect 62 478 66 482
rect 30 468 34 472
rect 70 468 74 472
rect 214 558 218 562
rect 118 548 122 552
rect 134 548 138 552
rect 150 548 154 552
rect 166 548 170 552
rect 182 548 186 552
rect 206 548 210 552
rect 222 538 226 542
rect 94 478 98 482
rect 6 458 10 462
rect 22 458 26 462
rect 46 438 50 442
rect 62 438 66 442
rect 6 338 10 342
rect 54 338 58 342
rect 118 458 122 462
rect 110 408 114 412
rect 102 368 106 372
rect 78 358 82 362
rect 94 338 98 342
rect 30 318 34 322
rect 54 318 58 322
rect 6 258 10 262
rect 70 288 74 292
rect 374 568 378 572
rect 366 558 370 562
rect 270 540 274 542
rect 270 538 274 540
rect 366 548 370 552
rect 382 548 386 552
rect 214 528 218 532
rect 238 528 242 532
rect 278 528 282 532
rect 302 528 306 532
rect 342 528 346 532
rect 366 528 370 532
rect 366 518 370 522
rect 150 478 154 482
rect 174 478 178 482
rect 222 478 226 482
rect 238 478 242 482
rect 254 478 258 482
rect 310 478 314 482
rect 342 478 346 482
rect 214 468 218 472
rect 174 448 178 452
rect 150 408 154 412
rect 126 358 130 362
rect 142 348 146 352
rect 110 338 114 342
rect 102 278 106 282
rect 198 458 202 462
rect 190 448 194 452
rect 182 368 186 372
rect 158 348 162 352
rect 134 318 138 322
rect 126 288 130 292
rect 46 258 50 262
rect 86 258 90 262
rect 110 258 114 262
rect 70 228 74 232
rect 102 168 106 172
rect 54 158 58 162
rect 62 158 66 162
rect 78 148 82 152
rect 6 138 10 142
rect 54 138 58 142
rect 70 128 74 132
rect 46 118 50 122
rect 62 118 66 122
rect 30 108 34 112
rect 6 88 10 92
rect 6 58 10 62
rect 54 108 58 112
rect 70 108 74 112
rect 62 68 66 72
rect 94 138 98 142
rect 86 88 90 92
rect 110 128 114 132
rect 94 78 98 82
rect 102 78 106 82
rect 182 298 186 302
rect 150 288 154 292
rect 222 418 226 422
rect 254 468 258 472
rect 262 468 266 472
rect 286 468 290 472
rect 310 468 314 472
rect 318 458 322 462
rect 334 458 338 462
rect 342 408 346 412
rect 342 388 346 392
rect 246 338 250 342
rect 278 338 282 342
rect 310 338 314 342
rect 326 338 330 342
rect 222 288 226 292
rect 166 278 170 282
rect 198 278 202 282
rect 214 278 218 282
rect 190 268 194 272
rect 166 258 170 262
rect 214 258 218 262
rect 158 248 162 252
rect 198 248 202 252
rect 182 228 186 232
rect 142 188 146 192
rect 174 188 178 192
rect 238 258 242 262
rect 262 288 266 292
rect 254 268 258 272
rect 230 238 234 242
rect 374 508 378 512
rect 430 648 434 652
rect 494 808 498 812
rect 454 758 458 762
rect 446 748 450 752
rect 510 748 514 752
rect 470 738 474 742
rect 486 738 490 742
rect 462 708 466 712
rect 454 678 458 682
rect 462 678 466 682
rect 454 658 458 662
rect 438 628 442 632
rect 398 558 402 562
rect 406 528 410 532
rect 406 428 410 432
rect 414 418 418 422
rect 454 548 458 552
rect 526 738 530 742
rect 550 738 554 742
rect 526 728 530 732
rect 550 688 554 692
rect 518 678 522 682
rect 574 758 578 762
rect 590 738 594 742
rect 582 678 586 682
rect 614 728 618 732
rect 662 938 666 942
rect 678 938 682 942
rect 718 940 722 942
rect 718 938 722 940
rect 646 928 650 932
rect 678 928 682 932
rect 726 928 730 932
rect 638 898 642 902
rect 654 868 658 872
rect 646 778 650 782
rect 750 1038 754 1042
rect 750 988 754 992
rect 750 928 754 932
rect 694 878 698 882
rect 726 878 730 882
rect 734 878 738 882
rect 710 868 714 872
rect 846 1138 850 1142
rect 806 1108 810 1112
rect 814 1108 818 1112
rect 814 1088 818 1092
rect 798 1068 802 1072
rect 790 998 794 1002
rect 798 998 802 1002
rect 766 938 770 942
rect 782 938 786 942
rect 758 908 762 912
rect 790 908 794 912
rect 758 888 762 892
rect 670 858 674 862
rect 686 858 690 862
rect 742 858 746 862
rect 702 848 706 852
rect 774 878 778 882
rect 750 838 754 842
rect 814 1058 818 1062
rect 814 998 818 1002
rect 846 1068 850 1072
rect 838 1058 842 1062
rect 830 1028 834 1032
rect 894 1138 898 1142
rect 910 1088 914 1092
rect 870 1078 874 1082
rect 934 1078 938 1082
rect 950 1078 954 1082
rect 966 1148 970 1152
rect 982 1148 986 1152
rect 1022 1158 1026 1162
rect 1118 1178 1122 1182
rect 1126 1168 1130 1172
rect 1142 1168 1146 1172
rect 1558 1168 1562 1172
rect 1422 1158 1426 1162
rect 1438 1158 1442 1162
rect 1038 1148 1042 1152
rect 1118 1148 1122 1152
rect 1214 1148 1218 1152
rect 1262 1148 1266 1152
rect 1366 1148 1370 1152
rect 1374 1148 1378 1152
rect 1406 1148 1410 1152
rect 990 1138 994 1142
rect 998 1138 1002 1142
rect 1006 1138 1010 1142
rect 974 1128 978 1132
rect 990 1108 994 1112
rect 1014 1108 1018 1112
rect 966 1068 970 1072
rect 974 1068 978 1072
rect 998 1098 1002 1102
rect 1006 1088 1010 1092
rect 870 1058 874 1062
rect 926 1058 930 1062
rect 886 1038 890 1042
rect 862 1028 866 1032
rect 902 1028 906 1032
rect 846 1008 850 1012
rect 894 1008 898 1012
rect 910 1008 914 1012
rect 862 958 866 962
rect 902 958 906 962
rect 822 938 826 942
rect 846 938 850 942
rect 958 1048 962 1052
rect 982 1018 986 1022
rect 1054 1078 1058 1082
rect 1086 1138 1090 1142
rect 1102 1118 1106 1122
rect 1078 1098 1082 1102
rect 1078 1078 1082 1082
rect 1062 1068 1066 1072
rect 1038 1058 1042 1062
rect 1054 1058 1058 1062
rect 1046 1038 1050 1042
rect 1038 1018 1042 1022
rect 1158 1128 1162 1132
rect 1174 1078 1178 1082
rect 1126 1068 1130 1072
rect 1142 1068 1146 1072
rect 1150 1068 1154 1072
rect 1166 1068 1170 1072
rect 1118 1058 1122 1062
rect 1134 1058 1138 1062
rect 1086 1048 1090 1052
rect 1150 1048 1154 1052
rect 1062 1038 1066 1042
rect 1110 1038 1114 1042
rect 1086 1008 1090 1012
rect 998 988 1002 992
rect 1102 978 1106 982
rect 998 958 1002 962
rect 1022 958 1026 962
rect 1118 958 1122 962
rect 934 948 938 952
rect 974 948 978 952
rect 1070 948 1074 952
rect 1150 948 1154 952
rect 1198 1068 1202 1072
rect 1190 1038 1194 1042
rect 1182 978 1186 982
rect 1230 1138 1234 1142
rect 1238 1108 1242 1112
rect 1254 1108 1258 1112
rect 1254 1098 1258 1102
rect 1222 1068 1226 1072
rect 1294 1138 1298 1142
rect 1318 1138 1322 1142
rect 1318 1128 1322 1132
rect 1278 1118 1282 1122
rect 1270 1098 1274 1102
rect 1262 1088 1266 1092
rect 1262 1068 1266 1072
rect 1334 1108 1338 1112
rect 1302 1068 1306 1072
rect 1310 1068 1314 1072
rect 1270 1058 1274 1062
rect 1262 1028 1266 1032
rect 1262 998 1266 1002
rect 1214 988 1218 992
rect 1238 988 1242 992
rect 1198 958 1202 962
rect 1206 958 1210 962
rect 1230 958 1234 962
rect 1206 948 1210 952
rect 838 908 842 912
rect 854 908 858 912
rect 846 898 850 902
rect 830 868 834 872
rect 822 858 826 862
rect 838 858 842 862
rect 790 828 794 832
rect 806 828 810 832
rect 686 808 690 812
rect 662 738 666 742
rect 686 738 690 742
rect 630 728 634 732
rect 638 728 642 732
rect 646 708 650 712
rect 614 678 618 682
rect 518 668 522 672
rect 558 668 562 672
rect 574 668 578 672
rect 494 658 498 662
rect 622 658 626 662
rect 542 648 546 652
rect 542 618 546 622
rect 494 588 498 592
rect 486 578 490 582
rect 478 568 482 572
rect 510 578 514 582
rect 518 548 522 552
rect 558 588 562 592
rect 606 578 610 582
rect 590 558 594 562
rect 558 548 562 552
rect 574 548 578 552
rect 638 648 642 652
rect 638 558 642 562
rect 502 538 506 542
rect 462 528 466 532
rect 446 518 450 522
rect 462 488 466 492
rect 438 468 442 472
rect 470 468 474 472
rect 406 408 410 412
rect 422 408 426 412
rect 382 378 386 382
rect 358 368 362 372
rect 382 368 386 372
rect 390 368 394 372
rect 374 338 378 342
rect 350 328 354 332
rect 366 328 370 332
rect 390 308 394 312
rect 414 378 418 382
rect 454 438 458 442
rect 438 368 442 372
rect 446 358 450 362
rect 422 348 426 352
rect 438 348 442 352
rect 526 518 530 522
rect 526 488 530 492
rect 502 468 506 472
rect 486 458 490 462
rect 502 458 506 462
rect 534 458 538 462
rect 518 448 522 452
rect 502 438 506 442
rect 502 408 506 412
rect 534 418 538 422
rect 518 388 522 392
rect 510 378 514 382
rect 510 368 514 372
rect 462 348 466 352
rect 342 278 346 282
rect 358 278 362 282
rect 270 268 274 272
rect 286 268 290 272
rect 302 268 306 272
rect 334 268 338 272
rect 406 268 410 272
rect 262 258 266 262
rect 230 168 234 172
rect 150 148 154 152
rect 134 128 138 132
rect 158 128 162 132
rect 166 128 170 132
rect 190 138 194 142
rect 174 118 178 122
rect 182 118 186 122
rect 142 98 146 102
rect 182 98 186 102
rect 198 98 202 102
rect 198 88 202 92
rect 222 158 226 162
rect 390 258 394 262
rect 414 258 418 262
rect 430 318 434 322
rect 446 308 450 312
rect 462 258 466 262
rect 358 248 362 252
rect 382 228 386 232
rect 310 218 314 222
rect 342 218 346 222
rect 334 208 338 212
rect 278 158 282 162
rect 286 138 290 142
rect 302 138 306 142
rect 246 128 250 132
rect 254 128 258 132
rect 246 108 250 112
rect 278 118 282 122
rect 246 98 250 102
rect 262 98 266 102
rect 190 68 194 72
rect 78 58 82 62
rect 150 58 154 62
rect 174 58 178 62
rect 214 78 218 82
rect 270 68 274 72
rect 118 48 122 52
rect 318 148 322 152
rect 310 108 314 112
rect 326 118 330 122
rect 398 228 402 232
rect 374 188 378 192
rect 342 168 346 172
rect 318 78 322 82
rect 318 58 322 62
rect 414 158 418 162
rect 350 148 354 152
rect 358 148 362 152
rect 382 148 386 152
rect 422 148 426 152
rect 350 118 354 122
rect 342 48 346 52
rect 382 138 386 142
rect 414 118 418 122
rect 374 98 378 102
rect 438 248 442 252
rect 462 248 466 252
rect 486 248 490 252
rect 502 348 506 352
rect 526 308 530 312
rect 494 238 498 242
rect 478 218 482 222
rect 446 198 450 202
rect 438 158 442 162
rect 446 148 450 152
rect 454 138 458 142
rect 430 118 434 122
rect 406 78 410 82
rect 422 78 426 82
rect 390 70 394 72
rect 390 68 394 70
rect 398 58 402 62
rect 366 48 370 52
rect 398 48 402 52
rect 446 58 450 62
rect 470 108 474 112
rect 462 98 466 102
rect 510 248 514 252
rect 518 228 522 232
rect 502 208 506 212
rect 526 198 530 202
rect 550 528 554 532
rect 582 518 586 522
rect 590 508 594 512
rect 558 468 562 472
rect 598 468 602 472
rect 606 458 610 462
rect 550 418 554 422
rect 574 428 578 432
rect 566 388 570 392
rect 542 368 546 372
rect 542 340 546 342
rect 542 338 546 340
rect 590 388 594 392
rect 542 308 546 312
rect 606 318 610 322
rect 574 268 578 272
rect 550 248 554 252
rect 566 218 570 222
rect 518 188 522 192
rect 670 698 674 702
rect 654 688 658 692
rect 662 658 666 662
rect 758 778 762 782
rect 750 738 754 742
rect 694 698 698 702
rect 734 718 738 722
rect 750 688 754 692
rect 694 678 698 682
rect 710 678 714 682
rect 814 748 818 752
rect 830 748 834 752
rect 790 738 794 742
rect 782 728 786 732
rect 806 728 810 732
rect 774 688 778 692
rect 702 668 706 672
rect 654 558 658 562
rect 854 888 858 892
rect 910 908 914 912
rect 926 908 930 912
rect 902 878 906 882
rect 902 868 906 872
rect 926 898 930 902
rect 958 938 962 942
rect 990 938 994 942
rect 1062 938 1066 942
rect 998 928 1002 932
rect 966 918 970 922
rect 950 908 954 912
rect 934 888 938 892
rect 1046 928 1050 932
rect 1038 918 1042 922
rect 926 878 930 882
rect 966 878 970 882
rect 958 868 962 872
rect 934 858 938 862
rect 862 828 866 832
rect 902 828 906 832
rect 942 778 946 782
rect 894 748 898 752
rect 910 748 914 752
rect 990 868 994 872
rect 1038 898 1042 902
rect 1030 888 1034 892
rect 1094 938 1098 942
rect 1166 938 1170 942
rect 1158 928 1162 932
rect 1190 928 1194 932
rect 1214 928 1218 932
rect 1230 928 1234 932
rect 1086 918 1090 922
rect 1182 908 1186 912
rect 1062 878 1066 882
rect 1070 878 1074 882
rect 1102 878 1106 882
rect 1158 878 1162 882
rect 1078 868 1082 872
rect 1094 868 1098 872
rect 1158 868 1162 872
rect 1126 858 1130 862
rect 1142 858 1146 862
rect 974 848 978 852
rect 1014 798 1018 802
rect 862 738 866 742
rect 886 740 890 742
rect 886 738 890 740
rect 894 738 898 742
rect 822 728 826 732
rect 822 708 826 712
rect 822 698 826 702
rect 838 718 842 722
rect 830 678 834 682
rect 678 628 682 632
rect 710 628 714 632
rect 670 568 674 572
rect 654 528 658 532
rect 622 508 626 512
rect 622 498 626 502
rect 622 448 626 452
rect 710 608 714 612
rect 694 568 698 572
rect 678 538 682 542
rect 670 498 674 502
rect 678 478 682 482
rect 670 458 674 462
rect 678 458 682 462
rect 702 548 706 552
rect 758 668 762 672
rect 798 668 802 672
rect 830 668 834 672
rect 790 658 794 662
rect 790 648 794 652
rect 734 538 738 542
rect 862 678 866 682
rect 854 648 858 652
rect 942 698 946 702
rect 910 688 914 692
rect 958 688 962 692
rect 910 678 914 682
rect 942 678 946 682
rect 950 678 954 682
rect 990 738 994 742
rect 982 728 986 732
rect 878 668 882 672
rect 934 668 938 672
rect 878 658 882 662
rect 902 648 906 652
rect 918 638 922 642
rect 894 628 898 632
rect 870 568 874 572
rect 822 548 826 552
rect 830 548 834 552
rect 718 518 722 522
rect 814 498 818 502
rect 766 488 770 492
rect 878 538 882 542
rect 862 528 866 532
rect 870 518 874 522
rect 846 488 850 492
rect 750 478 754 482
rect 766 478 770 482
rect 694 468 698 472
rect 670 398 674 402
rect 686 398 690 402
rect 710 468 714 472
rect 766 468 770 472
rect 726 458 730 462
rect 798 458 802 462
rect 742 448 746 452
rect 854 448 858 452
rect 638 378 642 382
rect 622 348 626 352
rect 622 318 626 322
rect 654 318 658 322
rect 614 218 618 222
rect 566 178 570 182
rect 598 178 602 182
rect 606 178 610 182
rect 518 158 522 162
rect 558 158 562 162
rect 486 148 490 152
rect 502 148 506 152
rect 502 138 506 142
rect 526 148 530 152
rect 518 128 522 132
rect 486 118 490 122
rect 502 78 506 82
rect 534 118 538 122
rect 542 88 546 92
rect 550 78 554 82
rect 494 68 498 72
rect 486 8 490 12
rect 694 338 698 342
rect 702 328 706 332
rect 670 318 674 322
rect 758 428 762 432
rect 814 418 818 422
rect 758 368 762 372
rect 766 368 770 372
rect 806 368 810 372
rect 726 348 730 352
rect 854 348 858 352
rect 726 338 730 342
rect 718 318 722 322
rect 662 288 666 292
rect 638 278 642 282
rect 646 258 650 262
rect 654 258 658 262
rect 678 258 682 262
rect 694 258 698 262
rect 686 248 690 252
rect 686 218 690 222
rect 758 328 762 332
rect 758 268 762 272
rect 838 338 842 342
rect 846 338 850 342
rect 838 328 842 332
rect 822 308 826 312
rect 846 288 850 292
rect 790 278 794 282
rect 806 278 810 282
rect 830 268 834 272
rect 926 608 930 612
rect 894 578 898 582
rect 934 548 938 552
rect 902 538 906 542
rect 974 668 978 672
rect 990 668 994 672
rect 966 658 970 662
rect 974 588 978 592
rect 966 528 970 532
rect 918 518 922 522
rect 910 508 914 512
rect 942 488 946 492
rect 982 568 986 572
rect 990 538 994 542
rect 990 528 994 532
rect 1062 828 1066 832
rect 1078 768 1082 772
rect 1070 758 1074 762
rect 1062 738 1066 742
rect 1046 718 1050 722
rect 1062 718 1066 722
rect 1046 678 1050 682
rect 1022 668 1026 672
rect 1014 658 1018 662
rect 1038 658 1042 662
rect 1022 648 1026 652
rect 1046 648 1050 652
rect 1030 558 1034 562
rect 1022 538 1026 542
rect 1022 528 1026 532
rect 982 518 986 522
rect 878 478 882 482
rect 886 478 890 482
rect 934 478 938 482
rect 958 478 962 482
rect 886 468 890 472
rect 878 458 882 462
rect 870 348 874 352
rect 958 448 962 452
rect 990 458 994 462
rect 974 428 978 432
rect 926 408 930 412
rect 902 398 906 402
rect 886 378 890 382
rect 958 378 962 382
rect 982 378 986 382
rect 1006 428 1010 432
rect 1014 428 1018 432
rect 998 398 1002 402
rect 990 358 994 362
rect 942 348 946 352
rect 958 348 962 352
rect 878 338 882 342
rect 934 338 938 342
rect 910 318 914 322
rect 878 278 882 282
rect 886 278 890 282
rect 902 278 906 282
rect 934 278 938 282
rect 966 338 970 342
rect 990 328 994 332
rect 1030 448 1034 452
rect 1022 398 1026 402
rect 1086 758 1090 762
rect 1102 758 1106 762
rect 1086 738 1090 742
rect 1102 738 1106 742
rect 1078 728 1082 732
rect 1078 698 1082 702
rect 1070 668 1074 672
rect 1054 638 1058 642
rect 1062 638 1066 642
rect 1046 618 1050 622
rect 1062 548 1066 552
rect 1094 658 1098 662
rect 1102 528 1106 532
rect 1086 518 1090 522
rect 1078 508 1082 512
rect 1062 498 1066 502
rect 1054 488 1058 492
rect 1086 498 1090 502
rect 1118 818 1122 822
rect 1126 778 1130 782
rect 1118 758 1122 762
rect 1118 718 1122 722
rect 1190 898 1194 902
rect 1222 878 1226 882
rect 1246 878 1250 882
rect 1254 878 1258 882
rect 1214 868 1218 872
rect 1222 868 1226 872
rect 1238 858 1242 862
rect 1254 858 1258 862
rect 1182 848 1186 852
rect 1254 788 1258 792
rect 1166 748 1170 752
rect 1198 748 1202 752
rect 1222 748 1226 752
rect 1238 748 1242 752
rect 1142 740 1146 742
rect 1142 738 1146 740
rect 1238 738 1242 742
rect 1246 738 1250 742
rect 1318 1058 1322 1062
rect 1334 1058 1338 1062
rect 1310 1048 1314 1052
rect 1302 968 1306 972
rect 1350 1098 1354 1102
rect 1366 1098 1370 1102
rect 1358 1088 1362 1092
rect 1638 1158 1642 1162
rect 1566 1148 1570 1152
rect 1630 1148 1634 1152
rect 1430 1128 1434 1132
rect 1414 1098 1418 1102
rect 1398 1088 1402 1092
rect 1390 1078 1394 1082
rect 1454 1128 1458 1132
rect 1462 1128 1466 1132
rect 1518 1128 1522 1132
rect 1486 1108 1490 1112
rect 1486 1088 1490 1092
rect 1454 1078 1458 1082
rect 1366 1068 1370 1072
rect 1446 1068 1450 1072
rect 1518 1088 1522 1092
rect 1582 1138 1586 1142
rect 1614 1140 1618 1142
rect 1614 1138 1618 1140
rect 1638 1138 1642 1142
rect 1590 1128 1594 1132
rect 1622 1128 1626 1132
rect 1662 1128 1666 1132
rect 1542 1118 1546 1122
rect 1654 1118 1658 1122
rect 1590 1098 1594 1102
rect 1582 1088 1586 1092
rect 1526 1078 1530 1082
rect 1542 1068 1546 1072
rect 1702 1140 1706 1142
rect 1702 1138 1706 1140
rect 1710 1128 1714 1132
rect 1710 1108 1714 1112
rect 1686 1098 1690 1102
rect 1702 1098 1706 1102
rect 1622 1088 1626 1092
rect 1614 1068 1618 1072
rect 1774 1138 1778 1142
rect 1814 1138 1818 1142
rect 1838 1138 1842 1142
rect 1782 1128 1786 1132
rect 1790 1118 1794 1122
rect 1814 1128 1818 1132
rect 1742 1078 1746 1082
rect 1766 1078 1770 1082
rect 1782 1068 1786 1072
rect 1822 1098 1826 1102
rect 1374 1058 1378 1062
rect 1406 1058 1410 1062
rect 1438 1058 1442 1062
rect 1462 1058 1466 1062
rect 1494 1058 1498 1062
rect 1526 1058 1530 1062
rect 1654 1058 1658 1062
rect 1342 1028 1346 1032
rect 1326 978 1330 982
rect 1270 928 1274 932
rect 1294 928 1298 932
rect 1286 918 1290 922
rect 1318 938 1322 942
rect 1278 908 1282 912
rect 1302 908 1306 912
rect 1342 968 1346 972
rect 1366 968 1370 972
rect 1334 948 1338 952
rect 1310 878 1314 882
rect 1278 868 1282 872
rect 1286 868 1290 872
rect 1270 768 1274 772
rect 1270 748 1274 752
rect 1158 728 1162 732
rect 1134 698 1138 702
rect 1182 698 1186 702
rect 1142 678 1146 682
rect 1198 678 1202 682
rect 1142 668 1146 672
rect 1142 648 1146 652
rect 1118 568 1122 572
rect 1126 538 1130 542
rect 1118 528 1122 532
rect 1086 478 1090 482
rect 1094 478 1098 482
rect 1110 468 1114 472
rect 1046 448 1050 452
rect 1086 428 1090 432
rect 1078 388 1082 392
rect 1014 348 1018 352
rect 1046 338 1050 342
rect 1070 338 1074 342
rect 1022 328 1026 332
rect 1102 368 1106 372
rect 1134 508 1138 512
rect 1126 498 1130 502
rect 1230 708 1234 712
rect 1230 668 1234 672
rect 1190 658 1194 662
rect 1174 638 1178 642
rect 1166 618 1170 622
rect 1262 668 1266 672
rect 1270 628 1274 632
rect 1254 608 1258 612
rect 1206 588 1210 592
rect 1246 588 1250 592
rect 1150 578 1154 582
rect 1206 568 1210 572
rect 1206 558 1210 562
rect 1254 558 1258 562
rect 1294 738 1298 742
rect 1302 718 1306 722
rect 1286 698 1290 702
rect 1294 698 1298 702
rect 1286 638 1290 642
rect 1198 548 1202 552
rect 1278 548 1282 552
rect 1326 858 1330 862
rect 1478 1048 1482 1052
rect 1414 978 1418 982
rect 1350 928 1354 932
rect 1406 928 1410 932
rect 1390 918 1394 922
rect 1374 908 1378 912
rect 1358 868 1362 872
rect 1390 898 1394 902
rect 1502 1028 1506 1032
rect 1510 1028 1514 1032
rect 1478 958 1482 962
rect 1382 878 1386 882
rect 1414 878 1418 882
rect 1454 928 1458 932
rect 1478 928 1482 932
rect 1494 928 1498 932
rect 1446 888 1450 892
rect 1454 878 1458 882
rect 1486 888 1490 892
rect 1382 868 1386 872
rect 1406 858 1410 862
rect 1350 848 1354 852
rect 1510 1018 1514 1022
rect 1638 1038 1642 1042
rect 1558 1018 1562 1022
rect 1550 988 1554 992
rect 1574 988 1578 992
rect 1630 988 1634 992
rect 1566 958 1570 962
rect 1654 968 1658 972
rect 1662 958 1666 962
rect 1598 948 1602 952
rect 1702 948 1706 952
rect 1590 938 1594 942
rect 1502 918 1506 922
rect 1550 908 1554 912
rect 1518 898 1522 902
rect 1542 878 1546 882
rect 1526 868 1530 872
rect 1518 848 1522 852
rect 1446 768 1450 772
rect 1342 758 1346 762
rect 1390 758 1394 762
rect 1406 758 1410 762
rect 1334 748 1338 752
rect 1366 748 1370 752
rect 1414 748 1418 752
rect 1446 748 1450 752
rect 1382 738 1386 742
rect 1318 728 1322 732
rect 1342 728 1346 732
rect 1406 698 1410 702
rect 1342 678 1346 682
rect 1350 668 1354 672
rect 1382 668 1386 672
rect 1350 648 1354 652
rect 1430 738 1434 742
rect 1454 738 1458 742
rect 1462 708 1466 712
rect 1502 728 1506 732
rect 1510 688 1514 692
rect 1494 678 1498 682
rect 1494 668 1498 672
rect 1510 668 1514 672
rect 1582 918 1586 922
rect 1582 908 1586 912
rect 1566 878 1570 882
rect 1574 868 1578 872
rect 1598 878 1602 882
rect 1590 858 1594 862
rect 1558 748 1562 752
rect 1582 748 1586 752
rect 1526 718 1530 722
rect 1422 658 1426 662
rect 1462 658 1466 662
rect 1470 658 1474 662
rect 1398 648 1402 652
rect 1414 648 1418 652
rect 1374 618 1378 622
rect 1326 578 1330 582
rect 1310 558 1314 562
rect 1342 548 1346 552
rect 1150 538 1154 542
rect 1190 528 1194 532
rect 1222 528 1226 532
rect 1230 518 1234 522
rect 1174 508 1178 512
rect 1214 498 1218 502
rect 1166 470 1170 472
rect 1166 468 1170 470
rect 1206 468 1210 472
rect 1174 458 1178 462
rect 1198 458 1202 462
rect 1118 428 1122 432
rect 1110 358 1114 362
rect 1182 398 1186 402
rect 1198 398 1202 402
rect 1142 388 1146 392
rect 1086 338 1090 342
rect 1118 338 1122 342
rect 1046 318 1050 322
rect 1150 318 1154 322
rect 1030 308 1034 312
rect 1054 288 1058 292
rect 1014 278 1018 282
rect 1022 268 1026 272
rect 774 258 778 262
rect 798 258 802 262
rect 830 258 834 262
rect 742 248 746 252
rect 774 248 778 252
rect 718 228 722 232
rect 838 228 842 232
rect 782 218 786 222
rect 814 218 818 222
rect 830 218 834 222
rect 742 208 746 212
rect 694 188 698 192
rect 622 168 626 172
rect 638 158 642 162
rect 670 148 674 152
rect 790 198 794 202
rect 758 168 762 172
rect 798 168 802 172
rect 766 158 770 162
rect 654 138 658 142
rect 614 128 618 132
rect 646 128 650 132
rect 662 128 666 132
rect 726 128 730 132
rect 750 128 754 132
rect 774 128 778 132
rect 782 128 786 132
rect 718 118 722 122
rect 638 98 642 102
rect 614 88 618 92
rect 766 108 770 112
rect 790 118 794 122
rect 806 138 810 142
rect 822 128 826 132
rect 798 108 802 112
rect 822 108 826 112
rect 670 78 674 82
rect 718 78 722 82
rect 694 68 698 72
rect 790 68 794 72
rect 662 58 666 62
rect 686 58 690 62
rect 710 58 714 62
rect 766 58 770 62
rect 598 48 602 52
rect 702 48 706 52
rect 526 8 530 12
rect 798 58 802 62
rect 1022 248 1026 252
rect 870 218 874 222
rect 910 218 914 222
rect 990 218 994 222
rect 886 208 890 212
rect 902 208 906 212
rect 1190 388 1194 392
rect 1190 378 1194 382
rect 1198 348 1202 352
rect 1278 538 1282 542
rect 1342 538 1346 542
rect 1366 538 1370 542
rect 1318 528 1322 532
rect 1278 478 1282 482
rect 1326 498 1330 502
rect 1334 498 1338 502
rect 1262 468 1266 472
rect 1294 468 1298 472
rect 1350 528 1354 532
rect 1366 528 1370 532
rect 1366 508 1370 512
rect 1230 458 1234 462
rect 1254 458 1258 462
rect 1294 458 1298 462
rect 1238 408 1242 412
rect 1246 408 1250 412
rect 1222 348 1226 352
rect 1206 338 1210 342
rect 1230 338 1234 342
rect 1246 338 1250 342
rect 1310 448 1314 452
rect 1334 358 1338 362
rect 1222 328 1226 332
rect 1270 328 1274 332
rect 1134 278 1138 282
rect 1174 278 1178 282
rect 1086 268 1090 272
rect 1102 268 1106 272
rect 1142 268 1146 272
rect 1166 268 1170 272
rect 1126 258 1130 262
rect 1086 248 1090 252
rect 1118 248 1122 252
rect 1062 228 1066 232
rect 1070 218 1074 222
rect 1054 198 1058 202
rect 998 188 1002 192
rect 1030 188 1034 192
rect 926 168 930 172
rect 918 148 922 152
rect 958 148 962 152
rect 982 148 986 152
rect 1014 158 1018 162
rect 1078 148 1082 152
rect 854 138 858 142
rect 902 140 906 142
rect 902 138 906 140
rect 934 138 938 142
rect 1094 138 1098 142
rect 1110 138 1114 142
rect 846 108 850 112
rect 838 98 842 102
rect 854 98 858 102
rect 846 88 850 92
rect 830 68 834 72
rect 822 48 826 52
rect 782 28 786 32
rect 902 108 906 112
rect 878 98 882 102
rect 894 98 898 102
rect 1006 118 1010 122
rect 966 78 970 82
rect 910 68 914 72
rect 926 68 930 72
rect 958 68 962 72
rect 1038 118 1042 122
rect 1062 118 1066 122
rect 1230 278 1234 282
rect 1278 308 1282 312
rect 1278 298 1282 302
rect 1302 288 1306 292
rect 1326 288 1330 292
rect 1302 278 1306 282
rect 1310 278 1314 282
rect 1238 268 1242 272
rect 1286 268 1290 272
rect 1302 268 1306 272
rect 1182 258 1186 262
rect 1214 258 1218 262
rect 1246 258 1250 262
rect 1262 258 1266 262
rect 1310 258 1314 262
rect 1166 248 1170 252
rect 1326 238 1330 242
rect 1142 198 1146 202
rect 1150 168 1154 172
rect 1190 168 1194 172
rect 1198 168 1202 172
rect 1134 158 1138 162
rect 1142 158 1146 162
rect 1126 128 1130 132
rect 1014 88 1018 92
rect 1038 88 1042 92
rect 1102 88 1106 92
rect 982 78 986 82
rect 998 78 1002 82
rect 1126 78 1130 82
rect 998 68 1002 72
rect 1214 168 1218 172
rect 1198 158 1202 162
rect 1206 158 1210 162
rect 1182 148 1186 152
rect 1190 108 1194 112
rect 1206 148 1210 152
rect 1230 138 1234 142
rect 1350 378 1354 382
rect 1398 598 1402 602
rect 1422 588 1426 592
rect 1382 578 1386 582
rect 1446 648 1450 652
rect 1398 568 1402 572
rect 1438 568 1442 572
rect 1454 568 1458 572
rect 1478 618 1482 622
rect 1518 558 1522 562
rect 1414 548 1418 552
rect 1462 548 1466 552
rect 1518 548 1522 552
rect 1438 538 1442 542
rect 1542 708 1546 712
rect 1542 668 1546 672
rect 1542 618 1546 622
rect 1542 608 1546 612
rect 1574 738 1578 742
rect 1598 838 1602 842
rect 1614 868 1618 872
rect 1606 768 1610 772
rect 1806 1048 1810 1052
rect 1782 1038 1786 1042
rect 1774 988 1778 992
rect 1830 1058 1834 1062
rect 1846 1058 1850 1062
rect 1838 1048 1842 1052
rect 1830 1038 1834 1042
rect 1798 968 1802 972
rect 1814 968 1818 972
rect 1678 938 1682 942
rect 1718 938 1722 942
rect 1654 918 1658 922
rect 1638 878 1642 882
rect 1630 868 1634 872
rect 1694 888 1698 892
rect 1662 868 1666 872
rect 1638 858 1642 862
rect 1646 858 1650 862
rect 1678 848 1682 852
rect 1710 928 1714 932
rect 1774 928 1778 932
rect 1790 928 1794 932
rect 1742 918 1746 922
rect 1806 928 1810 932
rect 1854 1008 1858 1012
rect 1854 998 1858 1002
rect 1822 918 1826 922
rect 1798 878 1802 882
rect 1718 868 1722 872
rect 1662 768 1666 772
rect 1734 768 1738 772
rect 1622 758 1626 762
rect 1654 758 1658 762
rect 1606 748 1610 752
rect 1622 748 1626 752
rect 1670 748 1674 752
rect 1558 728 1562 732
rect 1590 728 1594 732
rect 1598 728 1602 732
rect 1806 868 1810 872
rect 1814 868 1818 872
rect 1774 858 1778 862
rect 1750 838 1754 842
rect 1750 748 1754 752
rect 1742 738 1746 742
rect 1694 728 1698 732
rect 1686 718 1690 722
rect 1726 718 1730 722
rect 1718 698 1722 702
rect 1678 688 1682 692
rect 1590 678 1594 682
rect 1846 928 1850 932
rect 1862 978 1866 982
rect 1862 918 1866 922
rect 1846 878 1850 882
rect 1838 868 1842 872
rect 1830 858 1834 862
rect 1838 858 1842 862
rect 1830 748 1834 752
rect 1774 740 1778 742
rect 1774 738 1778 740
rect 1862 740 1866 742
rect 1862 738 1866 740
rect 1766 718 1770 722
rect 1774 718 1778 722
rect 1766 698 1770 702
rect 1662 678 1666 682
rect 1694 678 1698 682
rect 1726 678 1730 682
rect 1742 678 1746 682
rect 1566 668 1570 672
rect 1590 668 1594 672
rect 1574 658 1578 662
rect 1550 548 1554 552
rect 1494 538 1498 542
rect 1390 528 1394 532
rect 1446 528 1450 532
rect 1486 528 1490 532
rect 1526 528 1530 532
rect 1390 518 1394 522
rect 1462 508 1466 512
rect 1502 508 1506 512
rect 1406 468 1410 472
rect 1430 468 1434 472
rect 1470 478 1474 482
rect 1510 478 1514 482
rect 1494 470 1498 472
rect 1494 468 1498 470
rect 1526 470 1530 472
rect 1526 468 1530 470
rect 1390 458 1394 462
rect 1438 458 1442 462
rect 1478 458 1482 462
rect 1382 438 1386 442
rect 1358 368 1362 372
rect 1374 368 1378 372
rect 1358 358 1362 362
rect 1462 448 1466 452
rect 1502 448 1506 452
rect 1414 428 1418 432
rect 1446 418 1450 422
rect 1414 408 1418 412
rect 1390 378 1394 382
rect 1390 368 1394 372
rect 1366 338 1370 342
rect 1358 318 1362 322
rect 1350 308 1354 312
rect 1430 358 1434 362
rect 1398 318 1402 322
rect 1422 318 1426 322
rect 1398 308 1402 312
rect 1502 398 1506 402
rect 1526 358 1530 362
rect 1446 348 1450 352
rect 1542 508 1546 512
rect 1566 638 1570 642
rect 1598 628 1602 632
rect 1654 658 1658 662
rect 1638 648 1642 652
rect 1630 628 1634 632
rect 1686 668 1690 672
rect 1758 678 1762 682
rect 1718 668 1722 672
rect 1822 728 1826 732
rect 1854 728 1858 732
rect 1814 718 1818 722
rect 1790 678 1794 682
rect 1830 718 1834 722
rect 1854 718 1858 722
rect 1846 708 1850 712
rect 1702 658 1706 662
rect 1686 608 1690 612
rect 1870 678 1874 682
rect 1734 638 1738 642
rect 1814 628 1818 632
rect 1718 588 1722 592
rect 1766 588 1770 592
rect 1630 578 1634 582
rect 1622 558 1626 562
rect 1686 558 1690 562
rect 1734 558 1738 562
rect 1630 548 1634 552
rect 1574 528 1578 532
rect 1590 498 1594 502
rect 1558 488 1562 492
rect 1574 488 1578 492
rect 1622 538 1626 542
rect 1654 538 1658 542
rect 1678 528 1682 532
rect 1606 518 1610 522
rect 1566 478 1570 482
rect 1566 368 1570 372
rect 1558 358 1562 362
rect 1558 348 1562 352
rect 1494 338 1498 342
rect 1534 338 1538 342
rect 1446 318 1450 322
rect 1462 318 1466 322
rect 1390 278 1394 282
rect 1398 278 1402 282
rect 1406 268 1410 272
rect 1486 308 1490 312
rect 1486 298 1490 302
rect 1478 288 1482 292
rect 1534 308 1538 312
rect 1510 288 1514 292
rect 1510 278 1514 282
rect 1526 278 1530 282
rect 1382 218 1386 222
rect 1398 228 1402 232
rect 1350 188 1354 192
rect 1390 188 1394 192
rect 1342 168 1346 172
rect 1390 158 1394 162
rect 1318 148 1322 152
rect 1366 148 1370 152
rect 1222 128 1226 132
rect 1246 128 1250 132
rect 1278 138 1282 142
rect 1262 118 1266 122
rect 1310 138 1314 142
rect 1326 138 1330 142
rect 1342 138 1346 142
rect 1374 138 1378 142
rect 1318 128 1322 132
rect 1238 108 1242 112
rect 1254 108 1258 112
rect 1278 108 1282 112
rect 1294 108 1298 112
rect 1206 88 1210 92
rect 1150 68 1154 72
rect 1190 68 1194 72
rect 1030 58 1034 62
rect 1046 58 1050 62
rect 1054 58 1058 62
rect 1086 58 1090 62
rect 1150 58 1154 62
rect 886 48 890 52
rect 950 48 954 52
rect 862 38 866 42
rect 870 38 874 42
rect 878 38 882 42
rect 870 28 874 32
rect 966 8 970 12
rect 1054 8 1058 12
rect 1230 68 1234 72
rect 1246 70 1250 72
rect 1246 68 1250 70
rect 1294 78 1298 82
rect 1358 78 1362 82
rect 1342 68 1346 72
rect 1366 68 1370 72
rect 1454 258 1458 262
rect 1422 218 1426 222
rect 1446 218 1450 222
rect 1414 208 1418 212
rect 1446 178 1450 182
rect 1494 238 1498 242
rect 1478 198 1482 202
rect 1494 188 1498 192
rect 1430 148 1434 152
rect 1446 148 1450 152
rect 1510 148 1514 152
rect 1406 138 1410 142
rect 1470 138 1474 142
rect 1478 128 1482 132
rect 1438 108 1442 112
rect 1454 108 1458 112
rect 1438 88 1442 92
rect 1550 288 1554 292
rect 1550 278 1554 282
rect 1582 368 1586 372
rect 1646 508 1650 512
rect 1630 488 1634 492
rect 1694 548 1698 552
rect 1750 548 1754 552
rect 1782 548 1786 552
rect 1790 548 1794 552
rect 1686 468 1690 472
rect 1638 458 1642 462
rect 1614 368 1618 372
rect 1662 388 1666 392
rect 1686 358 1690 362
rect 1606 348 1610 352
rect 1622 348 1626 352
rect 1646 338 1650 342
rect 1646 328 1650 332
rect 1590 318 1594 322
rect 1606 318 1610 322
rect 1622 318 1626 322
rect 1574 298 1578 302
rect 1574 278 1578 282
rect 1622 308 1626 312
rect 1646 288 1650 292
rect 1614 278 1618 282
rect 1622 268 1626 272
rect 1702 538 1706 542
rect 1702 478 1706 482
rect 1726 478 1730 482
rect 1758 508 1762 512
rect 1822 568 1826 572
rect 1830 558 1834 562
rect 1862 558 1866 562
rect 1838 548 1842 552
rect 1870 548 1874 552
rect 1814 488 1818 492
rect 1750 478 1754 482
rect 1718 468 1722 472
rect 1702 388 1706 392
rect 1750 458 1754 462
rect 1798 458 1802 462
rect 1878 538 1882 542
rect 1878 528 1882 532
rect 1846 518 1850 522
rect 1838 498 1842 502
rect 1830 448 1834 452
rect 1710 338 1714 342
rect 1710 328 1714 332
rect 1742 328 1746 332
rect 1726 288 1730 292
rect 1702 278 1706 282
rect 1806 328 1810 332
rect 1798 318 1802 322
rect 1806 318 1810 322
rect 1798 308 1802 312
rect 1758 298 1762 302
rect 1750 278 1754 282
rect 1694 268 1698 272
rect 1710 268 1714 272
rect 1726 270 1730 272
rect 1726 268 1730 270
rect 1558 258 1562 262
rect 1590 248 1594 252
rect 1542 238 1546 242
rect 1574 218 1578 222
rect 1590 198 1594 202
rect 1598 198 1602 202
rect 1534 178 1538 182
rect 1550 168 1554 172
rect 1574 158 1578 162
rect 1558 148 1562 152
rect 1518 138 1522 142
rect 1534 128 1538 132
rect 1510 118 1514 122
rect 1534 98 1538 102
rect 1534 78 1538 82
rect 1414 68 1418 72
rect 1430 68 1434 72
rect 1462 68 1466 72
rect 1486 68 1490 72
rect 1278 58 1282 62
rect 1326 58 1330 62
rect 1222 38 1226 42
rect 1230 38 1234 42
rect 1214 28 1218 32
rect 1198 8 1202 12
rect 1214 8 1218 12
rect 1254 28 1258 32
rect 1350 58 1354 62
rect 1342 48 1346 52
rect 1390 48 1394 52
rect 1334 38 1338 42
rect 1254 8 1258 12
rect 1326 8 1330 12
rect 1486 58 1490 62
rect 1502 58 1506 62
rect 1694 258 1698 262
rect 1678 238 1682 242
rect 1646 218 1650 222
rect 1630 208 1634 212
rect 1606 158 1610 162
rect 1670 178 1674 182
rect 1622 148 1626 152
rect 1606 138 1610 142
rect 1622 128 1626 132
rect 1646 128 1650 132
rect 1662 118 1666 122
rect 1646 98 1650 102
rect 1670 98 1674 102
rect 1590 78 1594 82
rect 1622 78 1626 82
rect 1638 78 1642 82
rect 1526 58 1530 62
rect 1558 58 1562 62
rect 1670 88 1674 92
rect 1654 68 1658 72
rect 1702 148 1706 152
rect 1750 268 1754 272
rect 1766 268 1770 272
rect 1782 270 1786 272
rect 1782 268 1786 270
rect 1742 198 1746 202
rect 1742 188 1746 192
rect 1742 158 1746 162
rect 1718 138 1722 142
rect 1734 128 1738 132
rect 1694 68 1698 72
rect 1814 308 1818 312
rect 1766 188 1770 192
rect 1830 398 1834 402
rect 1862 468 1866 472
rect 1838 368 1842 372
rect 1854 368 1858 372
rect 1830 298 1834 302
rect 1830 278 1834 282
rect 1830 258 1834 262
rect 1846 258 1850 262
rect 1838 188 1842 192
rect 1846 168 1850 172
rect 1814 158 1818 162
rect 1822 158 1826 162
rect 1854 158 1858 162
rect 1782 148 1786 152
rect 1822 148 1826 152
rect 1758 138 1762 142
rect 1774 138 1778 142
rect 1766 98 1770 102
rect 1750 78 1754 82
rect 1758 78 1762 82
rect 1806 118 1810 122
rect 1806 88 1810 92
rect 1830 88 1834 92
rect 1782 78 1786 82
rect 1846 78 1850 82
rect 1774 68 1778 72
rect 1886 318 1890 322
rect 1886 258 1890 262
rect 1678 58 1682 62
rect 1702 58 1706 62
rect 1822 58 1826 62
rect 1878 58 1882 62
rect 1590 48 1594 52
<< metal3 >>
rect 866 1208 878 1211
rect 562 1178 614 1181
rect 954 1178 1118 1181
rect 354 1168 846 1171
rect 1130 1168 1142 1171
rect 1226 1168 1558 1171
rect -26 1158 6 1161
rect 338 1158 582 1161
rect 890 1158 934 1161
rect 938 1158 1022 1161
rect 1426 1158 1438 1161
rect 1442 1158 1638 1161
rect 210 1148 230 1151
rect 274 1148 278 1151
rect 290 1148 390 1151
rect 394 1148 414 1151
rect 426 1148 438 1151
rect 550 1148 558 1151
rect 586 1148 678 1151
rect 690 1148 702 1151
rect 858 1148 878 1151
rect 930 1148 942 1151
rect 970 1148 982 1151
rect 986 1148 1038 1151
rect 1122 1148 1214 1151
rect 1266 1148 1366 1151
rect 1378 1148 1406 1151
rect 1570 1148 1630 1151
rect 218 1138 270 1141
rect 282 1138 478 1141
rect 482 1138 582 1141
rect 586 1138 670 1141
rect 698 1138 750 1141
rect 850 1138 894 1141
rect 898 1138 990 1141
rect 994 1138 998 1141
rect 1010 1138 1086 1141
rect 1090 1138 1222 1141
rect 1234 1138 1294 1141
rect 1322 1138 1582 1141
rect 1586 1138 1614 1141
rect 1642 1138 1702 1141
rect 1778 1138 1814 1141
rect 1834 1138 1838 1141
rect 82 1128 150 1131
rect 154 1128 486 1131
rect 538 1128 566 1131
rect 570 1128 590 1131
rect 610 1128 758 1131
rect 978 1128 1158 1131
rect 1162 1128 1318 1131
rect 1434 1128 1454 1131
rect 1466 1128 1502 1131
rect 1522 1128 1590 1131
rect 1610 1128 1622 1131
rect 1646 1128 1662 1131
rect 1714 1128 1782 1131
rect 1786 1128 1814 1131
rect 138 1118 174 1121
rect 226 1118 246 1121
rect 250 1118 286 1121
rect 298 1118 382 1121
rect 450 1118 494 1121
rect 578 1118 630 1121
rect 634 1118 774 1121
rect 778 1118 1102 1121
rect 1106 1118 1278 1121
rect 1646 1121 1649 1128
rect 1546 1118 1649 1121
rect 1658 1118 1790 1121
rect 202 1108 310 1111
rect 354 1108 382 1111
rect 402 1108 430 1111
rect 434 1108 470 1111
rect 630 1108 806 1111
rect 810 1108 814 1111
rect 818 1108 990 1111
rect 994 1108 1014 1111
rect 1226 1108 1238 1111
rect 1258 1108 1334 1111
rect 1490 1108 1710 1111
rect 234 1098 270 1101
rect 274 1098 414 1101
rect 458 1098 478 1101
rect 514 1098 518 1101
rect 554 1098 566 1101
rect 630 1101 633 1108
rect 570 1098 633 1101
rect 674 1098 766 1101
rect 1002 1098 1078 1101
rect 1082 1098 1254 1101
rect 1266 1098 1270 1101
rect 1354 1098 1366 1101
rect 1378 1098 1414 1101
rect 1594 1098 1686 1101
rect 1706 1098 1822 1101
rect 50 1088 86 1091
rect 90 1088 334 1091
rect 346 1088 406 1091
rect 410 1088 558 1091
rect 562 1088 630 1091
rect 634 1088 766 1091
rect 770 1088 814 1091
rect 914 1088 1006 1091
rect 1010 1088 1262 1091
rect 1362 1088 1398 1091
rect 1402 1088 1486 1091
rect 1490 1088 1518 1091
rect 1586 1088 1622 1091
rect -26 1078 6 1081
rect 10 1078 46 1081
rect 250 1078 262 1081
rect 338 1078 870 1081
rect 938 1078 950 1081
rect 1058 1078 1078 1081
rect 1082 1078 1174 1081
rect 1178 1078 1390 1081
rect 1394 1078 1454 1081
rect 1458 1078 1526 1081
rect 1538 1078 1742 1081
rect 1754 1078 1766 1081
rect 178 1068 206 1071
rect 210 1068 254 1071
rect 266 1068 278 1071
rect 314 1068 350 1071
rect 362 1068 398 1071
rect 850 1068 966 1071
rect 978 1068 990 1071
rect 1002 1068 1062 1071
rect 1066 1068 1126 1071
rect 1138 1068 1142 1071
rect 1154 1068 1166 1071
rect 1202 1068 1222 1071
rect 1266 1068 1302 1071
rect 1306 1068 1310 1071
rect 1370 1068 1446 1071
rect 1450 1068 1542 1071
rect 1546 1068 1614 1071
rect 1618 1068 1782 1071
rect -26 1058 22 1061
rect 26 1058 38 1061
rect 42 1058 94 1061
rect 162 1058 182 1061
rect 258 1058 470 1061
rect 474 1058 606 1061
rect 610 1058 622 1061
rect 650 1058 654 1061
rect 670 1058 678 1061
rect 798 1061 801 1068
rect 798 1058 806 1061
rect 818 1058 838 1061
rect 874 1058 926 1061
rect 1042 1058 1054 1061
rect 1058 1058 1118 1061
rect 1138 1058 1270 1061
rect 1322 1058 1326 1061
rect 1338 1058 1374 1061
rect 1398 1058 1406 1061
rect 1450 1058 1462 1061
rect 1506 1058 1526 1061
rect 1834 1058 1846 1061
rect 122 1048 174 1051
rect 226 1048 262 1051
rect 266 1048 486 1051
rect 530 1048 742 1051
rect 746 1048 958 1051
rect 1090 1048 1150 1051
rect 1314 1048 1478 1051
rect 1494 1048 1497 1058
rect 1810 1048 1838 1051
rect 58 1038 286 1041
rect 378 1038 454 1041
rect 466 1038 486 1041
rect 658 1038 718 1041
rect 754 1038 886 1041
rect 1050 1038 1062 1041
rect 1114 1038 1190 1041
rect 1194 1038 1230 1041
rect 1234 1038 1638 1041
rect 1786 1038 1830 1041
rect 18 1028 62 1031
rect 66 1028 142 1031
rect 290 1028 502 1031
rect 834 1028 862 1031
rect 906 1028 1190 1031
rect 1266 1028 1342 1031
rect 1506 1028 1510 1031
rect 1514 1028 1534 1031
rect 50 1018 62 1021
rect 114 1018 166 1021
rect 266 1018 278 1021
rect 290 1018 414 1021
rect 418 1018 798 1021
rect 986 1018 1038 1021
rect 1514 1018 1558 1021
rect 178 1008 262 1011
rect 450 1008 462 1011
rect 466 1008 846 1011
rect 898 1008 910 1011
rect 914 1008 1086 1011
rect 1258 1008 1854 1011
rect 138 998 278 1001
rect 586 998 790 1001
rect 794 998 798 1001
rect 818 998 1262 1001
rect 1834 998 1854 1001
rect 602 988 646 991
rect 754 988 998 991
rect 1218 988 1238 991
rect 1554 988 1574 991
rect 1634 988 1774 991
rect 1778 988 1822 991
rect 482 978 534 981
rect 794 978 1102 981
rect 1186 978 1326 981
rect 1418 978 1862 981
rect 242 968 622 971
rect 626 968 1302 971
rect 1306 968 1342 971
rect 1370 968 1654 971
rect 1802 968 1814 971
rect -26 958 6 961
rect 186 958 254 961
rect 322 958 350 961
rect 466 958 494 961
rect 498 958 654 961
rect 866 958 902 961
rect 1002 958 1022 961
rect 1122 958 1198 961
rect 1210 958 1230 961
rect 1482 958 1566 961
rect 1570 958 1662 961
rect 178 948 190 951
rect 250 948 270 951
rect 298 948 318 951
rect 394 948 446 951
rect 506 948 542 951
rect 562 948 638 951
rect 674 948 702 951
rect 938 948 966 951
rect 970 948 974 951
rect 978 948 1070 951
rect 1154 948 1206 951
rect 1338 948 1590 951
rect 1602 948 1606 951
rect 1706 948 1734 951
rect 1590 942 1593 948
rect 106 938 206 941
rect 254 938 262 941
rect 354 938 382 941
rect 530 938 534 941
rect 610 938 662 941
rect 666 938 678 941
rect 722 938 766 941
rect 786 938 822 941
rect 826 938 846 941
rect 962 938 990 941
rect 1066 938 1094 941
rect 1098 938 1166 941
rect 1178 938 1318 941
rect 1682 938 1718 941
rect 254 932 257 938
rect 98 928 102 931
rect 162 928 190 931
rect 346 928 350 931
rect 354 928 566 931
rect 570 928 646 931
rect 666 928 678 931
rect 730 928 750 931
rect 762 928 998 931
rect 1050 928 1158 931
rect 1194 928 1214 931
rect 1226 928 1230 931
rect 1274 928 1294 931
rect 1298 928 1302 931
rect 1410 928 1454 931
rect 1458 928 1478 931
rect 1482 928 1494 931
rect 1498 928 1710 931
rect 1714 928 1774 931
rect 1778 928 1790 931
rect 1810 928 1846 931
rect 1350 922 1353 928
rect 66 918 70 921
rect 74 918 102 921
rect 130 918 294 921
rect 362 918 430 921
rect 498 918 518 921
rect 530 918 574 921
rect 634 918 966 921
rect 1042 918 1086 921
rect 1090 918 1174 921
rect 1290 918 1326 921
rect 1362 918 1390 921
rect 1394 918 1502 921
rect 1586 918 1654 921
rect 1746 918 1822 921
rect 1826 918 1862 921
rect 82 908 94 911
rect 338 908 366 911
rect 762 908 766 911
rect 794 908 838 911
rect 842 908 854 911
rect 858 908 910 911
rect 930 908 950 911
rect 954 908 1182 911
rect 1282 908 1302 911
rect 1306 908 1374 911
rect 1554 908 1582 911
rect 410 898 422 901
rect 434 898 582 901
rect 642 898 846 901
rect 930 898 1038 901
rect 1514 898 1518 901
rect 1190 892 1193 898
rect 66 888 78 891
rect 82 888 230 891
rect 266 888 438 891
rect 474 888 534 891
rect 586 888 758 891
rect 762 888 854 891
rect 858 888 934 891
rect 938 888 1030 891
rect 1390 891 1393 898
rect 1386 888 1393 891
rect 1450 888 1486 891
rect 1490 888 1694 891
rect -26 878 6 881
rect 90 878 166 881
rect 226 878 262 881
rect 410 878 446 881
rect 450 878 470 881
rect 474 878 582 881
rect 586 878 622 881
rect 698 878 726 881
rect 738 878 774 881
rect 906 878 926 881
rect 970 878 1062 881
rect 1074 878 1102 881
rect 1162 878 1214 881
rect 1218 878 1222 881
rect 1238 878 1246 881
rect 1258 878 1310 881
rect 1386 878 1414 881
rect 1418 878 1454 881
rect 1458 878 1542 881
rect 1570 878 1598 881
rect 1642 878 1798 881
rect 1826 878 1846 881
rect 162 868 190 871
rect 194 868 254 871
rect 314 868 342 871
rect 546 868 566 871
rect 594 868 614 871
rect 658 868 710 871
rect 834 868 902 871
rect 962 868 982 871
rect 994 868 1078 871
rect 1098 868 1110 871
rect 1162 868 1206 871
rect 1210 868 1214 871
rect 1226 868 1278 871
rect 1290 868 1358 871
rect 1386 868 1526 871
rect 1578 868 1614 871
rect 1634 868 1662 871
rect 1722 868 1806 871
rect 1818 868 1822 871
rect 1834 868 1838 871
rect -26 858 102 861
rect 218 858 230 861
rect 314 858 406 861
rect 418 858 470 861
rect 674 858 686 861
rect 746 858 750 861
rect 826 858 838 861
rect 850 858 934 861
rect 1130 858 1142 861
rect 1234 858 1238 861
rect 1258 858 1326 861
rect 1330 858 1406 861
rect 1594 858 1638 861
rect 1650 858 1774 861
rect 1778 858 1830 861
rect 1834 858 1838 861
rect 706 848 974 851
rect 1186 848 1350 851
rect 1354 848 1518 851
rect 1682 848 1822 851
rect 402 838 414 841
rect 418 838 502 841
rect 506 838 622 841
rect 722 838 750 841
rect 1602 838 1750 841
rect 442 828 454 831
rect 514 828 598 831
rect 602 828 790 831
rect 810 828 862 831
rect 866 828 902 831
rect 906 828 1062 831
rect 354 818 1118 821
rect 426 808 494 811
rect 690 808 1350 811
rect 1018 798 1262 801
rect 178 788 238 791
rect 274 788 334 791
rect 642 788 1254 791
rect -26 778 6 781
rect 346 778 350 781
rect 650 778 758 781
rect 946 778 1126 781
rect 362 768 374 771
rect 1082 768 1270 771
rect 1450 768 1502 771
rect 1610 768 1662 771
rect 1666 768 1734 771
rect 1738 768 1790 771
rect -26 758 190 761
rect 458 758 574 761
rect 1074 758 1086 761
rect 1094 758 1102 761
rect 1346 758 1390 761
rect 1410 758 1622 761
rect 1626 758 1654 761
rect 194 748 214 751
rect 258 748 270 751
rect 322 748 326 751
rect 386 748 430 751
rect 450 748 510 751
rect 818 748 830 751
rect 834 748 894 751
rect 914 748 1166 751
rect 1202 748 1222 751
rect 1242 748 1270 751
rect 1274 748 1334 751
rect 1370 748 1414 751
rect 1450 748 1454 751
rect 1562 748 1582 751
rect 1586 748 1606 751
rect 1626 748 1670 751
rect 1738 748 1750 751
rect 1818 748 1830 751
rect 170 738 222 741
rect 266 738 358 741
rect 370 738 470 741
rect 490 738 526 741
rect 554 738 590 741
rect 666 738 686 741
rect 690 738 750 741
rect 794 738 822 741
rect 866 738 886 741
rect 898 738 974 741
rect 986 738 990 741
rect 1066 738 1086 741
rect 1106 738 1110 741
rect 1146 738 1238 741
rect 1250 738 1294 741
rect 1306 738 1382 741
rect 1386 738 1430 741
rect 1450 738 1454 741
rect 1578 738 1742 741
rect 1746 738 1774 741
rect 1778 738 1862 741
rect 638 732 641 738
rect 822 732 825 738
rect 66 728 86 731
rect 170 728 198 731
rect 210 728 230 731
rect 250 728 526 731
rect 530 728 542 731
rect 618 728 630 731
rect 786 728 806 731
rect 986 728 1078 731
rect 1162 728 1318 731
rect 1322 728 1342 731
rect 1506 728 1558 731
rect 1562 728 1590 731
rect 1594 728 1598 731
rect 1658 728 1694 731
rect 1698 728 1822 731
rect 1842 728 1854 731
rect 738 718 838 721
rect 1050 718 1062 721
rect 1122 718 1302 721
rect 1530 718 1686 721
rect 1690 718 1718 721
rect 1730 718 1742 721
rect 1746 718 1766 721
rect 1770 718 1774 721
rect 1818 718 1830 721
rect 1850 718 1854 721
rect 458 708 462 711
rect 650 708 654 711
rect 826 708 1214 711
rect 1218 708 1230 711
rect 1466 708 1542 711
rect 1546 708 1590 711
rect 1594 708 1846 711
rect 418 698 670 701
rect 698 698 822 701
rect 946 698 1078 701
rect 1138 698 1182 701
rect 1290 698 1294 701
rect 1298 698 1406 701
rect 1586 698 1718 701
rect 1722 698 1766 701
rect 170 688 198 691
rect 298 688 414 691
rect 554 688 654 691
rect 754 688 774 691
rect 914 688 921 691
rect 1018 688 1510 691
rect 1514 688 1678 691
rect 114 678 206 681
rect 234 678 270 681
rect 394 678 406 681
rect 426 678 454 681
rect 466 678 518 681
rect 586 678 614 681
rect 618 678 694 681
rect 714 678 830 681
rect 834 678 862 681
rect 914 678 942 681
rect 958 681 961 688
rect 954 678 1046 681
rect 1146 678 1198 681
rect 1202 678 1342 681
rect 1594 678 1662 681
rect 1698 678 1726 681
rect 1730 678 1742 681
rect 1762 678 1790 681
rect 1858 678 1870 681
rect 878 672 881 678
rect 82 668 142 671
rect 170 668 190 671
rect 202 668 238 671
rect 522 668 558 671
rect 562 668 574 671
rect 706 668 750 671
rect 762 668 798 671
rect 802 668 830 671
rect 938 668 942 671
rect 978 668 985 671
rect 994 668 1001 671
rect 1010 668 1022 671
rect 1074 668 1142 671
rect 1154 668 1230 671
rect 1242 668 1262 671
rect 1354 668 1382 671
rect 1386 668 1481 671
rect 1498 668 1502 671
rect 1514 668 1542 671
rect 1570 668 1590 671
rect 1690 668 1718 671
rect 302 662 305 668
rect -26 658 6 661
rect 106 658 126 661
rect 226 658 238 661
rect 250 658 297 661
rect 354 658 390 661
rect 394 658 430 661
rect 458 658 494 661
rect 626 658 662 661
rect 666 658 718 661
rect 794 658 838 661
rect 882 658 966 661
rect 970 658 1014 661
rect 1026 658 1038 661
rect 1098 658 1118 661
rect 1426 658 1462 661
rect 1466 658 1470 661
rect 1478 661 1481 668
rect 1478 658 1574 661
rect 1658 658 1702 661
rect 266 648 286 651
rect 294 651 297 658
rect 294 648 334 651
rect 434 648 542 651
rect 642 648 790 651
rect 858 648 902 651
rect 1026 648 1030 651
rect 1042 648 1046 651
rect 1146 648 1350 651
rect 1402 648 1414 651
rect 1418 648 1446 651
rect 1466 648 1638 651
rect 418 638 918 641
rect 922 638 966 641
rect 970 638 1054 641
rect 1066 638 1174 641
rect 1178 638 1286 641
rect 1298 638 1566 641
rect 1570 638 1734 641
rect 122 628 438 631
rect 682 628 710 631
rect 898 628 1254 631
rect 1274 628 1598 631
rect 1634 628 1814 631
rect 42 618 310 621
rect 314 618 390 621
rect 394 618 542 621
rect 546 618 614 621
rect 834 618 1046 621
rect 1170 618 1374 621
rect 1482 618 1489 621
rect 1538 618 1542 621
rect 250 608 710 611
rect 930 608 1246 611
rect 1258 608 1542 611
rect 1546 608 1686 611
rect 82 598 1398 601
rect 498 588 558 591
rect 978 588 1206 591
rect 1250 588 1422 591
rect 1722 588 1766 591
rect 98 578 110 581
rect 490 578 510 581
rect 610 578 894 581
rect 1114 578 1150 581
rect 1158 578 1326 581
rect 1386 578 1630 581
rect 378 568 478 571
rect 674 568 694 571
rect 986 568 998 571
rect 1158 571 1161 578
rect 1822 572 1825 578
rect 1122 568 1161 571
rect 1210 568 1398 571
rect 1402 568 1438 571
rect 1442 568 1454 571
rect -26 558 6 561
rect 50 558 70 561
rect 106 558 214 561
rect 370 558 398 561
rect 410 558 590 561
rect 642 558 654 561
rect 658 558 1030 561
rect 1034 558 1206 561
rect 1258 558 1310 561
rect 1314 558 1518 561
rect 1626 558 1686 561
rect 1690 558 1734 561
rect 1834 558 1862 561
rect 66 548 118 551
rect 122 548 134 551
rect 154 548 166 551
rect 186 548 206 551
rect 370 548 382 551
rect 522 548 558 551
rect 578 548 694 551
rect 706 548 822 551
rect 834 548 934 551
rect 1066 548 1073 551
rect 1202 548 1206 551
rect 1282 548 1342 551
rect 1354 548 1414 551
rect 1418 548 1462 551
rect 1522 548 1550 551
rect 1562 548 1630 551
rect 1698 548 1750 551
rect 1754 548 1782 551
rect 1794 548 1822 551
rect 1826 548 1838 551
rect 1842 548 1870 551
rect 454 542 457 548
rect 90 538 94 541
rect 214 538 222 541
rect 274 538 446 541
rect 506 538 606 541
rect 646 538 678 541
rect 738 538 873 541
rect 882 538 902 541
rect 998 541 1001 548
rect 1654 542 1657 548
rect 994 538 1001 541
rect 1018 538 1022 541
rect 1154 538 1278 541
rect 1346 538 1366 541
rect 1370 538 1438 541
rect 1442 538 1494 541
rect 1626 538 1630 541
rect 1674 538 1702 541
rect 1730 538 1878 541
rect 218 528 238 531
rect 282 528 302 531
rect 346 528 366 531
rect 410 528 462 531
rect 466 528 550 531
rect 646 531 649 538
rect 554 528 649 531
rect 658 528 862 531
rect 870 531 873 538
rect 870 528 966 531
rect 994 528 1022 531
rect 1078 528 1102 531
rect 1126 531 1129 538
rect 1122 528 1129 531
rect 1194 528 1222 531
rect 1322 528 1350 531
rect 1370 528 1390 531
rect 1442 528 1446 531
rect 1490 528 1526 531
rect 1546 528 1574 531
rect 1578 528 1678 531
rect 1738 528 1878 531
rect 370 518 446 521
rect 450 518 526 521
rect 586 518 718 521
rect 874 518 918 521
rect 1078 521 1081 528
rect 986 518 1081 521
rect 1090 518 1230 521
rect 1394 518 1558 521
rect 1610 518 1846 521
rect 378 508 414 511
rect 594 508 622 511
rect 906 508 910 511
rect 1082 508 1134 511
rect 1146 508 1174 511
rect 1178 508 1366 511
rect 1466 508 1502 511
rect 1546 508 1646 511
rect 1650 508 1758 511
rect 1762 508 1814 511
rect 626 498 670 501
rect 818 498 1062 501
rect 1090 498 1126 501
rect 1134 498 1214 501
rect 1330 498 1334 501
rect 1338 498 1438 501
rect 1450 498 1590 501
rect 1722 498 1798 501
rect 1802 498 1838 501
rect 530 488 766 491
rect 850 488 942 491
rect 1134 491 1137 498
rect 1058 488 1137 491
rect 1154 488 1558 491
rect 1578 488 1582 491
rect 1634 488 1814 491
rect 462 482 465 488
rect -26 478 30 481
rect 66 478 94 481
rect 154 478 174 481
rect 178 478 222 481
rect 242 478 254 481
rect 314 478 342 481
rect 682 478 750 481
rect 770 478 846 481
rect 850 478 878 481
rect 938 478 958 481
rect 962 478 1014 481
rect 1018 478 1086 481
rect 1098 478 1278 481
rect 1474 478 1510 481
rect 1570 478 1670 481
rect 1706 478 1726 481
rect 1754 478 1758 481
rect 34 468 70 471
rect 218 468 254 471
rect 266 468 286 471
rect 306 468 310 471
rect 334 468 342 471
rect 442 468 470 471
rect 506 468 558 471
rect 602 468 694 471
rect 714 468 742 471
rect 758 468 766 471
rect 874 468 886 471
rect 898 468 1110 471
rect 1170 468 1206 471
rect 1266 468 1294 471
rect 1410 468 1430 471
rect 1498 468 1526 471
rect 1530 468 1686 471
rect 1722 468 1862 471
rect 334 462 337 468
rect -26 458 6 461
rect 26 458 118 461
rect 202 458 318 461
rect 490 458 502 461
rect 538 458 606 461
rect 626 458 670 461
rect 682 458 726 461
rect 794 458 798 461
rect 882 458 990 461
rect 1178 458 1198 461
rect 1234 458 1254 461
rect 1298 458 1390 461
rect 1442 458 1478 461
rect 1634 458 1638 461
rect 1754 458 1798 461
rect 1802 458 1806 461
rect 178 448 190 451
rect 522 448 622 451
rect 626 448 670 451
rect 746 448 854 451
rect 962 448 1030 451
rect 1050 448 1310 451
rect 1314 448 1454 451
rect 1458 448 1462 451
rect 1506 448 1558 451
rect 1562 448 1830 451
rect 50 438 62 441
rect 458 438 502 441
rect 842 438 1382 441
rect 410 428 574 431
rect 762 428 974 431
rect 978 428 1006 431
rect 1010 428 1014 431
rect 1018 428 1086 431
rect 1090 428 1110 431
rect 1122 428 1414 431
rect 90 418 174 421
rect 178 418 222 421
rect 226 418 414 421
rect 418 418 534 421
rect 554 418 678 421
rect 818 418 1190 421
rect 1194 418 1446 421
rect 114 408 150 411
rect 346 408 406 411
rect 426 408 502 411
rect 930 408 1238 411
rect 1250 408 1406 411
rect 1418 408 1542 411
rect 674 398 686 401
rect 906 398 998 401
rect 1026 398 1182 401
rect 1202 398 1502 401
rect 1830 392 1833 398
rect 162 388 342 391
rect 346 388 518 391
rect 570 388 590 391
rect 1082 388 1142 391
rect 1146 388 1150 391
rect 1194 388 1662 391
rect 1666 388 1702 391
rect 386 378 414 381
rect 514 378 638 381
rect 642 378 886 381
rect 962 378 982 381
rect 986 378 1190 381
rect 1354 378 1390 381
rect 106 368 182 371
rect 186 368 302 371
rect 362 368 382 371
rect 442 368 510 371
rect 546 368 758 371
rect 810 368 822 371
rect 826 368 1102 371
rect 1106 368 1358 371
rect 1362 368 1374 371
rect 1378 368 1390 371
rect 1570 368 1582 371
rect 1586 368 1614 371
rect 1842 368 1854 371
rect 450 358 761 361
rect 766 358 769 368
rect 994 358 1094 361
rect 1114 358 1278 361
rect 1290 358 1334 361
rect 1362 358 1430 361
rect 1434 358 1518 361
rect 1530 358 1558 361
rect 1570 358 1686 361
rect 146 348 158 351
rect 426 348 438 351
rect 466 348 502 351
rect 506 348 622 351
rect 678 348 726 351
rect 758 351 761 358
rect 758 348 854 351
rect 906 348 942 351
rect 946 348 950 351
rect 962 348 990 351
rect 1082 348 1198 351
rect 1226 348 1446 351
rect 1450 348 1545 351
rect 1610 348 1622 351
rect -26 338 6 341
rect 10 338 54 341
rect 98 338 110 341
rect 250 338 278 341
rect 314 338 326 341
rect 330 338 374 341
rect 678 341 681 348
rect 1014 342 1017 348
rect 546 338 681 341
rect 690 338 694 341
rect 730 338 838 341
rect 850 338 878 341
rect 938 338 966 341
rect 1050 338 1070 341
rect 1090 338 1118 341
rect 1210 338 1230 341
rect 1234 338 1246 341
rect 1250 338 1366 341
rect 1370 338 1494 341
rect 1498 338 1534 341
rect 1542 341 1545 348
rect 1542 338 1646 341
rect 1714 338 1721 341
rect 354 328 366 331
rect 698 328 702 331
rect 750 328 758 331
rect 842 328 990 331
rect 1026 328 1222 331
rect 1274 328 1646 331
rect 1714 328 1726 331
rect 1746 328 1806 331
rect 34 318 54 321
rect 138 318 430 321
rect 610 318 622 321
rect 658 318 670 321
rect 722 318 902 321
rect 914 318 1046 321
rect 1098 318 1150 321
rect 1362 318 1398 321
rect 1402 318 1422 321
rect 1450 318 1462 321
rect 1594 318 1606 321
rect 1626 318 1798 321
rect 1810 318 1886 321
rect 394 308 446 311
rect 498 308 526 311
rect 546 308 822 311
rect 826 308 1030 311
rect 1034 308 1278 311
rect 1354 308 1398 311
rect 1490 308 1534 311
rect 1538 308 1622 311
rect 1802 308 1814 311
rect 186 298 222 301
rect 226 298 1142 301
rect 1490 298 1574 301
rect 1762 298 1830 301
rect 74 288 126 291
rect 154 288 222 291
rect 226 288 254 291
rect 266 288 662 291
rect 858 288 1054 291
rect 1058 288 1302 291
rect 1330 288 1478 291
rect 1514 288 1534 291
rect 1538 288 1550 291
rect 1650 288 1726 291
rect 846 282 849 288
rect 106 278 166 281
rect 202 278 214 281
rect 362 278 638 281
rect 794 278 806 281
rect 850 278 878 281
rect 906 278 913 281
rect 1010 278 1014 281
rect 1138 278 1174 281
rect 1178 278 1230 281
rect 1234 278 1302 281
rect 1314 278 1390 281
rect 1402 278 1510 281
rect 1522 278 1526 281
rect 1554 278 1574 281
rect 1618 278 1702 281
rect 1706 278 1750 281
rect 1810 278 1830 281
rect 886 272 889 278
rect 194 268 254 271
rect 274 268 286 271
rect 306 268 334 271
rect 410 268 574 271
rect 578 268 758 271
rect 762 268 830 271
rect 934 271 937 278
rect 934 268 1022 271
rect 1090 268 1102 271
rect 1146 268 1166 271
rect 1242 268 1286 271
rect 1290 268 1297 271
rect 1306 268 1406 271
rect 1410 268 1622 271
rect 1698 268 1710 271
rect 1730 268 1742 271
rect 1770 268 1782 271
rect -26 258 6 261
rect 50 258 86 261
rect 114 258 126 261
rect 170 258 214 261
rect 242 258 262 261
rect 394 258 414 261
rect 466 258 561 261
rect 570 258 646 261
rect 682 258 694 261
rect 778 258 798 261
rect 802 258 806 261
rect 834 258 1126 261
rect 1130 258 1182 261
rect 1194 258 1214 261
rect 1226 258 1246 261
rect 1266 258 1310 261
rect 1330 258 1454 261
rect 1458 258 1558 261
rect 1562 258 1694 261
rect 1834 258 1846 261
rect 1890 258 1913 261
rect 162 248 198 251
rect 362 248 438 251
rect 442 248 462 251
rect 478 248 486 251
rect 514 248 550 251
rect 558 251 561 258
rect 558 248 686 251
rect 746 248 774 251
rect 1026 248 1086 251
rect 1090 248 1118 251
rect 1170 248 1590 251
rect 234 238 494 241
rect 498 238 1046 241
rect 1330 238 1494 241
rect 1546 238 1678 241
rect 74 228 182 231
rect 386 228 398 231
rect 522 228 718 231
rect 842 228 1062 231
rect 1066 228 1398 231
rect 1402 228 1758 231
rect 314 218 342 221
rect 346 218 478 221
rect 570 218 574 221
rect 618 218 686 221
rect 698 218 782 221
rect 818 218 830 221
rect 874 218 910 221
rect 994 218 1070 221
rect 1386 218 1422 221
rect 1426 218 1430 221
rect 1450 218 1574 221
rect 1578 218 1646 221
rect 338 208 502 211
rect 746 208 886 211
rect 906 208 1414 211
rect 450 198 526 201
rect 674 198 790 201
rect 1058 198 1142 201
rect 1482 198 1590 201
rect 1602 198 1742 201
rect 146 188 174 191
rect 378 188 518 191
rect 698 188 910 191
rect 914 188 998 191
rect 1002 188 1030 191
rect 1034 188 1086 191
rect 1098 188 1350 191
rect 1394 188 1494 191
rect 1746 188 1766 191
rect 1842 188 1854 191
rect 570 178 598 181
rect 610 178 718 181
rect 722 178 1446 181
rect 1538 178 1670 181
rect 82 168 102 171
rect 106 168 230 171
rect 346 168 622 171
rect 762 168 798 171
rect 930 168 1094 171
rect 1154 168 1190 171
rect 1202 168 1214 171
rect 1218 168 1342 171
rect 1410 168 1550 171
rect 1802 168 1846 171
rect -26 158 54 161
rect 282 158 414 161
rect 418 158 438 161
rect 522 158 558 161
rect 562 158 622 161
rect 642 158 766 161
rect 1018 158 1134 161
rect 1146 158 1198 161
rect 1210 158 1390 161
rect 1422 158 1574 161
rect 1610 158 1742 161
rect 1794 158 1814 161
rect 1826 158 1854 161
rect 222 152 225 158
rect 82 148 150 151
rect 322 148 350 151
rect 354 148 358 151
rect 362 148 382 151
rect 426 148 446 151
rect 490 148 502 151
rect 530 148 670 151
rect 682 148 918 151
rect 962 148 982 151
rect 1082 148 1182 151
rect 1186 148 1206 151
rect 1322 148 1358 151
rect 1422 151 1425 158
rect 1370 148 1425 151
rect 1434 148 1446 151
rect 1514 148 1558 151
rect 1626 148 1702 151
rect 1706 148 1782 151
rect 1818 148 1822 151
rect -26 138 6 141
rect 58 138 94 141
rect 194 138 286 141
rect 306 138 342 141
rect 386 138 454 141
rect 498 138 502 141
rect 658 138 806 141
rect 810 138 854 141
rect 906 138 934 141
rect 1098 138 1110 141
rect 1234 138 1278 141
rect 1314 138 1326 141
rect 1346 138 1374 141
rect 1410 138 1470 141
rect 1522 138 1606 141
rect 1610 138 1718 141
rect 1762 138 1774 141
rect 74 128 110 131
rect 138 128 158 131
rect 170 128 246 131
rect 258 128 518 131
rect 618 128 646 131
rect 666 128 726 131
rect 754 128 774 131
rect 786 128 822 131
rect 1130 128 1222 131
rect 1250 128 1318 131
rect 1362 128 1478 131
rect 1538 128 1622 131
rect 1650 128 1734 131
rect 50 118 62 121
rect 186 118 278 121
rect 282 118 326 121
rect 330 118 350 121
rect 418 118 430 121
rect 434 118 486 121
rect 538 118 654 121
rect 722 118 726 121
rect 794 118 985 121
rect 1010 118 1038 121
rect 1066 118 1262 121
rect 1266 118 1510 121
rect 1666 118 1806 121
rect 34 108 54 111
rect 250 108 310 111
rect 314 108 470 111
rect 474 108 766 111
rect 802 108 822 111
rect 850 108 902 111
rect 982 111 985 118
rect 982 108 1190 111
rect 1194 108 1238 111
rect 1242 108 1254 111
rect 1282 108 1294 111
rect 1442 108 1454 111
rect 146 98 182 101
rect 202 98 246 101
rect 266 98 374 101
rect 466 98 638 101
rect 658 98 838 101
rect 858 98 878 101
rect 882 98 894 101
rect 898 98 1534 101
rect 1650 98 1670 101
rect 1674 98 1766 101
rect 10 88 86 91
rect 90 88 198 91
rect 546 88 614 91
rect 618 88 846 91
rect 850 88 1014 91
rect 1018 88 1038 91
rect 1050 88 1102 91
rect 1106 88 1206 91
rect 1370 88 1438 91
rect 1562 88 1670 91
rect 1810 88 1822 91
rect 1834 88 1838 91
rect 98 78 102 81
rect 106 78 214 81
rect 322 78 406 81
rect 410 78 422 81
rect 426 78 502 81
rect 554 78 670 81
rect 730 78 966 81
rect 986 78 998 81
rect 1090 78 1126 81
rect 1298 78 1358 81
rect 1474 78 1534 81
rect 1594 78 1622 81
rect 1642 78 1750 81
rect 1762 78 1782 81
rect 214 72 217 78
rect 718 72 721 78
rect 1846 72 1849 78
rect 66 68 190 71
rect 226 68 270 71
rect 394 68 494 71
rect 674 68 694 71
rect 794 68 830 71
rect 930 68 958 71
rect 1002 68 1142 71
rect 1154 68 1190 71
rect 1250 68 1342 71
rect 1378 68 1414 71
rect 1466 68 1473 71
rect 1490 68 1654 71
rect 1698 68 1774 71
rect 910 62 913 68
rect -26 58 6 61
rect 82 58 150 61
rect 178 58 318 61
rect 402 58 446 61
rect 666 58 686 61
rect 690 58 710 61
rect 770 58 798 61
rect 1034 58 1046 61
rect 1058 58 1086 61
rect 1154 58 1278 61
rect 1330 58 1350 61
rect 1354 58 1486 61
rect 1506 58 1526 61
rect 1530 58 1558 61
rect 1562 58 1678 61
rect 1682 58 1702 61
rect 1826 58 1878 61
rect 122 48 342 51
rect 370 48 398 51
rect 602 48 702 51
rect 826 48 886 51
rect 954 48 1334 51
rect 1346 48 1390 51
rect 1594 48 1601 51
rect 866 38 870 41
rect 874 38 878 41
rect 1226 38 1230 41
rect 1234 38 1334 41
rect 786 28 870 31
rect 1210 28 1214 31
rect 1218 28 1254 31
rect 490 8 526 11
rect 954 8 966 11
rect 970 8 1054 11
rect 1202 8 1214 11
rect 1258 8 1326 11
<< m4contact >>
rect 622 1208 626 1212
rect 1222 1168 1226 1172
rect 582 1158 586 1162
rect 278 1148 282 1152
rect 414 1148 418 1152
rect 558 1148 562 1152
rect 582 1148 586 1152
rect 686 1148 690 1152
rect 278 1138 282 1142
rect 1222 1138 1226 1142
rect 1830 1138 1834 1142
rect 1502 1128 1506 1132
rect 1606 1128 1610 1132
rect 286 1118 290 1122
rect 542 1118 546 1122
rect 582 1108 586 1112
rect 622 1108 626 1112
rect 1222 1108 1226 1112
rect 518 1098 522 1102
rect 662 1098 666 1102
rect 1262 1098 1266 1102
rect 1374 1098 1378 1102
rect 1534 1078 1538 1082
rect 1750 1078 1754 1082
rect 254 1068 258 1072
rect 262 1068 266 1072
rect 990 1068 994 1072
rect 998 1068 1002 1072
rect 1134 1068 1138 1072
rect 622 1058 626 1062
rect 654 1058 658 1062
rect 678 1058 682 1062
rect 686 1058 690 1062
rect 806 1058 810 1062
rect 1118 1058 1122 1062
rect 1326 1058 1330 1062
rect 1406 1058 1410 1062
rect 1438 1058 1442 1062
rect 1446 1058 1450 1062
rect 1494 1058 1498 1062
rect 1502 1058 1506 1062
rect 1654 1058 1658 1062
rect 262 1048 266 1052
rect 1230 1038 1234 1042
rect 830 1028 834 1032
rect 1190 1028 1194 1032
rect 1534 1028 1538 1032
rect 286 1018 290 1022
rect 798 1018 802 1022
rect 462 1008 466 1012
rect 1254 1008 1258 1012
rect 278 998 282 1002
rect 582 998 586 1002
rect 1830 998 1834 1002
rect 1822 988 1826 992
rect 790 978 794 982
rect 654 958 658 962
rect 966 948 970 952
rect 1590 948 1594 952
rect 1606 948 1610 952
rect 1734 948 1738 952
rect 262 938 266 942
rect 526 938 530 942
rect 1174 938 1178 942
rect 94 928 98 932
rect 342 928 346 932
rect 662 928 666 932
rect 758 928 762 932
rect 1222 928 1226 932
rect 1302 928 1306 932
rect 614 918 618 922
rect 1174 918 1178 922
rect 1326 918 1330 922
rect 1350 918 1354 922
rect 1358 918 1362 922
rect 766 908 770 912
rect 1510 898 1514 902
rect 1190 888 1194 892
rect 1382 888 1386 892
rect 582 878 586 882
rect 1214 878 1218 882
rect 1246 878 1250 882
rect 1822 878 1826 882
rect 982 868 986 872
rect 1110 868 1114 872
rect 1206 868 1210 872
rect 1822 868 1826 872
rect 1830 868 1834 872
rect 406 858 410 862
rect 750 858 754 862
rect 846 858 850 862
rect 1230 858 1234 862
rect 1822 848 1826 852
rect 718 838 722 842
rect 1750 838 1754 842
rect 1350 808 1354 812
rect 1262 798 1266 802
rect 638 788 642 792
rect 342 778 346 782
rect 1502 768 1506 772
rect 1790 768 1794 772
rect 1102 758 1106 762
rect 1118 758 1122 762
rect 326 748 330 752
rect 1454 748 1458 752
rect 1734 748 1738 752
rect 1814 748 1818 752
rect 358 738 362 742
rect 638 738 642 742
rect 822 738 826 742
rect 974 738 978 742
rect 982 738 986 742
rect 1110 738 1114 742
rect 1302 738 1306 742
rect 1446 738 1450 742
rect 542 728 546 732
rect 1654 728 1658 732
rect 1838 728 1842 732
rect 1718 718 1722 722
rect 1742 718 1746 722
rect 1846 718 1850 722
rect 158 708 162 712
rect 454 708 458 712
rect 654 708 658 712
rect 1214 708 1218 712
rect 1590 708 1594 712
rect 414 698 418 702
rect 1582 698 1586 702
rect 414 688 418 692
rect 910 688 914 692
rect 1014 688 1018 692
rect 878 678 882 682
rect 1494 678 1498 682
rect 1854 678 1858 682
rect 302 668 306 672
rect 358 668 362 672
rect 750 668 754 672
rect 942 668 946 672
rect 974 668 978 672
rect 990 668 994 672
rect 1006 668 1010 672
rect 1150 668 1154 672
rect 1238 668 1242 672
rect 1502 668 1506 672
rect 238 658 242 662
rect 718 658 722 662
rect 838 658 842 662
rect 1022 658 1026 662
rect 1118 658 1122 662
rect 1190 658 1194 662
rect 1030 648 1034 652
rect 1038 648 1042 652
rect 1462 648 1466 652
rect 414 638 418 642
rect 966 638 970 642
rect 1294 638 1298 642
rect 1254 628 1258 632
rect 390 618 394 622
rect 614 618 618 622
rect 830 618 834 622
rect 1478 618 1482 622
rect 1534 618 1538 622
rect 1246 608 1250 612
rect 94 578 98 582
rect 1110 578 1114 582
rect 1822 578 1826 582
rect 870 568 874 572
rect 998 568 1002 572
rect 406 558 410 562
rect 694 548 698 552
rect 998 548 1002 552
rect 1062 548 1066 552
rect 1206 548 1210 552
rect 1350 548 1354 552
rect 1558 548 1562 552
rect 1654 548 1658 552
rect 1822 548 1826 552
rect 86 538 90 542
rect 222 538 226 542
rect 446 538 450 542
rect 454 538 458 542
rect 606 538 610 542
rect 1014 538 1018 542
rect 1630 538 1634 542
rect 1670 538 1674 542
rect 1726 538 1730 542
rect 1438 528 1442 532
rect 1542 528 1546 532
rect 1734 528 1738 532
rect 1558 518 1562 522
rect 414 508 418 512
rect 902 508 906 512
rect 1142 508 1146 512
rect 1814 508 1818 512
rect 1438 498 1442 502
rect 1446 498 1450 502
rect 1718 498 1722 502
rect 1798 498 1802 502
rect 1150 488 1154 492
rect 1582 488 1586 492
rect 462 478 466 482
rect 846 478 850 482
rect 886 478 890 482
rect 1014 478 1018 482
rect 1670 478 1674 482
rect 1758 478 1762 482
rect 302 468 306 472
rect 342 468 346 472
rect 694 468 698 472
rect 742 468 746 472
rect 766 468 770 472
rect 870 468 874 472
rect 894 468 898 472
rect 622 458 626 462
rect 790 458 794 462
rect 1630 458 1634 462
rect 1806 458 1810 462
rect 670 448 674 452
rect 1454 448 1458 452
rect 1558 448 1562 452
rect 838 438 842 442
rect 1110 428 1114 432
rect 86 418 90 422
rect 174 418 178 422
rect 678 418 682 422
rect 1190 418 1194 422
rect 1406 408 1410 412
rect 1542 408 1546 412
rect 158 388 162 392
rect 1150 388 1154 392
rect 1830 388 1834 392
rect 302 368 306 372
rect 390 368 394 372
rect 766 368 770 372
rect 822 368 826 372
rect 78 358 82 362
rect 126 358 130 362
rect 1094 358 1098 362
rect 1278 358 1282 362
rect 1286 358 1290 362
rect 1518 358 1522 362
rect 1566 358 1570 362
rect 870 348 874 352
rect 902 348 906 352
rect 950 348 954 352
rect 990 348 994 352
rect 1078 348 1082 352
rect 1558 348 1562 352
rect 686 338 690 342
rect 838 338 842 342
rect 1014 338 1018 342
rect 1710 338 1714 342
rect 694 328 698 332
rect 758 328 762 332
rect 1726 328 1730 332
rect 902 318 906 322
rect 1094 318 1098 322
rect 494 308 498 312
rect 222 298 226 302
rect 1142 298 1146 302
rect 1278 298 1282 302
rect 254 288 258 292
rect 854 288 858 292
rect 1534 288 1538 292
rect 342 278 346 282
rect 358 278 362 282
rect 846 278 850 282
rect 902 278 906 282
rect 1006 278 1010 282
rect 1518 278 1522 282
rect 1806 278 1810 282
rect 886 268 890 272
rect 1286 268 1290 272
rect 1742 268 1746 272
rect 1750 268 1754 272
rect 126 258 130 262
rect 566 258 570 262
rect 654 258 658 262
rect 806 258 810 262
rect 1190 258 1194 262
rect 1222 258 1226 262
rect 1326 258 1330 262
rect 486 248 490 252
rect 1046 238 1050 242
rect 70 228 74 232
rect 1758 228 1762 232
rect 574 218 578 222
rect 694 218 698 222
rect 1430 218 1434 222
rect 1630 208 1634 212
rect 670 198 674 202
rect 910 188 914 192
rect 1086 188 1090 192
rect 1094 188 1098 192
rect 1854 188 1858 192
rect 718 178 722 182
rect 78 168 82 172
rect 1094 168 1098 172
rect 1406 168 1410 172
rect 1798 168 1802 172
rect 62 158 66 162
rect 622 158 626 162
rect 1790 158 1794 162
rect 222 148 226 152
rect 678 148 682 152
rect 1358 148 1362 152
rect 1814 148 1818 152
rect 342 138 346 142
rect 494 138 498 142
rect 1358 128 1362 132
rect 174 118 178 122
rect 654 118 658 122
rect 726 118 730 122
rect 70 108 74 112
rect 654 98 658 102
rect 1046 88 1050 92
rect 1366 88 1370 92
rect 1558 88 1562 92
rect 1822 88 1826 92
rect 1838 88 1842 92
rect 726 78 730 82
rect 1086 78 1090 82
rect 1470 78 1474 82
rect 62 68 66 72
rect 214 68 218 72
rect 222 68 226 72
rect 670 68 674 72
rect 718 68 722 72
rect 1142 68 1146 72
rect 1230 68 1234 72
rect 1366 68 1370 72
rect 1374 68 1378 72
rect 1430 68 1434 72
rect 1462 68 1466 72
rect 1654 68 1658 72
rect 1846 68 1850 72
rect 910 58 914 62
rect 1150 58 1154 62
rect 1334 48 1338 52
rect 1590 48 1594 52
rect 1206 28 1210 32
rect 950 8 954 12
<< metal4 >>
rect 582 1152 585 1158
rect 554 1148 558 1151
rect 278 1142 281 1148
rect 254 1062 257 1068
rect 262 1052 265 1068
rect 278 1002 281 1138
rect 286 1022 289 1118
rect 258 938 262 941
rect 94 582 97 928
rect 342 782 345 928
rect 406 862 409 888
rect 322 748 326 751
rect 86 422 89 538
rect 158 392 161 708
rect 414 702 417 1148
rect 514 1098 518 1101
rect 218 538 222 541
rect 302 492 305 668
rect 302 472 305 488
rect 338 468 342 471
rect 62 72 65 158
rect 70 112 73 228
rect 78 172 81 358
rect 126 262 129 358
rect 174 122 177 418
rect 222 152 225 298
rect 214 72 217 88
rect 222 72 225 148
rect 254 102 257 288
rect 302 282 305 368
rect 358 282 361 668
rect 390 372 393 618
rect 406 542 409 558
rect 414 512 417 638
rect 454 542 457 708
rect 462 482 465 1008
rect 526 932 529 938
rect 542 732 545 1118
rect 582 1112 585 1148
rect 622 1112 625 1208
rect 1222 1142 1225 1168
rect 582 882 585 998
rect 614 622 617 918
rect 606 512 609 538
rect 622 462 625 1058
rect 654 962 657 1058
rect 638 742 641 788
rect 654 712 657 958
rect 662 932 665 1098
rect 686 1062 689 1078
rect 986 1068 990 1071
rect 998 1062 1001 1068
rect 674 1058 678 1061
rect 802 1058 806 1061
rect 798 1022 801 1058
rect 746 858 750 861
rect 718 662 721 838
rect 742 472 745 858
rect 766 482 769 908
rect 762 468 766 471
rect 342 142 345 278
rect 482 248 486 251
rect 494 142 497 308
rect 566 252 569 258
rect 570 218 574 221
rect 622 162 625 458
rect 654 262 657 268
rect 670 202 673 448
rect 622 62 625 158
rect 654 102 657 118
rect 670 72 673 198
rect 678 152 681 418
rect 686 342 689 348
rect 694 332 697 468
rect 790 462 793 978
rect 822 372 825 738
rect 830 622 833 1028
rect 846 862 849 938
rect 914 688 918 691
rect 838 442 841 658
rect 766 358 769 368
rect 834 338 838 341
rect 754 328 758 331
rect 846 282 849 478
rect 870 472 873 568
rect 870 352 873 358
rect 854 292 857 338
rect 878 332 881 678
rect 942 672 945 678
rect 966 642 969 948
rect 982 872 985 898
rect 974 742 977 758
rect 982 742 985 748
rect 978 668 982 671
rect 994 668 998 671
rect 906 508 910 511
rect 886 272 889 478
rect 990 352 993 638
rect 998 572 1001 608
rect 998 542 1001 548
rect 902 322 905 348
rect 906 278 910 281
rect 802 258 806 261
rect 718 72 721 178
rect 726 82 729 118
rect 910 62 913 188
rect 950 12 953 348
rect 1006 282 1009 668
rect 1014 542 1017 688
rect 1026 658 1030 661
rect 1038 652 1041 848
rect 1098 758 1102 761
rect 1110 742 1113 868
rect 1118 762 1121 1058
rect 1174 922 1177 938
rect 1190 892 1193 1028
rect 1222 932 1225 1108
rect 1206 872 1209 878
rect 1118 662 1121 758
rect 1214 712 1217 878
rect 1230 862 1233 1038
rect 1242 878 1246 881
rect 1150 672 1153 678
rect 1026 648 1030 651
rect 1066 548 1070 551
rect 1014 342 1017 478
rect 1110 432 1113 578
rect 1094 322 1097 358
rect 1142 302 1145 508
rect 1150 392 1153 488
rect 1190 422 1193 658
rect 1254 632 1257 1008
rect 1262 802 1265 1098
rect 1326 1062 1329 1068
rect 1502 1062 1505 1128
rect 1402 1058 1406 1061
rect 1438 1052 1441 1058
rect 1494 1052 1497 1058
rect 1534 1032 1537 1078
rect 1606 952 1609 1128
rect 1302 742 1305 928
rect 1326 862 1329 918
rect 1246 612 1249 618
rect 1294 612 1297 638
rect 1046 92 1049 238
rect 1086 82 1089 188
rect 1094 172 1097 188
rect 1154 58 1158 61
rect 1206 32 1209 548
rect 1278 302 1281 358
rect 1286 332 1289 358
rect 1290 268 1294 271
rect 1222 262 1225 268
rect 1326 262 1329 858
rect 1350 812 1353 918
rect 1358 852 1361 918
rect 1514 898 1518 901
rect 1386 888 1390 891
rect 1350 92 1353 548
rect 1442 528 1446 531
rect 1438 502 1441 528
rect 1446 492 1449 498
rect 1454 452 1457 748
rect 1494 642 1497 678
rect 1502 672 1505 768
rect 1590 712 1593 948
rect 1654 732 1657 1058
rect 1830 1002 1833 1138
rect 1734 752 1737 948
rect 1822 882 1825 988
rect 1822 852 1825 868
rect 1482 618 1486 621
rect 1406 172 1409 408
rect 1518 342 1521 358
rect 1534 292 1537 618
rect 1542 412 1545 528
rect 1558 522 1561 548
rect 1582 492 1585 698
rect 1630 532 1633 538
rect 1630 462 1633 528
rect 1558 352 1561 448
rect 1518 272 1521 278
rect 1358 132 1361 148
rect 1366 92 1369 98
rect 1366 72 1369 88
rect 1430 72 1433 218
rect 1558 92 1561 348
rect 1630 212 1633 458
rect 1470 72 1473 78
rect 1654 72 1657 548
rect 1670 482 1673 538
rect 1718 502 1721 718
rect 1714 338 1718 341
rect 1726 332 1729 538
rect 1734 532 1737 748
rect 1742 272 1745 718
rect 1750 272 1753 838
rect 1758 232 1761 478
rect 1790 162 1793 768
rect 1814 512 1817 748
rect 1822 582 1825 848
rect 1798 172 1801 498
rect 1806 282 1809 458
rect 1814 152 1817 508
rect 1822 92 1825 548
rect 1830 392 1833 868
rect 1838 92 1841 728
rect 1846 72 1849 718
rect 1854 192 1857 678
rect 1466 68 1470 71
rect 1230 62 1233 68
rect 1374 62 1377 68
rect 1594 48 1598 51
<< m5contact >>
rect 550 1148 554 1152
rect 254 1058 258 1062
rect 254 938 258 942
rect 406 888 410 892
rect 318 748 322 752
rect 358 738 362 742
rect 510 1098 514 1102
rect 414 688 418 692
rect 238 658 242 662
rect 214 538 218 542
rect 302 488 306 492
rect 334 468 338 472
rect 214 88 218 92
rect 406 538 410 542
rect 446 538 450 542
rect 526 928 530 932
rect 686 1148 690 1152
rect 606 508 610 512
rect 686 1078 690 1082
rect 982 1068 986 1072
rect 1134 1068 1138 1072
rect 670 1058 674 1062
rect 798 1058 802 1062
rect 998 1058 1002 1062
rect 758 928 762 932
rect 742 858 746 862
rect 694 548 698 552
rect 750 668 754 672
rect 766 478 770 482
rect 758 468 762 472
rect 302 278 306 282
rect 478 248 482 252
rect 566 248 570 252
rect 566 218 570 222
rect 654 268 658 272
rect 254 98 258 102
rect 686 348 690 352
rect 846 938 850 942
rect 918 688 922 692
rect 942 678 946 682
rect 766 368 770 372
rect 830 338 834 342
rect 750 328 754 332
rect 870 358 874 362
rect 854 338 858 342
rect 982 898 986 902
rect 1038 848 1042 852
rect 974 758 978 762
rect 982 748 986 752
rect 982 668 986 672
rect 998 668 1002 672
rect 990 638 994 642
rect 910 508 914 512
rect 878 328 882 332
rect 894 468 898 472
rect 998 608 1002 612
rect 998 538 1002 542
rect 910 278 914 282
rect 798 258 802 262
rect 694 218 698 222
rect 622 58 626 62
rect 1030 658 1034 662
rect 1094 758 1098 762
rect 1374 1098 1378 1102
rect 1206 878 1210 882
rect 1238 878 1242 882
rect 1150 678 1154 682
rect 1238 668 1242 672
rect 1022 648 1026 652
rect 1070 548 1074 552
rect 1078 348 1082 352
rect 1326 1068 1330 1072
rect 1398 1058 1402 1062
rect 1446 1058 1450 1062
rect 1438 1048 1442 1052
rect 1494 1048 1498 1052
rect 1750 1078 1754 1082
rect 1326 858 1330 862
rect 1246 618 1250 622
rect 1294 608 1298 612
rect 1190 258 1194 262
rect 1142 68 1146 72
rect 1158 58 1162 62
rect 1286 328 1290 332
rect 1222 268 1226 272
rect 1294 268 1298 272
rect 1518 898 1522 902
rect 1390 888 1394 892
rect 1358 848 1362 852
rect 1446 738 1450 742
rect 1446 528 1450 532
rect 1446 488 1450 492
rect 1462 648 1466 652
rect 1494 638 1498 642
rect 1486 618 1490 622
rect 1518 338 1522 342
rect 1630 528 1634 532
rect 1566 358 1570 362
rect 1518 268 1522 272
rect 1366 98 1370 102
rect 1350 88 1354 92
rect 1718 338 1722 342
rect 1470 68 1474 72
rect 1230 58 1234 62
rect 1374 58 1378 62
rect 1334 48 1338 52
rect 1598 48 1602 52
<< metal5 >>
rect 554 1148 686 1151
rect 514 1098 1374 1101
rect 690 1078 1750 1081
rect 986 1068 1134 1071
rect 1138 1068 1326 1071
rect 258 1058 670 1061
rect 802 1058 998 1061
rect 1402 1058 1446 1061
rect 1442 1048 1494 1051
rect 258 938 846 941
rect 530 928 758 931
rect 986 898 1518 901
rect 410 888 1390 891
rect 1210 878 1238 881
rect 746 858 1326 861
rect 1042 848 1358 851
rect 978 758 1094 761
rect 322 748 982 751
rect 362 738 1446 741
rect 418 688 918 691
rect 946 678 1150 681
rect 754 668 982 671
rect 1002 668 1238 671
rect 242 658 1030 661
rect 1026 648 1462 651
rect 994 638 1494 641
rect 1250 618 1486 621
rect 1002 608 1294 611
rect 698 548 1070 551
rect 218 538 406 541
rect 450 538 998 541
rect 1450 528 1630 531
rect 610 508 910 511
rect 306 488 1446 491
rect 338 468 758 471
rect 762 468 894 471
rect 766 362 769 368
rect 874 358 1566 361
rect 690 348 1078 351
rect 834 338 854 341
rect 1522 338 1718 341
rect 754 328 878 331
rect 882 328 1286 331
rect 306 278 910 281
rect 658 268 1222 271
rect 1298 268 1518 271
rect 802 258 1190 261
rect 482 248 566 251
rect 570 218 694 221
rect 258 98 1366 101
rect 218 88 1350 91
rect 1146 68 1470 71
rect 626 58 1158 61
rect 1234 58 1374 61
rect 1338 48 1598 51
<< m6contact >>
rect 765 478 766 482
rect 766 478 770 482
rect 765 477 770 478
rect 765 357 770 362
<< metal6 >>
rect 765 362 770 477
use BUFX2  BUFX2_70
timestamp 1514851247
transform -1 0 28 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_47
timestamp 1514851247
transform -1 0 52 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_68
timestamp 1514851247
transform -1 0 76 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_45
timestamp 1514851247
transform -1 0 100 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_53
timestamp 1514851247
transform -1 0 124 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_28
timestamp 1514851247
transform -1 0 148 0 1 1105
box 0 0 24 100
use XOR2X1  XOR2X1_5
timestamp 1514851247
transform 1 0 148 0 1 1105
box 0 0 56 100
use NAND2X1  NAND2X1_26
timestamp 1514851247
transform -1 0 228 0 1 1105
box 0 0 24 100
use NOR2X1  NOR2X1_4
timestamp 1514851247
transform -1 0 252 0 1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_8
timestamp 1514851247
transform -1 0 284 0 1 1105
box 0 0 32 100
use XOR2X1  XOR2X1_4
timestamp 1514851247
transform 1 0 284 0 1 1105
box 0 0 56 100
use BUFX2  BUFX2_54
timestamp 1514851247
transform -1 0 364 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_29
timestamp 1514851247
transform -1 0 388 0 1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_3
timestamp 1514851247
transform 1 0 388 0 1 1105
box 0 0 32 100
use AOI21X1  AOI21X1_4
timestamp 1514851247
transform 1 0 420 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_87
timestamp 1514851247
transform -1 0 484 0 1 1105
box 0 0 32 100
use XOR2X1  XOR2X1_1
timestamp 1514851247
transform 1 0 484 0 1 1105
box 0 0 56 100
use INVX1  INVX1_25
timestamp 1514851247
transform 1 0 540 0 1 1105
box 0 0 16 100
use NAND2X1  NAND2X1_31
timestamp 1514851247
transform -1 0 580 0 1 1105
box 0 0 24 100
use AOI21X1  AOI21X1_9
timestamp 1514851247
transform 1 0 580 0 1 1105
box 0 0 32 100
use NOR2X1  NOR2X1_5
timestamp 1514851247
transform -1 0 636 0 1 1105
box 0 0 24 100
use OR2X2  OR2X2_106
timestamp 1514851247
transform 1 0 636 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_67
timestamp 1514851247
transform 1 0 668 0 1 1105
box 0 0 32 100
use BUFX2  BUFX2_31
timestamp 1514851247
transform 1 0 700 0 1 1105
box 0 0 24 100
use BUFX2  BUFX2_56
timestamp 1514851247
transform 1 0 724 0 1 1105
box 0 0 24 100
use OAI21X1  OAI21X1_14
timestamp 1514851247
transform 1 0 748 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_27
timestamp 1514851247
transform -1 0 812 0 1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_33
timestamp 1514851247
transform -1 0 860 0 1 1105
box 0 0 48 100
use BUFX2  BUFX2_33
timestamp 1514851247
transform 1 0 860 0 1 1105
box 0 0 24 100
use MUX2X1  MUX2X1_9
timestamp 1514851247
transform 1 0 884 0 1 1105
box 0 0 48 100
use MUX2X1  MUX2X1_20
timestamp 1514851247
transform 1 0 932 0 1 1105
box 0 0 48 100
use MUX2X1  MUX2X1_19
timestamp 1514851247
transform -1 0 1028 0 1 1105
box 0 0 48 100
use MUX2X1  MUX2X1_11
timestamp 1514851247
transform 1 0 1028 0 1 1105
box 0 0 48 100
use OR2X2  OR2X2_25
timestamp 1514851247
transform 1 0 1076 0 1 1105
box 0 0 32 100
use NAND3X1  NAND3X1_11
timestamp 1514851247
transform 1 0 1108 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_26
timestamp 1514851247
transform -1 0 1172 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_65
timestamp 1514851247
transform 1 0 1172 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_102
timestamp 1514851247
transform 1 0 1204 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_34
timestamp 1514851247
transform -1 0 1268 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_103
timestamp 1514851247
transform -1 0 1300 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_64
timestamp 1514851247
transform -1 0 1332 0 1 1105
box 0 0 32 100
use BUFX2  BUFX2_23
timestamp 1514851247
transform -1 0 1356 0 1 1105
box 0 0 24 100
use MUX2X1  MUX2X1_30
timestamp 1514851247
transform -1 0 1404 0 1 1105
box 0 0 48 100
use AND2X2  AND2X2_74
timestamp 1514851247
transform 1 0 1404 0 1 1105
box 0 0 32 100
use INVX2  INVX2_1
timestamp 1514851247
transform -1 0 1452 0 1 1105
box 0 0 16 100
use OR2X2  OR2X2_38
timestamp 1514851247
transform 1 0 1452 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_39
timestamp 1514851247
transform 1 0 1484 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_117
timestamp 1514851247
transform 1 0 1516 0 1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_21
timestamp 1514851247
transform -1 0 1596 0 1 1105
box 0 0 48 100
use AND2X2  AND2X2_92
timestamp 1514851247
transform -1 0 1628 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_54
timestamp 1514851247
transform 1 0 1628 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_78
timestamp 1514851247
transform 1 0 1660 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_119
timestamp 1514851247
transform 1 0 1692 0 1 1105
box 0 0 32 100
use AND2X2  AND2X2_56
timestamp 1514851247
transform -1 0 1756 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_20
timestamp 1514851247
transform -1 0 1788 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_19
timestamp 1514851247
transform 1 0 1788 0 1 1105
box 0 0 32 100
use OR2X2  OR2X2_93
timestamp 1514851247
transform 1 0 1820 0 1 1105
box 0 0 32 100
use INVX1  INVX1_18
timestamp 1514851247
transform 1 0 1852 0 1 1105
box 0 0 16 100
use FILL  FILL_12_1
timestamp 1514851247
transform 1 0 1868 0 1 1105
box 0 0 8 100
use FILL  FILL_12_2
timestamp 1514851247
transform 1 0 1876 0 1 1105
box 0 0 8 100
use NAND2X1  NAND2X1_20
timestamp 1514851247
transform 1 0 4 0 -1 1105
box 0 0 24 100
use NAND3X1  NAND3X1_17
timestamp 1514851247
transform -1 0 60 0 -1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_21
timestamp 1514851247
transform -1 0 84 0 -1 1105
box 0 0 24 100
use OR2X2  OR2X2_74
timestamp 1514851247
transform 1 0 84 0 -1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_27
timestamp 1514851247
transform -1 0 140 0 -1 1105
box 0 0 24 100
use AND2X2  AND2X2_69
timestamp 1514851247
transform -1 0 172 0 -1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_17
timestamp 1514851247
transform -1 0 196 0 -1 1105
box 0 0 24 100
use AOI22X1  AOI22X1_3
timestamp 1514851247
transform 1 0 196 0 -1 1105
box 0 0 40 100
use OR2X2  OR2X2_97
timestamp 1514851247
transform 1 0 236 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_88
timestamp 1514851247
transform 1 0 268 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_36
timestamp 1514851247
transform -1 0 348 0 -1 1105
box 0 0 48 100
use OR2X2  OR2X2_50
timestamp 1514851247
transform 1 0 348 0 -1 1105
box 0 0 32 100
use NAND2X1  NAND2X1_18
timestamp 1514851247
transform 1 0 380 0 -1 1105
box 0 0 24 100
use MUX2X1  MUX2X1_39
timestamp 1514851247
transform 1 0 404 0 -1 1105
box 0 0 48 100
use OAI21X1  OAI21X1_4
timestamp 1514851247
transform -1 0 484 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_52
timestamp 1514851247
transform -1 0 516 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_28
timestamp 1514851247
transform -1 0 564 0 -1 1105
box 0 0 48 100
use NAND2X1  NAND2X1_16
timestamp 1514851247
transform 1 0 564 0 -1 1105
box 0 0 24 100
use MUX2X1  MUX2X1_1
timestamp 1514851247
transform -1 0 636 0 -1 1105
box 0 0 48 100
use NAND3X1  NAND3X1_13
timestamp 1514851247
transform -1 0 668 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_32
timestamp 1514851247
transform -1 0 700 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_31
timestamp 1514851247
transform -1 0 732 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_66
timestamp 1514851247
transform -1 0 764 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_41
timestamp 1514851247
transform 1 0 764 0 -1 1105
box 0 0 48 100
use BUFX2  BUFX2_48
timestamp 1514851247
transform -1 0 836 0 -1 1105
box 0 0 24 100
use MUX2X1  MUX2X1_37
timestamp 1514851247
transform 1 0 836 0 -1 1105
box 0 0 48 100
use AND2X2  AND2X2_65
timestamp 1514851247
transform -1 0 916 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_64
timestamp 1514851247
transform -1 0 948 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_8
timestamp 1514851247
transform 1 0 948 0 -1 1105
box 0 0 48 100
use OR2X2  OR2X2_44
timestamp 1514851247
transform 1 0 996 0 -1 1105
box 0 0 32 100
use NAND3X1  NAND3X1_14
timestamp 1514851247
transform 1 0 1028 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_45
timestamp 1514851247
transform -1 0 1092 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_22
timestamp 1514851247
transform -1 0 1140 0 -1 1105
box 0 0 48 100
use AND2X2  AND2X2_36
timestamp 1514851247
transform 1 0 1140 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_38
timestamp 1514851247
transform 1 0 1172 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_9
timestamp 1514851247
transform -1 0 1236 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_37
timestamp 1514851247
transform -1 0 1268 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_13
timestamp 1514851247
transform 1 0 1268 0 -1 1105
box 0 0 48 100
use MUX2X1  MUX2X1_10
timestamp 1514851247
transform -1 0 1364 0 -1 1105
box 0 0 48 100
use MUX2X1  MUX2X1_15
timestamp 1514851247
transform 1 0 1364 0 -1 1105
box 0 0 48 100
use AND2X2  AND2X2_77
timestamp 1514851247
transform -1 0 1444 0 -1 1105
box 0 0 32 100
use MUX2X1  MUX2X1_14
timestamp 1514851247
transform -1 0 1492 0 -1 1105
box 0 0 48 100
use AND2X2  AND2X2_76
timestamp 1514851247
transform -1 0 1524 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_75
timestamp 1514851247
transform -1 0 1556 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_56
timestamp 1514851247
transform -1 0 1588 0 -1 1105
box 0 0 32 100
use OR2X2  OR2X2_55
timestamp 1514851247
transform -1 0 1620 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_91
timestamp 1514851247
transform -1 0 1652 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_118
timestamp 1514851247
transform 1 0 1652 0 -1 1105
box 0 0 32 100
use BUFX2  BUFX2_12
timestamp 1514851247
transform -1 0 1708 0 -1 1105
box 0 0 24 100
use OR2X2  OR2X2_80
timestamp 1514851247
transform 1 0 1708 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_58
timestamp 1514851247
transform 1 0 1740 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_55
timestamp 1514851247
transform 1 0 1772 0 -1 1105
box 0 0 32 100
use NAND3X1  NAND3X1_24
timestamp 1514851247
transform 1 0 1804 0 -1 1105
box 0 0 32 100
use AND2X2  AND2X2_134
timestamp 1514851247
transform 1 0 1836 0 -1 1105
box 0 0 32 100
use FILL  FILL_11_1
timestamp 1514851247
transform -1 0 1876 0 -1 1105
box 0 0 8 100
use FILL  FILL_11_2
timestamp 1514851247
transform -1 0 1884 0 -1 1105
box 0 0 8 100
use BUFX2  BUFX2_57
timestamp 1514851247
transform -1 0 28 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_32
timestamp 1514851247
transform -1 0 52 0 1 905
box 0 0 24 100
use INVX1  INVX1_26
timestamp 1514851247
transform -1 0 68 0 1 905
box 0 0 16 100
use AOI21X1  AOI21X1_6
timestamp 1514851247
transform 1 0 68 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_143
timestamp 1514851247
transform -1 0 132 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_109
timestamp 1514851247
transform 1 0 132 0 1 905
box 0 0 32 100
use OAI21X1  OAI21X1_5
timestamp 1514851247
transform -1 0 196 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_110
timestamp 1514851247
transform 1 0 196 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_167
timestamp 1514851247
transform -1 0 260 0 1 905
box 0 0 32 100
use NAND2X1  NAND2X1_1
timestamp 1514851247
transform -1 0 284 0 1 905
box 0 0 24 100
use AND2X2  AND2X2_140
timestamp 1514851247
transform 1 0 284 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_100
timestamp 1514851247
transform -1 0 348 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_108
timestamp 1514851247
transform 1 0 348 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_137
timestamp 1514851247
transform 1 0 380 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_138
timestamp 1514851247
transform -1 0 444 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_200
timestamp 1514851247
transform 1 0 444 0 1 905
box 0 0 32 100
use NAND3X1  NAND3X1_16
timestamp 1514851247
transform -1 0 508 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_51
timestamp 1514851247
transform -1 0 540 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_49
timestamp 1514851247
transform -1 0 572 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_30
timestamp 1514851247
transform 1 0 572 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_191
timestamp 1514851247
transform 1 0 604 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_48
timestamp 1514851247
transform -1 0 668 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_145
timestamp 1514851247
transform 1 0 668 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_86
timestamp 1514851247
transform -1 0 732 0 1 905
box 0 0 32 100
use NAND3X1  NAND3X1_15
timestamp 1514851247
transform 1 0 732 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_47
timestamp 1514851247
transform -1 0 796 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_21
timestamp 1514851247
transform -1 0 820 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_25
timestamp 1514851247
transform 1 0 820 0 1 905
box 0 0 24 100
use AND2X2  AND2X2_127
timestamp 1514851247
transform 1 0 844 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_128
timestamp 1514851247
transform -1 0 908 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_2
timestamp 1514851247
transform -1 0 932 0 1 905
box 0 0 24 100
use BUFX2  BUFX2_51
timestamp 1514851247
transform -1 0 956 0 1 905
box 0 0 24 100
use AND2X2  AND2X2_83
timestamp 1514851247
transform -1 0 988 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_84
timestamp 1514851247
transform 1 0 988 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_43
timestamp 1514851247
transform -1 0 1052 0 1 905
box 0 0 32 100
use INVX1  INVX1_20
timestamp 1514851247
transform -1 0 1068 0 1 905
box 0 0 16 100
use OAI21X1  OAI21X1_6
timestamp 1514851247
transform -1 0 1100 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_39
timestamp 1514851247
transform -1 0 1132 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_10
timestamp 1514851247
transform -1 0 1164 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_7
timestamp 1514851247
transform 1 0 1164 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_8
timestamp 1514851247
transform -1 0 1228 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_122
timestamp 1514851247
transform 1 0 1228 0 1 905
box 0 0 32 100
use BUFX2  BUFX2_24
timestamp 1514851247
transform 1 0 1260 0 1 905
box 0 0 24 100
use INVX1  INVX1_16
timestamp 1514851247
transform -1 0 1300 0 1 905
box 0 0 16 100
use MUX2X1  MUX2X1_32
timestamp 1514851247
transform 1 0 1300 0 1 905
box 0 0 48 100
use OR2X2  OR2X2_82
timestamp 1514851247
transform -1 0 1380 0 1 905
box 0 0 32 100
use INVX1  INVX1_11
timestamp 1514851247
transform -1 0 1396 0 1 905
box 0 0 16 100
use AND2X2  AND2X2_26
timestamp 1514851247
transform 1 0 1396 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_37
timestamp 1514851247
transform -1 0 1460 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_96
timestamp 1514851247
transform -1 0 1492 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_95
timestamp 1514851247
transform -1 0 1524 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_59
timestamp 1514851247
transform -1 0 1556 0 1 905
box 0 0 32 100
use MUX2X1  MUX2X1_31
timestamp 1514851247
transform -1 0 1604 0 1 905
box 0 0 48 100
use MUX2X1  MUX2X1_25
timestamp 1514851247
transform 1 0 1604 0 1 905
box 0 0 48 100
use AND2X2  AND2X2_120
timestamp 1514851247
transform -1 0 1684 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_77
timestamp 1514851247
transform -1 0 1716 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_81
timestamp 1514851247
transform -1 0 1748 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_18
timestamp 1514851247
transform -1 0 1780 0 1 905
box 0 0 32 100
use OR2X2  OR2X2_17
timestamp 1514851247
transform -1 0 1812 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_52
timestamp 1514851247
transform -1 0 1844 0 1 905
box 0 0 32 100
use AND2X2  AND2X2_53
timestamp 1514851247
transform -1 0 1876 0 1 905
box 0 0 32 100
use FILL  FILL_10_1
timestamp 1514851247
transform 1 0 1876 0 1 905
box 0 0 8 100
use BUFX2  BUFX2_58
timestamp 1514851247
transform -1 0 28 0 -1 905
box 0 0 24 100
use BUFX2  BUFX2_34
timestamp 1514851247
transform -1 0 52 0 -1 905
box 0 0 24 100
use INVX1  INVX1_1
timestamp 1514851247
transform -1 0 68 0 -1 905
box 0 0 16 100
use AND2X2  AND2X2_230
timestamp 1514851247
transform 1 0 68 0 -1 905
box 0 0 32 100
use BUFX2  BUFX2_55
timestamp 1514851247
transform -1 0 124 0 -1 905
box 0 0 24 100
use BUFX2  BUFX2_30
timestamp 1514851247
transform -1 0 148 0 -1 905
box 0 0 24 100
use INVX1  INVX1_24
timestamp 1514851247
transform -1 0 164 0 -1 905
box 0 0 16 100
use OR2X2  OR2X2_75
timestamp 1514851247
transform 1 0 164 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_228
timestamp 1514851247
transform -1 0 228 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_227
timestamp 1514851247
transform -1 0 260 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_111
timestamp 1514851247
transform 1 0 260 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_142
timestamp 1514851247
transform -1 0 324 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_141
timestamp 1514851247
transform -1 0 356 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_71
timestamp 1514851247
transform -1 0 388 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_107
timestamp 1514851247
transform -1 0 420 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_98
timestamp 1514851247
transform 1 0 420 0 -1 905
box 0 0 32 100
use INVX1  INVX1_21
timestamp 1514851247
transform -1 0 468 0 -1 905
box 0 0 16 100
use OR2X2  OR2X2_28
timestamp 1514851247
transform 1 0 468 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_29
timestamp 1514851247
transform 1 0 500 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_142
timestamp 1514851247
transform 1 0 532 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_211
timestamp 1514851247
transform -1 0 596 0 -1 905
box 0 0 32 100
use INVX2  INVX2_3
timestamp 1514851247
transform -1 0 612 0 -1 905
box 0 0 16 100
use AND2X2  AND2X2_153
timestamp 1514851247
transform 1 0 612 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_1
timestamp 1514851247
transform 1 0 644 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_1
timestamp 1514851247
transform 1 0 676 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_108
timestamp 1514851247
transform -1 0 740 0 -1 905
box 0 0 32 100
use NAND3X1  NAND3X1_20
timestamp 1514851247
transform 1 0 740 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_149
timestamp 1514851247
transform -1 0 804 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_107
timestamp 1514851247
transform -1 0 836 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_148
timestamp 1514851247
transform -1 0 868 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_89
timestamp 1514851247
transform 1 0 868 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_147
timestamp 1514851247
transform -1 0 932 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_156
timestamp 1514851247
transform -1 0 964 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_112
timestamp 1514851247
transform -1 0 996 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_85
timestamp 1514851247
transform -1 0 1028 0 -1 905
box 0 0 32 100
use MUX2X1  MUX2X1_34
timestamp 1514851247
transform 1 0 1028 0 -1 905
box 0 0 48 100
use OR2X2  OR2X2_105
timestamp 1514851247
transform -1 0 1108 0 -1 905
box 0 0 32 100
use NAND3X1  NAND3X1_25
timestamp 1514851247
transform 1 0 1108 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_96
timestamp 1514851247
transform -1 0 1172 0 -1 905
box 0 0 32 100
use INVX2  INVX2_4
timestamp 1514851247
transform 1 0 1172 0 -1 905
box 0 0 16 100
use OR2X2  OR2X2_23
timestamp 1514851247
transform -1 0 1220 0 -1 905
box 0 0 32 100
use MUX2X1  MUX2X1_27
timestamp 1514851247
transform 1 0 1220 0 -1 905
box 0 0 48 100
use OR2X2  OR2X2_66
timestamp 1514851247
transform -1 0 1300 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_104
timestamp 1514851247
transform -1 0 1332 0 -1 905
box 0 0 32 100
use BUFX2  BUFX2_49
timestamp 1514851247
transform -1 0 1356 0 -1 905
box 0 0 24 100
use AND2X2  AND2X2_105
timestamp 1514851247
transform -1 0 1388 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_94
timestamp 1514851247
transform -1 0 1420 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_195
timestamp 1514851247
transform 1 0 1420 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_60
timestamp 1514851247
transform 1 0 1452 0 -1 905
box 0 0 32 100
use NAND3X1  NAND3X1_30
timestamp 1514851247
transform 1 0 1484 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_103
timestamp 1514851247
transform -1 0 1548 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_144
timestamp 1514851247
transform -1 0 1580 0 -1 905
box 0 0 32 100
use NAND3X1  NAND3X1_26
timestamp 1514851247
transform 1 0 1580 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_102
timestamp 1514851247
transform -1 0 1644 0 -1 905
box 0 0 32 100
use MUX2X1  MUX2X1_40
timestamp 1514851247
transform 1 0 1644 0 -1 905
box 0 0 48 100
use AND2X2  AND2X2_73
timestamp 1514851247
transform -1 0 1724 0 -1 905
box 0 0 32 100
use OR2X2  OR2X2_34
timestamp 1514851247
transform -1 0 1756 0 -1 905
box 0 0 32 100
use AND2X2  AND2X2_116
timestamp 1514851247
transform -1 0 1788 0 -1 905
box 0 0 32 100
use INVX1  INVX1_12
timestamp 1514851247
transform -1 0 1804 0 -1 905
box 0 0 16 100
use OR2X2  OR2X2_36
timestamp 1514851247
transform -1 0 1836 0 -1 905
box 0 0 32 100
use MUX2X1  MUX2X1_38
timestamp 1514851247
transform 1 0 1836 0 -1 905
box 0 0 48 100
use BUFX2  BUFX2_59
timestamp 1514851247
transform -1 0 28 0 1 705
box 0 0 24 100
use BUFX2  BUFX2_35
timestamp 1514851247
transform -1 0 52 0 1 705
box 0 0 24 100
use INVX1  INVX1_10
timestamp 1514851247
transform -1 0 68 0 1 705
box 0 0 16 100
use AND2X2  AND2X2_231
timestamp 1514851247
transform -1 0 100 0 1 705
box 0 0 32 100
use XOR2X1  XOR2X1_6
timestamp 1514851247
transform 1 0 100 0 1 705
box 0 0 56 100
use AOI21X1  AOI21X1_10
timestamp 1514851247
transform 1 0 156 0 1 705
box 0 0 32 100
use NOR2X1  NOR2X1_8
timestamp 1514851247
transform -1 0 212 0 1 705
box 0 0 24 100
use NAND2X1  NAND2X1_12
timestamp 1514851247
transform -1 0 236 0 1 705
box 0 0 24 100
use AND2X2  AND2X2_115
timestamp 1514851247
transform -1 0 268 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_114
timestamp 1514851247
transform -1 0 300 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_70
timestamp 1514851247
transform -1 0 332 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_73
timestamp 1514851247
transform -1 0 364 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_99
timestamp 1514851247
transform -1 0 396 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_136
timestamp 1514851247
transform -1 0 428 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_139
timestamp 1514851247
transform -1 0 460 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_157
timestamp 1514851247
transform -1 0 492 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_112
timestamp 1514851247
transform -1 0 524 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_155
timestamp 1514851247
transform -1 0 556 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_115
timestamp 1514851247
transform -1 0 588 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_114
timestamp 1514851247
transform -1 0 620 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_113
timestamp 1514851247
transform -1 0 652 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_132
timestamp 1514851247
transform -1 0 684 0 1 705
box 0 0 32 100
use NAND2X1  NAND2X1_14
timestamp 1514851247
transform 1 0 684 0 1 705
box 0 0 24 100
use OR2X2  OR2X2_156
timestamp 1514851247
transform 1 0 708 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_126
timestamp 1514851247
transform 1 0 740 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_91
timestamp 1514851247
transform 1 0 772 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_129
timestamp 1514851247
transform -1 0 836 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_122
timestamp 1514851247
transform 1 0 836 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_163
timestamp 1514851247
transform -1 0 900 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_79
timestamp 1514851247
transform 1 0 900 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_57
timestamp 1514851247
transform 1 0 932 0 1 705
box 0 0 32 100
use NOR2X1  NOR2X1_7
timestamp 1514851247
transform -1 0 988 0 1 705
box 0 0 24 100
use OR2X2  OR2X2_69
timestamp 1514851247
transform -1 0 1020 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_67
timestamp 1514851247
transform -1 0 1052 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_106
timestamp 1514851247
transform -1 0 1084 0 1 705
box 0 0 32 100
use AOI22X1  AOI22X1_1
timestamp 1514851247
transform -1 0 1124 0 1 705
box 0 0 40 100
use AND2X2  AND2X2_90
timestamp 1514851247
transform -1 0 1156 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_198
timestamp 1514851247
transform 1 0 1156 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_159
timestamp 1514851247
transform 1 0 1188 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_199
timestamp 1514851247
transform -1 0 1252 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_154
timestamp 1514851247
transform -1 0 1284 0 1 705
box 0 0 32 100
use MUX2X1  MUX2X1_43
timestamp 1514851247
transform -1 0 1332 0 1 705
box 0 0 48 100
use MUX2X1  MUX2X1_12
timestamp 1514851247
transform -1 0 1380 0 1 705
box 0 0 48 100
use MUX2X1  MUX2X1_24
timestamp 1514851247
transform 1 0 1380 0 1 705
box 0 0 48 100
use BUFX2  BUFX2_11
timestamp 1514851247
transform -1 0 1452 0 1 705
box 0 0 24 100
use OR2X2  OR2X2_61
timestamp 1514851247
transform -1 0 1484 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_89
timestamp 1514851247
transform -1 0 1516 0 1 705
box 0 0 32 100
use BUFX2  BUFX2_50
timestamp 1514851247
transform 1 0 1516 0 1 705
box 0 0 24 100
use AND2X2  AND2X2_32
timestamp 1514851247
transform 1 0 1540 0 1 705
box 0 0 32 100
use AOI21X1  AOI21X1_1
timestamp 1514851247
transform 1 0 1572 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_58
timestamp 1514851247
transform -1 0 1636 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_93
timestamp 1514851247
transform -1 0 1668 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_94
timestamp 1514851247
transform -1 0 1700 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_76
timestamp 1514851247
transform -1 0 1732 0 1 705
box 0 0 32 100
use BUFX2  BUFX2_13
timestamp 1514851247
transform -1 0 1756 0 1 705
box 0 0 24 100
use AND2X2  AND2X2_21
timestamp 1514851247
transform -1 0 1788 0 1 705
box 0 0 32 100
use OR2X2  OR2X2_189
timestamp 1514851247
transform -1 0 1820 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_151
timestamp 1514851247
transform 1 0 1820 0 1 705
box 0 0 32 100
use AND2X2  AND2X2_152
timestamp 1514851247
transform 1 0 1852 0 1 705
box 0 0 32 100
use BUFX2  BUFX2_69
timestamp 1514851247
transform -1 0 28 0 -1 705
box 0 0 24 100
use BUFX2  BUFX2_46
timestamp 1514851247
transform -1 0 52 0 -1 705
box 0 0 24 100
use AND2X2  AND2X2_232
timestamp 1514851247
transform -1 0 84 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_35
timestamp 1514851247
transform -1 0 116 0 -1 705
box 0 0 32 100
use NAND2X1  NAND2X1_23
timestamp 1514851247
transform -1 0 140 0 -1 705
box 0 0 24 100
use AND2X2  AND2X2_229
timestamp 1514851247
transform -1 0 172 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_131
timestamp 1514851247
transform 1 0 172 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_24
timestamp 1514851247
transform -1 0 236 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_2
timestamp 1514851247
transform 1 0 236 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_13
timestamp 1514851247
transform -1 0 300 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_100
timestamp 1514851247
transform 1 0 300 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_164
timestamp 1514851247
transform -1 0 364 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_72
timestamp 1514851247
transform -1 0 396 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_189
timestamp 1514851247
transform 1 0 396 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_153
timestamp 1514851247
transform -1 0 460 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_146
timestamp 1514851247
transform 1 0 460 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_222
timestamp 1514851247
transform -1 0 524 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_133
timestamp 1514851247
transform -1 0 556 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_132
timestamp 1514851247
transform -1 0 588 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_147
timestamp 1514851247
transform -1 0 620 0 -1 705
box 0 0 32 100
use BUFX2  BUFX2_8
timestamp 1514851247
transform -1 0 644 0 -1 705
box 0 0 24 100
use NAND3X1  NAND3X1_7
timestamp 1514851247
transform -1 0 676 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_131
timestamp 1514851247
transform -1 0 708 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_130
timestamp 1514851247
transform -1 0 740 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_92
timestamp 1514851247
transform -1 0 772 0 -1 705
box 0 0 32 100
use BUFX2  BUFX2_9
timestamp 1514851247
transform -1 0 796 0 -1 705
box 0 0 24 100
use OR2X2  OR2X2_35
timestamp 1514851247
transform -1 0 828 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_137
timestamp 1514851247
transform 1 0 828 0 -1 705
box 0 0 32 100
use NOR2X1  NOR2X1_1
timestamp 1514851247
transform -1 0 884 0 -1 705
box 0 0 24 100
use AND2X2  AND2X2_180
timestamp 1514851247
transform -1 0 916 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_7
timestamp 1514851247
transform -1 0 948 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_120
timestamp 1514851247
transform -1 0 980 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_86
timestamp 1514851247
transform -1 0 1012 0 -1 705
box 0 0 32 100
use OAI21X1  OAI21X1_1
timestamp 1514851247
transform 1 0 1012 0 -1 705
box 0 0 32 100
use INVX1  INVX1_30
timestamp 1514851247
transform 1 0 1044 0 -1 705
box 0 0 16 100
use AOI22X1  AOI22X1_2
timestamp 1514851247
transform -1 0 1100 0 -1 705
box 0 0 40 100
use NAND2X1  NAND2X1_30
timestamp 1514851247
transform -1 0 1124 0 -1 705
box 0 0 24 100
use NAND2X1  NAND2X1_29
timestamp 1514851247
transform -1 0 1148 0 -1 705
box 0 0 24 100
use NOR2X1  NOR2X1_2
timestamp 1514851247
transform -1 0 1172 0 -1 705
box 0 0 24 100
use AOI21X1  AOI21X1_7
timestamp 1514851247
transform -1 0 1204 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_160
timestamp 1514851247
transform -1 0 1236 0 -1 705
box 0 0 32 100
use NOR2X1  NOR2X1_6
timestamp 1514851247
transform -1 0 1260 0 -1 705
box 0 0 24 100
use OR2X2  OR2X2_85
timestamp 1514851247
transform -1 0 1292 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_84
timestamp 1514851247
transform -1 0 1324 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_123
timestamp 1514851247
transform -1 0 1356 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_33
timestamp 1514851247
transform -1 0 1388 0 -1 705
box 0 0 32 100
use MUX2X1  MUX2X1_23
timestamp 1514851247
transform -1 0 1436 0 -1 705
box 0 0 48 100
use MUX2X1  MUX2X1_6
timestamp 1514851247
transform 1 0 1436 0 -1 705
box 0 0 48 100
use OR2X2  OR2X2_196
timestamp 1514851247
transform -1 0 1516 0 -1 705
box 0 0 32 100
use BUFX2  BUFX2_1
timestamp 1514851247
transform 1 0 1516 0 -1 705
box 0 0 24 100
use AND2X2  AND2X2_22
timestamp 1514851247
transform -1 0 1572 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_4
timestamp 1514851247
transform -1 0 1604 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_31
timestamp 1514851247
transform -1 0 1636 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_178
timestamp 1514851247
transform -1 0 1668 0 -1 705
box 0 0 32 100
use AOI21X1  AOI21X1_5
timestamp 1514851247
transform -1 0 1700 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_109
timestamp 1514851247
transform -1 0 1732 0 -1 705
box 0 0 32 100
use OR2X2  OR2X2_190
timestamp 1514851247
transform -1 0 1764 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_18
timestamp 1514851247
transform 1 0 1764 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_20
timestamp 1514851247
transform -1 0 1828 0 -1 705
box 0 0 32 100
use AND2X2  AND2X2_19
timestamp 1514851247
transform -1 0 1860 0 -1 705
box 0 0 32 100
use FILL  FILL_7_1
timestamp 1514851247
transform -1 0 1868 0 -1 705
box 0 0 8 100
use FILL  FILL_7_2
timestamp 1514851247
transform -1 0 1876 0 -1 705
box 0 0 8 100
use FILL  FILL_7_3
timestamp 1514851247
transform -1 0 1884 0 -1 705
box 0 0 8 100
use BUFX2  BUFX2_60
timestamp 1514851247
transform -1 0 28 0 1 505
box 0 0 24 100
use BUFX2  BUFX2_36
timestamp 1514851247
transform -1 0 52 0 1 505
box 0 0 24 100
use INVX1  INVX1_19
timestamp 1514851247
transform -1 0 68 0 1 505
box 0 0 16 100
use NAND2X1  NAND2X1_34
timestamp 1514851247
transform -1 0 92 0 1 505
box 0 0 24 100
use OR2X2  OR2X2_90
timestamp 1514851247
transform 1 0 92 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_223
timestamp 1514851247
transform 1 0 124 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_225
timestamp 1514851247
transform 1 0 156 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_226
timestamp 1514851247
transform -1 0 220 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_135
timestamp 1514851247
transform -1 0 252 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_179
timestamp 1514851247
transform -1 0 284 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_177
timestamp 1514851247
transform -1 0 316 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_133
timestamp 1514851247
transform -1 0 348 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_173
timestamp 1514851247
transform -1 0 380 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_128
timestamp 1514851247
transform -1 0 412 0 1 505
box 0 0 32 100
use NAND3X1  NAND3X1_22
timestamp 1514851247
transform -1 0 444 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_116
timestamp 1514851247
transform 1 0 444 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_172
timestamp 1514851247
transform -1 0 508 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_190
timestamp 1514851247
transform 1 0 508 0 1 505
box 0 0 32 100
use INVX2  INVX2_2
timestamp 1514851247
transform 1 0 540 0 1 505
box 0 0 16 100
use AND2X2  AND2X2_188
timestamp 1514851247
transform -1 0 588 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_221
timestamp 1514851247
transform -1 0 620 0 1 505
box 0 0 32 100
use NAND2X1  NAND2X1_11
timestamp 1514851247
transform 1 0 620 0 1 505
box 0 0 24 100
use AOI21X1  AOI21X1_3
timestamp 1514851247
transform -1 0 676 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_46
timestamp 1514851247
transform 1 0 676 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_124
timestamp 1514851247
transform -1 0 740 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_79
timestamp 1514851247
transform -1 0 772 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_113
timestamp 1514851247
transform -1 0 804 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_101
timestamp 1514851247
transform -1 0 836 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_202
timestamp 1514851247
transform 1 0 836 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_14
timestamp 1514851247
transform 1 0 868 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_45
timestamp 1514851247
transform -1 0 932 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_68
timestamp 1514851247
transform -1 0 964 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_24
timestamp 1514851247
transform -1 0 996 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_127
timestamp 1514851247
transform -1 0 1028 0 1 505
box 0 0 32 100
use BUFX2  BUFX2_22
timestamp 1514851247
transform -1 0 1052 0 1 505
box 0 0 24 100
use INVX1  INVX1_14
timestamp 1514851247
transform 1 0 1052 0 1 505
box 0 0 16 100
use OR2X2  OR2X2_149
timestamp 1514851247
transform -1 0 1100 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_148
timestamp 1514851247
transform -1 0 1132 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_197
timestamp 1514851247
transform -1 0 1164 0 1 505
box 0 0 32 100
use MUX2X1  MUX2X1_45
timestamp 1514851247
transform -1 0 1212 0 1 505
box 0 0 48 100
use MUX2X1  MUX2X1_46
timestamp 1514851247
transform -1 0 1260 0 1 505
box 0 0 48 100
use AND2X2  AND2X2_170
timestamp 1514851247
transform -1 0 1292 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_171
timestamp 1514851247
transform -1 0 1324 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_187
timestamp 1514851247
transform -1 0 1356 0 1 505
box 0 0 32 100
use MUX2X1  MUX2X1_44
timestamp 1514851247
transform -1 0 1404 0 1 505
box 0 0 48 100
use MUX2X1  MUX2X1_42
timestamp 1514851247
transform -1 0 1452 0 1 505
box 0 0 48 100
use MUX2X1  MUX2X1_16
timestamp 1514851247
transform 1 0 1452 0 1 505
box 0 0 48 100
use AND2X2  AND2X2_62
timestamp 1514851247
transform -1 0 1532 0 1 505
box 0 0 32 100
use OR2X2  OR2X2_63
timestamp 1514851247
transform 1 0 1532 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_99
timestamp 1514851247
transform 1 0 1564 0 1 505
box 0 0 32 100
use BUFX2  BUFX2_20
timestamp 1514851247
transform 1 0 1596 0 1 505
box 0 0 24 100
use MUX2X1  MUX2X1_17
timestamp 1514851247
transform 1 0 1620 0 1 505
box 0 0 48 100
use INVX1  INVX1_23
timestamp 1514851247
transform -1 0 1684 0 1 505
box 0 0 16 100
use OR2X2  OR2X2_62
timestamp 1514851247
transform -1 0 1716 0 1 505
box 0 0 32 100
use AND2X2  AND2X2_97
timestamp 1514851247
transform -1 0 1748 0 1 505
box 0 0 32 100
use MUX2X1  MUX2X1_35
timestamp 1514851247
transform -1 0 1796 0 1 505
box 0 0 48 100
use MUX2X1  MUX2X1_29
timestamp 1514851247
transform -1 0 1844 0 1 505
box 0 0 48 100
use AND2X2  AND2X2_17
timestamp 1514851247
transform -1 0 1876 0 1 505
box 0 0 32 100
use FILL  FILL_6_1
timestamp 1514851247
transform 1 0 1876 0 1 505
box 0 0 8 100
use BUFX2  BUFX2_63
timestamp 1514851247
transform -1 0 28 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_33
timestamp 1514851247
transform 1 0 28 0 -1 505
box 0 0 24 100
use NAND3X1  NAND3X1_27
timestamp 1514851247
transform -1 0 84 0 -1 505
box 0 0 32 100
use AOI21X1  AOI21X1_11
timestamp 1514851247
transform 1 0 84 0 -1 505
box 0 0 32 100
use BUFX2  BUFX2_39
timestamp 1514851247
transform -1 0 140 0 -1 505
box 0 0 24 100
use INVX1  INVX1_29
timestamp 1514851247
transform -1 0 156 0 -1 505
box 0 0 16 100
use AND2X2  AND2X2_224
timestamp 1514851247
transform -1 0 188 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_68
timestamp 1514851247
transform 1 0 188 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_136
timestamp 1514851247
transform -1 0 252 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_176
timestamp 1514851247
transform 1 0 252 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_134
timestamp 1514851247
transform -1 0 316 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_175
timestamp 1514851247
transform -1 0 348 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_27
timestamp 1514851247
transform 1 0 348 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_170
timestamp 1514851247
transform 1 0 380 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_24
timestamp 1514851247
transform 1 0 412 0 -1 505
box 0 0 24 100
use NAND2X1  NAND2X1_22
timestamp 1514851247
transform -1 0 460 0 -1 505
box 0 0 24 100
use OR2X2  OR2X2_88
timestamp 1514851247
transform 1 0 460 0 -1 505
box 0 0 32 100
use NAND3X1  NAND3X1_19
timestamp 1514851247
transform -1 0 524 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_150
timestamp 1514851247
transform 1 0 524 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_125
timestamp 1514851247
transform 1 0 556 0 -1 505
box 0 0 32 100
use INVX1  INVX1_15
timestamp 1514851247
transform 1 0 588 0 -1 505
box 0 0 16 100
use NAND2X1  NAND2X1_13
timestamp 1514851247
transform 1 0 604 0 -1 505
box 0 0 24 100
use AND2X2  AND2X2_41
timestamp 1514851247
transform 1 0 628 0 -1 505
box 0 0 32 100
use OAI21X1  OAI21X1_12
timestamp 1514851247
transform 1 0 660 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_15
timestamp 1514851247
transform 1 0 692 0 -1 505
box 0 0 24 100
use AND2X2  AND2X2_43
timestamp 1514851247
transform 1 0 716 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_6
timestamp 1514851247
transform 1 0 748 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_40
timestamp 1514851247
transform 1 0 780 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_11
timestamp 1514851247
transform 1 0 812 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_44
timestamp 1514851247
transform 1 0 844 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_123
timestamp 1514851247
transform 1 0 876 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_130
timestamp 1514851247
transform -1 0 940 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_201
timestamp 1514851247
transform -1 0 972 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_28
timestamp 1514851247
transform 1 0 972 0 -1 505
box 0 0 24 100
use AND2X2  AND2X2_121
timestamp 1514851247
transform -1 0 1028 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_158
timestamp 1514851247
transform -1 0 1060 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_157
timestamp 1514851247
transform -1 0 1092 0 -1 505
box 0 0 32 100
use NAND2X1  NAND2X1_25
timestamp 1514851247
transform 1 0 1092 0 -1 505
box 0 0 24 100
use OR2X2  OR2X2_5
timestamp 1514851247
transform -1 0 1148 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_30
timestamp 1514851247
transform -1 0 1180 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_83
timestamp 1514851247
transform -1 0 1212 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_196
timestamp 1514851247
transform -1 0 1244 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_129
timestamp 1514851247
transform -1 0 1276 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_186
timestamp 1514851247
transform -1 0 1308 0 -1 505
box 0 0 32 100
use BUFX2  BUFX2_44
timestamp 1514851247
transform 1 0 1308 0 -1 505
box 0 0 24 100
use MUX2X1  MUX2X1_7
timestamp 1514851247
transform 1 0 1332 0 -1 505
box 0 0 48 100
use AND2X2  AND2X2_81
timestamp 1514851247
transform 1 0 1380 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_41
timestamp 1514851247
transform -1 0 1444 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_22
timestamp 1514851247
transform -1 0 1476 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_80
timestamp 1514851247
transform -1 0 1508 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_61
timestamp 1514851247
transform -1 0 1540 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_98
timestamp 1514851247
transform 1 0 1540 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_188
timestamp 1514851247
transform -1 0 1604 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_15
timestamp 1514851247
transform -1 0 1636 0 -1 505
box 0 0 32 100
use XNOR2X1  XNOR2X1_1
timestamp 1514851247
transform 1 0 1636 0 -1 505
box 0 0 56 100
use AND2X2  AND2X2_16
timestamp 1514851247
transform 1 0 1692 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_184
timestamp 1514851247
transform 1 0 1724 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_185
timestamp 1514851247
transform 1 0 1756 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_14
timestamp 1514851247
transform 1 0 1788 0 -1 505
box 0 0 32 100
use AND2X2  AND2X2_150
timestamp 1514851247
transform -1 0 1852 0 -1 505
box 0 0 32 100
use OR2X2  OR2X2_187
timestamp 1514851247
transform 1 0 1852 0 -1 505
box 0 0 32 100
use XOR2X1  XOR2X1_7
timestamp 1514851247
transform -1 0 60 0 1 305
box 0 0 56 100
use NOR2X1  NOR2X1_9
timestamp 1514851247
transform -1 0 84 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_186
timestamp 1514851247
transform 1 0 84 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_46
timestamp 1514851247
transform 1 0 116 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_57
timestamp 1514851247
transform 1 0 148 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_3
timestamp 1514851247
transform 1 0 180 0 1 305
box 0 0 24 100
use NAND2X1  NAND2X1_4
timestamp 1514851247
transform -1 0 228 0 1 305
box 0 0 24 100
use AOI21X1  AOI21X1_15
timestamp 1514851247
transform 1 0 228 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_181
timestamp 1514851247
transform -1 0 292 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_180
timestamp 1514851247
transform -1 0 324 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_179
timestamp 1514851247
transform -1 0 356 0 1 305
box 0 0 32 100
use NAND2X1  NAND2X1_32
timestamp 1514851247
transform 1 0 356 0 1 305
box 0 0 24 100
use NAND3X1  NAND3X1_6
timestamp 1514851247
transform 1 0 380 0 1 305
box 0 0 32 100
use INVX1  INVX1_13
timestamp 1514851247
transform -1 0 428 0 1 305
box 0 0 16 100
use AND2X2  AND2X2_162
timestamp 1514851247
transform -1 0 460 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_161
timestamp 1514851247
transform -1 0 492 0 1 305
box 0 0 32 100
use NAND3X1  NAND3X1_21
timestamp 1514851247
transform 1 0 492 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_216
timestamp 1514851247
transform -1 0 556 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_215
timestamp 1514851247
transform -1 0 588 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_87
timestamp 1514851247
transform -1 0 620 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_3
timestamp 1514851247
transform 1 0 620 0 1 305
box 0 0 24 100
use BUFX2  BUFX2_18
timestamp 1514851247
transform -1 0 668 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_12
timestamp 1514851247
transform -1 0 700 0 1 305
box 0 0 32 100
use BUFX2  BUFX2_3
timestamp 1514851247
transform -1 0 724 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_169
timestamp 1514851247
transform -1 0 756 0 1 305
box 0 0 32 100
use OAI21X1  OAI21X1_13
timestamp 1514851247
transform -1 0 788 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_63
timestamp 1514851247
transform -1 0 820 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_13
timestamp 1514851247
transform 1 0 820 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_111
timestamp 1514851247
transform -1 0 884 0 1 305
box 0 0 32 100
use XOR2X1  XOR2X1_3
timestamp 1514851247
transform 1 0 884 0 1 305
box 0 0 56 100
use BUFX2  BUFX2_4
timestamp 1514851247
transform 1 0 940 0 1 305
box 0 0 24 100
use AND2X2  AND2X2_23
timestamp 1514851247
transform -1 0 996 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_192
timestamp 1514851247
transform -1 0 1028 0 1 305
box 0 0 32 100
use NOR2X1  NOR2X1_12
timestamp 1514851247
transform 1 0 1028 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_2
timestamp 1514851247
transform -1 0 1084 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_82
timestamp 1514851247
transform -1 0 1116 0 1 305
box 0 0 32 100
use XOR2X1  XOR2X1_12
timestamp 1514851247
transform 1 0 1116 0 1 305
box 0 0 56 100
use AND2X2  AND2X2_11
timestamp 1514851247
transform -1 0 1204 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_183
timestamp 1514851247
transform -1 0 1236 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_213
timestamp 1514851247
transform 1 0 1236 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_139
timestamp 1514851247
transform 1 0 1268 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_140
timestamp 1514851247
transform 1 0 1300 0 1 305
box 0 0 32 100
use NAND3X1  NAND3X1_1
timestamp 1514851247
transform -1 0 1364 0 1 305
box 0 0 32 100
use BUFX2  BUFX2_7
timestamp 1514851247
transform -1 0 1388 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_54
timestamp 1514851247
transform 1 0 1388 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_53
timestamp 1514851247
transform -1 0 1452 0 1 305
box 0 0 32 100
use INVX1  INVX1_22
timestamp 1514851247
transform -1 0 1468 0 1 305
box 0 0 16 100
use BUFX4  BUFX4_1
timestamp 1514851247
transform 1 0 1468 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_3
timestamp 1514851247
transform -1 0 1532 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_28
timestamp 1514851247
transform -1 0 1564 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_29
timestamp 1514851247
transform -1 0 1596 0 1 305
box 0 0 32 100
use BUFX2  BUFX2_26
timestamp 1514851247
transform 1 0 1596 0 1 305
box 0 0 24 100
use OR2X2  OR2X2_182
timestamp 1514851247
transform 1 0 1620 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_12
timestamp 1514851247
transform 1 0 1652 0 1 305
box 0 0 32 100
use OR2X2  OR2X2_110
timestamp 1514851247
transform -1 0 1716 0 1 305
box 0 0 32 100
use AND2X2  AND2X2_48
timestamp 1514851247
transform 1 0 1716 0 1 305
box 0 0 32 100
use XOR2X1  XOR2X1_2
timestamp 1514851247
transform -1 0 1804 0 1 305
box 0 0 56 100
use OR2X2  OR2X2_16
timestamp 1514851247
transform 1 0 1804 0 1 305
box 0 0 32 100
use BUFX2  BUFX2_14
timestamp 1514851247
transform -1 0 1860 0 1 305
box 0 0 24 100
use FILL  FILL_4_1
timestamp 1514851247
transform 1 0 1860 0 1 305
box 0 0 8 100
use FILL  FILL_4_2
timestamp 1514851247
transform 1 0 1868 0 1 305
box 0 0 8 100
use FILL  FILL_4_3
timestamp 1514851247
transform 1 0 1876 0 1 305
box 0 0 8 100
use BUFX2  BUFX2_62
timestamp 1514851247
transform -1 0 28 0 -1 305
box 0 0 24 100
use BUFX2  BUFX2_38
timestamp 1514851247
transform -1 0 52 0 -1 305
box 0 0 24 100
use NAND3X1  NAND3X1_23
timestamp 1514851247
transform 1 0 52 0 -1 305
box 0 0 32 100
use INVX1  INVX1_28
timestamp 1514851247
transform -1 0 100 0 -1 305
box 0 0 16 100
use OR2X2  OR2X2_135
timestamp 1514851247
transform 1 0 100 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_174
timestamp 1514851247
transform 1 0 132 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_11
timestamp 1514851247
transform -1 0 188 0 -1 305
box 0 0 24 100
use AND2X2  AND2X2_175
timestamp 1514851247
transform 1 0 188 0 -1 305
box 0 0 32 100
use BUFX2  BUFX2_17
timestamp 1514851247
transform -1 0 244 0 -1 305
box 0 0 24 100
use BUFX2  BUFX2_16
timestamp 1514851247
transform -1 0 268 0 -1 305
box 0 0 24 100
use AND2X2  AND2X2_6
timestamp 1514851247
transform 1 0 268 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_178
timestamp 1514851247
transform 1 0 300 0 -1 305
box 0 0 32 100
use OAI21X1  OAI21X1_2
timestamp 1514851247
transform 1 0 332 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_9
timestamp 1514851247
transform -1 0 396 0 -1 305
box 0 0 32 100
use NAND3X1  NAND3X1_12
timestamp 1514851247
transform -1 0 428 0 -1 305
box 0 0 32 100
use NOR2X1  NOR2X1_13
timestamp 1514851247
transform -1 0 452 0 -1 305
box 0 0 24 100
use NAND3X1  NAND3X1_9
timestamp 1514851247
transform -1 0 484 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_160
timestamp 1514851247
transform -1 0 516 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_25
timestamp 1514851247
transform 1 0 516 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_118
timestamp 1514851247
transform -1 0 580 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_214
timestamp 1514851247
transform -1 0 612 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_174
timestamp 1514851247
transform -1 0 644 0 -1 305
box 0 0 32 100
use INVX1  INVX1_17
timestamp 1514851247
transform -1 0 660 0 -1 305
box 0 0 16 100
use BUFX2  BUFX2_19
timestamp 1514851247
transform 1 0 660 0 -1 305
box 0 0 24 100
use AND2X2  AND2X2_42
timestamp 1514851247
transform 1 0 684 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_168
timestamp 1514851247
transform 1 0 716 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_208
timestamp 1514851247
transform 1 0 748 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_117
timestamp 1514851247
transform -1 0 812 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_162
timestamp 1514851247
transform -1 0 844 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_161
timestamp 1514851247
transform 1 0 844 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_138
timestamp 1514851247
transform 1 0 876 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_126
timestamp 1514851247
transform -1 0 940 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_169
timestamp 1514851247
transform -1 0 972 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_168
timestamp 1514851247
transform -1 0 1004 0 -1 305
box 0 0 32 100
use NAND2X1  NAND2X1_19
timestamp 1514851247
transform 1 0 1004 0 -1 305
box 0 0 24 100
use AOI21X1  AOI21X1_14
timestamp 1514851247
transform -1 0 1060 0 -1 305
box 0 0 32 100
use NAND2X1  NAND2X1_2
timestamp 1514851247
transform 1 0 1060 0 -1 305
box 0 0 24 100
use OR2X2  OR2X2_42
timestamp 1514851247
transform -1 0 1116 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_78
timestamp 1514851247
transform -1 0 1148 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_104
timestamp 1514851247
transform -1 0 1180 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_143
timestamp 1514851247
transform 1 0 1180 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_60
timestamp 1514851247
transform -1 0 1244 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_173
timestamp 1514851247
transform -1 0 1276 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_95
timestamp 1514851247
transform -1 0 1308 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_212
timestamp 1514851247
transform -1 0 1340 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_210
timestamp 1514851247
transform -1 0 1372 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_172
timestamp 1514851247
transform -1 0 1404 0 -1 305
box 0 0 32 100
use BUFX2  BUFX2_10
timestamp 1514851247
transform -1 0 1428 0 -1 305
box 0 0 24 100
use AND2X2  AND2X2_47
timestamp 1514851247
transform -1 0 1460 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_141
timestamp 1514851247
transform -1 0 1492 0 -1 305
box 0 0 32 100
use AOI21X1  AOI21X1_2
timestamp 1514851247
transform -1 0 1524 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_59
timestamp 1514851247
transform -1 0 1556 0 -1 305
box 0 0 32 100
use NAND3X1  NAND3X1_10
timestamp 1514851247
transform 1 0 1556 0 -1 305
box 0 0 32 100
use OR2X2  OR2X2_40
timestamp 1514851247
transform -1 0 1620 0 -1 305
box 0 0 32 100
use XOR2X1  XOR2X1_13
timestamp 1514851247
transform 1 0 1620 0 -1 305
box 0 0 56 100
use OR2X2  OR2X2_21
timestamp 1514851247
transform -1 0 1708 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_146
timestamp 1514851247
transform -1 0 1740 0 -1 305
box 0 0 32 100
use AOI21X1  AOI21X1_12
timestamp 1514851247
transform -1 0 1772 0 -1 305
box 0 0 32 100
use AND2X2  AND2X2_51
timestamp 1514851247
transform 1 0 1772 0 -1 305
box 0 0 32 100
use BUFX2  BUFX2_27
timestamp 1514851247
transform 1 0 1804 0 -1 305
box 0 0 24 100
use INVX1  INVX1_9
timestamp 1514851247
transform 1 0 1828 0 -1 305
box 0 0 16 100
use BUFX2  BUFX2_52
timestamp 1514851247
transform 1 0 1844 0 -1 305
box 0 0 24 100
use FILL  FILL_3_1
timestamp 1514851247
transform -1 0 1876 0 -1 305
box 0 0 8 100
use FILL  FILL_3_2
timestamp 1514851247
transform -1 0 1884 0 -1 305
box 0 0 8 100
use XOR2X1  XOR2X1_8
timestamp 1514851247
transform -1 0 60 0 1 105
box 0 0 56 100
use INVX1  INVX1_27
timestamp 1514851247
transform -1 0 76 0 1 105
box 0 0 16 100
use NAND3X1  NAND3X1_29
timestamp 1514851247
transform -1 0 108 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_121
timestamp 1514851247
transform -1 0 140 0 1 105
box 0 0 32 100
use AOI21X1  AOI21X1_13
timestamp 1514851247
transform 1 0 140 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_32
timestamp 1514851247
transform -1 0 204 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_2
timestamp 1514851247
transform -1 0 236 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_177
timestamp 1514851247
transform -1 0 268 0 1 105
box 0 0 32 100
use INVX1  INVX1_8
timestamp 1514851247
transform -1 0 284 0 1 105
box 0 0 16 100
use AND2X2  AND2X2_5
timestamp 1514851247
transform -1 0 316 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_193
timestamp 1514851247
transform 1 0 316 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_194
timestamp 1514851247
transform 1 0 348 0 1 105
box 0 0 32 100
use INVX1  INVX1_6
timestamp 1514851247
transform 1 0 380 0 1 105
box 0 0 16 100
use AND2X2  AND2X2_8
timestamp 1514851247
transform -1 0 428 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_8
timestamp 1514851247
transform -1 0 460 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_176
timestamp 1514851247
transform 1 0 460 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_217
timestamp 1514851247
transform 1 0 492 0 1 105
box 0 0 32 100
use INVX4  INVX4_1
timestamp 1514851247
transform -1 0 548 0 1 105
box 0 0 24 100
use OAI21X1  OAI21X1_11
timestamp 1514851247
transform 1 0 548 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_171
timestamp 1514851247
transform -1 0 612 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_165
timestamp 1514851247
transform 1 0 612 0 1 105
box 0 0 32 100
use INVX1  INVX1_2
timestamp 1514851247
transform -1 0 660 0 1 105
box 0 0 16 100
use AND2X2  AND2X2_219
timestamp 1514851247
transform 1 0 660 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_220
timestamp 1514851247
transform -1 0 724 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_167
timestamp 1514851247
transform -1 0 756 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_203
timestamp 1514851247
transform 1 0 756 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_5
timestamp 1514851247
transform 1 0 788 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_204
timestamp 1514851247
transform 1 0 820 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_163
timestamp 1514851247
transform -1 0 884 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_207
timestamp 1514851247
transform -1 0 916 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_194
timestamp 1514851247
transform 1 0 916 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_195
timestamp 1514851247
transform 1 0 948 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_155
timestamp 1514851247
transform -1 0 1012 0 1 105
box 0 0 32 100
use XOR2X1  XOR2X1_10
timestamp 1514851247
transform 1 0 1012 0 1 105
box 0 0 56 100
use AND2X2  AND2X2_166
timestamp 1514851247
transform -1 0 1100 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_124
timestamp 1514851247
transform -1 0 1132 0 1 105
box 0 0 32 100
use NAND3X1  NAND3X1_31
timestamp 1514851247
transform 1 0 1132 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_164
timestamp 1514851247
transform -1 0 1196 0 1 105
box 0 0 32 100
use NAND2X1  NAND2X1_37
timestamp 1514851247
transform -1 0 1220 0 1 105
box 0 0 24 100
use OR2X2  OR2X2_151
timestamp 1514851247
transform 1 0 1220 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_191
timestamp 1514851247
transform 1 0 1252 0 1 105
box 0 0 32 100
use OAI21X1  OAI21X1_10
timestamp 1514851247
transform 1 0 1284 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_192
timestamp 1514851247
transform 1 0 1316 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_193
timestamp 1514851247
transform -1 0 1380 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_183
timestamp 1514851247
transform 1 0 1380 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_185
timestamp 1514851247
transform 1 0 1412 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_184
timestamp 1514851247
transform -1 0 1476 0 1 105
box 0 0 32 100
use MUX2X1  MUX2X1_2
timestamp 1514851247
transform -1 0 1524 0 1 105
box 0 0 48 100
use MUX2X1  MUX2X1_3
timestamp 1514851247
transform 1 0 1524 0 1 105
box 0 0 48 100
use OR2X2  OR2X2_154
timestamp 1514851247
transform -1 0 1604 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_50
timestamp 1514851247
transform -1 0 1636 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_71
timestamp 1514851247
transform 1 0 1636 0 1 105
box 0 0 32 100
use MUX2X1  MUX2X1_26
timestamp 1514851247
transform 1 0 1668 0 1 105
box 0 0 48 100
use OR2X2  OR2X2_15
timestamp 1514851247
transform 1 0 1716 0 1 105
box 0 0 32 100
use AND2X2  AND2X2_72
timestamp 1514851247
transform -1 0 1780 0 1 105
box 0 0 32 100
use OR2X2  OR2X2_33
timestamp 1514851247
transform -1 0 1812 0 1 105
box 0 0 32 100
use MUX2X1  MUX2X1_18
timestamp 1514851247
transform 1 0 1812 0 1 105
box 0 0 48 100
use FILL  FILL_2_1
timestamp 1514851247
transform 1 0 1860 0 1 105
box 0 0 8 100
use FILL  FILL_2_2
timestamp 1514851247
transform 1 0 1868 0 1 105
box 0 0 8 100
use FILL  FILL_2_3
timestamp 1514851247
transform 1 0 1876 0 1 105
box 0 0 8 100
use BUFX2  BUFX2_61
timestamp 1514851247
transform -1 0 28 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_37
timestamp 1514851247
transform -1 0 52 0 -1 105
box 0 0 24 100
use NAND3X1  NAND3X1_28
timestamp 1514851247
transform 1 0 52 0 -1 105
box 0 0 32 100
use NOR2X1  NOR2X1_10
timestamp 1514851247
transform -1 0 108 0 -1 105
box 0 0 24 100
use OR2X2  OR2X2_119
timestamp 1514851247
transform 1 0 108 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_158
timestamp 1514851247
transform 1 0 140 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_36
timestamp 1514851247
transform 1 0 172 0 -1 105
box 0 0 24 100
use NAND2X1  NAND2X1_35
timestamp 1514851247
transform -1 0 220 0 -1 105
box 0 0 24 100
use XOR2X1  XOR2X1_9
timestamp 1514851247
transform -1 0 276 0 -1 105
box 0 0 56 100
use AND2X2  AND2X2_10
timestamp 1514851247
transform 1 0 276 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_159
timestamp 1514851247
transform 1 0 308 0 -1 105
box 0 0 32 100
use NAND3X1  NAND3X1_18
timestamp 1514851247
transform -1 0 372 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_4
timestamp 1514851247
transform -1 0 404 0 -1 105
box 0 0 32 100
use INVX1  INVX1_7
timestamp 1514851247
transform 1 0 404 0 -1 105
box 0 0 16 100
use AND2X2  AND2X2_3
timestamp 1514851247
transform 1 0 420 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_7
timestamp 1514851247
transform 1 0 452 0 -1 105
box 0 0 32 100
use NOR3X1  NOR3X1_1
timestamp 1514851247
transform 1 0 484 0 -1 105
box 0 0 64 100
use INVX1  INVX1_5
timestamp 1514851247
transform 1 0 548 0 -1 105
box 0 0 16 100
use BUFX2  BUFX2_43
timestamp 1514851247
transform 1 0 564 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_67
timestamp 1514851247
transform 1 0 588 0 -1 105
box 0 0 24 100
use XOR2X1  XOR2X1_11
timestamp 1514851247
transform 1 0 612 0 -1 105
box 0 0 56 100
use AND2X2  AND2X2_209
timestamp 1514851247
transform -1 0 700 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_10
timestamp 1514851247
transform -1 0 724 0 -1 105
box 0 0 24 100
use INVX1  INVX1_4
timestamp 1514851247
transform 1 0 724 0 -1 105
box 0 0 16 100
use BUFX2  BUFX2_42
timestamp 1514851247
transform 1 0 740 0 -1 105
box 0 0 24 100
use AOI21X1  AOI21X1_17
timestamp 1514851247
transform -1 0 796 0 -1 105
box 0 0 32 100
use BUFX2  BUFX2_66
timestamp 1514851247
transform 1 0 796 0 -1 105
box 0 0 24 100
use NAND2X1  NAND2X1_9
timestamp 1514851247
transform -1 0 844 0 -1 105
box 0 0 24 100
use NAND3X1  NAND3X1_4
timestamp 1514851247
transform 1 0 844 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_8
timestamp 1514851247
transform -1 0 900 0 -1 105
box 0 0 24 100
use AND2X2  AND2X2_205
timestamp 1514851247
transform 1 0 900 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_206
timestamp 1514851247
transform -1 0 964 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_218
timestamp 1514851247
transform -1 0 996 0 -1 105
box 0 0 32 100
use INVX1  INVX1_32
timestamp 1514851247
transform 1 0 996 0 -1 105
box 0 0 16 100
use BUFX2  BUFX2_41
timestamp 1514851247
transform 1 0 1012 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_6
timestamp 1514851247
transform -1 0 1060 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_65
timestamp 1514851247
transform 1 0 1060 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_5
timestamp 1514851247
transform 1 0 1084 0 -1 105
box 0 0 24 100
use AND2X2  AND2X2_165
timestamp 1514851247
transform -1 0 1140 0 -1 105
box 0 0 32 100
use OAI21X1  OAI21X1_8
timestamp 1514851247
transform -1 0 1172 0 -1 105
box 0 0 32 100
use OR2X2  OR2X2_125
timestamp 1514851247
transform -1 0 1204 0 -1 105
box 0 0 32 100
use NAND3X1  NAND3X1_3
timestamp 1514851247
transform 1 0 1204 0 -1 105
box 0 0 32 100
use AND2X2  AND2X2_181
timestamp 1514851247
transform 1 0 1236 0 -1 105
box 0 0 32 100
use OAI21X1  OAI21X1_9
timestamp 1514851247
transform 1 0 1268 0 -1 105
box 0 0 32 100
use OR2X2  OR2X2_144
timestamp 1514851247
transform -1 0 1332 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_5
timestamp 1514851247
transform -1 0 1356 0 -1 105
box 0 0 24 100
use AND2X2  AND2X2_182
timestamp 1514851247
transform 1 0 1356 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_6
timestamp 1514851247
transform -1 0 1412 0 -1 105
box 0 0 24 100
use AOI21X1  AOI21X1_16
timestamp 1514851247
transform 1 0 1412 0 -1 105
box 0 0 32 100
use OR2X2  OR2X2_145
timestamp 1514851247
transform 1 0 1444 0 -1 105
box 0 0 32 100
use OR2X2  OR2X2_152
timestamp 1514851247
transform -1 0 1508 0 -1 105
box 0 0 32 100
use NAND2X1  NAND2X1_7
timestamp 1514851247
transform -1 0 1532 0 -1 105
box 0 0 24 100
use INVX1  INVX1_31
timestamp 1514851247
transform 1 0 1532 0 -1 105
box 0 0 16 100
use BUFX2  BUFX2_40
timestamp 1514851247
transform 1 0 1548 0 -1 105
box 0 0 24 100
use BUFX2  BUFX2_64
timestamp 1514851247
transform 1 0 1572 0 -1 105
box 0 0 24 100
use OR2X2  OR2X2_166
timestamp 1514851247
transform -1 0 1628 0 -1 105
box 0 0 32 100
use INVX1  INVX1_3
timestamp 1514851247
transform -1 0 1644 0 -1 105
box 0 0 16 100
use MUX2X1  MUX2X1_5
timestamp 1514851247
transform 1 0 1644 0 -1 105
box 0 0 48 100
use AND2X2  AND2X2_49
timestamp 1514851247
transform 1 0 1692 0 -1 105
box 0 0 32 100
use MUX2X1  MUX2X1_4
timestamp 1514851247
transform -1 0 1772 0 -1 105
box 0 0 48 100
use AND2X2  AND2X2_70
timestamp 1514851247
transform 1 0 1772 0 -1 105
box 0 0 32 100
use BUFX2  BUFX2_15
timestamp 1514851247
transform -1 0 1828 0 -1 105
box 0 0 24 100
use OR2X2  OR2X2_101
timestamp 1514851247
transform -1 0 1860 0 -1 105
box 0 0 32 100
use FILL  FILL_1_1
timestamp 1514851247
transform -1 0 1868 0 -1 105
box 0 0 8 100
use FILL  FILL_1_2
timestamp 1514851247
transform -1 0 1876 0 -1 105
box 0 0 8 100
use FILL  FILL_1_3
timestamp 1514851247
transform -1 0 1884 0 -1 105
box 0 0 8 100
<< labels >>
flabel metal2 960 1230 960 1230 3 FreeSans 24 90 0 0 ULA_A<0>
port 0 nsew
flabel metal2 824 1230 824 1230 3 FreeSans 24 90 0 0 ULA_A<1>
port 1 nsew
flabel metal2 1000 1230 1000 1230 3 FreeSans 24 90 0 0 ULA_A<2>
port 2 nsew
flabel metal3 -24 1080 -24 1080 7 FreeSans 24 0 0 0 ULA_A<3>
port 3 nsew
flabel metal2 984 1230 984 1230 3 FreeSans 24 90 0 0 ULA_A<4>
port 4 nsew
flabel metal2 1064 1230 1064 1230 3 FreeSans 24 90 0 0 ULA_A<5>
port 5 nsew
flabel metal2 584 1230 584 1230 3 FreeSans 24 90 0 0 ULA_A<6>
port 6 nsew
flabel metal2 624 1230 624 1230 3 FreeSans 24 90 0 0 ULA_A<7>
port 7 nsew
flabel metal3 -24 480 -24 480 7 FreeSans 24 0 0 0 ULA_A<8>
port 8 nsew
flabel metal3 -24 160 -24 160 7 FreeSans 24 0 0 0 ULA_A<9>
port 9 nsew
flabel metal2 1216 -20 1216 -20 7 FreeSans 24 270 0 0 ULA_A<10>
port 10 nsew
flabel metal2 272 -20 272 -20 7 FreeSans 24 270 0 0 ULA_A<11>
port 11 nsew
flabel metal2 1256 -20 1256 -20 7 FreeSans 24 270 0 0 ULA_A<12>
port 12 nsew
flabel metal2 1680 -20 1680 -20 7 FreeSans 24 270 0 0 ULA_A<13>
port 13 nsew
flabel metal2 856 -20 856 -20 7 FreeSans 24 270 0 0 ULA_A<14>
port 14 nsew
flabel metal2 1736 -20 1736 -20 7 FreeSans 24 270 0 0 ULA_A<15>
port 15 nsew
flabel metal2 880 1230 880 1230 3 FreeSans 24 90 0 0 ULA_B<0>
port 16 nsew
flabel metal2 1352 1230 1352 1230 3 FreeSans 24 90 0 0 ULA_B<1>
port 17 nsew
flabel metal2 1432 -20 1432 -20 7 FreeSans 24 270 0 0 ULA_B<2>
port 18 nsew
flabel metal3 -24 1060 -24 1060 7 FreeSans 24 0 0 0 ULA_B<3>
port 19 nsew
flabel metal2 432 -20 432 -20 7 FreeSans 24 270 0 0 ULA_B<4>
port 20 nsew
flabel metal2 208 1230 208 1230 3 FreeSans 24 90 0 0 ULA_B<5>
port 21 nsew
flabel metal2 560 1230 560 1230 3 FreeSans 24 90 0 0 ULA_B<6>
port 22 nsew
flabel metal3 -24 760 -24 760 7 FreeSans 24 0 0 0 ULA_B<7>
port 23 nsew
flabel metal3 -24 340 -24 340 7 FreeSans 24 0 0 0 ULA_B<8>
port 24 nsew
flabel metal3 -24 140 -24 140 7 FreeSans 24 0 0 0 ULA_B<9>
port 25 nsew
flabel metal2 1192 -20 1192 -20 7 FreeSans 24 270 0 0 ULA_B<10>
port 26 nsew
flabel metal2 224 -20 224 -20 7 FreeSans 24 270 0 0 ULA_B<11>
port 27 nsew
flabel metal2 1232 -20 1232 -20 7 FreeSans 24 270 0 0 ULA_B<12>
port 28 nsew
flabel metal2 1512 -20 1512 -20 7 FreeSans 24 270 0 0 ULA_B<13>
port 29 nsew
flabel metal2 880 -20 880 -20 7 FreeSans 24 270 0 0 ULA_B<14>
port 30 nsew
flabel metal2 704 -20 704 -20 7 FreeSans 24 270 0 0 ULA_B<15>
port 31 nsew
flabel metal2 968 -20 968 -20 7 FreeSans 24 270 0 0 ULA_ctrl<0>
port 32 nsew
flabel metal2 504 -20 504 -20 7 FreeSans 24 270 0 0 ULA_ctrl<1>
port 33 nsew
flabel metal2 352 -20 352 -20 7 FreeSans 24 270 0 0 ULA_ctrl<2>
port 34 nsew
flabel metal2 528 -20 528 -20 7 FreeSans 24 270 0 0 ULA_ctrl<3>
port 35 nsew
flabel metal3 1912 260 1912 260 3 FreeSans 24 0 0 0 ULA_OUT<0>
port 36 nsew
flabel metal2 104 1230 104 1230 3 FreeSans 24 90 0 0 ULA_OUT<1>
port 37 nsew
flabel metal2 344 1230 344 1230 3 FreeSans 24 90 0 0 ULA_OUT<2>
port 38 nsew
flabel metal3 -24 860 -24 860 7 FreeSans 24 0 0 0 ULA_OUT<3>
port 39 nsew
flabel metal2 744 1230 744 1230 3 FreeSans 24 90 0 0 ULA_OUT<4>
port 40 nsew
flabel metal3 -24 960 -24 960 7 FreeSans 24 0 0 0 ULA_OUT<5>
port 41 nsew
flabel metal3 -24 880 -24 880 7 FreeSans 24 0 0 0 ULA_OUT<6>
port 42 nsew
flabel metal3 -24 780 -24 780 7 FreeSans 24 0 0 0 ULA_OUT<7>
port 43 nsew
flabel metal3 -24 560 -24 560 7 FreeSans 24 0 0 0 ULA_OUT<8>
port 44 nsew
flabel metal3 -24 60 -24 60 7 FreeSans 24 270 0 0 ULA_OUT<9>
port 45 nsew
flabel metal3 -24 260 -24 260 7 FreeSans 24 0 0 0 ULA_OUT<10>
port 46 nsew
flabel metal3 -24 460 -24 460 7 FreeSans 24 0 0 0 ULA_OUT<11>
port 47 nsew
flabel metal2 1592 -20 1592 -20 7 FreeSans 24 270 0 0 ULA_OUT<12>
port 48 nsew
flabel metal2 1080 -20 1080 -20 7 FreeSans 24 270 0 0 ULA_OUT<13>
port 49 nsew
flabel metal2 816 -20 816 -20 7 FreeSans 24 270 0 0 ULA_OUT<14>
port 50 nsew
flabel metal2 608 -20 608 -20 7 FreeSans 24 270 0 0 ULA_OUT<15>
port 51 nsew
flabel metal2 56 1230 56 1230 7 FreeSans 24 90 0 0 ULA_flags<0>
port 52 nsew
flabel metal3 -24 660 -24 660 7 FreeSans 24 0 0 0 ULA_flags<1>
port 53 nsew
flabel metal3 -24 1160 -24 1160 7 FreeSans 24 90 0 0 ULA_flags<2>
port 54 nsew
<< end >>
