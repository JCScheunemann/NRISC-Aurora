module NRISC_ULA ( gnd, vdd, ULA_A, ULA_B, ULA_ctrl, ULA_OUT, ULA_flags);

input gnd, vdd;
input [15:0] ULA_A;
input [15:0] ULA_B;
input [3:0] ULA_ctrl;
output [15:0] ULA_OUT;
output [2:0] ULA_flags;

AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_322_), .Y(_323_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_350_), .Y(_351_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(ULA_ctrl[3]), .Y(_451_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_430_), .Y(_462_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .B(ULA_ctrl[1]), .Y(_494_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(ULA_ctrl[3]), .Y(_514_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(ULA_ctrl[2]), .Y(_515_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .B(ULA_ctrl[3]), .Y(_536_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_536_), .Y(_547_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_494_), .Y(_568_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(ULA_ctrl_0_bF_buf2), .Y(_603_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(ULA_ctrl_0_bF_buf2), .Y(_605_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_351_), .Y(_352_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_607_), .Y(_610_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_611_), .Y(_612_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(ULA_ctrl_0_bF_buf2), .Y(_615_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf0), .B(_617_), .Y(_618_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_606_), .Y(_620_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf0), .B(_622_), .Y(_623_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_624_), .Y(_0_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_621_), .Y(_2_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_604_), .Y(_4_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(ULA_ctrl_0_bF_buf2), .Y(_7_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_334_), .Y(_353_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_9_), .Y(_12_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_15_), .Y(_23_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_26_), .Y(_27_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_30__bF_buf1), .Y(_31_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(ULA_B_1_bF_buf0), .Y(_32_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(ULA_B_2_bF_buf3), .Y(_34_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(ULA_B_1_bF_buf5), .Y(_36_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_30__bF_buf3), .Y(_37_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_35_), .Y(_39_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(ULA_B_1_bF_buf3), .Y(_42_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_355_), .Y(_356_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_30__bF_buf0), .Y(_43_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(ULA_B_1_bF_buf3), .Y(_47_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_30__bF_buf4), .Y(_48_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_45_), .Y(_51_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_51_), .Y(_52_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_597_), .Y(_57_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_595__bF_buf0), .Y(_63_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_58_), .Y(_64_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_64_), .Y(_65_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_65_), .Y(_66_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_362_), .Y(_363_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(ULA_A[15]), .Y(_68_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(ULA_B_1_bF_buf5), .Y(_69_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(ULA_A[13]), .Y(_70_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(ULA_A[14]), .Y(_71_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf1), .B(_72_), .Y(_73_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_606_), .Y(_75_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_621_), .Y(_79_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_621_), .Y(_85_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_606_), .Y(_89_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_13_), .Y(_92_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_595__bF_buf2), .B(_363_), .Y(_364_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_81_), .Y(_93_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_96_), .Y(_97_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(ULA_B_2_bF_buf0), .Y(_98_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(ULA_B_1_bF_buf5), .Y(_99_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_30__bF_buf3), .Y(_100_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_35_), .Y(_102_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_27_), .Y(_110_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_105_), .Y(_111_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_111_), .Y(_112_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_114_), .Y(_115_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_358_), .Y(_365_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_127_), .Y(_625__1_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(ULA_A[14]), .Y(_131_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(ULA_A[15]), .Y(_132_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf1), .B(_133_), .Y(_134_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_135_), .Y(_138_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_621_), .Y(_141_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_606_), .Y(_143_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_13_), .Y(_146_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_139_), .Y(_147_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(ULA_B_2_bF_buf0), .Y(_149_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(ULA_B_1_bF_buf1), .Y(_372_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(ULA_B_1_bF_buf5), .Y(_150_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_30__bF_buf1), .Y(_151_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_35_), .Y(_153_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_27_), .Y(_161_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_157_), .Y(_162_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_162_), .Y(_163_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_165_), .Y(_167_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_128_), .Y(_171_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_175_), .Y(_625__2_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_604_), .Y(_182_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_30__bF_buf4), .Y(_374_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_86_), .Y(_183_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf2), .B(_83_), .Y(_184_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf2), .B(_87_), .Y(_187_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_76_), .Y(_188_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_186_), .Y(_191_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_15_), .Y(_192_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(ULA_B_1_bF_buf5), .Y(_195_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_30__bF_buf3), .Y(_196_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_178_), .Y(_199_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(ULA_B[3]), .Y(_200_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_371_), .Y(_377_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_106_), .Y(_203_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_201_), .Y(_204_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_30__bF_buf4), .Y(_206_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(ULA_B_1_bF_buf2), .Y(_207_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_205_), .Y(_209_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(ULA_B_1_bF_buf4), .Y(_213_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_30__bF_buf2), .Y(_215_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_220_), .Y(_221_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_595__bF_buf2), .Y(_223_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_218_), .Y(_224_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_323_), .Y(_324_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_370_), .Y(_378_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_224_), .Y(_225_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_225_), .Y(_226_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_606_), .Y(_233_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf3), .B(_19_), .Y(_234_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_20_), .Y(_235_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_621_), .Y(_237_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_232_), .Y(_240_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(ULA_B[3]), .Y(_243_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_106_), .Y(_244_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_205_), .Y(_245_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_379_), .Y(_380_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_251_), .Y(_255_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(ULA_B_2_bF_buf1), .Y(_257_) );
AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(ULA_B_1_bF_buf1), .Y(_258_) );
AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_30__bF_buf0), .Y(_260_) );
AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_35_), .Y(_262_) );
AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_255_), .Y(_265_) );
AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_265_), .Y(_266_) );
AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_266_), .Y(_267_) );
AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_270_), .Y(_271_) );
AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_272_), .Y(_275_) );
AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_365_), .Y(_381_) );
AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(ULA_B_2_bF_buf2), .Y(_286_) );
AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(ULA_B_1_bF_buf4), .Y(_287_) );
AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_30__bF_buf2), .Y(_289_) );
AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_35_), .Y(_291_) );
AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_293_), .Y(_294_) );
AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_294_), .Y(_295_) );
AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_276_), .Y(_296_) );
AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_298_), .Y(_299_) );
AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_300_), .Y(_303_) );
AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(ULA_B_2_bF_buf1), .Y(_315_) );
AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_606_), .Y(_388_) );
AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(ULA_B_1_bF_buf1), .Y(_316_) );
AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_30__bF_buf2), .Y(_318_) );
AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_35_), .Y(_320_) );
AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_616__bF_buf1), .B(_76_), .Y(_389_) );
AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_77_), .Y(_390_) );
AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_621_), .Y(_392_) );
AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(ULA_B_1_bF_buf4), .Y(_396_) );
AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_30__bF_buf4), .Y(_398_) );
AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_401_), .Y(_402_) );
AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_324_), .Y(_325_) );
AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_395_), .Y(_403_) );
AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_410_), .Y(_411_) );
AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_595__bF_buf3), .B(_411_), .Y(_412_) );
AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_412_), .Y(_413_) );
AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_404_), .Y(_414_) );
AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_394_), .Y(_415_) );
AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_422_), .Y(_427_) );
AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_432_), .Y(_433_) );
AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_595__bF_buf0), .Y(_435_) );
AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_429_), .Y(_436_) );
AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_327_), .Y(_328_) );
AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_436_), .Y(_437_) );
AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_421_), .Y(_438_) );
AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(ULA_B_1_bF_buf2), .Y(_445_) );
AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_30__bF_buf3), .Y(_447_) );
AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_452_), .Y(_453_) );
AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_444_), .Y(_454_) );
AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_460_), .Y(_461_) );
AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_595__bF_buf3), .B(_461_), .Y(_463_) );
AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_456_), .Y(_464_) );
AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_464_), .Y(_465_) );
AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_331_), .Y(_333_) );
AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_443_), .Y(_466_) );
AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_473_), .Y(_478_) );
AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_486_), .Y(_487_) );
AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_595__bF_buf2), .Y(_489_) );
AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_484_), .Y(_490_) );
AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_482_), .Y(_491_) );
AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_491_), .Y(_492_) );
AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_30__bF_buf1), .Y(_501_) );
AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(ULA_B_1_bF_buf2), .Y(_502_) );
AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_504_), .Y(_505_) );
AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(ULA_B_2_bF_buf2), .Y(_343_) );
AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_505_), .Y(_506_) );
AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_510_), .Y(_511_) );
AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_512_), .Y(_513_) );
AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_516_), .Y(_517_) );
AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_517_), .Y(_518_) );
AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_520_), .Y(_521_) );
AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_30__bF_buf3), .Y(_529_) );
AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(ULA_B_1_bF_buf2), .Y(_530_) );
AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(ULA_B_1_bF_buf1), .Y(_533_) );
AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_30__bF_buf4), .Y(_534_) );
AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(ULA_B_1_bF_buf4), .Y(_344_) );
AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_532_), .Y(_538_) );
AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_538_), .Y(_539_) );
AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_544_), .Y(_546_) );
AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_541_), .Y(_548_) );
AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_595__bF_buf0), .Y(_549_) );
AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_551_), .Y(_552_) );
AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_552_), .Y(_553_) );
AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_357_), .Y(_556_) );
AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_561_), .Y(_562_) );
AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_177_), .Y(_565_) );
AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_30__bF_buf2), .Y(_346_) );
AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_566_), .Y(_569_) );
AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(ULA_B_2_bF_buf3), .Y(_570_) );
AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_563_), .Y(_573_) );
AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_559_), .Y(_574_) );
AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_557_), .Y(_575_) );
AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_577_), .Y(_578_) );
AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_521_), .Y(_579_) );
AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_578_), .Y(_580_) );
AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_580_), .Y(_581_) );
AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_67_), .Y(_582_) );
AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_35_), .Y(_348_) );
AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_386_), .Y(_583_) );
AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_471_), .Y(_584_) );
AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_583_), .Y(_585_) );
AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_585_), .Y(_586_) );
AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_271_), .Y(_590_) );
AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_590_), .Y(_591_) );
AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_591_), .Y(_592_) );
AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_328_), .Y(_593_) );
AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_356_), .Y(_594_) );
AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_594_), .Y(zero) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_189_), .C(_604_), .Y(_332_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_30__bF_buf1), .C(ULA_B_2_bF_buf3), .Y(_566_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_599_), .C(_595__bF_buf1), .Y(_600_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(_128_), .C(_595__bF_buf1), .Y(_129_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_180_), .C(_179_), .Y(_181_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(_595__bF_buf2), .Y(_229_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_101_), .C(_28_), .Y(_280_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_283_), .C(_472_), .Y(_284_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_312_), .C(_472_), .Y(_313_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_340_), .C(_472_), .Y(_341_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_384_), .C(_595__bF_buf2), .Y(_385_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_616__bF_buf1), .C(_69_), .Y(_387_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_418_), .C(_595__bF_buf3), .Y(_419_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_440_), .C(_595__bF_buf0), .Y(_441_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_469_), .C(_595__bF_buf3), .Y(_470_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_495_), .C(_595__bF_buf2), .Y(_496_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_524_), .C(_595__bF_buf3), .Y(_526_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_425_), .C(_205_), .D(_423_), .Y(_426_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_476_), .C(_474_), .D(_205_), .Y(_477_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_124_), .C(_130_), .D(_175_), .Y(_587_) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf5) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf1) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf0) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf3) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf2) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf1) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf0) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf3) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf2) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf1) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf0) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf4) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_616_), .Y(_616__bF_buf3) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_616_), .Y(_616__bF_buf2) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_616_), .Y(_616__bF_buf1) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_616_), .Y(_616__bF_buf0) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_595_), .Y(_595__bF_buf3) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_595_), .Y(_595__bF_buf2) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_595_), .Y(_595__bF_buf1) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_595_), .Y(_595__bF_buf0) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf5) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf4) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf3) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf3) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf2) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf1) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf0) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_625__0_), .Y(_625__0_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_625__1_), .Y(_625__1_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_625__2_), .Y(_625__2_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_625__3_), .Y(_625__3_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_625__4_), .Y(_625__4_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_625__5_), .Y(_625__5_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf2) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_625__6_), .Y(_625__6_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_625__7_), .Y(_625__7_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_625__8_), .Y(_625__8_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_625__9_), .Y(_625__9_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_625__10_), .Y(_625__10_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_625__11_), .Y(_625__11_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_625__12_), .Y(_625__12_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_625__13_), .Y(_625__13_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_625__14_), .Y(_625__14_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_625__15_), .Y(_625__15_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf1) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_626__0_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(zero), .Y(_626__1_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(_626__2_) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf0) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf4) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf3) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_30__bF_buf2) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_328_), .Y(_625__6_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_542_), .Y(_543_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_550_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_554_), .Y(_625__14_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_625__15_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .Y(_430_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(_450_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[3]), .Y(_567_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .Y(_596_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_607_), .Y(_613_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_606_), .Y(_621_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_356_), .Y(_625__7_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_14_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_604_), .Y(_15_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[4]), .Y(_26_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(_29_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .Y(_35_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .Y(_54_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf4), .Y(_55_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(_60_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_625__0_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_386_), .Y(_625__8_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(_106_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_595__bF_buf1), .Y(_125_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .Y(_176_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_178_), .Y(_179_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_230_), .Y(_625__3_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_271_), .Y(_625__4_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_299_), .Y(_625__5_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_420_), .Y(_625__9_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_442_), .Y(_625__10_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_471_), .Y(_625__11_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_375_), .Y(_474_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_497_), .Y(_625__12_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_521_), .Y(_625__13_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf1), .Y(_30_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_A[7]), .S(ULA_B_0_bF_buf0), .Y(_345_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_A[13]), .S(ULA_B_0_bF_buf5), .Y(_500_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_A[14]), .S(ULA_B_0_bF_buf5), .Y(_528_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .B(ULA_A[14]), .S(ULA_B_0_bF_buf5), .Y(_611_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_A[12]), .S(ULA_B_0_bF_buf5), .Y(_617_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_A[8]), .S(ULA_B_0_bF_buf3), .Y(_622_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_A[10]), .S(ULA_B_0_bF_buf1), .Y(_624_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_A[0]), .S(ULA_B_0_bF_buf2), .Y(_16_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_A[2]), .S(ULA_B_0_bF_buf2), .Y(_17_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .S(_616__bF_buf3), .Y(_18_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_A[4]), .S(ULA_B_0_bF_buf2), .Y(_19_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_A[8]), .S(ULA_B_0_bF_buf4), .Y(_373_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_A[6]), .S(ULA_B_0_bF_buf4), .Y(_20_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_20_), .S(_616__bF_buf3), .Y(_21_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_18_), .S(_606_), .Y(_22_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_A[9]), .S(ULA_B_0_bF_buf3), .Y(_76_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_A[11]), .S(ULA_B_0_bF_buf1), .Y(_77_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .S(_616__bF_buf2), .Y(_78_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_A[1]), .S(ULA_B_0_bF_buf2), .Y(_82_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_A[3]), .S(ULA_B_0_bF_buf2), .Y(_83_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_83_), .S(_616__bF_buf3), .Y(_84_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_A[5]), .S(ULA_B_0_bF_buf4), .Y(_86_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_A[9]), .S(ULA_B_0_bF_buf4), .Y(_397_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_A[7]), .S(ULA_B_0_bF_buf4), .Y(_87_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .S(_616__bF_buf2), .Y(_88_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_A[13]), .S(ULA_B_0_bF_buf5), .Y(_95_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_86_), .S(ULA_B_1_bF_buf2), .Y(_104_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .B(ULA_A[1]), .S(ULA_B_0_bF_buf0), .Y(_117_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_617_), .S(_616__bF_buf0), .Y(_136_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_19_), .S(_616__bF_buf3), .Y(_140_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_622_), .S(_616__bF_buf2), .Y(_142_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_20_), .S(ULA_B_1_bF_buf2), .Y(_156_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_A[2]), .S(ULA_B_0_bF_buf2), .Y(_164_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_259_), .S(_30__bF_buf2), .Y(_423_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_95_), .S(_616__bF_buf0), .Y(_180_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_A[3]), .S(ULA_B_0_bF_buf0), .Y(_214_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_A[4]), .S(ULA_B_0_bF_buf0), .Y(_259_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_88_), .S(_606_), .Y(_273_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_A[5]), .S(ULA_B_0_bF_buf0), .Y(_288_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_142_), .S(_606_), .Y(_301_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_A[6]), .S(ULA_B_0_bF_buf0), .Y(_317_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_A[10]), .S(ULA_B_0_bF_buf1), .Y(_424_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_373_), .S(_30__bF_buf4), .Y(_425_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_A[11]), .S(ULA_B_0_bF_buf3), .Y(_446_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_A[12]), .S(ULA_B_0_bF_buf3), .Y(_475_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_424_), .S(_30__bF_buf3), .Y(_476_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_125_), .Y(_327_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_432_), .Y(_439_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_B[11]), .Y(_467_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_467_), .Y(_468_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_B[12]), .Y(_486_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_486_), .Y(_493_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_B[13]), .Y(_510_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_B[14]), .Y(_522_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_522_), .Y(_523_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .B(ULA_B[15]), .Y(_561_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .B(ULA_B_0_bF_buf3), .Y(_597_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_B[7]), .Y(_340_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_597_), .Y(_598_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .B(_29_), .Y(_46_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_55_), .Y(_56_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_B_1_bF_buf4), .Y(_114_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_125_), .Y(_127_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_B_2_bF_buf2), .Y(_128_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .B(_154_), .Y(_155_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_B[3]), .Y(_220_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_220_), .Y(_227_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_B[4]), .Y(_253_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_125_), .Y(_355_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_253_), .Y(_268_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .B(_277_), .Y(_278_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_B[5]), .Y(_283_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_125_), .Y(_298_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .B(_306_), .Y(_307_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_152_), .Y(_308_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_307_), .Y(_309_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_B[6]), .Y(_312_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_525_), .Y(_369_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_B[8]), .Y(_382_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_382_), .Y(_383_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_B[9]), .Y(_416_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_416_), .Y(_417_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_B[10]), .Y(_432_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_30__bF_buf1), .C(_35_), .Y(_329_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(ULA_A[11]), .C(ULA_B[11]), .Y(_469_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(ULA_A[12]), .C(ULA_B[12]), .Y(_495_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(ULA_A[14]), .C(ULA_B[14]), .Y(_524_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_522_), .C(_542_), .Y(_545_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(ULA_B[3]), .C(_26_), .Y(_558_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(ULA_A[0]), .C(ULA_B_0_bF_buf3), .Y(_599_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .B(ULA_ctrl[1]), .C(ULA_ctrl[3]), .Y(_9_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_515_), .C(_61_), .Y(_62_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(ULA_B_1_bF_buf0), .C(ULA_A[15]), .Y(_94_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_106_), .C(_108_), .Y(_109_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_430_), .C(_536_), .Y(_357_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_595__bF_buf1), .C(_121_), .Y(_122_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_106_), .C(_159_), .Y(_160_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(ULA_A[0]), .C(ULA_B_1_bF_buf3), .Y(_166_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_595__bF_buf1), .C(_172_), .Y(_173_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(ULA_A[3]), .C(ULA_B[3]), .Y(_228_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(ULA_ctrl[2]), .C(_567_), .Y(_249_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_252_), .C(_253_), .Y(_254_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(ULA_A[0]), .C(_30__bF_buf2), .Y(_256_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(ULA_A[4]), .C(ULA_B[4]), .Y(_269_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_268_), .C(_269_), .Y(_270_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_494_), .C(_567_), .Y(_362_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_604_), .C(_621_), .Y(_272_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_279_), .C(_280_), .Y(_281_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_604_), .C(_134_), .Y(_300_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(ULA_A[8]), .C(ULA_B[8]), .Y(_384_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_494_), .C(_567_), .Y(_410_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(ULA_A[9]), .C(ULA_B[9]), .Y(_418_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_15_), .C(_13_), .Y(_421_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(ULA_A[10]), .C(ULA_B[10]), .Y(_440_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_494_), .C(_567_), .Y(_460_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_29_), .Y(_330_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(ULA_B[3]), .Y(_205_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_B[4]), .Y(_250_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_B[5]), .Y(_282_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_B[6]), .Y(_311_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_46_), .Y(_335_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_5_), .Y(_336_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_B[7]), .Y(_339_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_B[8]), .Y(_359_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_B[9]), .Y(_407_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_B[11]), .Y(_457_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_8_), .Y(_13_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .B(ULA_B[4]), .Y(_61_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(ULA_ctrl[1]), .C(ULA_ctrl[3]), .Y(_472_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_333_), .C(_13_), .Y(_334_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_515_), .C(_61_), .Y(_120_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(_128_), .C(_129_), .Y(_130_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_472_), .C(_170_), .Y(_172_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_472_), .C(_219_), .Y(_222_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_156_), .C(_27_), .Y(_305_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_337_), .C(_27_), .Y(_338_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_472_), .C(_431_), .Y(_434_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_472_), .C(_485_), .Y(_488_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_472_), .C(_509_), .Y(_512_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_472_), .C(_560_), .Y(_563_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_472_), .C(_56_), .Y(_58_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_98_), .C(ULA_B[3]), .Y(_103_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_472_), .C(_113_), .Y(_116_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_321_), .Y(_322_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_8_), .Y(_366_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .Y(_33_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .Y(_38_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_39_), .Y(_40_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_40_), .Y(_41_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_43_), .Y(_44_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .Y(_45_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .Y(_49_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_49_), .Y(_50_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_52_), .Y(_53_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_602_), .Y(_59_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_366_), .Y(_367_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_66_), .Y(_67_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_70_), .Y(_72_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_73_), .Y(_74_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_75_), .Y(_80_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_80_), .Y(_81_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_89_), .Y(_90_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_90_), .Y(_91_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf0), .B(_95_), .Y(_96_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_101_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_104_), .Y(_105_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_3_), .Y(_368_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf3), .B(_82_), .Y(_107_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_30__bF_buf0), .B(_83_), .Y(_108_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_B_1_bF_buf4), .Y(_113_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf4), .B(_117_), .Y(_118_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf2), .B(_118_), .Y(_119_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_120_), .Y(_121_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_122_), .Y(_123_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_93_), .Y(_124_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_131_), .Y(_133_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_621_), .Y(_135_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_261_), .Y(_370_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_136_), .Y(_137_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_138_), .Y(_139_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .Y(_144_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_144_), .Y(_145_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf0), .B(_611_), .Y(_148_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .Y(_152_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_153_), .Y(_154_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_156_), .Y(_157_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf3), .B(_17_), .Y(_158_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_30__bF_buf0), .B(_19_), .Y(_159_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_59_), .Y(_371_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf1), .B(_164_), .Y(_165_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .B(_167_), .Y(_168_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_168_), .Y(_169_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_B_2_bF_buf2), .Y(_170_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_163_), .Y(_174_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_174_), .Y(_175_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_176_), .Y(_177_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_177_), .Y(_178_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_184_), .Y(_185_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_185_), .Y(_186_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_374_), .Y(_375_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .Y(_189_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_189_), .Y(_190_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_192_), .Y(_193_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_193_), .Y(_194_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .Y(_197_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf3), .B(_197_), .Y(_198_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf3), .B(_83_), .Y(_201_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_30__bF_buf0), .B(_86_), .Y(_202_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_207_), .Y(_208_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_209_), .Y(_210_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_375_), .Y(_376_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_210_), .Y(_211_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_211_), .Y(_212_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_215_), .Y(_216_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf2), .B(_216_), .Y(_217_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_120_), .Y(_218_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_B[3]), .Y(_219_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_226_), .Y(_230_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_619_), .Y(_231_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_231_), .Y(_232_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_235_), .Y(_236_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_378_), .Y(_379_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_237_), .Y(_238_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_238_), .Y(_239_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_240_), .Y(_241_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf3), .B(_33_), .Y(_242_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_245_), .Y(_246_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_246_), .Y(_247_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_247_), .Y(_248_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_249_), .Y(_251_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_B[4]), .Y(_252_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_260_), .Y(_261_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_381_), .Y(_386_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_262_), .Y(_263_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_263_), .Y(_264_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_273_), .Y(_274_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_275_), .Y(_276_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf0), .B(_97_), .Y(_277_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_104_), .Y(_279_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_284_), .Y(_285_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_289_), .Y(_290_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_291_), .Y(_292_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_292_), .Y(_293_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_390_), .Y(_391_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_301_), .Y(_302_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_303_), .Y(_304_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf0), .B(_148_), .Y(_306_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_309_), .Y(_310_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_313_), .Y(_314_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_318_), .Y(_319_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_315_), .Y(_321_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_180_), .Y(_331_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_388_), .Y(_393_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_393_), .Y(_394_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_119_), .Y(_395_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_398_), .Y(_399_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_399_), .Y(_400_) );
OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_290_), .Y(_401_) );
OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_403_), .Y(_404_) );
OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_98_), .Y(_405_) );
OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_405_), .Y(_406_) );
OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_249_), .Y(_408_) );
OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_330_), .Y(_337_) );
OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_415_), .Y(_420_) );
OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_168_), .Y(_422_) );
OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_427_), .Y(_428_) );
OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_154_), .Y(_429_) );
OR2X2 OR2X2_125 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_B[10]), .Y(_431_) );
OR2X2 OR2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_438_), .Y(_442_) );
OR2X2 OR2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_181_), .Y(_443_) );
OR2X2 OR2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_217_), .Y(_444_) );
OR2X2 OR2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_447_), .Y(_448_) );
OR2X2 OR2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_448_), .Y(_449_) );
OR2X2 OR2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_341_), .Y(_342_) );
OR2X2 OR2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_347_), .Y(_452_) );
OR2X2 OR2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_454_), .Y(_455_) );
OR2X2 OR2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_199_), .Y(_456_) );
OR2X2 OR2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_249_), .Y(_458_) );
OR2X2 OR2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_466_), .Y(_471_) );
OR2X2 OR2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_263_), .Y(_473_) );
OR2X2 OR2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_478_), .Y(_479_) );
OR2X2 OR2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_12_), .Y(_480_) );
OR2X2 OR2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_480_), .Y(_481_) );
OR2X2 OR2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_481_), .Y(_482_) );
OR2X2 OR2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_346_), .Y(_347_) );
OR2X2 OR2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_242_), .Y(_484_) );
OR2X2 OR2X2_144 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_B[12]), .Y(_485_) );
OR2X2 OR2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_492_), .Y(_497_) );
OR2X2 OR2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_292_), .Y(_498_) );
OR2X2 OR2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_399_), .Y(_499_) );
OR2X2 OR2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_502_), .Y(_503_) );
OR2X2 OR2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_503_), .Y(_504_) );
OR2X2 OR2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_506_), .Y(_507_) );
OR2X2 OR2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_277_), .Y(_508_) );
OR2X2 OR2X2_152 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_B[13]), .Y(_509_) );
OR2X2 OR2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_348_), .Y(_349_) );
OR2X2 OR2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_481_), .Y(_516_) );
OR2X2 OR2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_595__bF_buf0), .Y(_520_) );
OR2X2 OR2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_321_), .Y(_527_) );
OR2X2 OR2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_530_), .Y(_531_) );
OR2X2 OR2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_531_), .Y(_532_) );
OR2X2 OR2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_534_), .Y(_535_) );
OR2X2 OR2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_535_), .Y(_537_) );
OR2X2 OR2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_539_), .Y(_540_) );
OR2X2 OR2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_357_), .Y(_541_) );
OR2X2 OR2X2_163 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_B[14]), .Y(_542_) );
OR2X2 OR2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_349_), .Y(_350_) );
OR2X2 OR2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_249_), .Y(_544_) );
OR2X2 OR2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_550_), .Y(_551_) );
OR2X2 OR2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_553_), .Y(_554_) );
OR2X2 OR2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_366_), .Y(_555_) );
OR2X2 OR2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_556_), .Y(_557_) );
OR2X2 OR2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_558_), .Y(_559_) );
OR2X2 OR2X2_171 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .B(ULA_B[15]), .Y(_560_) );
OR2X2 OR2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_30__bF_buf1), .B(_500_), .Y(_564_) );
OR2X2 OR2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_569_), .Y(_571_) );
OR2X2 OR2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_571_), .Y(_572_) );
OR2X2 OR2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_40_), .Y(_358_) );
OR2X2 OR2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_595__bF_buf3), .Y(_577_) );
OR2X2 OR2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_472_), .Y(_483_) );
OR2X2 OR2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_515_), .Y(_525_) );
OR2X2 OR2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_568_), .Y(_588_) );
OR2X2 OR2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_525_), .Y(_589_) );
OR2X2 OR2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_483_), .Y(_595_) );
OR2X2 OR2X2_182 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf5), .B(ULA_B_1_bF_buf0), .Y(_601_) );
OR2X2 OR2X2_183 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf3), .B(_601_), .Y(_602_) );
OR2X2 OR2X2_184 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_B_1_bF_buf5), .Y(_607_) );
OR2X2 OR2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_608_), .Y(_609_) );
OR2X2 OR2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_249_), .Y(_360_) );
OR2X2 OR2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_615_), .Y(_616_) );
OR2X2 OR2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_612_), .Y(_619_) );
OR2X2 OR2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_0_), .Y(_1_) );
OR2X2 OR2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_2_), .Y(_3_) );
OR2X2 OR2X2_191 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .B(ULA_B[3]), .Y(_5_) );
OR2X2 OR2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_5_), .Y(_6_) );
OR2X2 OR2X2_193 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .B(_567_), .Y(_10_) );
OR2X2 OR2X2_194 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .B(_10_), .Y(_11_) );
OR2X2 OR2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_23_), .Y(_24_) );
OR2X2 OR2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_24_), .Y(_25_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(ULA_B_1_bF_buf5), .Y(_614_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_312_), .Y(_326_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf5), .B(ULA_B_1_bF_buf0), .Y(_608_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[4]), .B(_7_), .Y(_8_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(_114_), .Y(_126_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_283_), .Y(_297_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_340_), .Y(_354_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_B[8]), .Y(_361_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_B[9]), .Y(_409_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_B[11]), .Y(_459_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(_510_), .Y(_519_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(_561_), .Y(_576_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .B(_603_), .Y(_604_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf0), .B(_605_), .Y(_606_) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_625__0_), .Y(ULA_OUT[0]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_625__1_), .Y(ULA_OUT[1]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_625__2_), .Y(ULA_OUT[2]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_625__3_), .Y(ULA_OUT[3]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_625__4_), .Y(ULA_OUT[4]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_625__5_), .Y(ULA_OUT[5]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_625__6_), .Y(ULA_OUT[6]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_625__7_), .Y(ULA_OUT[7]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_625__8_), .Y(ULA_OUT[8]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_625__9_), .Y(ULA_OUT[9]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_625__10_), .Y(ULA_OUT[10]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_625__11_), .Y(ULA_OUT[11]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_625__12_), .Y(ULA_OUT[12]) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_625__13_), .Y(ULA_OUT[13]) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(_625__14_), .Y(ULA_OUT[14]) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_625__15_), .Y(ULA_OUT[15]) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(_626__0_), .Y(ULA_flags[0]) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(_626__1_), .Y(ULA_flags[1]) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(_626__2_), .Y(ULA_flags[2]) );
endmodule
