module NRISC_PC_ctrl (IDATA_CORE_out, CORE_PC_ctrl, CORE_STACK_ctrl, ULA_OUT, INTERRUPT_ch, INTERRUPT_flag, clk, rst, IDATA_CORE_addr, IDATA_clk, CORE_InstructionIN, REG_R0);

input INTERRUPT_flag;
input clk;
input rst;
output IDATA_clk;
input [15:0] IDATA_CORE_out;
input [1:0] CORE_PC_ctrl;
input [1:0] CORE_STACK_ctrl;
input [9:0] ULA_OUT;
input [7:0] INTERRUPT_ch;
output [9:0] IDATA_CORE_addr;
output [15:0] CORE_InstructionIN;
output [9:0] REG_R0;

wire vdd = 1'b1;
wire gnd = 1'b0;

AND2X2 AND2X2_1 ( .A(PC_pointer_0_), .B(PC_pointer_1_), .Y(_1012_) );
AND2X2 AND2X2_2 ( .A(_1314_), .B(_1308_), .Y(_1315_) );
AND2X2 AND2X2_3 ( .A(_1359_), .B(_1360_), .Y(_1361_) );
AND2X2 AND2X2_4 ( .A(_1363_), .B(_1362_), .Y(_1364_) );
AND2X2 AND2X2_5 ( .A(_1364_), .B(_1361_), .Y(_1365_) );
AND2X2 AND2X2_6 ( .A(_1274_), .B(_992__bF_buf0), .Y(_1420_) );
AND2X2 AND2X2_7 ( .A(_1434_), .B(_1430_), .Y(_1435_) );
AND2X2 AND2X2_8 ( .A(_1274_), .B(_1022_), .Y(_1494_) );
AND2X2 AND2X2_9 ( .A(_1508_), .B(_1505_), .Y(_1509_) );
AND2X2 AND2X2_10 ( .A(_1274_), .B(_1023_), .Y(_43_) );
AND2X2 AND2X2_11 ( .A(_55_), .B(_52_), .Y(_56_) );
AND2X2 AND2X2_12 ( .A(PC_pointer_2_), .B(PC_pointer_3_), .Y(_1079_) );
AND2X2 AND2X2_13 ( .A(_83_), .B(_86_), .Y(_87_) );
AND2X2 AND2X2_14 ( .A(_75_), .B(_1095__bF_buf2), .Y(_88_) );
AND2X2 AND2X2_15 ( .A(_89_), .B(_91_), .Y(_92_) );
AND2X2 AND2X2_16 ( .A(_1274_), .B(_1104_), .Y(_139_) );
AND2X2 AND2X2_17 ( .A(_151_), .B(_148_), .Y(_152_) );
AND2X2 AND2X2_18 ( .A(_1274_), .B(_1003_), .Y(_210_) );
AND2X2 AND2X2_19 ( .A(_222_), .B(_219_), .Y(_223_) );
AND2X2 AND2X2_20 ( .A(_1274_), .B(_997__bF_buf0), .Y(_282_) );
AND2X2 AND2X2_21 ( .A(_294_), .B(_291_), .Y(_295_) );
AND2X2 AND2X2_22 ( .A(_1274_), .B(_1000__bF_buf0), .Y(_355_) );
AND2X2 AND2X2_23 ( .A(_1192_), .B(_1193_), .Y(_1194_) );
AND2X2 AND2X2_24 ( .A(_367_), .B(_364_), .Y(_368_) );
AND2X2 AND2X2_25 ( .A(_1274_), .B(_1004__bF_buf1), .Y(_428_) );
AND2X2 AND2X2_26 ( .A(_440_), .B(_437_), .Y(_441_) );
AND2X2 AND2X2_27 ( .A(_1274_), .B(_1026_), .Y(_499_) );
AND2X2 AND2X2_28 ( .A(_511_), .B(_508_), .Y(_512_) );
AND2X2 AND2X2_29 ( .A(_1274_), .B(_987__bF_buf1), .Y(_572_) );
AND2X2 AND2X2_30 ( .A(_584_), .B(_581_), .Y(_585_) );
AND2X2 AND2X2_31 ( .A(_1274_), .B(_984_), .Y(_645_) );
AND2X2 AND2X2_32 ( .A(_657_), .B(_654_), .Y(_658_) );
AND2X2 AND2X2_33 ( .A(_1274_), .B(_1196_), .Y(_717_) );
AND2X2 AND2X2_34 ( .A(_1225_), .B(_1226_), .Y(_1227_) );
AND2X2 AND2X2_35 ( .A(_729_), .B(_726_), .Y(_730_) );
AND2X2 AND2X2_36 ( .A(_1274_), .B(_1191_), .Y(_791_) );
AND2X2 AND2X2_37 ( .A(_803_), .B(_800_), .Y(_804_) );
AND2X2 AND2X2_38 ( .A(_1274_), .B(_990__bF_buf1), .Y(_864_) );
AND2X2 AND2X2_39 ( .A(_876_), .B(_873_), .Y(_877_) );
AND2X2 AND2X2_40 ( .A(_1274_), .B(_1025_), .Y(_935_) );
AND2X2 AND2X2_41 ( .A(_947_), .B(_944_), .Y(_948_) );
AND2X2 AND2X2_42 ( .A(_1229_), .B(_1230_), .Y(_1231_) );
AND2X2 AND2X2_43 ( .A(_1274_), .B(_1102__bF_buf1), .Y(_1275_) );
AND2X2 AND2X2_44 ( .A(_1042_), .B(ULA_OUT[6]), .Y(_1280_) );
AND2X2 AND2X2_45 ( .A(_1297_), .B(_1296_), .Y(_1298_) );
AND2X2 AND2X2_46 ( .A(_1042_), .B(ULA_OUT[7]), .Y(_1313_) );
AOI21X1 AOI21X1_1 ( .A(_1212_), .B(_1211_), .C(rst_bF_buf0), .Y(_1213_) );
AOI21X1 AOI21X1_2 ( .A(_1430_), .B(_1431_), .C(_1307_), .Y(_1432_) );
AOI21X1 AOI21X1_3 ( .A(_1038__bF_buf2), .B(_1506_), .C(_1510_), .Y(_1511_) );
AOI21X1 AOI21X1_4 ( .A(_1040_), .B(_1022_), .C(_1037_), .Y(_1516_) );
AOI21X1 AOI21X1_5 ( .A(_1038__bF_buf2), .B(_53_), .C(_57_), .Y(_58_) );
AOI21X1 AOI21X1_6 ( .A(_1040_), .B(_1023_), .C(_1037_), .Y(_63_) );
AOI21X1 AOI21X1_7 ( .A(_1037_), .B(_70_), .C(_72_), .Y(_73_) );
AOI21X1 AOI21X1_8 ( .A(PC_pointer_2_), .B(_1012_), .C(_981_), .Y(_90_) );
AOI21X1 AOI21X1_9 ( .A(_1038__bF_buf4), .B(_131_), .C(_135_), .Y(_136_) );
AOI21X1 AOI21X1_10 ( .A(_1038__bF_buf9), .B(_149_), .C(_153_), .Y(_154_) );
AOI21X1 AOI21X1_11 ( .A(_1040_), .B(_1104_), .C(_1037_), .Y(_159_) );
AOI21X1 AOI21X1_12 ( .A(_1272_), .B(_1543__6_), .C(_1273_), .Y(_1274_) );
AOI21X1 AOI21X1_13 ( .A(_1038__bF_buf2), .B(_220_), .C(_224_), .Y(_225_) );
AOI21X1 AOI21X1_14 ( .A(_1038__bF_buf10), .B(_292_), .C(_296_), .Y(_297_) );
AOI21X1 AOI21X1_15 ( .A(_997__bF_buf0), .B(_1343_), .C(_299_), .Y(_300_) );
AOI21X1 AOI21X1_16 ( .A(_353_), .B(_359_), .C(_1311__bF_buf3), .Y(_360_) );
AOI21X1 AOI21X1_17 ( .A(_1038__bF_buf2), .B(_358_), .C(_360_), .Y(_361_) );
AOI21X1 AOI21X1_18 ( .A(_1038__bF_buf2), .B(_365_), .C(_369_), .Y(_370_) );
AOI21X1 AOI21X1_19 ( .A(_1000__bF_buf2), .B(_1343_), .C(_372_), .Y(_373_) );
AOI21X1 AOI21X1_20 ( .A(_1040_), .B(_1000__bF_buf0), .C(_1037_), .Y(_375_) );
AOI21X1 AOI21X1_21 ( .A(_1038__bF_buf3), .B(_420_), .C(_424_), .Y(_425_) );
AOI21X1 AOI21X1_22 ( .A(_1038__bF_buf2), .B(_438_), .C(_442_), .Y(_443_) );
AOI21X1 AOI21X1_23 ( .A(_1308_), .B(_1309_), .C(_1307_), .Y(_1310_) );
AOI21X1 AOI21X1_24 ( .A(_1004__bF_buf3), .B(_1343_), .C(_445_), .Y(_446_) );
AOI21X1 AOI21X1_25 ( .A(_1040_), .B(_1004__bF_buf3), .C(_1037_), .Y(_448_) );
AOI21X1 AOI21X1_26 ( .A(_1038__bF_buf2), .B(_509_), .C(_513_), .Y(_514_) );
AOI21X1 AOI21X1_27 ( .A(_1026_), .B(_1343_), .C(_516_), .Y(_517_) );
AOI21X1 AOI21X1_28 ( .A(_570_), .B(_576_), .C(_1311__bF_buf1), .Y(_577_) );
AOI21X1 AOI21X1_29 ( .A(_1038__bF_buf9), .B(_575_), .C(_577_), .Y(_578_) );
AOI21X1 AOI21X1_30 ( .A(_1038__bF_buf9), .B(_582_), .C(_586_), .Y(_587_) );
AOI21X1 AOI21X1_31 ( .A(_987__bF_buf0), .B(_1343_), .C(_589_), .Y(_590_) );
AOI21X1 AOI21X1_32 ( .A(_1038__bF_buf9), .B(_655_), .C(_659_), .Y(_660_) );
AOI21X1 AOI21X1_33 ( .A(_1038__bF_buf9), .B(_727_), .C(_731_), .Y(_732_) );
AOI21X1 AOI21X1_34 ( .A(PC_STACK_1__8_), .B(_990__bF_buf3), .C(_1330_), .Y(_1331_) );
AOI21X1 AOI21X1_35 ( .A(_1196_), .B(_1343_), .C(_734_), .Y(_735_) );
AOI21X1 AOI21X1_36 ( .A(_1038__bF_buf4), .B(_783_), .C(_787_), .Y(_788_) );
AOI21X1 AOI21X1_37 ( .A(_1038__bF_buf9), .B(_801_), .C(_805_), .Y(_806_) );
AOI21X1 AOI21X1_38 ( .A(_1040_), .B(_1191_), .C(_1037_), .Y(_811_) );
AOI21X1 AOI21X1_39 ( .A(_1038__bF_buf4), .B(_856_), .C(_860_), .Y(_861_) );
AOI21X1 AOI21X1_40 ( .A(_1038__bF_buf9), .B(_874_), .C(_878_), .Y(_879_) );
AOI21X1 AOI21X1_41 ( .A(_990__bF_buf3), .B(_1343_), .C(_881_), .Y(_882_) );
AOI21X1 AOI21X1_42 ( .A(_1040_), .B(_990__bF_buf3), .C(_1037_), .Y(_884_) );
AOI21X1 AOI21X1_43 ( .A(_1038__bF_buf5), .B(_945_), .C(_949_), .Y(_950_) );
AOI21X1 AOI21X1_44 ( .A(_1040_), .B(_1025_), .C(_1037_), .Y(_955_) );
AOI21X1 AOI21X1_45 ( .A(PC_STACK_6__8_), .B(_1102__bF_buf1), .C(_1334_), .Y(_1335_) );
AOI21X1 AOI21X1_46 ( .A(_1040_), .B(_963_), .C(rst_bF_buf0), .Y(_17_) );
AOI21X1 AOI21X1_47 ( .A(_1341_), .B(_1543__8_), .C(_1342_), .Y(_1343_) );
AOI21X1 AOI21X1_48 ( .A(_1102__bF_buf0), .B(_1343_), .C(_1340_), .Y(_1344_) );
AOI21X1 AOI21X1_49 ( .A(_1040_), .B(_1102__bF_buf0), .C(_1037_), .Y(_1347_) );
AOI21X1 AOI21X1_50 ( .A(_1367_), .B(_1368_), .C(rst_bF_buf1), .Y(_1369_) );
AOI22X1 AOI22X1_1 ( .A(_984_), .B(PC_STACK_4__0_), .C(PC_STACK_5__0_), .D(_987__bF_buf3), .Y(_988_) );
AOI22X1 AOI22X1_2 ( .A(_997__bF_buf2), .B(PC_STACK_9__1_), .C(PC_STACK_10__1_), .D(_1000__bF_buf1), .Y(_1050_) );
AOI22X1 AOI22X1_3 ( .A(PC_STACK_15__0_), .B(_1041__bF_buf2), .C(_171_), .D(_1045__bF_buf7), .Y(_172_) );
AOI22X1 AOI22X1_4 ( .A(PC_STACK_15__1_), .B(_1041__bF_buf7), .C(_178_), .D(_1038__bF_buf1), .Y(_179_) );
AOI22X1 AOI22X1_5 ( .A(PC_STACK_15__2_), .B(_1041__bF_buf7), .C(_185_), .D(_1038__bF_buf1), .Y(_186_) );
AOI22X1 AOI22X1_6 ( .A(PC_STACK_15__3_), .B(_1041__bF_buf8), .C(_192_), .D(_1045__bF_buf0), .Y(_193_) );
AOI22X1 AOI22X1_7 ( .A(PC_STACK_15__4_), .B(_1041__bF_buf7), .C(_199_), .D(_1045__bF_buf8), .Y(_200_) );
AOI22X1 AOI22X1_8 ( .A(PC_STACK_15__5_), .B(_1041__bF_buf7), .C(_206_), .D(_1045__bF_buf8), .Y(_207_) );
AOI22X1 AOI22X1_9 ( .A(_213_), .B(_1038__bF_buf10), .C(_1045__bF_buf2), .D(_215_), .Y(_216_) );
AOI22X1 AOI22X1_10 ( .A(_1045__bF_buf1), .B(_229_), .C(_231_), .D(PC_STACK_15__8_), .Y(_232_) );
AOI22X1 AOI22X1_11 ( .A(_1045__bF_buf1), .B(_236_), .C(_231_), .D(PC_STACK_15__9_), .Y(_237_) );
AOI22X1 AOI22X1_12 ( .A(PC_STACK_9__0_), .B(_1041__bF_buf5), .C(_243_), .D(_1045__bF_buf3), .Y(_244_) );
AOI22X1 AOI22X1_13 ( .A(PC_STACK_15__1_), .B(_1003_), .C(_1004__bF_buf0), .D(PC_STACK_8__1_), .Y(_1051_) );
AOI22X1 AOI22X1_14 ( .A(PC_STACK_9__1_), .B(_1041__bF_buf2), .C(_250_), .D(_1038__bF_buf0), .Y(_251_) );
AOI22X1 AOI22X1_15 ( .A(PC_STACK_9__2_), .B(_1041__bF_buf0), .C(_257_), .D(_1038__bF_buf10), .Y(_258_) );
AOI22X1 AOI22X1_16 ( .A(PC_STACK_9__3_), .B(_1041__bF_buf2), .C(_264_), .D(_1045__bF_buf7), .Y(_265_) );
AOI22X1 AOI22X1_17 ( .A(PC_STACK_9__4_), .B(_1041__bF_buf2), .C(_271_), .D(_1045__bF_buf7), .Y(_272_) );
AOI22X1 AOI22X1_18 ( .A(PC_STACK_9__5_), .B(_1041__bF_buf5), .C(_278_), .D(_1045__bF_buf3), .Y(_279_) );
AOI22X1 AOI22X1_19 ( .A(_285_), .B(_1038__bF_buf6), .C(_1045__bF_buf3), .D(_287_), .Y(_288_) );
AOI22X1 AOI22X1_20 ( .A(_1045__bF_buf2), .B(_301_), .C(_303_), .D(PC_STACK_9__8_), .Y(_304_) );
AOI22X1 AOI22X1_21 ( .A(_1045__bF_buf2), .B(_308_), .C(_303_), .D(PC_STACK_9__9_), .Y(_309_) );
AOI22X1 AOI22X1_22 ( .A(PC_STACK_10__0_), .B(_1041__bF_buf5), .C(_316_), .D(_1045__bF_buf3), .Y(_317_) );
AOI22X1 AOI22X1_23 ( .A(PC_STACK_10__1_), .B(_1041__bF_buf5), .C(_323_), .D(_1038__bF_buf0), .Y(_324_) );
AOI22X1 AOI22X1_24 ( .A(_1022_), .B(PC_STACK_13__1_), .C(PC_STACK_14__1_), .D(_1023_), .Y(_1060_) );
AOI22X1 AOI22X1_25 ( .A(PC_STACK_10__2_), .B(_1041__bF_buf5), .C(_330_), .D(_1038__bF_buf6), .Y(_331_) );
AOI22X1 AOI22X1_26 ( .A(PC_STACK_10__3_), .B(_1041__bF_buf0), .C(_337_), .D(_1045__bF_buf1), .Y(_338_) );
AOI22X1 AOI22X1_27 ( .A(PC_STACK_10__4_), .B(_1041__bF_buf5), .C(_344_), .D(_1045__bF_buf3), .Y(_345_) );
AOI22X1 AOI22X1_28 ( .A(PC_STACK_10__5_), .B(_1041__bF_buf5), .C(_351_), .D(_1045__bF_buf3), .Y(_352_) );
AOI22X1 AOI22X1_29 ( .A(PC_STACK_10__8_), .B(_375_), .C(_374_), .D(_1045__bF_buf2), .Y(_376_) );
AOI22X1 AOI22X1_30 ( .A(PC_STACK_10__9_), .B(_375_), .C(_380_), .D(_1045__bF_buf2), .Y(_381_) );
AOI22X1 AOI22X1_31 ( .A(PC_STACK_8__0_), .B(_1041__bF_buf7), .C(_387_), .D(_1045__bF_buf7), .Y(_388_) );
AOI22X1 AOI22X1_32 ( .A(PC_STACK_8__1_), .B(_1041__bF_buf2), .C(_394_), .D(_1038__bF_buf0), .Y(_395_) );
AOI22X1 AOI22X1_33 ( .A(PC_STACK_8__2_), .B(_1041__bF_buf7), .C(_401_), .D(_1038__bF_buf1), .Y(_402_) );
AOI22X1 AOI22X1_34 ( .A(PC_STACK_8__3_), .B(_1041__bF_buf2), .C(_408_), .D(_1045__bF_buf7), .Y(_409_) );
AOI22X1 AOI22X1_35 ( .A(PC_STACK_11__1_), .B(_1026_), .C(_1025_), .D(PC_STACK_0__1_), .Y(_1061_) );
AOI22X1 AOI22X1_36 ( .A(PC_STACK_8__4_), .B(_1041__bF_buf5), .C(_415_), .D(_1045__bF_buf3), .Y(_416_) );
AOI22X1 AOI22X1_37 ( .A(_431_), .B(_1038__bF_buf6), .C(_1045__bF_buf2), .D(_433_), .Y(_434_) );
AOI22X1 AOI22X1_38 ( .A(_1045__bF_buf2), .B(_447_), .C(_448_), .D(PC_STACK_8__8_), .Y(_449_) );
AOI22X1 AOI22X1_39 ( .A(_1045__bF_buf2), .B(_453_), .C(_448_), .D(PC_STACK_8__9_), .Y(_454_) );
AOI22X1 AOI22X1_40 ( .A(PC_STACK_11__0_), .B(_1041__bF_buf7), .C(_460_), .D(_1045__bF_buf7), .Y(_461_) );
AOI22X1 AOI22X1_41 ( .A(PC_STACK_11__1_), .B(_1041__bF_buf7), .C(_467_), .D(_1038__bF_buf1), .Y(_468_) );
AOI22X1 AOI22X1_42 ( .A(PC_STACK_11__2_), .B(_1041__bF_buf2), .C(_474_), .D(_1038__bF_buf0), .Y(_475_) );
AOI22X1 AOI22X1_43 ( .A(PC_STACK_11__3_), .B(_1041__bF_buf7), .C(_481_), .D(_1045__bF_buf8), .Y(_482_) );
AOI22X1 AOI22X1_44 ( .A(PC_STACK_11__4_), .B(_1041__bF_buf5), .C(_488_), .D(_1045__bF_buf3), .Y(_489_) );
AOI22X1 AOI22X1_45 ( .A(PC_STACK_11__5_), .B(_1041__bF_buf7), .C(_495_), .D(_1045__bF_buf7), .Y(_496_) );
AOI22X1 AOI22X1_46 ( .A(_1007_), .B(_1029_), .C(_1053_), .D(_1063_), .Y(_1065_) );
AOI22X1 AOI22X1_47 ( .A(_502_), .B(_1038__bF_buf6), .C(_1045__bF_buf3), .D(_504_), .Y(_505_) );
AOI22X1 AOI22X1_48 ( .A(_1045__bF_buf2), .B(_518_), .C(_520_), .D(PC_STACK_11__8_), .Y(_521_) );
AOI22X1 AOI22X1_49 ( .A(_1045__bF_buf2), .B(_525_), .C(_520_), .D(PC_STACK_11__9_), .Y(_526_) );
AOI22X1 AOI22X1_50 ( .A(PC_STACK_5__0_), .B(_1041__bF_buf4), .C(_533_), .D(_1045__bF_buf1), .Y(_534_) );
AOI22X1 AOI22X1_51 ( .A(PC_STACK_5__1_), .B(_1041__bF_buf4), .C(_540_), .D(_1038__bF_buf10), .Y(_541_) );
AOI22X1 AOI22X1_52 ( .A(PC_STACK_5__2_), .B(_1041__bF_buf0), .C(_547_), .D(_1038__bF_buf10), .Y(_548_) );
AOI22X1 AOI22X1_53 ( .A(PC_STACK_5__3_), .B(_1041__bF_buf4), .C(_554_), .D(_1045__bF_buf0), .Y(_555_) );
AOI22X1 AOI22X1_54 ( .A(PC_STACK_5__4_), .B(_1041__bF_buf3), .C(_561_), .D(_1045__bF_buf0), .Y(_562_) );
AOI22X1 AOI22X1_55 ( .A(PC_STACK_5__5_), .B(_1041__bF_buf3), .C(_568_), .D(_1045__bF_buf0), .Y(_569_) );
AOI22X1 AOI22X1_56 ( .A(_1045__bF_buf0), .B(_591_), .C(_593_), .D(PC_STACK_5__8_), .Y(_594_) );
AOI22X1 AOI22X1_57 ( .A(PC_STACK_6__1_), .B(_1041__bF_buf1), .C(_1074_), .D(_1038__bF_buf8), .Y(_1075_) );
AOI22X1 AOI22X1_58 ( .A(_1045__bF_buf0), .B(_599_), .C(_593_), .D(PC_STACK_5__9_), .Y(_600_) );
AOI22X1 AOI22X1_59 ( .A(PC_STACK_4__0_), .B(_1041__bF_buf9), .C(_606_), .D(_1045__bF_buf6), .Y(_607_) );
AOI22X1 AOI22X1_60 ( .A(PC_STACK_4__1_), .B(_1041__bF_buf4), .C(_613_), .D(_1038__bF_buf10), .Y(_614_) );
AOI22X1 AOI22X1_61 ( .A(PC_STACK_4__2_), .B(_1041__bF_buf1), .C(_620_), .D(_1038__bF_buf7), .Y(_621_) );
AOI22X1 AOI22X1_62 ( .A(PC_STACK_4__3_), .B(_1041__bF_buf2), .C(_627_), .D(_1045__bF_buf6), .Y(_628_) );
AOI22X1 AOI22X1_63 ( .A(PC_STACK_4__4_), .B(_1041__bF_buf1), .C(_634_), .D(_1045__bF_buf4), .Y(_635_) );
AOI22X1 AOI22X1_64 ( .A(PC_STACK_4__5_), .B(_1041__bF_buf9), .C(_641_), .D(_1045__bF_buf5), .Y(_642_) );
AOI22X1 AOI22X1_65 ( .A(_648_), .B(_1038__bF_buf5), .C(_1045__bF_buf0), .D(_650_), .Y(_651_) );
AOI22X1 AOI22X1_66 ( .A(_1045__bF_buf5), .B(_664_), .C(_666_), .D(PC_STACK_4__8_), .Y(_667_) );
AOI22X1 AOI22X1_67 ( .A(_1045__bF_buf5), .B(_671_), .C(_666_), .D(PC_STACK_4__9_), .Y(_672_) );
AOI22X1 AOI22X1_68 ( .A(_984_), .B(PC_STACK_4__2_), .C(PC_STACK_9__2_), .D(_997__bF_buf2), .Y(_1088_) );
AOI22X1 AOI22X1_69 ( .A(PC_STACK_3__0_), .B(_1041__bF_buf1), .C(_678_), .D(_1045__bF_buf9), .Y(_679_) );
AOI22X1 AOI22X1_70 ( .A(PC_STACK_3__1_), .B(_1041__bF_buf1), .C(_685_), .D(_1038__bF_buf8), .Y(_686_) );
AOI22X1 AOI22X1_71 ( .A(PC_STACK_3__2_), .B(_1041__bF_buf6), .C(_692_), .D(_1038__bF_buf1), .Y(_693_) );
AOI22X1 AOI22X1_72 ( .A(PC_STACK_3__3_), .B(_1041__bF_buf10), .C(_699_), .D(_1045__bF_buf9), .Y(_700_) );
AOI22X1 AOI22X1_73 ( .A(PC_STACK_3__4_), .B(_1041__bF_buf10), .C(_706_), .D(_1045__bF_buf9), .Y(_707_) );
AOI22X1 AOI22X1_74 ( .A(PC_STACK_3__5_), .B(_1041__bF_buf1), .C(_713_), .D(_1045__bF_buf9), .Y(_714_) );
AOI22X1 AOI22X1_75 ( .A(_720_), .B(_1038__bF_buf9), .C(_1045__bF_buf0), .D(_722_), .Y(_723_) );
AOI22X1 AOI22X1_76 ( .A(_1045__bF_buf5), .B(_736_), .C(_738_), .D(PC_STACK_3__8_), .Y(_739_) );
AOI22X1 AOI22X1_77 ( .A(_1045__bF_buf10), .B(_743_), .C(_738_), .D(PC_STACK_3__9_), .Y(_744_) );
AOI22X1 AOI22X1_78 ( .A(PC_STACK_2__0_), .B(_1041__bF_buf1), .C(_750_), .D(_1045__bF_buf4), .Y(_751_) );
AOI22X1 AOI22X1_79 ( .A(PC_STACK_12__2_), .B(_992__bF_buf2), .C(_987__bF_buf3), .D(PC_STACK_5__2_), .Y(_1089_) );
AOI22X1 AOI22X1_80 ( .A(PC_STACK_2__1_), .B(_1041__bF_buf6), .C(_757_), .D(_1038__bF_buf7), .Y(_758_) );
AOI22X1 AOI22X1_81 ( .A(PC_STACK_2__2_), .B(_1041__bF_buf6), .C(_764_), .D(_1038__bF_buf7), .Y(_765_) );
AOI22X1 AOI22X1_82 ( .A(PC_STACK_2__3_), .B(_1041__bF_buf1), .C(_771_), .D(_1045__bF_buf4), .Y(_772_) );
AOI22X1 AOI22X1_83 ( .A(PC_STACK_2__4_), .B(_1041__bF_buf1), .C(_778_), .D(_1045__bF_buf4), .Y(_779_) );
AOI22X1 AOI22X1_84 ( .A(_794_), .B(_1038__bF_buf9), .C(_1045__bF_buf5), .D(_796_), .Y(_797_) );
AOI22X1 AOI22X1_85 ( .A(_1045__bF_buf10), .B(_810_), .C(_811_), .D(PC_STACK_2__8_), .Y(_812_) );
AOI22X1 AOI22X1_86 ( .A(_1045__bF_buf10), .B(_816_), .C(_811_), .D(PC_STACK_2__9_), .Y(_817_) );
AOI22X1 AOI22X1_87 ( .A(PC_STACK_1__0_), .B(_1041__bF_buf9), .C(_823_), .D(_1045__bF_buf6), .Y(_824_) );
AOI22X1 AOI22X1_88 ( .A(PC_STACK_1__1_), .B(_1041__bF_buf9), .C(_830_), .D(_1038__bF_buf8), .Y(_831_) );
AOI22X1 AOI22X1_89 ( .A(PC_STACK_1__2_), .B(_1041__bF_buf9), .C(_837_), .D(_1038__bF_buf3), .Y(_838_) );
AOI22X1 AOI22X1_90 ( .A(_1000__bF_buf1), .B(PC_STACK_10__2_), .C(PC_STACK_6__2_), .D(_1102__bF_buf3), .Y(_1103_) );
AOI22X1 AOI22X1_91 ( .A(PC_STACK_1__3_), .B(_1041__bF_buf10), .C(_844_), .D(_1045__bF_buf10), .Y(_845_) );
AOI22X1 AOI22X1_92 ( .A(PC_STACK_1__4_), .B(_1041__bF_buf10), .C(_851_), .D(_1045__bF_buf10), .Y(_852_) );
AOI22X1 AOI22X1_93 ( .A(_867_), .B(_1038__bF_buf5), .C(_1045__bF_buf5), .D(_869_), .Y(_870_) );
AOI22X1 AOI22X1_94 ( .A(_1045__bF_buf10), .B(_883_), .C(_884_), .D(PC_STACK_1__8_), .Y(_885_) );
AOI22X1 AOI22X1_95 ( .A(_1045__bF_buf10), .B(_889_), .C(_884_), .D(PC_STACK_1__9_), .Y(_890_) );
AOI22X1 AOI22X1_96 ( .A(PC_STACK_0__0_), .B(_1041__bF_buf6), .C(_896_), .D(_1045__bF_buf8), .Y(_897_) );
AOI22X1 AOI22X1_97 ( .A(PC_STACK_0__1_), .B(_1041__bF_buf6), .C(_903_), .D(_1038__bF_buf7), .Y(_904_) );
AOI22X1 AOI22X1_98 ( .A(PC_STACK_0__2_), .B(_1041__bF_buf6), .C(_910_), .D(_1038__bF_buf7), .Y(_911_) );
AOI22X1 AOI22X1_99 ( .A(PC_STACK_0__3_), .B(_1041__bF_buf6), .C(_917_), .D(_1045__bF_buf4), .Y(_918_) );
AOI22X1 AOI22X1_100 ( .A(PC_STACK_0__4_), .B(_1041__bF_buf6), .C(_924_), .D(_1045__bF_buf8), .Y(_925_) );
AOI22X1 AOI22X1_101 ( .A(PC_STACK_1__2_), .B(_990__bF_buf1), .C(_1104_), .D(PC_STACK_7__2_), .Y(_1105_) );
AOI22X1 AOI22X1_102 ( .A(PC_STACK_0__5_), .B(_1041__bF_buf6), .C(_931_), .D(_1045__bF_buf8), .Y(_932_) );
AOI22X1 AOI22X1_103 ( .A(_938_), .B(_1038__bF_buf2), .C(_1045__bF_buf0), .D(_940_), .Y(_941_) );
AOI22X1 AOI22X1_104 ( .A(_954_), .B(_1045__bF_buf6), .C(_955_), .D(PC_STACK_0__8_), .Y(_956_) );
AOI22X1 AOI22X1_105 ( .A(_960_), .B(_1045__bF_buf6), .C(_955_), .D(PC_STACK_0__9_), .Y(_961_) );
AOI22X1 AOI22X1_106 ( .A(PC_STACK_12__0_), .B(_992__bF_buf1), .C(_990__bF_buf1), .D(PC_STACK_1__0_), .Y(_993_) );
AOI22X1 AOI22X1_107 ( .A(PC_STACK_6__0_), .B(_1102__bF_buf3), .C(_1104_), .D(PC_STACK_7__0_), .Y(_1113_) );
AOI22X1 AOI22X1_108 ( .A(PC_STACK_6__1_), .B(_1102__bF_buf3), .C(_1104_), .D(PC_STACK_7__1_), .Y(_1129_) );
AOI22X1 AOI22X1_109 ( .A(PC_STACK_6__2_), .B(_1041__bF_buf2), .C(_1149_), .D(_1038__bF_buf3), .Y(_1150_) );
AOI22X1 AOI22X1_110 ( .A(_984_), .B(PC_STACK_4__3_), .C(PC_STACK_9__3_), .D(_997__bF_buf2), .Y(_1158_) );
AOI22X1 AOI22X1_111 ( .A(PC_STACK_12__3_), .B(_992__bF_buf2), .C(_987__bF_buf3), .D(PC_STACK_5__3_), .Y(_1159_) );
AOI22X1 AOI22X1_112 ( .A(PC_STACK_6__3_), .B(_1041__bF_buf10), .C(_1189_), .D(_1045__bF_buf9), .Y(_1190_) );
AOI22X1 AOI22X1_113 ( .A(PC_STACK_4__4_), .B(_984_), .C(_1191_), .D(PC_STACK_2__4_), .Y(_1192_) );
AOI22X1 AOI22X1_114 ( .A(PC_STACK_14__4_), .B(_1023_), .C(_1025_), .D(PC_STACK_0__4_), .Y(_1193_) );
AOI22X1 AOI22X1_115 ( .A(PC_STACK_6__4_), .B(_1102__bF_buf3), .C(_1104_), .D(PC_STACK_7__4_), .Y(_1195_) );
AOI22X1 AOI22X1_116 ( .A(PC_STACK_3__4_), .B(_1196_), .C(_990__bF_buf0), .D(PC_STACK_1__4_), .Y(_1197_) );
AOI22X1 AOI22X1_117 ( .A(_997__bF_buf1), .B(PC_STACK_9__0_), .C(PC_STACK_10__0_), .D(_1000__bF_buf1), .Y(_1001_) );
AOI22X1 AOI22X1_118 ( .A(PC_STACK_11__4_), .B(_1026_), .C(_1000__bF_buf2), .D(PC_STACK_10__4_), .Y(_1207_) );
AOI22X1 AOI22X1_119 ( .A(PC_STACK_12__4_), .B(_992__bF_buf2), .C(_987__bF_buf3), .D(PC_STACK_5__4_), .Y(_1208_) );
AOI22X1 AOI22X1_120 ( .A(PC_STACK_6__4_), .B(_1041__bF_buf10), .C(_1221_), .D(_1045__bF_buf9), .Y(_1222_) );
AOI22X1 AOI22X1_121 ( .A(PC_STACK_13__5_), .B(_1022_), .C(_997__bF_buf2), .D(PC_STACK_9__5_), .Y(_1223_) );
AOI22X1 AOI22X1_122 ( .A(PC_STACK_12__5_), .B(_992__bF_buf1), .C(_1102__bF_buf3), .D(PC_STACK_6__5_), .Y(_1224_) );
AOI22X1 AOI22X1_123 ( .A(PC_STACK_11__5_), .B(_1026_), .C(_1000__bF_buf1), .D(PC_STACK_10__5_), .Y(_1225_) );
AOI22X1 AOI22X1_124 ( .A(PC_STACK_15__5_), .B(_1003_), .C(_1004__bF_buf0), .D(PC_STACK_8__5_), .Y(_1226_) );
AOI22X1 AOI22X1_125 ( .A(PC_STACK_3__5_), .B(_1196_), .C(_1191_), .D(PC_STACK_2__5_), .Y(_1229_) );
AOI22X1 AOI22X1_126 ( .A(_984_), .B(PC_STACK_4__5_), .C(PC_STACK_1__5_), .D(_990__bF_buf0), .Y(_1230_) );
AOI22X1 AOI22X1_127 ( .A(PC_STACK_14__5_), .B(_1023_), .C(_1025_), .D(PC_STACK_0__5_), .Y(_1232_) );
AOI22X1 AOI22X1_128 ( .A(PC_STACK_15__0_), .B(_1003_), .C(_1004__bF_buf0), .D(PC_STACK_8__0_), .Y(_1005_) );
AOI22X1 AOI22X1_129 ( .A(PC_STACK_5__5_), .B(_987__bF_buf2), .C(_1104_), .D(PC_STACK_7__5_), .Y(_1233_) );
AOI22X1 AOI22X1_130 ( .A(PC_STACK_6__5_), .B(_1041__bF_buf10), .C(_1246_), .D(_1045__bF_buf9), .Y(_1247_) );
AOI22X1 AOI22X1_131 ( .A(PC_STACK_5__6_), .B(_987__bF_buf1), .C(_1104_), .D(PC_STACK_7__6_), .Y(_1256_) );
AOI22X1 AOI22X1_132 ( .A(PC_STACK_12__6_), .B(_992__bF_buf0), .C(_1102__bF_buf1), .D(PC_STACK_6__6_), .Y(_1257_) );
AOI22X1 AOI22X1_133 ( .A(PC_STACK_3__6_), .B(_1196_), .C(_990__bF_buf2), .D(PC_STACK_1__6_), .Y(_1266_) );
AOI22X1 AOI22X1_134 ( .A(PC_STACK_0__6_), .B(_1025_), .C(_1000__bF_buf3), .D(PC_STACK_10__6_), .Y(_1267_) );
AOI22X1 AOI22X1_135 ( .A(_1279_), .B(_1038__bF_buf5), .C(_1045__bF_buf10), .D(_1282_), .Y(_1283_) );
AOI22X1 AOI22X1_136 ( .A(PC_STACK_11__7_), .B(_1026_), .C(_1000__bF_buf3), .D(PC_STACK_10__7_), .Y(_1291_) );
AOI22X1 AOI22X1_137 ( .A(PC_STACK_14__7_), .B(_1023_), .C(_1004__bF_buf2), .D(PC_STACK_8__7_), .Y(_1292_) );
AOI22X1 AOI22X1_138 ( .A(PC_STACK_12__7_), .B(_992__bF_buf3), .C(_984_), .D(PC_STACK_4__7_), .Y(_1294_) );
AOI22X1 AOI22X1_139 ( .A(_1022_), .B(PC_STACK_13__0_), .C(PC_STACK_14__0_), .D(_1023_), .Y(_1024_) );
AOI22X1 AOI22X1_140 ( .A(PC_STACK_6__7_), .B(_1102__bF_buf2), .C(_1191_), .D(PC_STACK_2__7_), .Y(_1295_) );
AOI22X1 AOI22X1_141 ( .A(PC_STACK_15__7_), .B(_1003_), .C(_1025_), .D(PC_STACK_0__7_), .Y(_1296_) );
AOI22X1 AOI22X1_142 ( .A(_990__bF_buf2), .B(PC_STACK_1__7_), .C(PC_STACK_5__7_), .D(_987__bF_buf2), .Y(_1297_) );
AOI22X1 AOI22X1_143 ( .A(_1004__bF_buf3), .B(PC_STACK_8__8_), .C(PC_STACK_9__8_), .D(_997__bF_buf0), .Y(_1318_) );
AOI22X1 AOI22X1_144 ( .A(PC_STACK_11__8_), .B(_1026_), .C(_1000__bF_buf2), .D(PC_STACK_10__8_), .Y(_1319_) );
AOI22X1 AOI22X1_145 ( .A(PC_STACK_3__8_), .B(_1196_), .C(_987__bF_buf2), .D(PC_STACK_5__8_), .Y(_1336_) );
AOI22X1 AOI22X1_146 ( .A(_1347_), .B(PC_STACK_6__8_), .C(_1045__bF_buf10), .D(_1346_), .Y(_1348_) );
AOI22X1 AOI22X1_147 ( .A(_1023_), .B(PC_STACK_14__9_), .C(PC_STACK_11__9_), .D(_1026_), .Y(_1350_) );
AOI22X1 AOI22X1_148 ( .A(PC_STACK_15__9_), .B(_1003_), .C(_997__bF_buf3), .D(PC_STACK_9__9_), .Y(_1351_) );
AOI22X1 AOI22X1_149 ( .A(_990__bF_buf2), .B(PC_STACK_1__9_), .C(PC_STACK_5__9_), .D(_987__bF_buf2), .Y(_1359_) );
AOI22X1 AOI22X1_150 ( .A(PC_STACK_11__0_), .B(_1026_), .C(_1025_), .D(PC_STACK_0__0_), .Y(_1027_) );
AOI22X1 AOI22X1_151 ( .A(_1004__bF_buf3), .B(PC_STACK_8__9_), .C(PC_STACK_10__9_), .D(_1000__bF_buf0), .Y(_1360_) );
AOI22X1 AOI22X1_152 ( .A(PC_STACK_3__9_), .B(_1196_), .C(_1102__bF_buf0), .D(PC_STACK_6__9_), .Y(_1362_) );
AOI22X1 AOI22X1_153 ( .A(PC_STACK_12__9_), .B(_992__bF_buf1), .C(_1191_), .D(PC_STACK_2__9_), .Y(_1363_) );
AOI22X1 AOI22X1_154 ( .A(_1349_), .B(_1025_), .C(_1365_), .D(_1358_), .Y(_1543__9_) );
AOI22X1 AOI22X1_155 ( .A(_1347_), .B(PC_STACK_6__9_), .C(_1045__bF_buf10), .D(_1374_), .Y(_1375_) );
AOI22X1 AOI22X1_156 ( .A(PC_STACK_12__0_), .B(_1041__bF_buf9), .C(_1381_), .D(_1045__bF_buf6), .Y(_1382_) );
AOI22X1 AOI22X1_157 ( .A(PC_STACK_12__1_), .B(_1041__bF_buf9), .C(_1388_), .D(_1038__bF_buf5), .Y(_1389_) );
AOI22X1 AOI22X1_158 ( .A(PC_STACK_12__2_), .B(_1041__bF_buf4), .C(_1395_), .D(_1038__bF_buf10), .Y(_1396_) );
AOI22X1 AOI22X1_159 ( .A(PC_STACK_12__3_), .B(_1041__bF_buf9), .C(_1402_), .D(_1045__bF_buf6), .Y(_1403_) );
AOI22X1 AOI22X1_160 ( .A(PC_STACK_12__4_), .B(_1041__bF_buf9), .C(_1409_), .D(_1045__bF_buf5), .Y(_1410_) );
AOI22X1 AOI22X1_161 ( .A(PC_STACK_6__0_), .B(_1041__bF_buf6), .C(_1044_), .D(_1045__bF_buf4), .Y(_1046_) );
AOI22X1 AOI22X1_162 ( .A(PC_STACK_12__5_), .B(_1041__bF_buf9), .C(_1416_), .D(_1045__bF_buf5), .Y(_1417_) );
AOI22X1 AOI22X1_163 ( .A(_1424_), .B(_1038__bF_buf5), .C(_1045__bF_buf5), .D(_1426_), .Y(_1427_) );
AOI22X1 AOI22X1_164 ( .A(_1045__bF_buf0), .B(_1441_), .C(_1443_), .D(PC_STACK_12__8_), .Y(_1444_) );
AOI22X1 AOI22X1_165 ( .A(_1045__bF_buf5), .B(_1448_), .C(_1443_), .D(PC_STACK_12__9_), .Y(_1449_) );
AOI22X1 AOI22X1_166 ( .A(PC_STACK_13__0_), .B(_1041__bF_buf0), .C(_1455_), .D(_1045__bF_buf6), .Y(_1456_) );
AOI22X1 AOI22X1_167 ( .A(PC_STACK_13__1_), .B(_1041__bF_buf2), .C(_1462_), .D(_1038__bF_buf0), .Y(_1463_) );
AOI22X1 AOI22X1_168 ( .A(PC_STACK_13__2_), .B(_1041__bF_buf7), .C(_1469_), .D(_1038__bF_buf0), .Y(_1470_) );
AOI22X1 AOI22X1_169 ( .A(PC_STACK_13__3_), .B(_1041__bF_buf2), .C(_1476_), .D(_1045__bF_buf6), .Y(_1477_) );
AOI22X1 AOI22X1_170 ( .A(PC_STACK_13__4_), .B(_1041__bF_buf5), .C(_1483_), .D(_1045__bF_buf3), .Y(_1484_) );
AOI22X1 AOI22X1_171 ( .A(PC_STACK_13__5_), .B(_1041__bF_buf0), .C(_1490_), .D(_1045__bF_buf2), .Y(_1491_) );
AOI22X1 AOI22X1_172 ( .A(_984_), .B(PC_STACK_4__1_), .C(PC_STACK_5__1_), .D(_987__bF_buf3), .Y(_1047_) );
AOI22X1 AOI22X1_173 ( .A(_1498_), .B(_1038__bF_buf10), .C(_1045__bF_buf2), .D(_1500_), .Y(_1501_) );
AOI22X1 AOI22X1_174 ( .A(PC_STACK_13__8_), .B(_1516_), .C(_1515_), .D(_1045__bF_buf1), .Y(_1517_) );
AOI22X1 AOI22X1_175 ( .A(PC_STACK_13__9_), .B(_1516_), .C(_1521_), .D(_1045__bF_buf1), .Y(_1522_) );
AOI22X1 AOI22X1_176 ( .A(PC_STACK_14__0_), .B(_1041__bF_buf0), .C(_1528_), .D(_1045__bF_buf1), .Y(_1529_) );
AOI22X1 AOI22X1_177 ( .A(PC_STACK_14__1_), .B(_1041__bF_buf4), .C(_1535_), .D(_1038__bF_buf10), .Y(_1536_) );
AOI22X1 AOI22X1_178 ( .A(PC_STACK_14__2_), .B(_1041__bF_buf0), .C(_18_), .D(_1038__bF_buf2), .Y(_19_) );
AOI22X1 AOI22X1_179 ( .A(PC_STACK_14__3_), .B(_1041__bF_buf8), .C(_25_), .D(_1045__bF_buf0), .Y(_26_) );
AOI22X1 AOI22X1_180 ( .A(PC_STACK_14__4_), .B(_1041__bF_buf6), .C(_32_), .D(_1045__bF_buf4), .Y(_33_) );
AOI22X1 AOI22X1_181 ( .A(PC_STACK_14__5_), .B(_1041__bF_buf6), .C(_39_), .D(_1045__bF_buf4), .Y(_40_) );
AOI22X1 AOI22X1_182 ( .A(_46_), .B(_1038__bF_buf2), .C(_1045__bF_buf1), .D(_48_), .Y(_49_) );
AOI22X1 AOI22X1_183 ( .A(PC_STACK_12__1_), .B(_992__bF_buf1), .C(_990__bF_buf1), .D(PC_STACK_1__1_), .Y(_1048_) );
AOI22X1 AOI22X1_184 ( .A(PC_STACK_14__8_), .B(_63_), .C(_62_), .D(_1045__bF_buf1), .Y(_64_) );
AOI22X1 AOI22X1_185 ( .A(PC_STACK_14__9_), .B(_63_), .C(_68_), .D(_1045__bF_buf1), .Y(_69_) );
AOI22X1 AOI22X1_186 ( .A(PC_STACK_7__0_), .B(_1041__bF_buf1), .C(_98_), .D(_1045__bF_buf4), .Y(_99_) );
AOI22X1 AOI22X1_187 ( .A(PC_STACK_7__1_), .B(_1041__bF_buf1), .C(_105_), .D(_1038__bF_buf8), .Y(_106_) );
AOI22X1 AOI22X1_188 ( .A(PC_STACK_7__2_), .B(_1041__bF_buf9), .C(_112_), .D(_1038__bF_buf8), .Y(_113_) );
AOI22X1 AOI22X1_189 ( .A(PC_STACK_7__3_), .B(_1041__bF_buf10), .C(_119_), .D(_1045__bF_buf9), .Y(_120_) );
AOI22X1 AOI22X1_190 ( .A(PC_STACK_7__4_), .B(_1041__bF_buf10), .C(_126_), .D(_1045__bF_buf9), .Y(_127_) );
AOI22X1 AOI22X1_191 ( .A(_142_), .B(_1038__bF_buf9), .C(_1045__bF_buf0), .D(_144_), .Y(_145_) );
AOI22X1 AOI22X1_192 ( .A(_1045__bF_buf10), .B(_158_), .C(_159_), .D(PC_STACK_7__8_), .Y(_160_) );
AOI22X1 AOI22X1_193 ( .A(_1045__bF_buf10), .B(_164_), .C(_159_), .D(PC_STACK_7__9_), .Y(_165_) );
BUFX2 BUFX2_1 ( .A(_1542__0_), .Y(_0__0_) );
BUFX2 BUFX2_2 ( .A(_1542__9_), .Y(_0__9_) );
BUFX2 BUFX2_3 ( .A(_1542__10_), .Y(_0__10_) );
BUFX2 BUFX2_4 ( .A(_1542__11_), .Y(_0__11_) );
BUFX2 BUFX2_5 ( .A(_1542__12_), .Y(_0__12_) );
BUFX2 BUFX2_6 ( .A(_1542__13_), .Y(_0__13_) );
BUFX2 BUFX2_7 ( .A(_1542__14_), .Y(_0__14_) );
BUFX2 BUFX2_8 ( .A(IDATA_CORE_out[15]), .Y(_0__15_) );
BUFX2 BUFX2_9 ( .A(_1543__0_), .Y(_1__0_) );
BUFX2 BUFX2_10 ( .A(_1543__1_), .Y(_1__1_) );
BUFX2 BUFX2_11 ( .A(_1543__2_), .Y(_1__2_) );
BUFX2 BUFX2_12 ( .A(_1542__1_), .Y(_0__1_) );
BUFX2 BUFX2_13 ( .A(_1543__3_), .Y(_1__3_) );
BUFX2 BUFX2_14 ( .A(_1543__4_), .Y(_1__4_) );
BUFX2 BUFX2_15 ( .A(_1543__5_), .Y(_1__5_) );
BUFX2 BUFX2_16 ( .A(_1543__6_), .Y(_1__6_) );
BUFX2 BUFX2_17 ( .A(_1543__7_), .Y(_1__7_) );
BUFX2 BUFX2_18 ( .A(_1543__8_), .Y(_1__8_) );
BUFX2 BUFX2_19 ( .A(_1543__9_), .Y(_1__9_) );
BUFX2 BUFX2_20 ( .A(_1544_), .Y(_2_) );
BUFX2 BUFX2_21 ( .A(_1545__0_), .Y(_3__0_) );
BUFX2 BUFX2_22 ( .A(_1545__1_), .Y(_3__1_) );
BUFX2 BUFX2_23 ( .A(_1542__2_), .Y(_0__2_) );
BUFX2 BUFX2_24 ( .A(_1545__2_), .Y(_3__2_) );
BUFX2 BUFX2_25 ( .A(_1545__3_), .Y(_3__3_) );
BUFX2 BUFX2_26 ( .A(_1545__4_), .Y(_3__4_) );
BUFX2 BUFX2_27 ( .A(_1545__5_), .Y(_3__5_) );
BUFX2 BUFX2_28 ( .A(_1545__6_), .Y(_3__6_) );
BUFX2 BUFX2_29 ( .A(_1545__7_), .Y(_3__7_) );
BUFX2 BUFX2_30 ( .A(_1545__8_), .Y(_3__8_) );
BUFX2 BUFX2_31 ( .A(_1545__9_), .Y(_3__9_) );
BUFX2 BUFX2_32 ( .A(_1542__3_), .Y(_0__3_) );
BUFX2 BUFX2_33 ( .A(_1542__4_), .Y(_0__4_) );
BUFX2 BUFX2_34 ( .A(_1542__5_), .Y(_0__5_) );
BUFX2 BUFX2_35 ( .A(_1542__6_), .Y(_0__6_) );
BUFX2 BUFX2_36 ( .A(_1542__7_), .Y(_0__7_) );
BUFX2 BUFX2_37 ( .A(_1542__8_), .Y(_0__8_) );
BUFX4 BUFX4_1 ( .A(_1116_), .Y(_1116__bF_buf4) );
BUFX4 BUFX4_2 ( .A(_999_), .Y(_999__bF_buf5) );
BUFX4 BUFX4_3 ( .A(rst), .Y(rst_bF_buf3) );
BUFX4 BUFX4_4 ( .A(rst), .Y(rst_bF_buf2) );
BUFX4 BUFX4_5 ( .A(rst), .Y(rst_bF_buf1) );
BUFX4 BUFX4_6 ( .A(rst), .Y(rst_bF_buf0) );
BUFX4 BUFX4_7 ( .A(_1109_), .Y(_1109__bF_buf4) );
BUFX4 BUFX4_8 ( .A(_1109_), .Y(_1109__bF_buf3) );
BUFX4 BUFX4_9 ( .A(_1109_), .Y(_1109__bF_buf2) );
BUFX4 BUFX4_10 ( .A(_1109_), .Y(_1109__bF_buf1) );
BUFX4 BUFX4_11 ( .A(_1109_), .Y(_1109__bF_buf0) );
BUFX4 BUFX4_12 ( .A(_992_), .Y(_992__bF_buf3) );
BUFX4 BUFX4_13 ( .A(_999_), .Y(_999__bF_buf4) );
BUFX4 BUFX4_14 ( .A(_992_), .Y(_992__bF_buf2) );
BUFX4 BUFX4_15 ( .A(_992_), .Y(_992__bF_buf1) );
BUFX4 BUFX4_16 ( .A(_992_), .Y(_992__bF_buf0) );
BUFX4 BUFX4_17 ( .A(_989_), .Y(_989__bF_buf5) );
BUFX4 BUFX4_18 ( .A(_989_), .Y(_989__bF_buf4) );
BUFX4 BUFX4_19 ( .A(_989_), .Y(_989__bF_buf3) );
BUFX4 BUFX4_20 ( .A(_989_), .Y(_989__bF_buf2) );
BUFX4 BUFX4_21 ( .A(_989_), .Y(_989__bF_buf1) );
BUFX4 BUFX4_22 ( .A(_989_), .Y(_989__bF_buf0) );
BUFX4 BUFX4_23 ( .A(_1085_), .Y(_1085__bF_buf4) );
BUFX4 BUFX4_24 ( .A(_999_), .Y(_999__bF_buf3) );
BUFX4 BUFX4_25 ( .A(_1085_), .Y(_1085__bF_buf3) );
BUFX4 BUFX4_26 ( .A(_1085_), .Y(_1085__bF_buf2) );
BUFX4 BUFX4_27 ( .A(_1085_), .Y(_1085__bF_buf1) );
BUFX4 BUFX4_28 ( .A(_1085_), .Y(_1085__bF_buf0) );
BUFX4 BUFX4_29 ( .A(_986_), .Y(_986__bF_buf5) );
BUFX4 BUFX4_30 ( .A(_986_), .Y(_986__bF_buf4) );
BUFX4 BUFX4_31 ( .A(_986_), .Y(_986__bF_buf3) );
BUFX4 BUFX4_32 ( .A(_986_), .Y(_986__bF_buf2) );
BUFX4 BUFX4_33 ( .A(_986_), .Y(_986__bF_buf1) );
BUFX4 BUFX4_34 ( .A(_986_), .Y(_986__bF_buf0) );
BUFX4 BUFX4_35 ( .A(_999_), .Y(_999__bF_buf2) );
BUFX4 BUFX4_36 ( .A(_983_), .Y(_983__bF_buf6) );
BUFX4 BUFX4_37 ( .A(_983_), .Y(_983__bF_buf5) );
BUFX4 BUFX4_38 ( .A(_983_), .Y(_983__bF_buf4) );
BUFX4 BUFX4_39 ( .A(_983_), .Y(_983__bF_buf3) );
BUFX4 BUFX4_40 ( .A(_983_), .Y(_983__bF_buf2) );
BUFX4 BUFX4_41 ( .A(_983_), .Y(_983__bF_buf1) );
BUFX4 BUFX4_42 ( .A(_983_), .Y(_983__bF_buf0) );
BUFX4 BUFX4_43 ( .A(_1041_), .Y(_1041__bF_buf10) );
BUFX4 BUFX4_44 ( .A(_1041_), .Y(_1041__bF_buf9) );
BUFX4 BUFX4_45 ( .A(_1041_), .Y(_1041__bF_buf8) );
BUFX4 BUFX4_46 ( .A(_999_), .Y(_999__bF_buf1) );
BUFX4 BUFX4_47 ( .A(_1041_), .Y(_1041__bF_buf7) );
BUFX4 BUFX4_48 ( .A(_1041_), .Y(_1041__bF_buf6) );
BUFX4 BUFX4_49 ( .A(_1041_), .Y(_1041__bF_buf5) );
BUFX4 BUFX4_50 ( .A(_1041_), .Y(_1041__bF_buf4) );
BUFX4 BUFX4_51 ( .A(_1041_), .Y(_1041__bF_buf3) );
BUFX4 BUFX4_52 ( .A(_1041_), .Y(_1041__bF_buf2) );
BUFX4 BUFX4_53 ( .A(_1041_), .Y(_1041__bF_buf1) );
BUFX4 BUFX4_54 ( .A(_1041_), .Y(_1041__bF_buf0) );
BUFX4 BUFX4_55 ( .A(_1038_), .Y(_1038__bF_buf10) );
BUFX4 BUFX4_56 ( .A(_1038_), .Y(_1038__bF_buf9) );
BUFX4 BUFX4_57 ( .A(_999_), .Y(_999__bF_buf0) );
BUFX4 BUFX4_58 ( .A(_1038_), .Y(_1038__bF_buf8) );
BUFX4 BUFX4_59 ( .A(_1038_), .Y(_1038__bF_buf7) );
BUFX4 BUFX4_60 ( .A(_1038_), .Y(_1038__bF_buf6) );
BUFX4 BUFX4_61 ( .A(_1038_), .Y(_1038__bF_buf5) );
BUFX4 BUFX4_62 ( .A(_1038_), .Y(_1038__bF_buf4) );
BUFX4 BUFX4_63 ( .A(_1038_), .Y(_1038__bF_buf3) );
BUFX4 BUFX4_64 ( .A(_1038_), .Y(_1038__bF_buf2) );
BUFX4 BUFX4_65 ( .A(_1038_), .Y(_1038__bF_buf1) );
BUFX4 BUFX4_66 ( .A(_1038_), .Y(_1038__bF_buf0) );
BUFX4 BUFX4_67 ( .A(_1000_), .Y(_1000__bF_buf3) );
BUFX4 BUFX4_68 ( .A(_1095_), .Y(_1095__bF_buf4) );
BUFX4 BUFX4_69 ( .A(_1000_), .Y(_1000__bF_buf2) );
BUFX4 BUFX4_70 ( .A(_1000_), .Y(_1000__bF_buf1) );
BUFX4 BUFX4_71 ( .A(_1000_), .Y(_1000__bF_buf0) );
BUFX4 BUFX4_72 ( .A(_1099_), .Y(_1099__bF_buf4) );
BUFX4 BUFX4_73 ( .A(_1099_), .Y(_1099__bF_buf3) );
BUFX4 BUFX4_74 ( .A(_1099_), .Y(_1099__bF_buf2) );
BUFX4 BUFX4_75 ( .A(_1099_), .Y(_1099__bF_buf1) );
BUFX4 BUFX4_76 ( .A(_1099_), .Y(_1099__bF_buf0) );
BUFX4 BUFX4_77 ( .A(_1311_), .Y(_1311__bF_buf3) );
BUFX4 BUFX4_78 ( .A(_1311_), .Y(_1311__bF_buf2) );
BUFX4 BUFX4_79 ( .A(_1095_), .Y(_1095__bF_buf3) );
BUFX4 BUFX4_80 ( .A(_1311_), .Y(_1311__bF_buf1) );
BUFX4 BUFX4_81 ( .A(_1311_), .Y(_1311__bF_buf0) );
BUFX4 BUFX4_82 ( .A(_1117_), .Y(_1117__bF_buf4) );
BUFX4 BUFX4_83 ( .A(_1117_), .Y(_1117__bF_buf3) );
BUFX4 BUFX4_84 ( .A(_1117_), .Y(_1117__bF_buf2) );
BUFX4 BUFX4_85 ( .A(_1117_), .Y(_1117__bF_buf1) );
BUFX4 BUFX4_86 ( .A(_1117_), .Y(_1117__bF_buf0) );
BUFX4 BUFX4_87 ( .A(_1020_), .Y(_1020__bF_buf4) );
BUFX4 BUFX4_88 ( .A(_1020_), .Y(_1020__bF_buf3) );
BUFX4 BUFX4_89 ( .A(_1020_), .Y(_1020__bF_buf2) );
BUFX4 BUFX4_90 ( .A(_1095_), .Y(_1095__bF_buf2) );
BUFX4 BUFX4_91 ( .A(_1020_), .Y(_1020__bF_buf1) );
BUFX4 BUFX4_92 ( .A(_1020_), .Y(_1020__bF_buf0) );
BUFX4 BUFX4_93 ( .A(_997_), .Y(_997__bF_buf3) );
BUFX4 BUFX4_94 ( .A(_997_), .Y(_997__bF_buf2) );
BUFX4 BUFX4_95 ( .A(_997_), .Y(_997__bF_buf1) );
BUFX4 BUFX4_96 ( .A(_997_), .Y(_997__bF_buf0) );
BUFX4 BUFX4_97 ( .A(_310_), .Y(_310__bF_buf3) );
BUFX4 BUFX4_98 ( .A(_310_), .Y(_310__bF_buf2) );
BUFX4 BUFX4_99 ( .A(_310_), .Y(_310__bF_buf1) );
BUFX4 BUFX4_100 ( .A(_310_), .Y(_310__bF_buf0) );
BUFX4 BUFX4_101 ( .A(_1095_), .Y(_1095__bF_buf1) );
BUFX4 BUFX4_102 ( .A(_1011_), .Y(_1011__bF_buf4) );
BUFX4 BUFX4_103 ( .A(_1011_), .Y(_1011__bF_buf3) );
BUFX4 BUFX4_104 ( .A(_1011_), .Y(_1011__bF_buf2) );
BUFX4 BUFX4_105 ( .A(_1011_), .Y(_1011__bF_buf1) );
BUFX4 BUFX4_106 ( .A(_1011_), .Y(_1011__bF_buf0) );
BUFX4 BUFX4_107 ( .A(_991_), .Y(_991__bF_buf6) );
BUFX4 BUFX4_108 ( .A(_991_), .Y(_991__bF_buf5) );
BUFX4 BUFX4_109 ( .A(_991_), .Y(_991__bF_buf4) );
BUFX4 BUFX4_110 ( .A(_991_), .Y(_991__bF_buf3) );
BUFX4 BUFX4_111 ( .A(_991_), .Y(_991__bF_buf2) );
BUFX4 BUFX4_112 ( .A(_1116_), .Y(_1116__bF_buf3) );
BUFX4 BUFX4_113 ( .A(_1095_), .Y(_1095__bF_buf0) );
BUFX4 BUFX4_114 ( .A(_991_), .Y(_991__bF_buf1) );
BUFX4 BUFX4_115 ( .A(_991_), .Y(_991__bF_buf0) );
BUFX4 BUFX4_116 ( .A(_1084_), .Y(_1084__bF_buf4) );
BUFX4 BUFX4_117 ( .A(_1084_), .Y(_1084__bF_buf3) );
BUFX4 BUFX4_118 ( .A(_1084_), .Y(_1084__bF_buf2) );
BUFX4 BUFX4_119 ( .A(_1084_), .Y(_1084__bF_buf1) );
BUFX4 BUFX4_120 ( .A(_1084_), .Y(_1084__bF_buf0) );
BUFX4 BUFX4_121 ( .A(_1102_), .Y(_1102__bF_buf3) );
BUFX4 BUFX4_122 ( .A(_1102_), .Y(_1102__bF_buf2) );
BUFX4 BUFX4_123 ( .A(_1102_), .Y(_1102__bF_buf1) );
BUFX4 BUFX4_124 ( .A(_996_), .Y(_996__bF_buf5) );
BUFX4 BUFX4_125 ( .A(_1102_), .Y(_1102__bF_buf0) );
BUFX4 BUFX4_126 ( .A(_527_), .Y(_527__bF_buf3) );
BUFX4 BUFX4_127 ( .A(_527_), .Y(_527__bF_buf2) );
BUFX4 BUFX4_128 ( .A(_527_), .Y(_527__bF_buf1) );
BUFX4 BUFX4_129 ( .A(_527_), .Y(_527__bF_buf0) );
BUFX4 BUFX4_130 ( .A(_1002_), .Y(_1002__bF_buf5) );
BUFX4 BUFX4_131 ( .A(_1002_), .Y(_1002__bF_buf4) );
BUFX4 BUFX4_132 ( .A(_1002_), .Y(_1002__bF_buf3) );
BUFX4 BUFX4_133 ( .A(_1002_), .Y(_1002__bF_buf2) );
BUFX4 BUFX4_134 ( .A(_1002_), .Y(_1002__bF_buf1) );
BUFX4 BUFX4_135 ( .A(_996_), .Y(_996__bF_buf4) );
BUFX4 BUFX4_136 ( .A(_1002_), .Y(_1002__bF_buf0) );
BUFX4 BUFX4_137 ( .A(_982_), .Y(_982__bF_buf6) );
BUFX4 BUFX4_138 ( .A(_982_), .Y(_982__bF_buf5) );
BUFX4 BUFX4_139 ( .A(_982_), .Y(_982__bF_buf4) );
BUFX4 BUFX4_140 ( .A(_982_), .Y(_982__bF_buf3) );
BUFX4 BUFX4_141 ( .A(_982_), .Y(_982__bF_buf2) );
BUFX4 BUFX4_142 ( .A(_982_), .Y(_982__bF_buf1) );
BUFX4 BUFX4_143 ( .A(_982_), .Y(_982__bF_buf0) );
BUFX4 BUFX4_144 ( .A(_996_), .Y(_996__bF_buf3) );
BUFX4 BUFX4_145 ( .A(_996_), .Y(_996__bF_buf2) );
BUFX4 BUFX4_146 ( .A(_996_), .Y(_996__bF_buf1) );
BUFX4 BUFX4_147 ( .A(_996_), .Y(_996__bF_buf0) );
BUFX4 BUFX4_148 ( .A(_1301_), .Y(_1301__bF_buf6) );
BUFX4 BUFX4_149 ( .A(_1301_), .Y(_1301__bF_buf5) );
BUFX4 BUFX4_150 ( .A(_1301_), .Y(_1301__bF_buf4) );
BUFX4 BUFX4_151 ( .A(_1116_), .Y(_1116__bF_buf2) );
BUFX4 BUFX4_152 ( .A(_1301_), .Y(_1301__bF_buf3) );
BUFX4 BUFX4_153 ( .A(_1301_), .Y(_1301__bF_buf2) );
BUFX4 BUFX4_154 ( .A(_1301_), .Y(_1301__bF_buf1) );
BUFX4 BUFX4_155 ( .A(_1301_), .Y(_1301__bF_buf0) );
BUFX4 BUFX4_156 ( .A(_1013_), .Y(_1013__bF_buf4) );
BUFX4 BUFX4_157 ( .A(_1013_), .Y(_1013__bF_buf3) );
BUFX4 BUFX4_158 ( .A(_1013_), .Y(_1013__bF_buf2) );
BUFX4 BUFX4_159 ( .A(_1013_), .Y(_1013__bF_buf1) );
BUFX4 BUFX4_160 ( .A(_1013_), .Y(_1013__bF_buf0) );
BUFX4 BUFX4_161 ( .A(_1201_), .Y(_1201__bF_buf4) );
BUFX4 BUFX4_162 ( .A(_1116_), .Y(_1116__bF_buf1) );
BUFX4 BUFX4_163 ( .A(_1201_), .Y(_1201__bF_buf3) );
BUFX4 BUFX4_164 ( .A(_1201_), .Y(_1201__bF_buf2) );
BUFX4 BUFX4_165 ( .A(_1201_), .Y(_1201__bF_buf1) );
BUFX4 BUFX4_166 ( .A(_1201_), .Y(_1201__bF_buf0) );
BUFX4 BUFX4_167 ( .A(clk), .Y(clk_bF_buf12) );
BUFX4 BUFX4_168 ( .A(clk), .Y(clk_bF_buf11) );
BUFX4 BUFX4_169 ( .A(clk), .Y(clk_bF_buf10) );
BUFX4 BUFX4_170 ( .A(clk), .Y(clk_bF_buf9) );
BUFX4 BUFX4_171 ( .A(clk), .Y(clk_bF_buf8) );
BUFX4 BUFX4_172 ( .A(clk), .Y(clk_bF_buf7) );
BUFX4 BUFX4_173 ( .A(_1116_), .Y(_1116__bF_buf0) );
BUFX4 BUFX4_174 ( .A(clk), .Y(clk_bF_buf6) );
BUFX4 BUFX4_175 ( .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_176 ( .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_177 ( .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_178 ( .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_179 ( .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_180 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_181 ( .A(_990_), .Y(_990__bF_buf3) );
BUFX4 BUFX4_182 ( .A(_990_), .Y(_990__bF_buf2) );
BUFX4 BUFX4_183 ( .A(_990_), .Y(_990__bF_buf1) );
BUFX4 BUFX4_184 ( .A(_1019_), .Y(_1019__bF_buf3) );
BUFX4 BUFX4_185 ( .A(_990_), .Y(_990__bF_buf0) );
BUFX4 BUFX4_186 ( .A(_987_), .Y(_987__bF_buf3) );
BUFX4 BUFX4_187 ( .A(_987_), .Y(_987__bF_buf2) );
BUFX4 BUFX4_188 ( .A(_987_), .Y(_987__bF_buf1) );
BUFX4 BUFX4_189 ( .A(_987_), .Y(_987__bF_buf0) );
BUFX4 BUFX4_190 ( .A(_1045_), .Y(_1045__bF_buf10) );
BUFX4 BUFX4_191 ( .A(_1045_), .Y(_1045__bF_buf9) );
BUFX4 BUFX4_192 ( .A(_1045_), .Y(_1045__bF_buf8) );
BUFX4 BUFX4_193 ( .A(_1045_), .Y(_1045__bF_buf7) );
BUFX4 BUFX4_194 ( .A(_1045_), .Y(_1045__bF_buf6) );
BUFX4 BUFX4_195 ( .A(_1019_), .Y(_1019__bF_buf2) );
BUFX4 BUFX4_196 ( .A(_1045_), .Y(_1045__bF_buf5) );
BUFX4 BUFX4_197 ( .A(_1045_), .Y(_1045__bF_buf4) );
BUFX4 BUFX4_198 ( .A(_1045_), .Y(_1045__bF_buf3) );
BUFX4 BUFX4_199 ( .A(_1045_), .Y(_1045__bF_buf2) );
BUFX4 BUFX4_200 ( .A(_1045_), .Y(_1045__bF_buf1) );
BUFX4 BUFX4_201 ( .A(_1045_), .Y(_1045__bF_buf0) );
BUFX4 BUFX4_202 ( .A(_1004_), .Y(_1004__bF_buf3) );
BUFX4 BUFX4_203 ( .A(_1004_), .Y(_1004__bF_buf2) );
BUFX4 BUFX4_204 ( .A(_1004_), .Y(_1004__bF_buf1) );
BUFX4 BUFX4_205 ( .A(_1004_), .Y(_1004__bF_buf0) );
BUFX4 BUFX4_206 ( .A(_1019_), .Y(_1019__bF_buf1) );
BUFX4 BUFX4_207 ( .A(_1080_), .Y(_1080__bF_buf4) );
BUFX4 BUFX4_208 ( .A(_1080_), .Y(_1080__bF_buf3) );
BUFX4 BUFX4_209 ( .A(_1080_), .Y(_1080__bF_buf2) );
BUFX4 BUFX4_210 ( .A(_1080_), .Y(_1080__bF_buf1) );
BUFX4 BUFX4_211 ( .A(_1080_), .Y(_1080__bF_buf0) );
BUFX4 BUFX4_212 ( .A(_1030_), .Y(_1030__bF_buf9) );
BUFX4 BUFX4_213 ( .A(_1030_), .Y(_1030__bF_buf8) );
BUFX4 BUFX4_214 ( .A(_1030_), .Y(_1030__bF_buf7) );
BUFX4 BUFX4_215 ( .A(_1030_), .Y(_1030__bF_buf6) );
BUFX4 BUFX4_216 ( .A(_1030_), .Y(_1030__bF_buf5) );
BUFX4 BUFX4_217 ( .A(_1019_), .Y(_1019__bF_buf0) );
BUFX4 BUFX4_218 ( .A(_1030_), .Y(_1030__bF_buf4) );
BUFX4 BUFX4_219 ( .A(_1030_), .Y(_1030__bF_buf3) );
BUFX4 BUFX4_220 ( .A(_1030_), .Y(_1030__bF_buf2) );
BUFX4 BUFX4_221 ( .A(_1030_), .Y(_1030__bF_buf1) );
BUFX4 BUFX4_222 ( .A(_1030_), .Y(_1030__bF_buf0) );
BUFX4 BUFX4_223 ( .A(_1250_), .Y(_1250__bF_buf4) );
BUFX4 BUFX4_224 ( .A(_1250_), .Y(_1250__bF_buf3) );
BUFX4 BUFX4_225 ( .A(_1250_), .Y(_1250__bF_buf2) );
BUFX4 BUFX4_226 ( .A(_1250_), .Y(_1250__bF_buf1) );
BUFX4 BUFX4_227 ( .A(_1250_), .Y(_1250__bF_buf0) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf9), .D(_17_), .Q(delay) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf9), .D(_1543__4_), .Q(ADDR_stack_0__4_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf0), .D(_13__4_), .Q(PC_STACK_7__4_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf11), .D(_13__5_), .Q(PC_STACK_7__5_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf6), .D(_13__6_), .Q(PC_STACK_7__6_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf9), .D(_13__7_), .Q(PC_STACK_7__7_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf0), .D(_13__8_), .Q(PC_STACK_7__8_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf0), .D(_13__9_), .Q(PC_STACK_7__9_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf8), .D(_14__0_), .Q(PC_STACK_8__0_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf7), .D(_14__1_), .Q(PC_STACK_8__1_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf5), .D(_14__2_), .Q(PC_STACK_8__2_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf1), .D(_14__3_), .Q(PC_STACK_8__3_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf9), .D(_1543__5_), .Q(ADDR_stack_0__5_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf1), .D(_14__4_), .Q(PC_STACK_8__4_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf7), .D(_14__5_), .Q(PC_STACK_8__5_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf1), .D(_14__6_), .Q(PC_STACK_8__6_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf2), .D(_14__7_), .Q(PC_STACK_8__7_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf10), .D(_14__8_), .Q(PC_STACK_8__8_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf10), .D(_14__9_), .Q(PC_STACK_8__9_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf7), .D(_15__0_), .Q(PC_STACK_9__0_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf8), .D(_15__1_), .Q(PC_STACK_9__1_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf10), .D(_15__2_), .Q(PC_STACK_9__2_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf7), .D(_15__3_), .Q(PC_STACK_9__3_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf9), .D(_1543__6_), .Q(ADDR_stack_0__6_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf8), .D(_15__4_), .Q(PC_STACK_9__4_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf1), .D(_15__5_), .Q(PC_STACK_9__5_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf7), .D(_15__6_), .Q(PC_STACK_9__6_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf10), .D(_15__7_), .Q(PC_STACK_9__7_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf10), .D(_15__8_), .Q(PC_STACK_9__8_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf10), .D(_15__9_), .Q(PC_STACK_9__9_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf1), .D(_1__0_), .Q(PC_STACK_10__0_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf1), .D(_1__1_), .Q(PC_STACK_10__1_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf1), .D(_1__2_), .Q(PC_STACK_10__2_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf7), .D(_1__3_), .Q(PC_STACK_10__3_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf9), .D(_1543__7_), .Q(ADDR_stack_0__7_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf1), .D(_1__4_), .Q(PC_STACK_10__4_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf1), .D(_1__5_), .Q(PC_STACK_10__5_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf10), .D(_1__6_), .Q(PC_STACK_10__6_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf2), .D(_1__7_), .Q(PC_STACK_10__7_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf1), .D(_1__8_), .Q(PC_STACK_10__8_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf10), .D(_1__9_), .Q(PC_STACK_10__9_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf8), .D(_2__0_), .Q(PC_STACK_11__0_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf8), .D(_2__1_), .Q(PC_STACK_11__1_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf8), .D(_2__2_), .Q(PC_STACK_11__2_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf8), .D(_2__3_), .Q(PC_STACK_11__3_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf9), .D(_1543__8_), .Q(ADDR_stack_0__8_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf1), .D(_2__4_), .Q(PC_STACK_11__4_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf8), .D(_2__5_), .Q(PC_STACK_11__5_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf1), .D(_2__6_), .Q(PC_STACK_11__6_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf2), .D(_2__7_), .Q(PC_STACK_11__7_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf10), .D(_2__8_), .Q(PC_STACK_11__8_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf10), .D(_2__9_), .Q(PC_STACK_11__9_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf4), .D(_3__0_), .Q(PC_STACK_12__0_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf11), .D(_3__1_), .Q(PC_STACK_12__1_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf4), .D(_3__2_), .Q(PC_STACK_12__2_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf4), .D(_3__3_), .Q(PC_STACK_12__3_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf1), .D(_1543__9_), .Q(ADDR_stack_0__9_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf11), .D(_3__4_), .Q(PC_STACK_12__4_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf11), .D(_3__5_), .Q(PC_STACK_12__5_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf11), .D(_3__6_), .Q(PC_STACK_12__6_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf6), .D(_3__7_), .Q(PC_STACK_12__7_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf2), .D(_3__8_), .Q(PC_STACK_12__8_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf11), .D(_3__9_), .Q(PC_STACK_12__9_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf7), .D(_4__0_), .Q(PC_STACK_13__0_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf8), .D(_4__1_), .Q(PC_STACK_13__1_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf8), .D(_4__2_), .Q(PC_STACK_13__2_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf7), .D(_4__3_), .Q(PC_STACK_13__3_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf5), .D(ADDR_stack_0__0_), .Q(_1545__0_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf7), .D(_4__4_), .Q(PC_STACK_13__4_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf7), .D(_4__5_), .Q(PC_STACK_13__5_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf10), .D(_4__6_), .Q(PC_STACK_13__6_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf10), .D(_4__7_), .Q(PC_STACK_13__7_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf10), .D(_4__8_), .Q(PC_STACK_13__8_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf4), .D(_4__9_), .Q(PC_STACK_13__9_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf4), .D(_5__0_), .Q(PC_STACK_14__0_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf4), .D(_5__1_), .Q(PC_STACK_14__1_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf10), .D(_5__2_), .Q(PC_STACK_14__2_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf2), .D(_5__3_), .Q(PC_STACK_14__3_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf12), .D(ADDR_stack_0__1_), .Q(_1545__1_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf3), .D(_5__4_), .Q(PC_STACK_14__4_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf3), .D(_5__5_), .Q(PC_STACK_14__5_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf4), .D(_5__6_), .Q(PC_STACK_14__6_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf2), .D(_5__7_), .Q(PC_STACK_14__7_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf2), .D(_5__8_), .Q(PC_STACK_14__8_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf2), .D(_5__9_), .Q(PC_STACK_14__9_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf8), .D(_6__0_), .Q(PC_STACK_15__0_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf8), .D(_6__1_), .Q(PC_STACK_15__1_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf8), .D(_6__2_), .Q(PC_STACK_15__2_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf6), .D(_6__3_), .Q(PC_STACK_15__3_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf5), .D(ADDR_stack_0__2_), .Q(_1545__2_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf8), .D(_6__4_), .Q(PC_STACK_15__4_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf5), .D(_6__5_), .Q(PC_STACK_15__5_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf7), .D(_6__6_), .Q(PC_STACK_15__6_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf2), .D(_6__7_), .Q(PC_STACK_15__7_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf2), .D(_6__8_), .Q(PC_STACK_15__8_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf10), .D(_6__9_), .Q(PC_STACK_15__9_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf5), .D(ADDR_stack_0__3_), .Q(_1545__3_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf5), .D(_16__0_), .Q(PC_pointer_0_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf9), .D(ADDR_stack_0__4_), .Q(_1545__4_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf9), .D(ADDR_stack_0__5_), .Q(_1545__5_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf9), .D(ADDR_stack_0__6_), .Q(_1545__6_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf9), .D(ADDR_stack_0__7_), .Q(_1545__7_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf9), .D(ADDR_stack_0__8_), .Q(_1545__8_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf1), .D(ADDR_stack_0__9_), .Q(_1545__9_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf5), .D(_0__0_), .Q(PC_STACK_0__0_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf5), .D(_0__1_), .Q(PC_STACK_0__1_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf5), .D(_0__2_), .Q(PC_STACK_0__2_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf3), .D(_0__3_), .Q(PC_STACK_0__3_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf3), .D(_16__1_), .Q(PC_pointer_1_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf3), .D(_0__4_), .Q(PC_STACK_0__4_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf5), .D(_0__5_), .Q(PC_STACK_0__5_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf2), .D(_0__6_), .Q(PC_STACK_0__6_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf6), .D(_0__7_), .Q(PC_STACK_0__7_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf7), .D(_0__8_), .Q(PC_STACK_0__8_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf3), .D(_0__9_), .Q(PC_STACK_0__9_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf4), .D(_7__0_), .Q(PC_STACK_1__0_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf12), .D(_7__1_), .Q(PC_STACK_1__1_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf3), .D(_7__2_), .Q(PC_STACK_1__2_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf0), .D(_7__3_), .Q(PC_STACK_1__3_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf3), .D(_16__2_), .Q(PC_pointer_2_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf0), .D(_7__4_), .Q(PC_STACK_1__4_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf11), .D(_7__5_), .Q(PC_STACK_1__5_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf2), .D(_7__6_), .Q(PC_STACK_1__6_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf6), .D(_7__7_), .Q(PC_STACK_1__7_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf11), .D(_7__8_), .Q(PC_STACK_1__8_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf11), .D(_7__9_), .Q(PC_STACK_1__9_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf12), .D(_8__0_), .Q(PC_STACK_2__0_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf3), .D(_8__1_), .Q(PC_STACK_2__1_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf3), .D(_8__2_), .Q(PC_STACK_2__2_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf12), .D(_8__3_), .Q(PC_STACK_2__3_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf3), .D(_16__3_), .Q(PC_pointer_3_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf3), .D(_8__4_), .Q(PC_STACK_2__4_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf12), .D(_8__5_), .Q(PC_STACK_2__5_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf11), .D(_8__6_), .Q(PC_STACK_2__6_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf6), .D(_8__7_), .Q(PC_STACK_2__7_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf11), .D(_8__8_), .Q(PC_STACK_2__8_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf0), .D(_8__9_), .Q(PC_STACK_2__9_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf12), .D(_9__0_), .Q(PC_STACK_3__0_) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf12), .D(_9__1_), .Q(PC_STACK_3__1_) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf5), .D(_9__2_), .Q(PC_STACK_3__2_) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf12), .D(_9__3_), .Q(PC_STACK_3__3_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf5), .D(_1543__0_), .Q(ADDR_stack_0__0_) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf0), .D(_9__4_), .Q(PC_STACK_3__4_) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf12), .D(_9__5_), .Q(PC_STACK_3__5_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf6), .D(_9__6_), .Q(PC_STACK_3__6_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf9), .D(_9__7_), .Q(PC_STACK_3__7_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf11), .D(_9__8_), .Q(PC_STACK_3__8_) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf0), .D(_9__9_), .Q(PC_STACK_3__9_) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf4), .D(_10__0_), .Q(PC_STACK_4__0_) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf4), .D(_10__1_), .Q(PC_STACK_4__1_) );
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf3), .D(_10__2_), .Q(PC_STACK_4__2_) );
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf7), .D(_10__3_), .Q(PC_STACK_4__3_) );
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf12), .D(_1543__1_), .Q(ADDR_stack_0__1_) );
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf12), .D(_10__4_), .Q(PC_STACK_4__4_) );
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf11), .D(_10__5_), .Q(PC_STACK_4__5_) );
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf6), .D(_10__6_), .Q(PC_STACK_4__6_) );
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf6), .D(_10__7_), .Q(PC_STACK_4__7_) );
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf11), .D(_10__8_), .Q(PC_STACK_4__8_) );
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf11), .D(_10__9_), .Q(PC_STACK_4__9_) );
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf4), .D(_11__0_), .Q(PC_STACK_5__0_) );
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf4), .D(_11__1_), .Q(PC_STACK_5__1_) );
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf4), .D(_11__2_), .Q(PC_STACK_5__2_) );
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf2), .D(_11__3_), .Q(PC_STACK_5__3_) );
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf5), .D(_1543__2_), .Q(ADDR_stack_0__2_) );
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf2), .D(_11__4_), .Q(PC_STACK_5__4_) );
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf6), .D(_11__5_), .Q(PC_STACK_5__5_) );
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf6), .D(_11__6_), .Q(PC_STACK_5__6_) );
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf6), .D(_11__7_), .Q(PC_STACK_5__7_) );
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf9), .D(_11__8_), .Q(PC_STACK_5__8_) );
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf6), .D(_11__9_), .Q(PC_STACK_5__9_) );
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf3), .D(_12__0_), .Q(PC_STACK_6__0_) );
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf12), .D(_12__1_), .Q(PC_STACK_6__1_) );
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf7), .D(_12__2_), .Q(PC_STACK_6__2_) );
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf0), .D(_12__3_), .Q(PC_STACK_6__3_) );
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf5), .D(_1543__3_), .Q(ADDR_stack_0__3_) );
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf12), .D(_12__4_), .Q(PC_STACK_6__4_) );
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf0), .D(_12__5_), .Q(PC_STACK_6__5_) );
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf0), .D(_12__6_), .Q(PC_STACK_6__6_) );
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf6), .D(_12__7_), .Q(PC_STACK_6__7_) );
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf0), .D(_12__8_), .Q(PC_STACK_6__8_) );
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf0), .D(_12__9_), .Q(PC_STACK_6__9_) );
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf12), .D(_13__0_), .Q(PC_STACK_7__0_) );
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf12), .D(_13__1_), .Q(PC_STACK_7__1_) );
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf4), .D(_13__2_), .Q(PC_STACK_7__2_) );
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf0), .D(_13__3_), .Q(PC_STACK_7__3_) );
INVX1 INVX1_1 ( .A(PC_STACK_2__0_), .Y(_1008_) );
INVX1 INVX1_2 ( .A(PC_STACK_2__2_), .Y(_1078_) );
INVX1 INVX1_3 ( .A(_862_), .Y(_863_) );
INVX1 INVX1_4 ( .A(_880_), .Y(_881_) );
INVX1 INVX1_5 ( .A(_933_), .Y(_934_) );
INVX1 INVX1_6 ( .A(clk_bF_buf9), .Y(_962_) );
INVX1 INVX1_7 ( .A(CORE_PC_ctrl[1]), .Y(_963_) );
INVX1 INVX1_8 ( .A(IDATA_CORE_out[0]), .Y(_966_) );
INVX1 INVX1_9 ( .A(IDATA_CORE_out[1]), .Y(_967_) );
INVX1 INVX1_10 ( .A(IDATA_CORE_out[2]), .Y(_968_) );
INVX1 INVX1_11 ( .A(IDATA_CORE_out[3]), .Y(_969_) );
INVX1 INVX1_12 ( .A(IDATA_CORE_out[4]), .Y(_970_) );
INVX1 INVX1_13 ( .A(PC_STACK_11__2_), .Y(_1082_) );
INVX1 INVX1_14 ( .A(IDATA_CORE_out[5]), .Y(_971_) );
INVX1 INVX1_15 ( .A(IDATA_CORE_out[6]), .Y(_972_) );
INVX1 INVX1_16 ( .A(IDATA_CORE_out[7]), .Y(_973_) );
INVX1 INVX1_17 ( .A(IDATA_CORE_out[8]), .Y(_974_) );
INVX1 INVX1_18 ( .A(IDATA_CORE_out[9]), .Y(_975_) );
INVX1 INVX1_19 ( .A(IDATA_CORE_out[10]), .Y(_976_) );
INVX1 INVX1_20 ( .A(IDATA_CORE_out[11]), .Y(_977_) );
INVX1 INVX1_21 ( .A(IDATA_CORE_out[12]), .Y(_978_) );
INVX1 INVX1_22 ( .A(IDATA_CORE_out[13]), .Y(_979_) );
INVX1 INVX1_23 ( .A(IDATA_CORE_out[14]), .Y(_980_) );
INVX1 INVX1_24 ( .A(PC_STACK_15__2_), .Y(_1083_) );
INVX1 INVX1_25 ( .A(PC_STACK_14__2_), .Y(_1091_) );
INVX1 INVX1_26 ( .A(PC_STACK_8__2_), .Y(_1093_) );
INVX1 INVX1_27 ( .A(PC_STACK_0__2_), .Y(_1097_) );
INVX1 INVX1_28 ( .A(PC_STACK_3__2_), .Y(_1098_) );
INVX1 INVX1_29 ( .A(PC_STACK_14__0_), .Y(_1107_) );
INVX1 INVX1_30 ( .A(PC_STACK_13__0_), .Y(_1108_) );
INVX1 INVX1_31 ( .A(PC_STACK_12__0_), .Y(_1114_) );
INVX1 INVX1_32 ( .A(PC_STACK_3__0_), .Y(_1009_) );
INVX1 INVX1_33 ( .A(PC_STACK_1__0_), .Y(_1115_) );
INVX1 INVX1_34 ( .A(PC_STACK_8__0_), .Y(_1119_) );
INVX1 INVX1_35 ( .A(PC_STACK_15__0_), .Y(_1120_) );
INVX1 INVX1_36 ( .A(PC_STACK_14__1_), .Y(_1124_) );
INVX1 INVX1_37 ( .A(PC_STACK_13__1_), .Y(_1125_) );
INVX1 INVX1_38 ( .A(PC_STACK_12__1_), .Y(_1130_) );
INVX1 INVX1_39 ( .A(PC_STACK_1__1_), .Y(_1131_) );
INVX1 INVX1_40 ( .A(PC_STACK_8__1_), .Y(_1133_) );
INVX1 INVX1_41 ( .A(PC_STACK_15__1_), .Y(_1134_) );
INVX1 INVX1_42 ( .A(PC_STACK_13__3_), .Y(_1151_) );
INVX1 INVX1_43 ( .A(PC_STACK_6__0_), .Y(_1015_) );
INVX1 INVX1_44 ( .A(PC_STACK_2__3_), .Y(_1152_) );
INVX1 INVX1_45 ( .A(PC_STACK_11__3_), .Y(_1154_) );
INVX1 INVX1_46 ( .A(PC_STACK_8__3_), .Y(_1155_) );
INVX1 INVX1_47 ( .A(PC_STACK_15__3_), .Y(_1161_) );
INVX1 INVX1_48 ( .A(PC_STACK_14__3_), .Y(_1162_) );
INVX1 INVX1_49 ( .A(PC_STACK_0__3_), .Y(_1164_) );
INVX1 INVX1_50 ( .A(PC_STACK_6__3_), .Y(_1166_) );
INVX1 INVX1_51 ( .A(PC_STACK_3__3_), .Y(_1169_) );
INVX1 INVX1_52 ( .A(PC_STACK_1__3_), .Y(_1173_) );
INVX1 INVX1_53 ( .A(PC_STACK_7__3_), .Y(_1174_) );
INVX1 INVX1_54 ( .A(PC_STACK_7__0_), .Y(_1016_) );
INVX1 INVX1_55 ( .A(PC_STACK_9__4_), .Y(_1199_) );
INVX1 INVX1_56 ( .A(PC_STACK_15__4_), .Y(_1200_) );
INVX1 INVX1_57 ( .A(PC_STACK_8__4_), .Y(_1203_) );
INVX1 INVX1_58 ( .A(PC_STACK_13__4_), .Y(_1204_) );
INVX1 INVX1_59 ( .A(_1235_), .Y(_1543__5_) );
INVX1 INVX1_60 ( .A(PC_STACK_2__6_), .Y(_1248_) );
INVX1 INVX1_61 ( .A(PC_STACK_4__6_), .Y(_1249_) );
INVX1 INVX1_62 ( .A(PC_STACK_11__6_), .Y(_1252_) );
INVX1 INVX1_63 ( .A(PC_STACK_14__6_), .Y(_1253_) );
INVX1 INVX1_64 ( .A(PC_STACK_9__6_), .Y(_1259_) );
INVX1 INVX1_65 ( .A(PC_STACK_2__1_), .Y(_1054_) );
INVX1 INVX1_66 ( .A(PC_STACK_8__6_), .Y(_1260_) );
INVX1 INVX1_67 ( .A(PC_STACK_15__6_), .Y(_1262_) );
INVX1 INVX1_68 ( .A(PC_STACK_13__6_), .Y(_1263_) );
INVX1 INVX1_69 ( .A(_1270_), .Y(_1271_) );
INVX1 INVX1_70 ( .A(PC_STACK_13__7_), .Y(_1284_) );
INVX1 INVX1_71 ( .A(PC_STACK_3__7_), .Y(_1287_) );
INVX1 INVX1_72 ( .A(PC_STACK_7__7_), .Y(_1288_) );
INVX1 INVX1_73 ( .A(_1300_), .Y(_1543__7_) );
INVX1 INVX1_74 ( .A(_1038__bF_buf9), .Y(_1307_) );
INVX1 INVX1_75 ( .A(PC_STACK_13__8_), .Y(_1320_) );
INVX1 INVX1_76 ( .A(PC_STACK_3__1_), .Y(_1055_) );
INVX1 INVX1_77 ( .A(PC_STACK_12__8_), .Y(_1321_) );
INVX1 INVX1_78 ( .A(PC_STACK_15__8_), .Y(_1323_) );
INVX1 INVX1_79 ( .A(PC_STACK_14__8_), .Y(_1324_) );
INVX1 INVX1_80 ( .A(PC_STACK_2__8_), .Y(_1328_) );
INVX1 INVX1_81 ( .A(PC_STACK_7__8_), .Y(_1329_) );
INVX1 INVX1_82 ( .A(PC_STACK_4__8_), .Y(_1332_) );
INVX1 INVX1_83 ( .A(PC_STACK_0__8_), .Y(_1333_) );
INVX1 INVX1_84 ( .A(_1339_), .Y(_1340_) );
INVX1 INVX1_85 ( .A(PC_STACK_0__9_), .Y(_1349_) );
INVX1 INVX1_86 ( .A(PC_STACK_7__9_), .Y(_1353_) );
INVX1 INVX1_87 ( .A(PC_STACK_6__1_), .Y(_1057_) );
INVX1 INVX1_88 ( .A(PC_STACK_13__9_), .Y(_1355_) );
INVX1 INVX1_89 ( .A(PC_STACK_4__9_), .Y(_1356_) );
INVX1 INVX1_90 ( .A(_1543__9_), .Y(_1366_) );
INVX1 INVX1_91 ( .A(_1418_), .Y(_1419_) );
INVX1 INVX1_92 ( .A(_1442_), .Y(_1443_) );
INVX1 INVX1_93 ( .A(_1492_), .Y(_1493_) );
INVX1 INVX1_94 ( .A(_41_), .Y(_42_) );
INVX1 INVX1_95 ( .A(_137_), .Y(_138_) );
INVX1 INVX1_96 ( .A(_208_), .Y(_209_) );
INVX1 INVX1_97 ( .A(_230_), .Y(_231_) );
INVX1 INVX1_98 ( .A(PC_STACK_7__1_), .Y(_1058_) );
INVX1 INVX1_99 ( .A(_280_), .Y(_281_) );
INVX1 INVX1_100 ( .A(_298_), .Y(_299_) );
INVX1 INVX1_101 ( .A(_302_), .Y(_303_) );
INVX1 INVX1_102 ( .A(_353_), .Y(_354_) );
INVX1 INVX1_103 ( .A(_371_), .Y(_372_) );
INVX1 INVX1_104 ( .A(_426_), .Y(_427_) );
INVX1 INVX1_105 ( .A(_444_), .Y(_445_) );
INVX1 INVX1_106 ( .A(_497_), .Y(_498_) );
INVX1 INVX1_107 ( .A(_515_), .Y(_516_) );
INVX1 INVX1_108 ( .A(_519_), .Y(_520_) );
INVX1 INVX1_109 ( .A(PC_STACK_13__2_), .Y(_1077_) );
INVX1 INVX1_110 ( .A(_570_), .Y(_571_) );
INVX1 INVX1_111 ( .A(_588_), .Y(_589_) );
INVX1 INVX1_112 ( .A(_592_), .Y(_593_) );
INVX1 INVX1_113 ( .A(PC_STACK_5__9_), .Y(_595_) );
INVX1 INVX1_114 ( .A(_643_), .Y(_644_) );
INVX1 INVX1_115 ( .A(_665_), .Y(_666_) );
INVX1 INVX1_116 ( .A(_715_), .Y(_716_) );
INVX1 INVX1_117 ( .A(_733_), .Y(_734_) );
INVX1 INVX1_118 ( .A(_737_), .Y(_738_) );
INVX1 INVX1_119 ( .A(_789_), .Y(_790_) );
INVX2 INVX2_1 ( .A(_1269_), .Y(_1543__6_) );
INVX2 INVX2_2 ( .A(_1338_), .Y(_1543__8_) );
INVX2 INVX2_3 ( .A(CORE_STACK_ctrl[0]), .Y(_70_) );
INVX2 INVX2_4 ( .A(CORE_STACK_ctrl[1]), .Y(_71_) );
INVX2 INVX2_5 ( .A(_76_), .Y(_77_) );
INVX4 INVX4_1 ( .A(PC_pointer_3_), .Y(_981_) );
INVX4 INVX4_2 ( .A(PC_pointer_1_), .Y(_985_) );
INVX4 INVX4_3 ( .A(PC_pointer_2_), .Y(_995_) );
INVX4 INVX4_4 ( .A(PC_pointer_0_), .Y(_998_) );
INVX8 INVX8_1 ( .A(INTERRUPT_ch[0]), .Y(_1035_) );
INVX8 INVX8_2 ( .A(_997__bF_buf1), .Y(_1201_) );
INVX8 INVX8_3 ( .A(INTERRUPT_ch[4]), .Y(_1217_) );
INVX8 INVX8_4 ( .A(INTERRUPT_ch[5]), .Y(_1242_) );
INVX8 INVX8_5 ( .A(_1030__bF_buf9), .Y(_1301_) );
INVX8 INVX8_6 ( .A(_1045__bF_buf0), .Y(_1311_) );
INVX8 INVX8_7 ( .A(INTERRUPT_ch[6]), .Y(_1497_) );
INVX8 INVX8_8 ( .A(INTERRUPT_ch[7]), .Y(_1504_) );
INVX8 INVX8_9 ( .A(_1000__bF_buf2), .Y(_310_) );
INVX8 INVX8_10 ( .A(_987__bF_buf1), .Y(_527_) );
INVX8 INVX8_11 ( .A(INTERRUPT_flag), .Y(_1037_) );
INVX8 INVX8_12 ( .A(CORE_PC_ctrl[0]), .Y(_1040_) );
INVX8 INVX8_13 ( .A(rst_bF_buf0), .Y(_1042_) );
INVX8 INVX8_14 ( .A(INTERRUPT_ch[1]), .Y(_1073_) );
INVX8 INVX8_15 ( .A(_1020__bF_buf1), .Y(_1104_) );
INVX8 INVX8_16 ( .A(INTERRUPT_ch[2]), .Y(_1148_) );
INVX8 INVX8_17 ( .A(INTERRUPT_ch[3]), .Y(_1185_) );
INVX8 INVX8_18 ( .A(_1011__bF_buf2), .Y(_1191_) );
NAND2X1 NAND2X1_1 ( .A(PC_pointer_2_), .B(_981_), .Y(_982_) );
NAND2X1 NAND2X1_2 ( .A(_1017_), .B(_1018_), .Y(_1019_) );
NAND2X1 NAND2X1_3 ( .A(_1038__bF_buf7), .B(_37_), .Y(_38_) );
NAND2X1 NAND2X1_4 ( .A(PC_STACK_14__6_), .B(_1041__bF_buf4), .Y(_45_) );
NAND2X1 NAND2X1_5 ( .A(_1280_), .B(_1023_), .Y(_47_) );
NAND2X1 NAND2X1_6 ( .A(PC_STACK_14__7_), .B(_1041__bF_buf3), .Y(_54_) );
NAND2X1 NAND2X1_7 ( .A(_1313_), .B(_1023_), .Y(_55_) );
NAND2X1 NAND2X1_8 ( .A(_1037_), .B(_70_), .Y(_74_) );
NAND2X1 NAND2X1_9 ( .A(_1002__bF_buf2), .B(_983__bF_buf1), .Y(_78_) );
NAND2X1 NAND2X1_10 ( .A(PC_pointer_2_), .B(_1012_), .Y(_81_) );
NAND2X1 NAND2X1_11 ( .A(_1030__bF_buf3), .B(_94_), .Y(_95_) );
NAND2X1 NAND2X1_12 ( .A(_1038__bF_buf8), .B(_96_), .Y(_97_) );
NAND2X1 NAND2X1_13 ( .A(_1024_), .B(_1027_), .Y(_1028_) );
NAND2X1 NAND2X1_14 ( .A(_1030__bF_buf3), .B(_101_), .Y(_102_) );
NAND2X1 NAND2X1_15 ( .A(_1045__bF_buf4), .B(_103_), .Y(_104_) );
NAND2X1 NAND2X1_16 ( .A(_1030__bF_buf4), .B(_108_), .Y(_109_) );
NAND2X1 NAND2X1_17 ( .A(_1045__bF_buf4), .B(_110_), .Y(_111_) );
NAND2X1 NAND2X1_18 ( .A(_1030__bF_buf3), .B(_115_), .Y(_116_) );
NAND2X1 NAND2X1_19 ( .A(_1038__bF_buf4), .B(_117_), .Y(_118_) );
NAND2X1 NAND2X1_20 ( .A(_1030__bF_buf3), .B(_122_), .Y(_123_) );
NAND2X1 NAND2X1_21 ( .A(_1038__bF_buf4), .B(_124_), .Y(_125_) );
NAND2X1 NAND2X1_22 ( .A(_1104_), .B(_1239_), .Y(_128_) );
NAND2X1 NAND2X1_23 ( .A(PC_STACK_7__5_), .B(_1041__bF_buf10), .Y(_132_) );
NAND2X1 NAND2X1_24 ( .A(_1029_), .B(_1007_), .Y(_1543__0_) );
NAND2X1 NAND2X1_25 ( .A(_1045__bF_buf10), .B(_133_), .Y(_134_) );
NAND2X1 NAND2X1_26 ( .A(_132_), .B(_134_), .Y(_135_) );
NAND2X1 NAND2X1_27 ( .A(PC_STACK_7__6_), .B(_1041__bF_buf3), .Y(_141_) );
NAND2X1 NAND2X1_28 ( .A(_1280_), .B(_1104_), .Y(_143_) );
NAND2X1 NAND2X1_29 ( .A(_137_), .B(_143_), .Y(_144_) );
NAND2X1 NAND2X1_30 ( .A(PC_STACK_7__7_), .B(_1041__bF_buf3), .Y(_150_) );
NAND2X1 NAND2X1_31 ( .A(_1313_), .B(_1104_), .Y(_151_) );
NAND2X1 NAND2X1_32 ( .A(_1030__bF_buf8), .B(_167_), .Y(_168_) );
NAND2X1 NAND2X1_33 ( .A(_1038__bF_buf0), .B(_169_), .Y(_170_) );
NAND2X1 NAND2X1_34 ( .A(_1030__bF_buf2), .B(_174_), .Y(_175_) );
NAND2X1 NAND2X1_35 ( .A(_1030__bF_buf1), .B(_1033_), .Y(_1034_) );
NAND2X1 NAND2X1_36 ( .A(_1045__bF_buf8), .B(_176_), .Y(_177_) );
NAND2X1 NAND2X1_37 ( .A(_1030__bF_buf2), .B(_181_), .Y(_182_) );
NAND2X1 NAND2X1_38 ( .A(_1045__bF_buf8), .B(_183_), .Y(_184_) );
NAND2X1 NAND2X1_39 ( .A(_1030__bF_buf5), .B(_188_), .Y(_189_) );
NAND2X1 NAND2X1_40 ( .A(_1038__bF_buf5), .B(_190_), .Y(_191_) );
NAND2X1 NAND2X1_41 ( .A(_1030__bF_buf2), .B(_195_), .Y(_196_) );
NAND2X1 NAND2X1_42 ( .A(_1038__bF_buf1), .B(_197_), .Y(_198_) );
NAND2X1 NAND2X1_43 ( .A(_1030__bF_buf2), .B(_202_), .Y(_203_) );
NAND2X1 NAND2X1_44 ( .A(_1038__bF_buf1), .B(_204_), .Y(_205_) );
NAND2X1 NAND2X1_45 ( .A(PC_STACK_15__6_), .B(_1041__bF_buf0), .Y(_212_) );
NAND2X1 NAND2X1_46 ( .A(_1038__bF_buf7), .B(_1036_), .Y(_1039_) );
NAND2X1 NAND2X1_47 ( .A(_1280_), .B(_1003_), .Y(_214_) );
NAND2X1 NAND2X1_48 ( .A(PC_STACK_15__7_), .B(_1041__bF_buf3), .Y(_221_) );
NAND2X1 NAND2X1_49 ( .A(_1313_), .B(_1003_), .Y(_222_) );
NAND2X1 NAND2X1_50 ( .A(_1030__bF_buf6), .B(_239_), .Y(_240_) );
NAND2X1 NAND2X1_51 ( .A(_1038__bF_buf6), .B(_241_), .Y(_242_) );
NAND2X1 NAND2X1_52 ( .A(_1030__bF_buf6), .B(_246_), .Y(_247_) );
NAND2X1 NAND2X1_53 ( .A(_1045__bF_buf7), .B(_248_), .Y(_249_) );
NAND2X1 NAND2X1_54 ( .A(_1030__bF_buf9), .B(_253_), .Y(_254_) );
NAND2X1 NAND2X1_55 ( .A(_1045__bF_buf2), .B(_255_), .Y(_256_) );
NAND2X1 NAND2X1_56 ( .A(_1030__bF_buf6), .B(_260_), .Y(_261_) );
NAND2X1 NAND2X1_57 ( .A(ULA_OUT[0]), .B(_1042_), .Y(_1043_) );
NAND2X1 NAND2X1_58 ( .A(_1038__bF_buf3), .B(_262_), .Y(_263_) );
NAND2X1 NAND2X1_59 ( .A(_1030__bF_buf6), .B(_267_), .Y(_268_) );
NAND2X1 NAND2X1_60 ( .A(_1038__bF_buf0), .B(_269_), .Y(_270_) );
NAND2X1 NAND2X1_61 ( .A(_1030__bF_buf6), .B(_274_), .Y(_275_) );
NAND2X1 NAND2X1_62 ( .A(_1038__bF_buf0), .B(_276_), .Y(_277_) );
NAND2X1 NAND2X1_63 ( .A(PC_STACK_9__6_), .B(_1041__bF_buf0), .Y(_284_) );
NAND2X1 NAND2X1_64 ( .A(_1280_), .B(_997__bF_buf1), .Y(_286_) );
NAND2X1 NAND2X1_65 ( .A(PC_STACK_9__7_), .B(_1041__bF_buf0), .Y(_293_) );
NAND2X1 NAND2X1_66 ( .A(_1313_), .B(_997__bF_buf3), .Y(_294_) );
NAND2X1 NAND2X1_67 ( .A(_1030__bF_buf6), .B(_312_), .Y(_313_) );
NAND2X1 NAND2X1_68 ( .A(_1048_), .B(_1047_), .Y(_1049_) );
NAND2X1 NAND2X1_69 ( .A(_1038__bF_buf6), .B(_314_), .Y(_315_) );
NAND2X1 NAND2X1_70 ( .A(_1030__bF_buf6), .B(_319_), .Y(_320_) );
NAND2X1 NAND2X1_71 ( .A(_1045__bF_buf3), .B(_321_), .Y(_322_) );
NAND2X1 NAND2X1_72 ( .A(_1030__bF_buf0), .B(_326_), .Y(_327_) );
NAND2X1 NAND2X1_73 ( .A(_1045__bF_buf3), .B(_328_), .Y(_329_) );
NAND2X1 NAND2X1_74 ( .A(_1030__bF_buf9), .B(_333_), .Y(_334_) );
NAND2X1 NAND2X1_75 ( .A(_1038__bF_buf10), .B(_335_), .Y(_336_) );
NAND2X1 NAND2X1_76 ( .A(_1030__bF_buf0), .B(_340_), .Y(_341_) );
NAND2X1 NAND2X1_77 ( .A(_1038__bF_buf6), .B(_342_), .Y(_343_) );
NAND2X1 NAND2X1_78 ( .A(_1030__bF_buf0), .B(_347_), .Y(_348_) );
NAND2X1 NAND2X1_79 ( .A(_1051_), .B(_1050_), .Y(_1052_) );
NAND2X1 NAND2X1_80 ( .A(_1038__bF_buf6), .B(_349_), .Y(_350_) );
NAND2X1 NAND2X1_81 ( .A(PC_STACK_10__6_), .B(_1041__bF_buf4), .Y(_357_) );
NAND2X1 NAND2X1_82 ( .A(_1280_), .B(_1000__bF_buf0), .Y(_359_) );
NAND2X1 NAND2X1_83 ( .A(PC_STACK_10__7_), .B(_1041__bF_buf4), .Y(_366_) );
NAND2X1 NAND2X1_84 ( .A(_1313_), .B(_1000__bF_buf3), .Y(_367_) );
NAND2X1 NAND2X1_85 ( .A(_1030__bF_buf8), .B(_383_), .Y(_384_) );
NAND2X1 NAND2X1_86 ( .A(_1038__bF_buf3), .B(_385_), .Y(_386_) );
NAND2X1 NAND2X1_87 ( .A(_1030__bF_buf8), .B(_390_), .Y(_391_) );
NAND2X1 NAND2X1_88 ( .A(_1045__bF_buf3), .B(_392_), .Y(_393_) );
NAND2X1 NAND2X1_89 ( .A(_1030__bF_buf8), .B(_397_), .Y(_398_) );
NAND2X1 NAND2X1_90 ( .A(_1060_), .B(_1061_), .Y(_1062_) );
NAND2X1 NAND2X1_91 ( .A(_1045__bF_buf8), .B(_399_), .Y(_400_) );
NAND2X1 NAND2X1_92 ( .A(_1030__bF_buf8), .B(_404_), .Y(_405_) );
NAND2X1 NAND2X1_93 ( .A(_1038__bF_buf0), .B(_406_), .Y(_407_) );
NAND2X1 NAND2X1_94 ( .A(_1030__bF_buf0), .B(_411_), .Y(_412_) );
NAND2X1 NAND2X1_95 ( .A(_1038__bF_buf6), .B(_413_), .Y(_414_) );
NAND2X1 NAND2X1_96 ( .A(_1004__bF_buf1), .B(_1239_), .Y(_417_) );
NAND2X1 NAND2X1_97 ( .A(PC_STACK_8__5_), .B(_1041__bF_buf7), .Y(_421_) );
NAND2X1 NAND2X1_98 ( .A(_1045__bF_buf7), .B(_422_), .Y(_423_) );
NAND2X1 NAND2X1_99 ( .A(_421_), .B(_423_), .Y(_424_) );
NAND2X1 NAND2X1_100 ( .A(PC_STACK_8__6_), .B(_1041__bF_buf5), .Y(_430_) );
NAND2X1 NAND2X1_101 ( .A(_1063_), .B(_1053_), .Y(_1543__1_) );
NAND2X1 NAND2X1_102 ( .A(_1280_), .B(_1004__bF_buf1), .Y(_432_) );
NAND2X1 NAND2X1_103 ( .A(PC_STACK_8__7_), .B(_1041__bF_buf4), .Y(_439_) );
NAND2X1 NAND2X1_104 ( .A(_1313_), .B(_1004__bF_buf2), .Y(_440_) );
NAND2X1 NAND2X1_105 ( .A(_1030__bF_buf8), .B(_456_), .Y(_457_) );
NAND2X1 NAND2X1_106 ( .A(_1038__bF_buf0), .B(_458_), .Y(_459_) );
NAND2X1 NAND2X1_107 ( .A(_1030__bF_buf8), .B(_463_), .Y(_464_) );
NAND2X1 NAND2X1_108 ( .A(_1045__bF_buf7), .B(_465_), .Y(_466_) );
NAND2X1 NAND2X1_109 ( .A(_1030__bF_buf6), .B(_470_), .Y(_471_) );
NAND2X1 NAND2X1_110 ( .A(_1045__bF_buf7), .B(_472_), .Y(_473_) );
NAND2X1 NAND2X1_111 ( .A(_1030__bF_buf2), .B(_477_), .Y(_478_) );
NAND2X1 NAND2X1_112 ( .A(PC_pointer_0_), .B(_985_), .Y(_986_) );
NAND2X1 NAND2X1_113 ( .A(_1030__bF_buf3), .B(_1068_), .Y(_1069_) );
NAND2X1 NAND2X1_114 ( .A(_1038__bF_buf1), .B(_479_), .Y(_480_) );
NAND2X1 NAND2X1_115 ( .A(_1030__bF_buf0), .B(_484_), .Y(_485_) );
NAND2X1 NAND2X1_116 ( .A(_1038__bF_buf6), .B(_486_), .Y(_487_) );
NAND2X1 NAND2X1_117 ( .A(_1030__bF_buf8), .B(_491_), .Y(_492_) );
NAND2X1 NAND2X1_118 ( .A(_1038__bF_buf1), .B(_493_), .Y(_494_) );
NAND2X1 NAND2X1_119 ( .A(PC_STACK_11__6_), .B(_1041__bF_buf5), .Y(_501_) );
NAND2X1 NAND2X1_120 ( .A(_1280_), .B(_1026_), .Y(_503_) );
NAND2X1 NAND2X1_121 ( .A(PC_STACK_11__7_), .B(_1041__bF_buf4), .Y(_510_) );
NAND2X1 NAND2X1_122 ( .A(_1313_), .B(_1026_), .Y(_511_) );
NAND2X1 NAND2X1_123 ( .A(_1030__bF_buf9), .B(_529_), .Y(_530_) );
NAND2X1 NAND2X1_124 ( .A(ULA_OUT[1]), .B(_1042_), .Y(_1070_) );
NAND2X1 NAND2X1_125 ( .A(_1038__bF_buf10), .B(_531_), .Y(_532_) );
NAND2X1 NAND2X1_126 ( .A(_1030__bF_buf9), .B(_536_), .Y(_537_) );
NAND2X1 NAND2X1_127 ( .A(_1045__bF_buf1), .B(_538_), .Y(_539_) );
NAND2X1 NAND2X1_128 ( .A(_1030__bF_buf9), .B(_543_), .Y(_544_) );
NAND2X1 NAND2X1_129 ( .A(_1045__bF_buf1), .B(_545_), .Y(_546_) );
NAND2X1 NAND2X1_130 ( .A(_1030__bF_buf5), .B(_550_), .Y(_551_) );
NAND2X1 NAND2X1_131 ( .A(_1038__bF_buf10), .B(_552_), .Y(_553_) );
NAND2X1 NAND2X1_132 ( .A(_1030__bF_buf5), .B(_557_), .Y(_558_) );
NAND2X1 NAND2X1_133 ( .A(_1038__bF_buf2), .B(_559_), .Y(_560_) );
NAND2X1 NAND2X1_134 ( .A(_1030__bF_buf5), .B(_564_), .Y(_565_) );
NAND2X1 NAND2X1_135 ( .A(_1045__bF_buf9), .B(_1071_), .Y(_1072_) );
NAND2X1 NAND2X1_136 ( .A(_1038__bF_buf9), .B(_566_), .Y(_567_) );
NAND2X1 NAND2X1_137 ( .A(PC_STACK_5__6_), .B(_1041__bF_buf3), .Y(_574_) );
NAND2X1 NAND2X1_138 ( .A(_1280_), .B(_987__bF_buf1), .Y(_576_) );
NAND2X1 NAND2X1_139 ( .A(PC_STACK_5__7_), .B(_1041__bF_buf3), .Y(_583_) );
NAND2X1 NAND2X1_140 ( .A(_1313_), .B(_987__bF_buf0), .Y(_584_) );
NAND2X1 NAND2X1_141 ( .A(_1030__bF_buf4), .B(_602_), .Y(_603_) );
NAND2X1 NAND2X1_142 ( .A(_1038__bF_buf5), .B(_604_), .Y(_605_) );
NAND2X1 NAND2X1_143 ( .A(_1030__bF_buf4), .B(_609_), .Y(_610_) );
NAND2X1 NAND2X1_144 ( .A(_1045__bF_buf5), .B(_611_), .Y(_612_) );
NAND2X1 NAND2X1_145 ( .A(_1030__bF_buf1), .B(_616_), .Y(_617_) );
NAND2X1 NAND2X1_146 ( .A(_1012_), .B(_1079_), .Y(_1085_) );
NAND2X1 NAND2X1_147 ( .A(_1045__bF_buf4), .B(_618_), .Y(_619_) );
NAND2X1 NAND2X1_148 ( .A(_1030__bF_buf8), .B(_623_), .Y(_624_) );
NAND2X1 NAND2X1_149 ( .A(_1038__bF_buf3), .B(_625_), .Y(_626_) );
NAND2X1 NAND2X1_150 ( .A(_1030__bF_buf1), .B(_630_), .Y(_631_) );
NAND2X1 NAND2X1_151 ( .A(_1038__bF_buf7), .B(_632_), .Y(_633_) );
NAND2X1 NAND2X1_152 ( .A(_1030__bF_buf7), .B(_637_), .Y(_638_) );
NAND2X1 NAND2X1_153 ( .A(_1038__bF_buf5), .B(_639_), .Y(_640_) );
NAND2X1 NAND2X1_154 ( .A(PC_STACK_4__6_), .B(_1041__bF_buf8), .Y(_647_) );
NAND2X1 NAND2X1_155 ( .A(_1280_), .B(_984_), .Y(_649_) );
NAND2X1 NAND2X1_156 ( .A(PC_STACK_4__7_), .B(_1041__bF_buf3), .Y(_656_) );
NAND2X1 NAND2X1_157 ( .A(_1010_), .B(_1094_), .Y(_1099_) );
NAND2X1 NAND2X1_158 ( .A(_1313_), .B(_984_), .Y(_657_) );
NAND2X1 NAND2X1_159 ( .A(_1030__bF_buf3), .B(_674_), .Y(_675_) );
NAND2X1 NAND2X1_160 ( .A(_1038__bF_buf8), .B(_676_), .Y(_677_) );
NAND2X1 NAND2X1_161 ( .A(_1030__bF_buf3), .B(_681_), .Y(_682_) );
NAND2X1 NAND2X1_162 ( .A(_1045__bF_buf9), .B(_683_), .Y(_684_) );
NAND2X1 NAND2X1_163 ( .A(_1030__bF_buf2), .B(_688_), .Y(_689_) );
NAND2X1 NAND2X1_164 ( .A(_1045__bF_buf8), .B(_690_), .Y(_691_) );
NAND2X1 NAND2X1_165 ( .A(_1030__bF_buf3), .B(_695_), .Y(_696_) );
NAND2X1 NAND2X1_166 ( .A(_1038__bF_buf8), .B(_697_), .Y(_698_) );
NAND2X1 NAND2X1_167 ( .A(_1030__bF_buf7), .B(_702_), .Y(_703_) );
NAND2X1 NAND2X1_168 ( .A(_1094_), .B(_1079_), .Y(_1117_) );
NAND2X1 NAND2X1_169 ( .A(_1038__bF_buf4), .B(_704_), .Y(_705_) );
NAND2X1 NAND2X1_170 ( .A(_1030__bF_buf7), .B(_709_), .Y(_710_) );
NAND2X1 NAND2X1_171 ( .A(_1038__bF_buf8), .B(_711_), .Y(_712_) );
NAND2X1 NAND2X1_172 ( .A(PC_STACK_3__6_), .B(_1041__bF_buf8), .Y(_719_) );
NAND2X1 NAND2X1_173 ( .A(_1280_), .B(_1196_), .Y(_721_) );
NAND2X1 NAND2X1_174 ( .A(_715_), .B(_721_), .Y(_722_) );
NAND2X1 NAND2X1_175 ( .A(PC_STACK_3__7_), .B(_1041__bF_buf3), .Y(_728_) );
NAND2X1 NAND2X1_176 ( .A(_1313_), .B(_1196_), .Y(_729_) );
NAND2X1 NAND2X1_177 ( .A(_1030__bF_buf1), .B(_746_), .Y(_747_) );
NAND2X1 NAND2X1_178 ( .A(_1038__bF_buf8), .B(_748_), .Y(_749_) );
NAND2X1 NAND2X1_179 ( .A(_1030__bF_buf8), .B(_1143_), .Y(_1144_) );
NAND2X1 NAND2X1_180 ( .A(_1030__bF_buf1), .B(_753_), .Y(_754_) );
NAND2X1 NAND2X1_181 ( .A(_1045__bF_buf4), .B(_755_), .Y(_756_) );
NAND2X1 NAND2X1_182 ( .A(_1030__bF_buf2), .B(_760_), .Y(_761_) );
NAND2X1 NAND2X1_183 ( .A(_1045__bF_buf8), .B(_762_), .Y(_763_) );
NAND2X1 NAND2X1_184 ( .A(_1030__bF_buf1), .B(_767_), .Y(_768_) );
NAND2X1 NAND2X1_185 ( .A(_1038__bF_buf7), .B(_769_), .Y(_770_) );
NAND2X1 NAND2X1_186 ( .A(_1030__bF_buf1), .B(_774_), .Y(_775_) );
NAND2X1 NAND2X1_187 ( .A(_1038__bF_buf8), .B(_776_), .Y(_777_) );
NAND2X1 NAND2X1_188 ( .A(_1191_), .B(_1239_), .Y(_780_) );
NAND2X1 NAND2X1_189 ( .A(PC_STACK_2__5_), .B(_1041__bF_buf10), .Y(_784_) );
NAND2X1 NAND2X1_190 ( .A(ULA_OUT[2]), .B(_1042_), .Y(_1145_) );
NAND2X1 NAND2X1_191 ( .A(_1045__bF_buf9), .B(_785_), .Y(_786_) );
NAND2X1 NAND2X1_192 ( .A(_784_), .B(_786_), .Y(_787_) );
NAND2X1 NAND2X1_193 ( .A(PC_STACK_2__6_), .B(_1041__bF_buf8), .Y(_793_) );
NAND2X1 NAND2X1_194 ( .A(_1280_), .B(_1191_), .Y(_795_) );
NAND2X1 NAND2X1_195 ( .A(PC_STACK_2__7_), .B(_1041__bF_buf8), .Y(_802_) );
NAND2X1 NAND2X1_196 ( .A(_1313_), .B(_1191_), .Y(_803_) );
NAND2X1 NAND2X1_197 ( .A(_1030__bF_buf4), .B(_819_), .Y(_820_) );
NAND2X1 NAND2X1_198 ( .A(_1038__bF_buf8), .B(_821_), .Y(_822_) );
NAND2X1 NAND2X1_199 ( .A(_1030__bF_buf7), .B(_826_), .Y(_827_) );
NAND2X1 NAND2X1_200 ( .A(_1045__bF_buf5), .B(_828_), .Y(_829_) );
NAND2X1 NAND2X1_201 ( .A(_1045__bF_buf6), .B(_1146_), .Y(_1147_) );
NAND2X1 NAND2X1_202 ( .A(_1030__bF_buf4), .B(_833_), .Y(_834_) );
NAND2X1 NAND2X1_203 ( .A(_1045__bF_buf6), .B(_835_), .Y(_836_) );
NAND2X1 NAND2X1_204 ( .A(_1030__bF_buf7), .B(_840_), .Y(_841_) );
NAND2X1 NAND2X1_205 ( .A(_1038__bF_buf4), .B(_842_), .Y(_843_) );
NAND2X1 NAND2X1_206 ( .A(_1030__bF_buf7), .B(_847_), .Y(_848_) );
NAND2X1 NAND2X1_207 ( .A(_1038__bF_buf4), .B(_849_), .Y(_850_) );
NAND2X1 NAND2X1_208 ( .A(_990__bF_buf0), .B(_1239_), .Y(_853_) );
NAND2X1 NAND2X1_209 ( .A(PC_STACK_1__5_), .B(_1041__bF_buf9), .Y(_857_) );
NAND2X1 NAND2X1_210 ( .A(_1045__bF_buf9), .B(_858_), .Y(_859_) );
NAND2X1 NAND2X1_211 ( .A(_857_), .B(_859_), .Y(_860_) );
NAND2X1 NAND2X1_212 ( .A(_1168_), .B(_1176_), .Y(_1177_) );
NAND2X1 NAND2X1_213 ( .A(PC_STACK_1__6_), .B(_1041__bF_buf8), .Y(_866_) );
NAND2X1 NAND2X1_214 ( .A(_1280_), .B(_990__bF_buf1), .Y(_868_) );
NAND2X1 NAND2X1_215 ( .A(_862_), .B(_868_), .Y(_869_) );
NAND2X1 NAND2X1_216 ( .A(PC_STACK_1__7_), .B(_1041__bF_buf8), .Y(_875_) );
NAND2X1 NAND2X1_217 ( .A(_1313_), .B(_990__bF_buf3), .Y(_876_) );
NAND2X1 NAND2X1_218 ( .A(_1030__bF_buf2), .B(_892_), .Y(_893_) );
NAND2X1 NAND2X1_219 ( .A(_1038__bF_buf1), .B(_894_), .Y(_895_) );
NAND2X1 NAND2X1_220 ( .A(_1030__bF_buf2), .B(_899_), .Y(_900_) );
NAND2X1 NAND2X1_221 ( .A(_1045__bF_buf8), .B(_901_), .Y(_902_) );
NAND2X1 NAND2X1_222 ( .A(_1030__bF_buf2), .B(_906_), .Y(_907_) );
NAND2X1 NAND2X1_223 ( .A(PC_pointer_2_), .B(PC_pointer_3_), .Y(_991_) );
NAND2X1 NAND2X1_224 ( .A(_1030__bF_buf3), .B(_1183_), .Y(_1184_) );
NAND2X1 NAND2X1_225 ( .A(_1045__bF_buf8), .B(_908_), .Y(_909_) );
NAND2X1 NAND2X1_226 ( .A(_1030__bF_buf1), .B(_913_), .Y(_914_) );
NAND2X1 NAND2X1_227 ( .A(_1038__bF_buf7), .B(_915_), .Y(_916_) );
NAND2X1 NAND2X1_228 ( .A(_1030__bF_buf1), .B(_920_), .Y(_921_) );
NAND2X1 NAND2X1_229 ( .A(_1038__bF_buf7), .B(_922_), .Y(_923_) );
NAND2X1 NAND2X1_230 ( .A(_1030__bF_buf2), .B(_927_), .Y(_928_) );
NAND2X1 NAND2X1_231 ( .A(_1038__bF_buf1), .B(_929_), .Y(_930_) );
NAND2X1 NAND2X1_232 ( .A(PC_STACK_0__6_), .B(_1041__bF_buf3), .Y(_937_) );
NAND2X1 NAND2X1_233 ( .A(_1280_), .B(_1025_), .Y(_939_) );
NAND2X1 NAND2X1_234 ( .A(_933_), .B(_939_), .Y(_940_) );
NAND2X1 NAND2X1_235 ( .A(_1038__bF_buf4), .B(_1186_), .Y(_1187_) );
NAND2X1 NAND2X1_236 ( .A(PC_STACK_0__7_), .B(_1041__bF_buf8), .Y(_946_) );
NAND2X1 NAND2X1_237 ( .A(_1313_), .B(_1025_), .Y(_947_) );
NAND2X1 NAND2X1_238 ( .A(_963_), .B(_964_), .Y(_965_) );
NAND2X1 NAND2X1_239 ( .A(ULA_OUT[3]), .B(_1042_), .Y(_1188_) );
NAND2X1 NAND2X1_240 ( .A(_1030__bF_buf3), .B(_1215_), .Y(_1216_) );
NAND2X1 NAND2X1_241 ( .A(_1038__bF_buf4), .B(_1218_), .Y(_1219_) );
NAND2X1 NAND2X1_242 ( .A(ULA_OUT[4]), .B(_1042_), .Y(_1220_) );
NAND2X1 NAND2X1_243 ( .A(_1030__bF_buf3), .B(_1240_), .Y(_1241_) );
NAND2X1 NAND2X1_244 ( .A(_1038__bF_buf4), .B(_1243_), .Y(_1244_) );
NAND2X1 NAND2X1_245 ( .A(ULA_OUT[5]), .B(_1042_), .Y(_1245_) );
NAND2X1 NAND2X1_246 ( .A(_1094_), .B(_1018_), .Y(_1250_) );
NAND2X1 NAND2X1_247 ( .A(_993_), .B(_988_), .Y(_994_) );
NAND2X1 NAND2X1_248 ( .A(PC_STACK_6__6_), .B(_1041__bF_buf10), .Y(_1277_) );
NAND2X1 NAND2X1_249 ( .A(INTERRUPT_ch[6]), .B(_1102__bF_buf1), .Y(_1278_) );
NAND2X1 NAND2X1_250 ( .A(_1270_), .B(_1278_), .Y(_1279_) );
NAND2X1 NAND2X1_251 ( .A(_1280_), .B(_1102__bF_buf1), .Y(_1281_) );
NAND2X1 NAND2X1_252 ( .A(_1270_), .B(_1281_), .Y(_1282_) );
NAND2X1 NAND2X1_253 ( .A(PC_STACK_9__7_), .B(_997__bF_buf3), .Y(_1285_) );
NAND2X1 NAND2X1_254 ( .A(_1303_), .B(_1302_), .Y(_1304_) );
NAND2X1 NAND2X1_255 ( .A(INTERRUPT_ch[7]), .B(_1102__bF_buf2), .Y(_1309_) );
NAND2X1 NAND2X1_256 ( .A(PC_STACK_6__7_), .B(_1041__bF_buf8), .Y(_1312_) );
NAND2X1 NAND2X1_257 ( .A(_1313_), .B(_1102__bF_buf2), .Y(_1314_) );
NAND2X1 NAND2X1_258 ( .A(PC_pointer_3_), .B(_995_), .Y(_996_) );
NAND2X1 NAND2X1_259 ( .A(ULA_OUT[8]), .B(_1042_), .Y(_1345_) );
NAND2X1 NAND2X1_260 ( .A(_1350_), .B(_1351_), .Y(_1352_) );
NAND2X1 NAND2X1_261 ( .A(ULA_OUT[9]), .B(_1042_), .Y(_1373_) );
NAND2X1 NAND2X1_262 ( .A(_1030__bF_buf4), .B(_1377_), .Y(_1378_) );
NAND2X1 NAND2X1_263 ( .A(_1038__bF_buf3), .B(_1379_), .Y(_1380_) );
NAND2X1 NAND2X1_264 ( .A(_1030__bF_buf7), .B(_1384_), .Y(_1385_) );
NAND2X1 NAND2X1_265 ( .A(_1045__bF_buf5), .B(_1386_), .Y(_1387_) );
NAND2X1 NAND2X1_266 ( .A(_1030__bF_buf4), .B(_1391_), .Y(_1392_) );
NAND2X1 NAND2X1_267 ( .A(_1045__bF_buf6), .B(_1393_), .Y(_1394_) );
NAND2X1 NAND2X1_268 ( .A(_1030__bF_buf4), .B(_1398_), .Y(_1399_) );
NAND2X1 NAND2X1_269 ( .A(PC_pointer_1_), .B(_998_), .Y(_999_) );
NAND2X1 NAND2X1_270 ( .A(_1038__bF_buf3), .B(_1400_), .Y(_1401_) );
NAND2X1 NAND2X1_271 ( .A(_1030__bF_buf7), .B(_1405_), .Y(_1406_) );
NAND2X1 NAND2X1_272 ( .A(_1038__bF_buf5), .B(_1407_), .Y(_1408_) );
NAND2X1 NAND2X1_273 ( .A(_1030__bF_buf4), .B(_1412_), .Y(_1413_) );
NAND2X1 NAND2X1_274 ( .A(_1038__bF_buf5), .B(_1414_), .Y(_1415_) );
NAND2X1 NAND2X1_275 ( .A(PC_STACK_12__6_), .B(_1041__bF_buf8), .Y(_1422_) );
NAND2X1 NAND2X1_276 ( .A(INTERRUPT_ch[6]), .B(_992__bF_buf0), .Y(_1423_) );
NAND2X1 NAND2X1_277 ( .A(_1418_), .B(_1423_), .Y(_1424_) );
NAND2X1 NAND2X1_278 ( .A(_1280_), .B(_992__bF_buf0), .Y(_1425_) );
NAND2X1 NAND2X1_279 ( .A(_1418_), .B(_1425_), .Y(_1426_) );
NAND2X1 NAND2X1_280 ( .A(PC_pointer_0_), .B(PC_pointer_1_), .Y(_1002_) );
NAND2X1 NAND2X1_281 ( .A(INTERRUPT_ch[7]), .B(_992__bF_buf3), .Y(_1431_) );
NAND2X1 NAND2X1_282 ( .A(PC_STACK_12__7_), .B(_1041__bF_buf8), .Y(_1433_) );
NAND2X1 NAND2X1_283 ( .A(_1313_), .B(_992__bF_buf3), .Y(_1434_) );
NAND2X1 NAND2X1_284 ( .A(_1030__bF_buf8), .B(_1451_), .Y(_1452_) );
NAND2X1 NAND2X1_285 ( .A(_1038__bF_buf3), .B(_1453_), .Y(_1454_) );
NAND2X1 NAND2X1_286 ( .A(_1030__bF_buf6), .B(_1458_), .Y(_1459_) );
NAND2X1 NAND2X1_287 ( .A(_1045__bF_buf7), .B(_1460_), .Y(_1461_) );
NAND2X1 NAND2X1_288 ( .A(_1030__bF_buf6), .B(_1465_), .Y(_1466_) );
NAND2X1 NAND2X1_289 ( .A(_1045__bF_buf7), .B(_1467_), .Y(_1468_) );
NAND2X1 NAND2X1_290 ( .A(_1030__bF_buf6), .B(_1472_), .Y(_1473_) );
NAND2X1 NAND2X1_291 ( .A(_1005_), .B(_1001_), .Y(_1006_) );
NAND2X1 NAND2X1_292 ( .A(_1038__bF_buf3), .B(_1474_), .Y(_1475_) );
NAND2X1 NAND2X1_293 ( .A(_1030__bF_buf0), .B(_1479_), .Y(_1480_) );
NAND2X1 NAND2X1_294 ( .A(_1038__bF_buf6), .B(_1481_), .Y(_1482_) );
NAND2X1 NAND2X1_295 ( .A(_1030__bF_buf0), .B(_1486_), .Y(_1487_) );
NAND2X1 NAND2X1_296 ( .A(_1038__bF_buf6), .B(_1488_), .Y(_1489_) );
NAND2X1 NAND2X1_297 ( .A(PC_STACK_13__6_), .B(_1041__bF_buf0), .Y(_1496_) );
NAND2X1 NAND2X1_298 ( .A(_1280_), .B(_1022_), .Y(_1499_) );
NAND2X1 NAND2X1_299 ( .A(PC_STACK_13__7_), .B(_1041__bF_buf4), .Y(_1507_) );
NAND2X1 NAND2X1_300 ( .A(_1313_), .B(_1022_), .Y(_1508_) );
NAND2X1 NAND2X1_301 ( .A(_1030__bF_buf4), .B(_1524_), .Y(_1525_) );
NAND2X1 NAND2X1_302 ( .A(_1010_), .B(_1012_), .Y(_1013_) );
NAND2X1 NAND2X1_303 ( .A(_1038__bF_buf3), .B(_1526_), .Y(_1527_) );
NAND2X1 NAND2X1_304 ( .A(_1030__bF_buf4), .B(_1531_), .Y(_1532_) );
NAND2X1 NAND2X1_305 ( .A(_1045__bF_buf6), .B(_1533_), .Y(_1534_) );
NAND2X1 NAND2X1_306 ( .A(_1030__bF_buf9), .B(_1538_), .Y(_1539_) );
NAND2X1 NAND2X1_307 ( .A(_1045__bF_buf1), .B(_1540_), .Y(_1541_) );
NAND2X1 NAND2X1_308 ( .A(_1030__bF_buf5), .B(_21_), .Y(_22_) );
NAND2X1 NAND2X1_309 ( .A(_1038__bF_buf5), .B(_23_), .Y(_24_) );
NAND2X1 NAND2X1_310 ( .A(_1030__bF_buf1), .B(_28_), .Y(_29_) );
NAND2X1 NAND2X1_311 ( .A(_1038__bF_buf7), .B(_30_), .Y(_31_) );
NAND2X1 NAND2X1_312 ( .A(_1030__bF_buf1), .B(_35_), .Y(_36_) );
NAND3X1 NAND3X1_1 ( .A(_998_), .B(PC_pointer_1_), .C(_1010_), .Y(_1011_) );
NAND3X1 NAND3X1_2 ( .A(_998_), .B(PC_pointer_1_), .C(_1079_), .Y(_1109_) );
NAND3X1 NAND3X1_3 ( .A(_532_), .B(_534_), .C(_530_), .Y(_11__0_) );
NAND3X1 NAND3X1_4 ( .A(_539_), .B(_541_), .C(_537_), .Y(_11__1_) );
NAND3X1 NAND3X1_5 ( .A(_546_), .B(_548_), .C(_544_), .Y(_11__2_) );
NAND3X1 NAND3X1_6 ( .A(_553_), .B(_555_), .C(_551_), .Y(_11__3_) );
NAND3X1 NAND3X1_7 ( .A(_560_), .B(_562_), .C(_558_), .Y(_11__4_) );
NAND3X1 NAND3X1_8 ( .A(_567_), .B(_569_), .C(_565_), .Y(_11__5_) );
NAND3X1 NAND3X1_9 ( .A(_574_), .B(_578_), .C(_573_), .Y(_11__6_) );
NAND3X1 NAND3X1_10 ( .A(_605_), .B(_607_), .C(_603_), .Y(_10__0_) );
NAND3X1 NAND3X1_11 ( .A(_612_), .B(_614_), .C(_610_), .Y(_10__1_) );
NAND3X1 NAND3X1_12 ( .A(_619_), .B(_621_), .C(_617_), .Y(_10__2_) );
NAND3X1 NAND3X1_13 ( .A(_988_), .B(_1001_), .C(_1111_), .Y(_1112_) );
NAND3X1 NAND3X1_14 ( .A(_626_), .B(_628_), .C(_624_), .Y(_10__3_) );
NAND3X1 NAND3X1_15 ( .A(_633_), .B(_635_), .C(_631_), .Y(_10__4_) );
NAND3X1 NAND3X1_16 ( .A(_640_), .B(_642_), .C(_638_), .Y(_10__5_) );
NAND3X1 NAND3X1_17 ( .A(_647_), .B(_651_), .C(_646_), .Y(_10__6_) );
NAND3X1 NAND3X1_18 ( .A(_677_), .B(_679_), .C(_675_), .Y(_9__0_) );
NAND3X1 NAND3X1_19 ( .A(_684_), .B(_686_), .C(_682_), .Y(_9__1_) );
NAND3X1 NAND3X1_20 ( .A(_691_), .B(_693_), .C(_689_), .Y(_9__2_) );
NAND3X1 NAND3X1_21 ( .A(_698_), .B(_700_), .C(_696_), .Y(_9__3_) );
NAND3X1 NAND3X1_22 ( .A(_705_), .B(_707_), .C(_703_), .Y(_9__4_) );
NAND3X1 NAND3X1_23 ( .A(_712_), .B(_714_), .C(_710_), .Y(_9__5_) );
NAND3X1 NAND3X1_24 ( .A(PC_pointer_0_), .B(_985_), .C(_1010_), .Y(_1116_) );
NAND3X1 NAND3X1_25 ( .A(_719_), .B(_723_), .C(_718_), .Y(_9__6_) );
NAND3X1 NAND3X1_26 ( .A(_749_), .B(_751_), .C(_747_), .Y(_8__0_) );
NAND3X1 NAND3X1_27 ( .A(_756_), .B(_758_), .C(_754_), .Y(_8__1_) );
NAND3X1 NAND3X1_28 ( .A(_763_), .B(_765_), .C(_761_), .Y(_8__2_) );
NAND3X1 NAND3X1_29 ( .A(_770_), .B(_772_), .C(_768_), .Y(_8__3_) );
NAND3X1 NAND3X1_30 ( .A(_777_), .B(_779_), .C(_775_), .Y(_8__4_) );
NAND3X1 NAND3X1_31 ( .A(_793_), .B(_797_), .C(_792_), .Y(_8__6_) );
NAND3X1 NAND3X1_32 ( .A(_822_), .B(_824_), .C(_820_), .Y(_7__0_) );
NAND3X1 NAND3X1_33 ( .A(_829_), .B(_831_), .C(_827_), .Y(_7__1_) );
NAND3X1 NAND3X1_34 ( .A(_836_), .B(_838_), .C(_834_), .Y(_7__2_) );
NAND3X1 NAND3X1_35 ( .A(_1113_), .B(_1027_), .C(_1122_), .Y(_1123_) );
NAND3X1 NAND3X1_36 ( .A(_843_), .B(_845_), .C(_841_), .Y(_7__3_) );
NAND3X1 NAND3X1_37 ( .A(_850_), .B(_852_), .C(_848_), .Y(_7__4_) );
NAND3X1 NAND3X1_38 ( .A(_866_), .B(_870_), .C(_865_), .Y(_7__6_) );
NAND3X1 NAND3X1_39 ( .A(_895_), .B(_897_), .C(_893_), .Y(_0__0_) );
NAND3X1 NAND3X1_40 ( .A(_902_), .B(_904_), .C(_900_), .Y(_0__1_) );
NAND3X1 NAND3X1_41 ( .A(_909_), .B(_911_), .C(_907_), .Y(_0__2_) );
NAND3X1 NAND3X1_42 ( .A(_916_), .B(_918_), .C(_914_), .Y(_0__3_) );
NAND3X1 NAND3X1_43 ( .A(_923_), .B(_925_), .C(_921_), .Y(_0__4_) );
NAND3X1 NAND3X1_44 ( .A(_930_), .B(_932_), .C(_928_), .Y(_0__5_) );
NAND3X1 NAND3X1_45 ( .A(_937_), .B(_941_), .C(_936_), .Y(_0__6_) );
NAND3X1 NAND3X1_46 ( .A(_1047_), .B(_1050_), .C(_1127_), .Y(_1128_) );
NAND3X1 NAND3X1_47 ( .A(_1129_), .B(_1061_), .C(_1136_), .Y(_1137_) );
NAND3X1 NAND3X1_48 ( .A(_1147_), .B(_1150_), .C(_1144_), .Y(_12__2_) );
NAND3X1 NAND3X1_49 ( .A(_1158_), .B(_1159_), .C(_1157_), .Y(_1160_) );
NAND3X1 NAND3X1_50 ( .A(PC_STACK_10__3_), .B(_1017_), .C(_1170_), .Y(_1171_) );
NAND3X1 NAND3X1_51 ( .A(_1187_), .B(_1190_), .C(_1184_), .Y(_12__3_) );
NAND3X1 NAND3X1_52 ( .A(PC_pointer_2_), .B(_981_), .C(_1012_), .Y(_1020_) );
NAND3X1 NAND3X1_53 ( .A(_1195_), .B(_1197_), .C(_1194_), .Y(_1198_) );
NAND3X1 NAND3X1_54 ( .A(_1207_), .B(_1208_), .C(_1206_), .Y(_1209_) );
NAND3X1 NAND3X1_55 ( .A(_1543__2_), .B(_1543__3_), .C(_1065_), .Y(_1211_) );
NAND3X1 NAND3X1_56 ( .A(_1219_), .B(_1222_), .C(_1216_), .Y(_12__4_) );
NAND3X1 NAND3X1_57 ( .A(_1223_), .B(_1224_), .C(_1227_), .Y(_1228_) );
NAND3X1 NAND3X1_58 ( .A(_1232_), .B(_1233_), .C(_1231_), .Y(_1234_) );
NAND3X1 NAND3X1_59 ( .A(_1543__4_), .B(_1543__5_), .C(_1180_), .Y(_1237_) );
NAND3X1 NAND3X1_60 ( .A(_1042_), .B(_1237_), .C(_1238_), .Y(_1239_) );
NAND3X1 NAND3X1_61 ( .A(_1244_), .B(_1247_), .C(_1241_), .Y(_12__5_) );
NAND3X1 NAND3X1_62 ( .A(_1256_), .B(_1257_), .C(_1255_), .Y(_1258_) );
NAND3X1 NAND3X1_63 ( .A(_1039_), .B(_1046_), .C(_1034_), .Y(_12__0_) );
NAND3X1 NAND3X1_64 ( .A(_1266_), .B(_1267_), .C(_1265_), .Y(_1268_) );
NAND3X1 NAND3X1_65 ( .A(_1277_), .B(_1283_), .C(_1276_), .Y(_12__6_) );
NAND3X1 NAND3X1_66 ( .A(_1291_), .B(_1292_), .C(_1290_), .Y(_1293_) );
NAND3X1 NAND3X1_67 ( .A(_1294_), .B(_1295_), .C(_1298_), .Y(_1299_) );
NAND3X1 NAND3X1_68 ( .A(_1543__6_), .B(_1543__7_), .C(_1272_), .Y(_1302_) );
NAND3X1 NAND3X1_69 ( .A(_1318_), .B(_1319_), .C(_1326_), .Y(_1327_) );
NAND3X1 NAND3X1_70 ( .A(_1331_), .B(_1336_), .C(_1335_), .Y(_1337_) );
NAND3X1 NAND3X1_71 ( .A(_1543__8_), .B(_1366_), .C(_1341_), .Y(_1367_) );
NAND3X1 NAND3X1_72 ( .A(_1380_), .B(_1382_), .C(_1378_), .Y(_3__0_) );
NAND3X1 NAND3X1_73 ( .A(_1387_), .B(_1389_), .C(_1385_), .Y(_3__1_) );
NAND3X1 NAND3X1_74 ( .A(_1072_), .B(_1075_), .C(_1069_), .Y(_12__1_) );
NAND3X1 NAND3X1_75 ( .A(_1394_), .B(_1396_), .C(_1392_), .Y(_3__2_) );
NAND3X1 NAND3X1_76 ( .A(_1401_), .B(_1403_), .C(_1399_), .Y(_3__3_) );
NAND3X1 NAND3X1_77 ( .A(_1408_), .B(_1410_), .C(_1406_), .Y(_3__4_) );
NAND3X1 NAND3X1_78 ( .A(_1415_), .B(_1417_), .C(_1413_), .Y(_3__5_) );
NAND3X1 NAND3X1_79 ( .A(_1422_), .B(_1427_), .C(_1421_), .Y(_3__6_) );
NAND3X1 NAND3X1_80 ( .A(_1454_), .B(_1456_), .C(_1452_), .Y(_4__0_) );
NAND3X1 NAND3X1_81 ( .A(_1461_), .B(_1463_), .C(_1459_), .Y(_4__1_) );
NAND3X1 NAND3X1_82 ( .A(_1468_), .B(_1470_), .C(_1466_), .Y(_4__2_) );
NAND3X1 NAND3X1_83 ( .A(_1475_), .B(_1477_), .C(_1473_), .Y(_4__3_) );
NAND3X1 NAND3X1_84 ( .A(_1482_), .B(_1484_), .C(_1480_), .Y(_4__4_) );
NAND3X1 NAND3X1_85 ( .A(PC_pointer_0_), .B(_985_), .C(_1079_), .Y(_1080_) );
NAND3X1 NAND3X1_86 ( .A(_1489_), .B(_1491_), .C(_1487_), .Y(_4__5_) );
NAND3X1 NAND3X1_87 ( .A(_1496_), .B(_1501_), .C(_1495_), .Y(_4__6_) );
NAND3X1 NAND3X1_88 ( .A(_1527_), .B(_1529_), .C(_1525_), .Y(_5__0_) );
NAND3X1 NAND3X1_89 ( .A(_1534_), .B(_1536_), .C(_1532_), .Y(_5__1_) );
NAND3X1 NAND3X1_90 ( .A(_1541_), .B(_19_), .C(_1539_), .Y(_5__2_) );
NAND3X1 NAND3X1_91 ( .A(_24_), .B(_26_), .C(_22_), .Y(_5__3_) );
NAND3X1 NAND3X1_92 ( .A(_31_), .B(_33_), .C(_29_), .Y(_5__4_) );
NAND3X1 NAND3X1_93 ( .A(_38_), .B(_40_), .C(_36_), .Y(_5__5_) );
NAND3X1 NAND3X1_94 ( .A(_45_), .B(_49_), .C(_44_), .Y(_5__6_) );
NAND3X1 NAND3X1_95 ( .A(_81_), .B(_82_), .C(_73_), .Y(_83_) );
NAND3X1 NAND3X1_96 ( .A(_995_), .B(PC_pointer_3_), .C(_1012_), .Y(_1084_) );
NAND3X1 NAND3X1_97 ( .A(_97_), .B(_99_), .C(_95_), .Y(_13__0_) );
NAND3X1 NAND3X1_98 ( .A(_104_), .B(_106_), .C(_102_), .Y(_13__1_) );
NAND3X1 NAND3X1_99 ( .A(_111_), .B(_113_), .C(_109_), .Y(_13__2_) );
NAND3X1 NAND3X1_100 ( .A(_118_), .B(_120_), .C(_116_), .Y(_13__3_) );
NAND3X1 NAND3X1_101 ( .A(_125_), .B(_127_), .C(_123_), .Y(_13__4_) );
NAND3X1 NAND3X1_102 ( .A(_141_), .B(_145_), .C(_140_), .Y(_13__6_) );
NAND3X1 NAND3X1_103 ( .A(_170_), .B(_172_), .C(_168_), .Y(_6__0_) );
NAND3X1 NAND3X1_104 ( .A(_177_), .B(_179_), .C(_175_), .Y(_6__1_) );
NAND3X1 NAND3X1_105 ( .A(_184_), .B(_186_), .C(_182_), .Y(_6__2_) );
NAND3X1 NAND3X1_106 ( .A(_191_), .B(_193_), .C(_189_), .Y(_6__3_) );
NAND3X1 NAND3X1_107 ( .A(_1088_), .B(_1089_), .C(_1087_), .Y(_1090_) );
NAND3X1 NAND3X1_108 ( .A(_198_), .B(_200_), .C(_196_), .Y(_6__4_) );
NAND3X1 NAND3X1_109 ( .A(_205_), .B(_207_), .C(_203_), .Y(_6__5_) );
NAND3X1 NAND3X1_110 ( .A(_212_), .B(_216_), .C(_211_), .Y(_6__6_) );
NAND3X1 NAND3X1_111 ( .A(_242_), .B(_244_), .C(_240_), .Y(_15__0_) );
NAND3X1 NAND3X1_112 ( .A(_249_), .B(_251_), .C(_247_), .Y(_15__1_) );
NAND3X1 NAND3X1_113 ( .A(_256_), .B(_258_), .C(_254_), .Y(_15__2_) );
NAND3X1 NAND3X1_114 ( .A(_263_), .B(_265_), .C(_261_), .Y(_15__3_) );
NAND3X1 NAND3X1_115 ( .A(_270_), .B(_272_), .C(_268_), .Y(_15__4_) );
NAND3X1 NAND3X1_116 ( .A(_277_), .B(_279_), .C(_275_), .Y(_15__5_) );
NAND3X1 NAND3X1_117 ( .A(_284_), .B(_288_), .C(_283_), .Y(_15__6_) );
NAND3X1 NAND3X1_118 ( .A(_995_), .B(PC_pointer_3_), .C(_1094_), .Y(_1095_) );
NAND3X1 NAND3X1_119 ( .A(_315_), .B(_317_), .C(_313_), .Y(_1__0_) );
NAND3X1 NAND3X1_120 ( .A(_322_), .B(_324_), .C(_320_), .Y(_1__1_) );
NAND3X1 NAND3X1_121 ( .A(_329_), .B(_331_), .C(_327_), .Y(_1__2_) );
NAND3X1 NAND3X1_122 ( .A(_336_), .B(_338_), .C(_334_), .Y(_1__3_) );
NAND3X1 NAND3X1_123 ( .A(_343_), .B(_345_), .C(_341_), .Y(_1__4_) );
NAND3X1 NAND3X1_124 ( .A(_350_), .B(_352_), .C(_348_), .Y(_1__5_) );
NAND3X1 NAND3X1_125 ( .A(_357_), .B(_361_), .C(_356_), .Y(_1__6_) );
NAND3X1 NAND3X1_126 ( .A(_386_), .B(_388_), .C(_384_), .Y(_14__0_) );
NAND3X1 NAND3X1_127 ( .A(_393_), .B(_395_), .C(_391_), .Y(_14__1_) );
NAND3X1 NAND3X1_128 ( .A(_400_), .B(_402_), .C(_398_), .Y(_14__2_) );
NAND3X1 NAND3X1_129 ( .A(_1103_), .B(_1105_), .C(_1101_), .Y(_1106_) );
NAND3X1 NAND3X1_130 ( .A(_407_), .B(_409_), .C(_405_), .Y(_14__3_) );
NAND3X1 NAND3X1_131 ( .A(_414_), .B(_416_), .C(_412_), .Y(_14__4_) );
NAND3X1 NAND3X1_132 ( .A(_430_), .B(_434_), .C(_429_), .Y(_14__6_) );
NAND3X1 NAND3X1_133 ( .A(_459_), .B(_461_), .C(_457_), .Y(_2__0_) );
NAND3X1 NAND3X1_134 ( .A(_466_), .B(_468_), .C(_464_), .Y(_2__1_) );
NAND3X1 NAND3X1_135 ( .A(_473_), .B(_475_), .C(_471_), .Y(_2__2_) );
NAND3X1 NAND3X1_136 ( .A(_480_), .B(_482_), .C(_478_), .Y(_2__3_) );
NAND3X1 NAND3X1_137 ( .A(_487_), .B(_489_), .C(_485_), .Y(_2__4_) );
NAND3X1 NAND3X1_138 ( .A(_494_), .B(_496_), .C(_492_), .Y(_2__5_) );
NAND3X1 NAND3X1_139 ( .A(_501_), .B(_505_), .C(_500_), .Y(_2__6_) );
NOR2X1 NOR2X1_1 ( .A(_983__bF_buf0), .B(_982__bF_buf2), .Y(_984_) );
NOR2X1 NOR2X1_2 ( .A(PC_pointer_2_), .B(PC_pointer_3_), .Y(_1010_) );
NOR2X1 NOR2X1_3 ( .A(PC_pointer_0_), .B(_985_), .Y(_1017_) );
NOR2X1 NOR2X1_4 ( .A(PC_pointer_3_), .B(_995_), .Y(_1018_) );
NOR2X1 NOR2X1_5 ( .A(_989__bF_buf3), .B(_983__bF_buf5), .Y(_1025_) );
NOR2X1 NOR2X1_6 ( .A(CORE_PC_ctrl[0]), .B(INTERRUPT_flag), .Y(_1030_) );
NOR2X1 NOR2X1_7 ( .A(CORE_PC_ctrl[0]), .B(_1037_), .Y(_1038_) );
NOR2X1 NOR2X1_8 ( .A(_1040_), .B(_1037_), .Y(_1041_) );
NOR2X1 NOR2X1_9 ( .A(INTERRUPT_flag), .B(_1040_), .Y(_1045_) );
NOR2X1 NOR2X1_10 ( .A(_1049_), .B(_1052_), .Y(_1053_) );
NOR2X1 NOR2X1_11 ( .A(_1086_), .B(_1081_), .Y(_1087_) );
NOR2X1 NOR2X1_12 ( .A(_986__bF_buf3), .B(_982__bF_buf2), .Y(_987_) );
NOR2X1 NOR2X1_13 ( .A(PC_pointer_0_), .B(PC_pointer_1_), .Y(_1094_) );
NOR2X1 NOR2X1_14 ( .A(_1093_), .B(_1095__bF_buf2), .Y(_1096_) );
NOR2X1 NOR2X1_15 ( .A(_999__bF_buf2), .B(_982__bF_buf1), .Y(_1102_) );
NOR2X1 NOR2X1_16 ( .A(_1014_), .B(_1110_), .Y(_1111_) );
NOR2X1 NOR2X1_17 ( .A(_1118_), .B(_1121_), .Y(_1122_) );
NOR2X1 NOR2X1_18 ( .A(_1056_), .B(_1126_), .Y(_1127_) );
NOR2X1 NOR2X1_19 ( .A(_1132_), .B(_1135_), .Y(_1136_) );
NOR2X1 NOR2X1_20 ( .A(_1090_), .B(_1106_), .Y(_1139_) );
NOR2X1 NOR2X1_21 ( .A(_1139_), .B(_1138_), .Y(_1140_) );
NOR2X1 NOR2X1_22 ( .A(rst_bF_buf2), .B(_1140_), .Y(_1141_) );
NOR2X1 NOR2X1_23 ( .A(_989__bF_buf4), .B(_986__bF_buf3), .Y(_990_) );
NOR2X1 NOR2X1_24 ( .A(_1153_), .B(_1156_), .Y(_1157_) );
NOR2X1 NOR2X1_25 ( .A(_1164_), .B(_1099__bF_buf4), .Y(_1165_) );
NOR2X1 NOR2X1_26 ( .A(PC_pointer_2_), .B(_981_), .Y(_1170_) );
NOR2X1 NOR2X1_27 ( .A(_1175_), .B(_1172_), .Y(_1176_) );
NOR2X1 NOR2X1_28 ( .A(_1160_), .B(_1177_), .Y(_1179_) );
NOR2X1 NOR2X1_29 ( .A(_1002__bF_buf5), .B(_989__bF_buf5), .Y(_1196_) );
NOR2X1 NOR2X1_30 ( .A(_1205_), .B(_1202_), .Y(_1206_) );
NOR2X1 NOR2X1_31 ( .A(_1198_), .B(_1209_), .Y(_1212_) );
NOR2X1 NOR2X1_32 ( .A(_1228_), .B(_1234_), .Y(_1235_) );
NOR2X1 NOR2X1_33 ( .A(_1254_), .B(_1251_), .Y(_1255_) );
NOR2X1 NOR2X1_34 ( .A(_991__bF_buf6), .B(_983__bF_buf0), .Y(_992_) );
NOR2X1 NOR2X1_35 ( .A(_1264_), .B(_1261_), .Y(_1265_) );
NOR2X1 NOR2X1_36 ( .A(_1258_), .B(_1268_), .Y(_1269_) );
NOR2X1 NOR2X1_37 ( .A(_1289_), .B(_1286_), .Y(_1290_) );
NOR2X1 NOR2X1_38 ( .A(_1299_), .B(_1293_), .Y(_1300_) );
NOR2X1 NOR2X1_39 ( .A(_1310_), .B(_1316_), .Y(_1317_) );
NOR2X1 NOR2X1_40 ( .A(_1325_), .B(_1322_), .Y(_1326_) );
NOR2X1 NOR2X1_41 ( .A(_1327_), .B(_1337_), .Y(_1338_) );
NOR2X1 NOR2X1_42 ( .A(_1432_), .B(_1436_), .Y(_1437_) );
NOR2X1 NOR2X1_43 ( .A(_71_), .B(_74_), .Y(_75_) );
NOR2X1 NOR2X1_44 ( .A(_75_), .B(_73_), .Y(_76_) );
NOR2X1 NOR2X1_45 ( .A(_986__bF_buf4), .B(_996__bF_buf2), .Y(_997_) );
NOR2X1 NOR2X1_46 ( .A(PC_pointer_2_), .B(_983__bF_buf4), .Y(_84_) );
NOR2X1 NOR2X1_47 ( .A(_995_), .B(_1094_), .Y(_85_) );
NOR2X1 NOR2X1_48 ( .A(CORE_PC_ctrl[0]), .B(delay), .Y(_964_) );
NOR2X1 NOR2X1_49 ( .A(_962_), .B(_965_), .Y(_1544_) );
NOR2X1 NOR2X1_50 ( .A(_966_), .B(_965_), .Y(_1542__0_) );
NOR2X1 NOR2X1_51 ( .A(_967_), .B(_965_), .Y(_1542__1_) );
NOR2X1 NOR2X1_52 ( .A(_968_), .B(_965_), .Y(_1542__2_) );
NOR2X1 NOR2X1_53 ( .A(_969_), .B(_965_), .Y(_1542__3_) );
NOR2X1 NOR2X1_54 ( .A(_970_), .B(_965_), .Y(_1542__4_) );
NOR2X1 NOR2X1_55 ( .A(_971_), .B(_965_), .Y(_1542__5_) );
NOR2X1 NOR2X1_56 ( .A(_999__bF_buf4), .B(_996__bF_buf2), .Y(_1000_) );
NOR2X1 NOR2X1_57 ( .A(_972_), .B(_965_), .Y(_1542__6_) );
NOR2X1 NOR2X1_58 ( .A(_973_), .B(_965_), .Y(_1542__7_) );
NOR2X1 NOR2X1_59 ( .A(_974_), .B(_965_), .Y(_1542__8_) );
NOR2X1 NOR2X1_60 ( .A(_975_), .B(_965_), .Y(_1542__9_) );
NOR2X1 NOR2X1_61 ( .A(_976_), .B(_965_), .Y(_1542__10_) );
NOR2X1 NOR2X1_62 ( .A(_977_), .B(_965_), .Y(_1542__11_) );
NOR2X1 NOR2X1_63 ( .A(_978_), .B(_965_), .Y(_1542__12_) );
NOR2X1 NOR2X1_64 ( .A(_979_), .B(_965_), .Y(_1542__13_) );
NOR2X1 NOR2X1_65 ( .A(_980_), .B(_965_), .Y(_1542__14_) );
NOR2X1 NOR2X1_66 ( .A(_1002__bF_buf1), .B(_991__bF_buf5), .Y(_1003_) );
NOR2X1 NOR2X1_67 ( .A(_983__bF_buf2), .B(_996__bF_buf0), .Y(_1004_) );
NOR2X1 NOR2X1_68 ( .A(_994_), .B(_1006_), .Y(_1007_) );
NOR3X1 NOR3X1_1 ( .A(_998_), .B(PC_pointer_1_), .C(_991__bF_buf1), .Y(_1022_) );
NOR3X1 NOR3X1_2 ( .A(_1139_), .B(_1179_), .C(_1138_), .Y(_1180_) );
NOR3X1 NOR3X1_3 ( .A(_1212_), .B(_1235_), .C(_1211_), .Y(_1272_) );
NOR3X1 NOR3X1_4 ( .A(_1269_), .B(_1300_), .C(_1237_), .Y(_1341_) );
NOR3X1 NOR3X1_5 ( .A(_1354_), .B(_1357_), .C(_1352_), .Y(_1358_) );
NOR3X1 NOR3X1_6 ( .A(PC_pointer_0_), .B(_985_), .C(_991__bF_buf1), .Y(_1023_) );
NOR3X1 NOR3X1_7 ( .A(PC_pointer_2_), .B(_981_), .C(_1002__bF_buf1), .Y(_1026_) );
NOR3X1 NOR3X1_8 ( .A(_1014_), .B(_1021_), .C(_1028_), .Y(_1029_) );
NOR3X1 NOR3X1_9 ( .A(_1056_), .B(_1059_), .C(_1062_), .Y(_1063_) );
NOR3X1 NOR3X1_10 ( .A(_1091_), .B(_991__bF_buf1), .C(_999__bF_buf1), .Y(_1092_) );
NOR3X1 NOR3X1_11 ( .A(_1096_), .B(_1092_), .C(_1100_), .Y(_1101_) );
NOR3X1 NOR3X1_12 ( .A(_999__bF_buf5), .B(_1166_), .C(_982__bF_buf0), .Y(_1167_) );
NOR3X1 NOR3X1_13 ( .A(_1165_), .B(_1167_), .C(_1163_), .Y(_1168_) );
OAI21X1 OAI21X1_1 ( .A(_999__bF_buf3), .B(_982__bF_buf5), .C(PC_STACK_6__0_), .Y(_1031_) );
OAI21X1 OAI21X1_2 ( .A(_999__bF_buf1), .B(_982__bF_buf6), .C(PC_STACK_6__2_), .Y(_1076_) );
OAI21X1 OAI21X1_3 ( .A(_986__bF_buf5), .B(_991__bF_buf2), .C(PC_STACK_13__2_), .Y(_1464_) );
OAI21X1 OAI21X1_4 ( .A(_1142_), .B(_1080__bF_buf1), .C(_1464_), .Y(_1465_) );
OAI21X1 OAI21X1_5 ( .A(_1080__bF_buf1), .B(_1145_), .C(_1464_), .Y(_1467_) );
OAI21X1 OAI21X1_6 ( .A(_1148_), .B(_1080__bF_buf1), .C(_1464_), .Y(_1469_) );
OAI21X1 OAI21X1_7 ( .A(_986__bF_buf4), .B(_991__bF_buf4), .C(PC_STACK_13__3_), .Y(_1471_) );
OAI21X1 OAI21X1_8 ( .A(_1182_), .B(_1080__bF_buf3), .C(_1471_), .Y(_1472_) );
OAI21X1 OAI21X1_9 ( .A(_1185_), .B(_1080__bF_buf3), .C(_1471_), .Y(_1474_) );
OAI21X1 OAI21X1_10 ( .A(_1080__bF_buf3), .B(_1188_), .C(_1471_), .Y(_1476_) );
OAI21X1 OAI21X1_11 ( .A(_986__bF_buf5), .B(_991__bF_buf4), .C(PC_STACK_13__4_), .Y(_1478_) );
OAI21X1 OAI21X1_12 ( .A(_1214_), .B(_1080__bF_buf0), .C(_1478_), .Y(_1479_) );
OAI21X1 OAI21X1_13 ( .A(_1065_), .B(_1543__2_), .C(_1141_), .Y(_1142_) );
OAI21X1 OAI21X1_14 ( .A(_1217_), .B(_1080__bF_buf0), .C(_1478_), .Y(_1481_) );
OAI21X1 OAI21X1_15 ( .A(_1080__bF_buf0), .B(_1220_), .C(_1478_), .Y(_1483_) );
OAI21X1 OAI21X1_16 ( .A(_986__bF_buf4), .B(_991__bF_buf4), .C(PC_STACK_13__5_), .Y(_1485_) );
OAI21X1 OAI21X1_17 ( .A(_1239_), .B(_1080__bF_buf0), .C(_1485_), .Y(_1486_) );
OAI21X1 OAI21X1_18 ( .A(_1242_), .B(_1080__bF_buf0), .C(_1485_), .Y(_1488_) );
OAI21X1 OAI21X1_19 ( .A(_1080__bF_buf3), .B(_1245_), .C(_1485_), .Y(_1490_) );
OAI21X1 OAI21X1_20 ( .A(_986__bF_buf4), .B(_991__bF_buf4), .C(PC_STACK_13__6_), .Y(_1492_) );
OAI21X1 OAI21X1_21 ( .A(_1494_), .B(_1493_), .C(_1030__bF_buf9), .Y(_1495_) );
OAI21X1 OAI21X1_22 ( .A(_1497_), .B(_1080__bF_buf4), .C(_1492_), .Y(_1498_) );
OAI21X1 OAI21X1_23 ( .A(_1263_), .B(_1022_), .C(_1499_), .Y(_1500_) );
OAI21X1 OAI21X1_24 ( .A(_1142_), .B(_1019__bF_buf2), .C(_1076_), .Y(_1143_) );
OAI21X1 OAI21X1_25 ( .A(_1304_), .B(rst_bF_buf2), .C(_1022_), .Y(_1502_) );
OAI21X1 OAI21X1_26 ( .A(PC_STACK_13__7_), .B(_1022_), .C(_1502_), .Y(_1503_) );
OAI21X1 OAI21X1_27 ( .A(_986__bF_buf0), .B(_991__bF_buf3), .C(PC_STACK_13__7_), .Y(_1505_) );
OAI21X1 OAI21X1_28 ( .A(_1504_), .B(_1080__bF_buf4), .C(_1505_), .Y(_1506_) );
OAI21X1 OAI21X1_29 ( .A(_1509_), .B(_1311__bF_buf3), .C(_1507_), .Y(_1510_) );
OAI21X1 OAI21X1_30 ( .A(_1503_), .B(_1301__bF_buf4), .C(_1511_), .Y(_4__7_) );
OAI21X1 OAI21X1_31 ( .A(_986__bF_buf0), .B(_991__bF_buf3), .C(_1320_), .Y(_1512_) );
OAI21X1 OAI21X1_32 ( .A(_1343_), .B(_1080__bF_buf4), .C(_1512_), .Y(_1513_) );
OAI21X1 OAI21X1_33 ( .A(_986__bF_buf0), .B(_991__bF_buf4), .C(PC_STACK_13__8_), .Y(_1514_) );
OAI21X1 OAI21X1_34 ( .A(_1080__bF_buf4), .B(_1345_), .C(_1514_), .Y(_1515_) );
OAI21X1 OAI21X1_35 ( .A(_1019__bF_buf2), .B(_1145_), .C(_1076_), .Y(_1146_) );
OAI21X1 OAI21X1_36 ( .A(_1513_), .B(_1301__bF_buf1), .C(_1517_), .Y(_4__8_) );
OAI21X1 OAI21X1_37 ( .A(_986__bF_buf4), .B(_991__bF_buf5), .C(_1355_), .Y(_1518_) );
OAI21X1 OAI21X1_38 ( .A(_1369_), .B(_1080__bF_buf2), .C(_1518_), .Y(_1519_) );
OAI21X1 OAI21X1_39 ( .A(_986__bF_buf0), .B(_991__bF_buf4), .C(PC_STACK_13__9_), .Y(_1520_) );
OAI21X1 OAI21X1_40 ( .A(_1080__bF_buf4), .B(_1373_), .C(_1520_), .Y(_1521_) );
OAI21X1 OAI21X1_41 ( .A(_1519_), .B(_1301__bF_buf1), .C(_1522_), .Y(_4__9_) );
OAI21X1 OAI21X1_42 ( .A(_999__bF_buf1), .B(_991__bF_buf5), .C(PC_STACK_14__0_), .Y(_1523_) );
OAI21X1 OAI21X1_43 ( .A(_1032_), .B(_1109__bF_buf3), .C(_1523_), .Y(_1524_) );
OAI21X1 OAI21X1_44 ( .A(_1035_), .B(_1109__bF_buf3), .C(_1523_), .Y(_1526_) );
OAI21X1 OAI21X1_45 ( .A(_1109__bF_buf3), .B(_1043_), .C(_1523_), .Y(_1528_) );
OAI21X1 OAI21X1_46 ( .A(_1019__bF_buf2), .B(_1148_), .C(_1076_), .Y(_1149_) );
OAI21X1 OAI21X1_47 ( .A(_999__bF_buf1), .B(_991__bF_buf5), .C(PC_STACK_14__1_), .Y(_1530_) );
OAI21X1 OAI21X1_48 ( .A(_1067_), .B(_1109__bF_buf1), .C(_1530_), .Y(_1531_) );
OAI21X1 OAI21X1_49 ( .A(_1109__bF_buf1), .B(_1070_), .C(_1530_), .Y(_1533_) );
OAI21X1 OAI21X1_50 ( .A(_1073_), .B(_1109__bF_buf3), .C(_1530_), .Y(_1535_) );
OAI21X1 OAI21X1_51 ( .A(_999__bF_buf1), .B(_991__bF_buf3), .C(PC_STACK_14__2_), .Y(_1537_) );
OAI21X1 OAI21X1_52 ( .A(_1142_), .B(_1109__bF_buf4), .C(_1537_), .Y(_1538_) );
OAI21X1 OAI21X1_53 ( .A(_1109__bF_buf4), .B(_1145_), .C(_1537_), .Y(_1540_) );
OAI21X1 OAI21X1_54 ( .A(_1148_), .B(_1109__bF_buf4), .C(_1537_), .Y(_18_) );
OAI21X1 OAI21X1_55 ( .A(_999__bF_buf0), .B(_991__bF_buf6), .C(PC_STACK_14__3_), .Y(_20_) );
OAI21X1 OAI21X1_56 ( .A(_1182_), .B(_1109__bF_buf1), .C(_20_), .Y(_21_) );
OAI21X1 OAI21X1_57 ( .A(_1169_), .B(_1013__bF_buf2), .C(_1171_), .Y(_1172_) );
OAI21X1 OAI21X1_58 ( .A(_1185_), .B(_1109__bF_buf1), .C(_20_), .Y(_23_) );
OAI21X1 OAI21X1_59 ( .A(_1109__bF_buf1), .B(_1188_), .C(_20_), .Y(_25_) );
OAI21X1 OAI21X1_60 ( .A(_999__bF_buf3), .B(_991__bF_buf1), .C(PC_STACK_14__4_), .Y(_27_) );
OAI21X1 OAI21X1_61 ( .A(_1214_), .B(_1109__bF_buf2), .C(_27_), .Y(_28_) );
OAI21X1 OAI21X1_62 ( .A(_1217_), .B(_1109__bF_buf2), .C(_27_), .Y(_30_) );
OAI21X1 OAI21X1_63 ( .A(_1109__bF_buf2), .B(_1220_), .C(_27_), .Y(_32_) );
OAI21X1 OAI21X1_64 ( .A(_999__bF_buf3), .B(_991__bF_buf1), .C(PC_STACK_14__5_), .Y(_34_) );
OAI21X1 OAI21X1_65 ( .A(_1239_), .B(_1109__bF_buf2), .C(_34_), .Y(_35_) );
OAI21X1 OAI21X1_66 ( .A(_1242_), .B(_1109__bF_buf2), .C(_34_), .Y(_37_) );
OAI21X1 OAI21X1_67 ( .A(_1109__bF_buf2), .B(_1245_), .C(_34_), .Y(_39_) );
OAI21X1 OAI21X1_68 ( .A(_999__bF_buf5), .B(_982__bF_buf0), .C(PC_STACK_6__3_), .Y(_1178_) );
OAI21X1 OAI21X1_69 ( .A(_999__bF_buf1), .B(_991__bF_buf3), .C(PC_STACK_14__6_), .Y(_41_) );
OAI21X1 OAI21X1_70 ( .A(_43_), .B(_42_), .C(_1030__bF_buf9), .Y(_44_) );
OAI21X1 OAI21X1_71 ( .A(_1497_), .B(_1109__bF_buf4), .C(_41_), .Y(_46_) );
OAI21X1 OAI21X1_72 ( .A(_1253_), .B(_1023_), .C(_47_), .Y(_48_) );
OAI21X1 OAI21X1_73 ( .A(_1304_), .B(rst_bF_buf1), .C(_1023_), .Y(_50_) );
OAI21X1 OAI21X1_74 ( .A(PC_STACK_14__7_), .B(_1023_), .C(_50_), .Y(_51_) );
OAI21X1 OAI21X1_75 ( .A(_999__bF_buf0), .B(_991__bF_buf0), .C(PC_STACK_14__7_), .Y(_52_) );
OAI21X1 OAI21X1_76 ( .A(_1504_), .B(_1109__bF_buf0), .C(_52_), .Y(_53_) );
OAI21X1 OAI21X1_77 ( .A(_56_), .B(_1311__bF_buf0), .C(_54_), .Y(_57_) );
OAI21X1 OAI21X1_78 ( .A(_51_), .B(_1301__bF_buf6), .C(_58_), .Y(_5__7_) );
OAI21X1 OAI21X1_79 ( .A(_1140_), .B(_1543__3_), .C(_1042_), .Y(_1181_) );
OAI21X1 OAI21X1_80 ( .A(_999__bF_buf0), .B(_991__bF_buf3), .C(_1324_), .Y(_59_) );
OAI21X1 OAI21X1_81 ( .A(_1343_), .B(_1109__bF_buf0), .C(_59_), .Y(_60_) );
OAI21X1 OAI21X1_82 ( .A(_999__bF_buf0), .B(_991__bF_buf3), .C(PC_STACK_14__8_), .Y(_61_) );
OAI21X1 OAI21X1_83 ( .A(_1109__bF_buf0), .B(_1345_), .C(_61_), .Y(_62_) );
OAI21X1 OAI21X1_84 ( .A(_60_), .B(_1301__bF_buf4), .C(_64_), .Y(_5__8_) );
OAI21X1 OAI21X1_85 ( .A(_1369_), .B(_1109__bF_buf0), .C(_65_), .Y(_66_) );
OAI21X1 OAI21X1_86 ( .A(_999__bF_buf0), .B(_991__bF_buf0), .C(PC_STACK_14__9_), .Y(_67_) );
OAI21X1 OAI21X1_87 ( .A(_1109__bF_buf0), .B(_1373_), .C(_67_), .Y(_68_) );
OAI21X1 OAI21X1_88 ( .A(_66_), .B(_1301__bF_buf4), .C(_69_), .Y(_5__9_) );
OAI21X1 OAI21X1_89 ( .A(_1037_), .B(_70_), .C(_71_), .Y(_72_) );
OAI21X1 OAI21X1_90 ( .A(_1182_), .B(_1019__bF_buf0), .C(_1178_), .Y(_1183_) );
OAI21X1 OAI21X1_91 ( .A(_71_), .B(_74_), .C(_78_), .Y(_79_) );
OAI21X1 OAI21X1_92 ( .A(_73_), .B(_78_), .C(_79_), .Y(_80_) );
OAI21X1 OAI21X1_93 ( .A(_77_), .B(_985_), .C(_80_), .Y(_16__1_) );
OAI21X1 OAI21X1_94 ( .A(_998_), .B(_985_), .C(_995_), .Y(_82_) );
OAI21X1 OAI21X1_95 ( .A(_84_), .B(_85_), .C(_75_), .Y(_86_) );
OAI21X1 OAI21X1_96 ( .A(_995_), .B(_77_), .C(_87_), .Y(_16__2_) );
OAI21X1 OAI21X1_97 ( .A(PC_pointer_3_), .B(_84_), .C(_88_), .Y(_89_) );
OAI21X1 OAI21X1_98 ( .A(_1104_), .B(_90_), .C(_73_), .Y(_91_) );
OAI21X1 OAI21X1_99 ( .A(_981_), .B(_77_), .C(_92_), .Y(_16__3_) );
OAI21X1 OAI21X1_100 ( .A(_982__bF_buf5), .B(_1002__bF_buf4), .C(PC_STACK_7__0_), .Y(_93_) );
OAI21X1 OAI21X1_101 ( .A(_1019__bF_buf0), .B(_1185_), .C(_1178_), .Y(_1186_) );
OAI21X1 OAI21X1_102 ( .A(_1032_), .B(_1020__bF_buf3), .C(_93_), .Y(_94_) );
OAI21X1 OAI21X1_103 ( .A(_1035_), .B(_1020__bF_buf3), .C(_93_), .Y(_96_) );
OAI21X1 OAI21X1_104 ( .A(_1020__bF_buf3), .B(_1043_), .C(_93_), .Y(_98_) );
OAI21X1 OAI21X1_105 ( .A(_982__bF_buf5), .B(_1002__bF_buf4), .C(PC_STACK_7__1_), .Y(_100_) );
OAI21X1 OAI21X1_106 ( .A(_1067_), .B(_1020__bF_buf3), .C(_100_), .Y(_101_) );
OAI21X1 OAI21X1_107 ( .A(_1020__bF_buf3), .B(_1070_), .C(_100_), .Y(_103_) );
OAI21X1 OAI21X1_108 ( .A(_1073_), .B(_1020__bF_buf3), .C(_100_), .Y(_105_) );
OAI21X1 OAI21X1_109 ( .A(_982__bF_buf5), .B(_1002__bF_buf1), .C(PC_STACK_7__2_), .Y(_107_) );
OAI21X1 OAI21X1_110 ( .A(_1142_), .B(_1020__bF_buf2), .C(_107_), .Y(_108_) );
OAI21X1 OAI21X1_111 ( .A(_1020__bF_buf2), .B(_1145_), .C(_107_), .Y(_110_) );
OAI21X1 OAI21X1_112 ( .A(_1032_), .B(_1019__bF_buf2), .C(_1031_), .Y(_1033_) );
OAI21X1 OAI21X1_113 ( .A(_1019__bF_buf0), .B(_1188_), .C(_1178_), .Y(_1189_) );
OAI21X1 OAI21X1_114 ( .A(_1148_), .B(_1020__bF_buf2), .C(_107_), .Y(_112_) );
OAI21X1 OAI21X1_115 ( .A(_982__bF_buf0), .B(_1002__bF_buf4), .C(PC_STACK_7__3_), .Y(_114_) );
OAI21X1 OAI21X1_116 ( .A(_1182_), .B(_1020__bF_buf0), .C(_114_), .Y(_115_) );
OAI21X1 OAI21X1_117 ( .A(_1185_), .B(_1020__bF_buf0), .C(_114_), .Y(_117_) );
OAI21X1 OAI21X1_118 ( .A(_1020__bF_buf0), .B(_1188_), .C(_114_), .Y(_119_) );
OAI21X1 OAI21X1_119 ( .A(_982__bF_buf0), .B(_1002__bF_buf5), .C(PC_STACK_7__4_), .Y(_121_) );
OAI21X1 OAI21X1_120 ( .A(_1214_), .B(_1020__bF_buf0), .C(_121_), .Y(_122_) );
OAI21X1 OAI21X1_121 ( .A(_1217_), .B(_1020__bF_buf1), .C(_121_), .Y(_124_) );
OAI21X1 OAI21X1_122 ( .A(_1020__bF_buf0), .B(_1220_), .C(_121_), .Y(_126_) );
OAI21X1 OAI21X1_123 ( .A(PC_STACK_7__5_), .B(_1104_), .C(_128_), .Y(_129_) );
OAI21X1 OAI21X1_124 ( .A(_999__bF_buf5), .B(_982__bF_buf0), .C(PC_STACK_6__4_), .Y(_1210_) );
OAI21X1 OAI21X1_125 ( .A(_982__bF_buf3), .B(_1002__bF_buf5), .C(PC_STACK_7__5_), .Y(_130_) );
OAI21X1 OAI21X1_126 ( .A(_1242_), .B(_1020__bF_buf4), .C(_130_), .Y(_131_) );
OAI21X1 OAI21X1_127 ( .A(_1020__bF_buf4), .B(_1245_), .C(_130_), .Y(_133_) );
OAI21X1 OAI21X1_128 ( .A(_129_), .B(_1301__bF_buf0), .C(_136_), .Y(_13__5_) );
OAI21X1 OAI21X1_129 ( .A(_982__bF_buf2), .B(_1002__bF_buf3), .C(PC_STACK_7__6_), .Y(_137_) );
OAI21X1 OAI21X1_130 ( .A(_139_), .B(_138_), .C(_1030__bF_buf5), .Y(_140_) );
OAI21X1 OAI21X1_131 ( .A(_1497_), .B(_1020__bF_buf4), .C(_137_), .Y(_142_) );
OAI21X1 OAI21X1_132 ( .A(_1304_), .B(rst_bF_buf0), .C(_1104_), .Y(_146_) );
OAI21X1 OAI21X1_133 ( .A(PC_STACK_7__7_), .B(_1104_), .C(_146_), .Y(_147_) );
OAI21X1 OAI21X1_134 ( .A(_982__bF_buf4), .B(_1002__bF_buf3), .C(PC_STACK_7__7_), .Y(_148_) );
OAI21X1 OAI21X1_135 ( .A(_1211_), .B(_1212_), .C(_1213_), .Y(_1214_) );
OAI21X1 OAI21X1_136 ( .A(_1504_), .B(_1020__bF_buf4), .C(_148_), .Y(_149_) );
OAI21X1 OAI21X1_137 ( .A(_152_), .B(_1311__bF_buf0), .C(_150_), .Y(_153_) );
OAI21X1 OAI21X1_138 ( .A(_147_), .B(_1301__bF_buf6), .C(_154_), .Y(_13__7_) );
OAI21X1 OAI21X1_139 ( .A(_982__bF_buf3), .B(_1002__bF_buf5), .C(_1329_), .Y(_155_) );
OAI21X1 OAI21X1_140 ( .A(_1343_), .B(_1020__bF_buf1), .C(_155_), .Y(_156_) );
OAI21X1 OAI21X1_141 ( .A(_982__bF_buf3), .B(_1002__bF_buf5), .C(PC_STACK_7__8_), .Y(_157_) );
OAI21X1 OAI21X1_142 ( .A(_1020__bF_buf1), .B(_1345_), .C(_157_), .Y(_158_) );
OAI21X1 OAI21X1_143 ( .A(_156_), .B(_1301__bF_buf5), .C(_160_), .Y(_13__8_) );
OAI21X1 OAI21X1_144 ( .A(_982__bF_buf3), .B(_1002__bF_buf5), .C(_1353_), .Y(_161_) );
OAI21X1 OAI21X1_145 ( .A(_1369_), .B(_1020__bF_buf1), .C(_161_), .Y(_162_) );
OAI21X1 OAI21X1_146 ( .A(_1214_), .B(_1019__bF_buf3), .C(_1210_), .Y(_1215_) );
OAI21X1 OAI21X1_147 ( .A(_982__bF_buf3), .B(_1002__bF_buf5), .C(PC_STACK_7__9_), .Y(_163_) );
OAI21X1 OAI21X1_148 ( .A(_1020__bF_buf1), .B(_1373_), .C(_163_), .Y(_164_) );
OAI21X1 OAI21X1_149 ( .A(_162_), .B(_1301__bF_buf5), .C(_165_), .Y(_13__9_) );
OAI21X1 OAI21X1_150 ( .A(_1002__bF_buf0), .B(_991__bF_buf2), .C(PC_STACK_15__0_), .Y(_166_) );
OAI21X1 OAI21X1_151 ( .A(_1032_), .B(_1085__bF_buf0), .C(_166_), .Y(_167_) );
OAI21X1 OAI21X1_152 ( .A(_1085__bF_buf0), .B(_1035_), .C(_166_), .Y(_169_) );
OAI21X1 OAI21X1_153 ( .A(_1085__bF_buf0), .B(_1043_), .C(_166_), .Y(_171_) );
OAI21X1 OAI21X1_154 ( .A(_1002__bF_buf2), .B(_991__bF_buf2), .C(PC_STACK_15__1_), .Y(_173_) );
OAI21X1 OAI21X1_155 ( .A(_1067_), .B(_1085__bF_buf2), .C(_173_), .Y(_174_) );
OAI21X1 OAI21X1_156 ( .A(_1085__bF_buf2), .B(_1070_), .C(_173_), .Y(_176_) );
OAI21X1 OAI21X1_157 ( .A(_1019__bF_buf1), .B(_1217_), .C(_1210_), .Y(_1218_) );
OAI21X1 OAI21X1_158 ( .A(_1085__bF_buf2), .B(_1073_), .C(_173_), .Y(_178_) );
OAI21X1 OAI21X1_159 ( .A(_1002__bF_buf2), .B(_991__bF_buf2), .C(PC_STACK_15__2_), .Y(_180_) );
OAI21X1 OAI21X1_160 ( .A(_1142_), .B(_1085__bF_buf1), .C(_180_), .Y(_181_) );
OAI21X1 OAI21X1_161 ( .A(_1085__bF_buf1), .B(_1145_), .C(_180_), .Y(_183_) );
OAI21X1 OAI21X1_162 ( .A(_1085__bF_buf1), .B(_1148_), .C(_180_), .Y(_185_) );
OAI21X1 OAI21X1_163 ( .A(_1002__bF_buf3), .B(_991__bF_buf6), .C(PC_STACK_15__3_), .Y(_187_) );
OAI21X1 OAI21X1_164 ( .A(_1182_), .B(_1085__bF_buf4), .C(_187_), .Y(_188_) );
OAI21X1 OAI21X1_165 ( .A(_1085__bF_buf4), .B(_1185_), .C(_187_), .Y(_190_) );
OAI21X1 OAI21X1_166 ( .A(_1085__bF_buf4), .B(_1188_), .C(_187_), .Y(_192_) );
OAI21X1 OAI21X1_167 ( .A(_1002__bF_buf2), .B(_991__bF_buf2), .C(PC_STACK_15__4_), .Y(_194_) );
OAI21X1 OAI21X1_168 ( .A(_1019__bF_buf3), .B(_1220_), .C(_1210_), .Y(_1221_) );
OAI21X1 OAI21X1_169 ( .A(_1214_), .B(_1085__bF_buf1), .C(_194_), .Y(_195_) );
OAI21X1 OAI21X1_170 ( .A(_1085__bF_buf1), .B(_1217_), .C(_194_), .Y(_197_) );
OAI21X1 OAI21X1_171 ( .A(_1085__bF_buf1), .B(_1220_), .C(_194_), .Y(_199_) );
OAI21X1 OAI21X1_172 ( .A(_1002__bF_buf2), .B(_991__bF_buf2), .C(PC_STACK_15__5_), .Y(_201_) );
OAI21X1 OAI21X1_173 ( .A(_1239_), .B(_1085__bF_buf2), .C(_201_), .Y(_202_) );
OAI21X1 OAI21X1_174 ( .A(_1085__bF_buf2), .B(_1242_), .C(_201_), .Y(_204_) );
OAI21X1 OAI21X1_175 ( .A(_1085__bF_buf2), .B(_1245_), .C(_201_), .Y(_206_) );
OAI21X1 OAI21X1_176 ( .A(_1002__bF_buf1), .B(_991__bF_buf4), .C(PC_STACK_15__6_), .Y(_208_) );
OAI21X1 OAI21X1_177 ( .A(_210_), .B(_209_), .C(_1030__bF_buf9), .Y(_211_) );
OAI21X1 OAI21X1_178 ( .A(_1085__bF_buf4), .B(_1497_), .C(_208_), .Y(_213_) );
OAI21X1 OAI21X1_179 ( .A(_999__bF_buf5), .B(_982__bF_buf0), .C(PC_STACK_6__5_), .Y(_1236_) );
OAI21X1 OAI21X1_180 ( .A(_1262_), .B(_1003_), .C(_214_), .Y(_215_) );
OAI21X1 OAI21X1_181 ( .A(_1304_), .B(rst_bF_buf2), .C(_1003_), .Y(_217_) );
OAI21X1 OAI21X1_182 ( .A(PC_STACK_15__7_), .B(_1003_), .C(_217_), .Y(_218_) );
OAI21X1 OAI21X1_183 ( .A(_1002__bF_buf3), .B(_991__bF_buf0), .C(PC_STACK_15__7_), .Y(_219_) );
OAI21X1 OAI21X1_184 ( .A(_1085__bF_buf3), .B(_1504_), .C(_219_), .Y(_220_) );
OAI21X1 OAI21X1_185 ( .A(_223_), .B(_1311__bF_buf0), .C(_221_), .Y(_224_) );
OAI21X1 OAI21X1_186 ( .A(_218_), .B(_1301__bF_buf6), .C(_225_), .Y(_6__7_) );
OAI21X1 OAI21X1_187 ( .A(_1002__bF_buf1), .B(_991__bF_buf0), .C(_1323_), .Y(_226_) );
OAI21X1 OAI21X1_188 ( .A(_1343_), .B(_1085__bF_buf3), .C(_226_), .Y(_227_) );
OAI21X1 OAI21X1_189 ( .A(_1002__bF_buf3), .B(_991__bF_buf0), .C(PC_STACK_15__8_), .Y(_228_) );
OAI21X1 OAI21X1_190 ( .A(_1211_), .B(_1212_), .C(_1235_), .Y(_1238_) );
OAI21X1 OAI21X1_191 ( .A(_1085__bF_buf3), .B(_1345_), .C(_228_), .Y(_229_) );
OAI21X1 OAI21X1_192 ( .A(_1085__bF_buf3), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_230_) );
OAI21X1 OAI21X1_193 ( .A(_227_), .B(_1301__bF_buf4), .C(_232_), .Y(_6__8_) );
OAI21X1 OAI21X1_194 ( .A(_1369_), .B(_1085__bF_buf3), .C(_233_), .Y(_234_) );
OAI21X1 OAI21X1_195 ( .A(_1002__bF_buf1), .B(_991__bF_buf3), .C(PC_STACK_15__9_), .Y(_235_) );
OAI21X1 OAI21X1_196 ( .A(_1085__bF_buf3), .B(_1373_), .C(_235_), .Y(_236_) );
OAI21X1 OAI21X1_197 ( .A(_234_), .B(_1301__bF_buf4), .C(_237_), .Y(_6__9_) );
OAI21X1 OAI21X1_198 ( .A(_986__bF_buf5), .B(_996__bF_buf5), .C(PC_STACK_9__0_), .Y(_238_) );
OAI21X1 OAI21X1_199 ( .A(_1032_), .B(_1201__bF_buf1), .C(_238_), .Y(_239_) );
OAI21X1 OAI21X1_200 ( .A(_1201__bF_buf2), .B(_1035_), .C(_238_), .Y(_241_) );
OAI21X1 OAI21X1_201 ( .A(_1239_), .B(_1019__bF_buf3), .C(_1236_), .Y(_1240_) );
OAI21X1 OAI21X1_202 ( .A(_1201__bF_buf1), .B(_1043_), .C(_238_), .Y(_243_) );
OAI21X1 OAI21X1_203 ( .A(_986__bF_buf5), .B(_996__bF_buf5), .C(PC_STACK_9__1_), .Y(_245_) );
OAI21X1 OAI21X1_204 ( .A(_1067_), .B(_1201__bF_buf3), .C(_245_), .Y(_246_) );
OAI21X1 OAI21X1_205 ( .A(_1201__bF_buf3), .B(_1070_), .C(_245_), .Y(_248_) );
OAI21X1 OAI21X1_206 ( .A(_1201__bF_buf3), .B(_1073_), .C(_245_), .Y(_250_) );
OAI21X1 OAI21X1_207 ( .A(_986__bF_buf4), .B(_996__bF_buf2), .C(PC_STACK_9__2_), .Y(_252_) );
OAI21X1 OAI21X1_208 ( .A(_1142_), .B(_1201__bF_buf2), .C(_252_), .Y(_253_) );
OAI21X1 OAI21X1_209 ( .A(_1201__bF_buf4), .B(_1145_), .C(_252_), .Y(_255_) );
OAI21X1 OAI21X1_210 ( .A(_1201__bF_buf2), .B(_1148_), .C(_252_), .Y(_257_) );
OAI21X1 OAI21X1_211 ( .A(_986__bF_buf5), .B(_996__bF_buf5), .C(PC_STACK_9__3_), .Y(_259_) );
OAI21X1 OAI21X1_212 ( .A(_1019__bF_buf0), .B(_1242_), .C(_1236_), .Y(_1243_) );
OAI21X1 OAI21X1_213 ( .A(_1182_), .B(_1201__bF_buf1), .C(_259_), .Y(_260_) );
OAI21X1 OAI21X1_214 ( .A(_1201__bF_buf1), .B(_1185_), .C(_259_), .Y(_262_) );
OAI21X1 OAI21X1_215 ( .A(_1201__bF_buf1), .B(_1188_), .C(_259_), .Y(_264_) );
OAI21X1 OAI21X1_216 ( .A(_986__bF_buf5), .B(_996__bF_buf5), .C(PC_STACK_9__4_), .Y(_266_) );
OAI21X1 OAI21X1_217 ( .A(_1214_), .B(_1201__bF_buf3), .C(_266_), .Y(_267_) );
OAI21X1 OAI21X1_218 ( .A(_1201__bF_buf0), .B(_1217_), .C(_266_), .Y(_269_) );
OAI21X1 OAI21X1_219 ( .A(_1201__bF_buf0), .B(_1220_), .C(_266_), .Y(_271_) );
OAI21X1 OAI21X1_220 ( .A(_986__bF_buf5), .B(_996__bF_buf3), .C(PC_STACK_9__5_), .Y(_273_) );
OAI21X1 OAI21X1_221 ( .A(_1239_), .B(_1201__bF_buf3), .C(_273_), .Y(_274_) );
OAI21X1 OAI21X1_222 ( .A(_1201__bF_buf0), .B(_1242_), .C(_273_), .Y(_276_) );
OAI21X1 OAI21X1_223 ( .A(_1019__bF_buf2), .B(_1035_), .C(_1031_), .Y(_1036_) );
OAI21X1 OAI21X1_224 ( .A(_1019__bF_buf0), .B(_1245_), .C(_1236_), .Y(_1246_) );
OAI21X1 OAI21X1_225 ( .A(_1201__bF_buf0), .B(_1245_), .C(_273_), .Y(_278_) );
OAI21X1 OAI21X1_226 ( .A(_986__bF_buf4), .B(_996__bF_buf2), .C(PC_STACK_9__6_), .Y(_280_) );
OAI21X1 OAI21X1_227 ( .A(_282_), .B(_281_), .C(_1030__bF_buf0), .Y(_283_) );
OAI21X1 OAI21X1_228 ( .A(_1201__bF_buf2), .B(_1497_), .C(_280_), .Y(_285_) );
OAI21X1 OAI21X1_229 ( .A(_1259_), .B(_997__bF_buf1), .C(_286_), .Y(_287_) );
OAI21X1 OAI21X1_230 ( .A(_1304_), .B(rst_bF_buf2), .C(_997__bF_buf3), .Y(_289_) );
OAI21X1 OAI21X1_231 ( .A(PC_STACK_9__7_), .B(_997__bF_buf3), .C(_289_), .Y(_290_) );
OAI21X1 OAI21X1_232 ( .A(_986__bF_buf0), .B(_996__bF_buf4), .C(PC_STACK_9__7_), .Y(_291_) );
OAI21X1 OAI21X1_233 ( .A(_1201__bF_buf4), .B(_1504_), .C(_291_), .Y(_292_) );
OAI21X1 OAI21X1_234 ( .A(_295_), .B(_1311__bF_buf3), .C(_293_), .Y(_296_) );
OAI21X1 OAI21X1_235 ( .A(_999__bF_buf2), .B(_982__bF_buf1), .C(PC_STACK_6__6_), .Y(_1270_) );
OAI21X1 OAI21X1_236 ( .A(_290_), .B(_1301__bF_buf1), .C(_297_), .Y(_15__7_) );
OAI21X1 OAI21X1_237 ( .A(_986__bF_buf0), .B(_996__bF_buf4), .C(PC_STACK_9__8_), .Y(_298_) );
OAI21X1 OAI21X1_238 ( .A(_1201__bF_buf4), .B(_1345_), .C(_298_), .Y(_301_) );
OAI21X1 OAI21X1_239 ( .A(_1201__bF_buf4), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_302_) );
OAI21X1 OAI21X1_240 ( .A(_300_), .B(_1301__bF_buf3), .C(_304_), .Y(_15__8_) );
OAI21X1 OAI21X1_241 ( .A(_1369_), .B(_1201__bF_buf4), .C(_305_), .Y(_306_) );
OAI21X1 OAI21X1_242 ( .A(_986__bF_buf0), .B(_996__bF_buf2), .C(PC_STACK_9__9_), .Y(_307_) );
OAI21X1 OAI21X1_243 ( .A(_1201__bF_buf4), .B(_1373_), .C(_307_), .Y(_308_) );
OAI21X1 OAI21X1_244 ( .A(_306_), .B(_1301__bF_buf3), .C(_309_), .Y(_15__9_) );
OAI21X1 OAI21X1_245 ( .A(_999__bF_buf4), .B(_996__bF_buf3), .C(PC_STACK_10__0_), .Y(_311_) );
OAI21X1 OAI21X1_246 ( .A(_1272_), .B(_1543__6_), .C(_1042_), .Y(_1273_) );
OAI21X1 OAI21X1_247 ( .A(_1032_), .B(_310__bF_buf2), .C(_311_), .Y(_312_) );
OAI21X1 OAI21X1_248 ( .A(_310__bF_buf2), .B(_1035_), .C(_311_), .Y(_314_) );
OAI21X1 OAI21X1_249 ( .A(_310__bF_buf2), .B(_1043_), .C(_311_), .Y(_316_) );
OAI21X1 OAI21X1_250 ( .A(_999__bF_buf4), .B(_996__bF_buf5), .C(PC_STACK_10__1_), .Y(_318_) );
OAI21X1 OAI21X1_251 ( .A(_1067_), .B(_310__bF_buf2), .C(_318_), .Y(_319_) );
OAI21X1 OAI21X1_252 ( .A(_310__bF_buf2), .B(_1070_), .C(_318_), .Y(_321_) );
OAI21X1 OAI21X1_253 ( .A(_310__bF_buf2), .B(_1073_), .C(_318_), .Y(_323_) );
OAI21X1 OAI21X1_254 ( .A(_999__bF_buf4), .B(_996__bF_buf3), .C(PC_STACK_10__2_), .Y(_325_) );
OAI21X1 OAI21X1_255 ( .A(_1142_), .B(_310__bF_buf0), .C(_325_), .Y(_326_) );
OAI21X1 OAI21X1_256 ( .A(_310__bF_buf0), .B(_1145_), .C(_325_), .Y(_328_) );
OAI21X1 OAI21X1_257 ( .A(_1275_), .B(_1271_), .C(_1030__bF_buf7), .Y(_1276_) );
OAI21X1 OAI21X1_258 ( .A(_310__bF_buf0), .B(_1148_), .C(_325_), .Y(_330_) );
OAI21X1 OAI21X1_259 ( .A(_999__bF_buf1), .B(_996__bF_buf2), .C(PC_STACK_10__3_), .Y(_332_) );
OAI21X1 OAI21X1_260 ( .A(_1182_), .B(_310__bF_buf3), .C(_332_), .Y(_333_) );
OAI21X1 OAI21X1_261 ( .A(_310__bF_buf3), .B(_1185_), .C(_332_), .Y(_335_) );
OAI21X1 OAI21X1_262 ( .A(_310__bF_buf3), .B(_1188_), .C(_332_), .Y(_337_) );
OAI21X1 OAI21X1_263 ( .A(_999__bF_buf4), .B(_996__bF_buf3), .C(PC_STACK_10__4_), .Y(_339_) );
OAI21X1 OAI21X1_264 ( .A(_1214_), .B(_310__bF_buf1), .C(_339_), .Y(_340_) );
OAI21X1 OAI21X1_265 ( .A(_310__bF_buf1), .B(_1217_), .C(_339_), .Y(_342_) );
OAI21X1 OAI21X1_266 ( .A(_310__bF_buf1), .B(_1220_), .C(_339_), .Y(_344_) );
OAI21X1 OAI21X1_267 ( .A(_999__bF_buf4), .B(_996__bF_buf3), .C(PC_STACK_10__5_), .Y(_346_) );
OAI21X1 OAI21X1_268 ( .A(_1284_), .B(_1080__bF_buf4), .C(_1285_), .Y(_1286_) );
OAI21X1 OAI21X1_269 ( .A(_1239_), .B(_310__bF_buf1), .C(_346_), .Y(_347_) );
OAI21X1 OAI21X1_270 ( .A(_310__bF_buf0), .B(_1242_), .C(_346_), .Y(_349_) );
OAI21X1 OAI21X1_271 ( .A(_310__bF_buf0), .B(_1245_), .C(_346_), .Y(_351_) );
OAI21X1 OAI21X1_272 ( .A(_999__bF_buf0), .B(_996__bF_buf4), .C(PC_STACK_10__6_), .Y(_353_) );
OAI21X1 OAI21X1_273 ( .A(_355_), .B(_354_), .C(_1030__bF_buf9), .Y(_356_) );
OAI21X1 OAI21X1_274 ( .A(_310__bF_buf3), .B(_1497_), .C(_353_), .Y(_358_) );
OAI21X1 OAI21X1_275 ( .A(_1304_), .B(rst_bF_buf1), .C(_1000__bF_buf3), .Y(_362_) );
OAI21X1 OAI21X1_276 ( .A(PC_STACK_10__7_), .B(_1000__bF_buf3), .C(_362_), .Y(_363_) );
OAI21X1 OAI21X1_277 ( .A(_999__bF_buf0), .B(_996__bF_buf4), .C(PC_STACK_10__7_), .Y(_364_) );
OAI21X1 OAI21X1_278 ( .A(_310__bF_buf3), .B(_1504_), .C(_364_), .Y(_365_) );
OAI21X1 OAI21X1_279 ( .A(_1237_), .B(_1269_), .C(_1300_), .Y(_1303_) );
OAI21X1 OAI21X1_280 ( .A(_368_), .B(_1311__bF_buf3), .C(_366_), .Y(_369_) );
OAI21X1 OAI21X1_281 ( .A(_363_), .B(_1301__bF_buf4), .C(_370_), .Y(_1__7_) );
OAI21X1 OAI21X1_282 ( .A(_999__bF_buf4), .B(_996__bF_buf0), .C(PC_STACK_10__8_), .Y(_371_) );
OAI21X1 OAI21X1_283 ( .A(_310__bF_buf1), .B(_1345_), .C(_371_), .Y(_374_) );
OAI21X1 OAI21X1_284 ( .A(_373_), .B(_1301__bF_buf3), .C(_376_), .Y(_1__8_) );
OAI21X1 OAI21X1_285 ( .A(_1369_), .B(_310__bF_buf1), .C(_377_), .Y(_378_) );
OAI21X1 OAI21X1_286 ( .A(_999__bF_buf4), .B(_996__bF_buf0), .C(PC_STACK_10__9_), .Y(_379_) );
OAI21X1 OAI21X1_287 ( .A(_310__bF_buf3), .B(_1373_), .C(_379_), .Y(_380_) );
OAI21X1 OAI21X1_288 ( .A(_378_), .B(_1301__bF_buf3), .C(_381_), .Y(_1__9_) );
OAI21X1 OAI21X1_289 ( .A(_996__bF_buf1), .B(_983__bF_buf3), .C(PC_STACK_8__0_), .Y(_382_) );
OAI21X1 OAI21X1_290 ( .A(_1304_), .B(rst_bF_buf3), .C(_1102__bF_buf2), .Y(_1305_) );
OAI21X1 OAI21X1_291 ( .A(_1032_), .B(_1095__bF_buf1), .C(_382_), .Y(_383_) );
OAI21X1 OAI21X1_292 ( .A(_1035_), .B(_1095__bF_buf2), .C(_382_), .Y(_385_) );
OAI21X1 OAI21X1_293 ( .A(_1095__bF_buf1), .B(_1043_), .C(_382_), .Y(_387_) );
OAI21X1 OAI21X1_294 ( .A(_996__bF_buf5), .B(_983__bF_buf2), .C(PC_STACK_8__1_), .Y(_389_) );
OAI21X1 OAI21X1_295 ( .A(_1067_), .B(_1095__bF_buf0), .C(_389_), .Y(_390_) );
OAI21X1 OAI21X1_296 ( .A(_1095__bF_buf3), .B(_1070_), .C(_389_), .Y(_392_) );
OAI21X1 OAI21X1_297 ( .A(_1073_), .B(_1095__bF_buf3), .C(_389_), .Y(_394_) );
OAI21X1 OAI21X1_298 ( .A(_996__bF_buf1), .B(_983__bF_buf3), .C(PC_STACK_8__2_), .Y(_396_) );
OAI21X1 OAI21X1_299 ( .A(_1142_), .B(_1095__bF_buf2), .C(_396_), .Y(_397_) );
OAI21X1 OAI21X1_300 ( .A(_1095__bF_buf2), .B(_1145_), .C(_396_), .Y(_399_) );
OAI21X1 OAI21X1_301 ( .A(PC_STACK_6__7_), .B(_1102__bF_buf2), .C(_1305_), .Y(_1306_) );
OAI21X1 OAI21X1_302 ( .A(_1148_), .B(_1095__bF_buf2), .C(_396_), .Y(_401_) );
OAI21X1 OAI21X1_303 ( .A(_996__bF_buf5), .B(_983__bF_buf2), .C(PC_STACK_8__3_), .Y(_403_) );
OAI21X1 OAI21X1_304 ( .A(_1182_), .B(_1095__bF_buf0), .C(_403_), .Y(_404_) );
OAI21X1 OAI21X1_305 ( .A(_1185_), .B(_1095__bF_buf0), .C(_403_), .Y(_406_) );
OAI21X1 OAI21X1_306 ( .A(_1095__bF_buf0), .B(_1188_), .C(_403_), .Y(_408_) );
OAI21X1 OAI21X1_307 ( .A(_996__bF_buf3), .B(_983__bF_buf2), .C(PC_STACK_8__4_), .Y(_410_) );
OAI21X1 OAI21X1_308 ( .A(_1214_), .B(_1095__bF_buf3), .C(_410_), .Y(_411_) );
OAI21X1 OAI21X1_309 ( .A(_1217_), .B(_1095__bF_buf3), .C(_410_), .Y(_413_) );
OAI21X1 OAI21X1_310 ( .A(_1095__bF_buf3), .B(_1220_), .C(_410_), .Y(_415_) );
OAI21X1 OAI21X1_311 ( .A(PC_STACK_8__5_), .B(_1004__bF_buf0), .C(_417_), .Y(_418_) );
OAI21X1 OAI21X1_312 ( .A(_999__bF_buf2), .B(_982__bF_buf2), .C(PC_STACK_6__7_), .Y(_1308_) );
OAI21X1 OAI21X1_313 ( .A(_996__bF_buf5), .B(_983__bF_buf3), .C(PC_STACK_8__5_), .Y(_419_) );
OAI21X1 OAI21X1_314 ( .A(_1242_), .B(_1095__bF_buf1), .C(_419_), .Y(_420_) );
OAI21X1 OAI21X1_315 ( .A(_1095__bF_buf1), .B(_1245_), .C(_419_), .Y(_422_) );
OAI21X1 OAI21X1_316 ( .A(_418_), .B(_1301__bF_buf1), .C(_425_), .Y(_14__5_) );
OAI21X1 OAI21X1_317 ( .A(_996__bF_buf0), .B(_983__bF_buf2), .C(PC_STACK_8__6_), .Y(_426_) );
OAI21X1 OAI21X1_318 ( .A(_428_), .B(_427_), .C(_1030__bF_buf0), .Y(_429_) );
OAI21X1 OAI21X1_319 ( .A(_1497_), .B(_1095__bF_buf4), .C(_426_), .Y(_431_) );
OAI21X1 OAI21X1_320 ( .A(_1260_), .B(_1004__bF_buf1), .C(_432_), .Y(_433_) );
OAI21X1 OAI21X1_321 ( .A(_1304_), .B(rst_bF_buf1), .C(_1004__bF_buf2), .Y(_435_) );
OAI21X1 OAI21X1_322 ( .A(PC_STACK_8__7_), .B(_1004__bF_buf2), .C(_435_), .Y(_436_) );
OAI21X1 OAI21X1_323 ( .A(_1315_), .B(_1311__bF_buf2), .C(_1312_), .Y(_1316_) );
OAI21X1 OAI21X1_324 ( .A(_996__bF_buf4), .B(_983__bF_buf6), .C(PC_STACK_8__7_), .Y(_437_) );
OAI21X1 OAI21X1_325 ( .A(_1504_), .B(_1095__bF_buf4), .C(_437_), .Y(_438_) );
OAI21X1 OAI21X1_326 ( .A(_441_), .B(_1311__bF_buf3), .C(_439_), .Y(_442_) );
OAI21X1 OAI21X1_327 ( .A(_436_), .B(_1301__bF_buf4), .C(_443_), .Y(_14__7_) );
OAI21X1 OAI21X1_328 ( .A(_996__bF_buf0), .B(_983__bF_buf2), .C(PC_STACK_8__8_), .Y(_444_) );
OAI21X1 OAI21X1_329 ( .A(_1095__bF_buf4), .B(_1345_), .C(_444_), .Y(_447_) );
OAI21X1 OAI21X1_330 ( .A(_446_), .B(_1301__bF_buf3), .C(_449_), .Y(_14__8_) );
OAI21X1 OAI21X1_331 ( .A(_1369_), .B(_1095__bF_buf4), .C(_450_), .Y(_451_) );
OAI21X1 OAI21X1_332 ( .A(_996__bF_buf2), .B(_983__bF_buf2), .C(PC_STACK_8__9_), .Y(_452_) );
OAI21X1 OAI21X1_333 ( .A(_1095__bF_buf4), .B(_1373_), .C(_452_), .Y(_453_) );
OAI21X1 OAI21X1_334 ( .A(_1019__bF_buf2), .B(_1043_), .C(_1031_), .Y(_1044_) );
OAI21X1 OAI21X1_335 ( .A(_1306_), .B(_1301__bF_buf2), .C(_1317_), .Y(_12__7_) );
OAI21X1 OAI21X1_336 ( .A(_451_), .B(_1301__bF_buf1), .C(_454_), .Y(_14__9_) );
OAI21X1 OAI21X1_337 ( .A(_996__bF_buf1), .B(_1002__bF_buf0), .C(PC_STACK_11__0_), .Y(_455_) );
OAI21X1 OAI21X1_338 ( .A(_1032_), .B(_1084__bF_buf1), .C(_455_), .Y(_456_) );
OAI21X1 OAI21X1_339 ( .A(_1035_), .B(_1084__bF_buf3), .C(_455_), .Y(_458_) );
OAI21X1 OAI21X1_340 ( .A(_1084__bF_buf3), .B(_1043_), .C(_455_), .Y(_460_) );
OAI21X1 OAI21X1_341 ( .A(_996__bF_buf1), .B(_1002__bF_buf2), .C(PC_STACK_11__1_), .Y(_462_) );
OAI21X1 OAI21X1_342 ( .A(_1067_), .B(_1084__bF_buf0), .C(_462_), .Y(_463_) );
OAI21X1 OAI21X1_343 ( .A(_1084__bF_buf1), .B(_1070_), .C(_462_), .Y(_465_) );
OAI21X1 OAI21X1_344 ( .A(_1073_), .B(_1084__bF_buf0), .C(_462_), .Y(_467_) );
OAI21X1 OAI21X1_345 ( .A(_996__bF_buf1), .B(_1002__bF_buf0), .C(PC_STACK_11__2_), .Y(_469_) );
OAI21X1 OAI21X1_346 ( .A(_999__bF_buf2), .B(_982__bF_buf3), .C(PC_STACK_6__8_), .Y(_1339_) );
OAI21X1 OAI21X1_347 ( .A(_1142_), .B(_1084__bF_buf3), .C(_469_), .Y(_470_) );
OAI21X1 OAI21X1_348 ( .A(_1084__bF_buf3), .B(_1145_), .C(_469_), .Y(_472_) );
OAI21X1 OAI21X1_349 ( .A(_1148_), .B(_1084__bF_buf3), .C(_469_), .Y(_474_) );
OAI21X1 OAI21X1_350 ( .A(_996__bF_buf1), .B(_1002__bF_buf2), .C(PC_STACK_11__3_), .Y(_476_) );
OAI21X1 OAI21X1_351 ( .A(_1182_), .B(_1084__bF_buf0), .C(_476_), .Y(_477_) );
OAI21X1 OAI21X1_352 ( .A(_1185_), .B(_1084__bF_buf0), .C(_476_), .Y(_479_) );
OAI21X1 OAI21X1_353 ( .A(_1084__bF_buf0), .B(_1188_), .C(_476_), .Y(_481_) );
OAI21X1 OAI21X1_354 ( .A(_996__bF_buf3), .B(_1002__bF_buf0), .C(PC_STACK_11__4_), .Y(_483_) );
OAI21X1 OAI21X1_355 ( .A(_1214_), .B(_1084__bF_buf2), .C(_483_), .Y(_484_) );
OAI21X1 OAI21X1_356 ( .A(_1217_), .B(_1084__bF_buf2), .C(_483_), .Y(_486_) );
OAI21X1 OAI21X1_357 ( .A(_1341_), .B(_1543__8_), .C(_1042_), .Y(_1342_) );
OAI21X1 OAI21X1_358 ( .A(_1084__bF_buf2), .B(_1220_), .C(_483_), .Y(_488_) );
OAI21X1 OAI21X1_359 ( .A(_996__bF_buf1), .B(_1002__bF_buf0), .C(PC_STACK_11__5_), .Y(_490_) );
OAI21X1 OAI21X1_360 ( .A(_1239_), .B(_1084__bF_buf1), .C(_490_), .Y(_491_) );
OAI21X1 OAI21X1_361 ( .A(_1242_), .B(_1084__bF_buf1), .C(_490_), .Y(_493_) );
OAI21X1 OAI21X1_362 ( .A(_1084__bF_buf1), .B(_1245_), .C(_490_), .Y(_495_) );
OAI21X1 OAI21X1_363 ( .A(_996__bF_buf0), .B(_1002__bF_buf0), .C(PC_STACK_11__6_), .Y(_497_) );
OAI21X1 OAI21X1_364 ( .A(_499_), .B(_498_), .C(_1030__bF_buf0), .Y(_500_) );
OAI21X1 OAI21X1_365 ( .A(_1497_), .B(_1084__bF_buf2), .C(_497_), .Y(_502_) );
OAI21X1 OAI21X1_366 ( .A(_1252_), .B(_1026_), .C(_503_), .Y(_504_) );
OAI21X1 OAI21X1_367 ( .A(_1304_), .B(rst_bF_buf1), .C(_1026_), .Y(_506_) );
OAI21X1 OAI21X1_368 ( .A(_1019__bF_buf3), .B(_1345_), .C(_1339_), .Y(_1346_) );
OAI21X1 OAI21X1_369 ( .A(PC_STACK_11__7_), .B(_1026_), .C(_506_), .Y(_507_) );
OAI21X1 OAI21X1_370 ( .A(_996__bF_buf4), .B(_1002__bF_buf1), .C(PC_STACK_11__7_), .Y(_508_) );
OAI21X1 OAI21X1_371 ( .A(_1504_), .B(_1084__bF_buf4), .C(_508_), .Y(_509_) );
OAI21X1 OAI21X1_372 ( .A(_512_), .B(_1311__bF_buf0), .C(_510_), .Y(_513_) );
OAI21X1 OAI21X1_373 ( .A(_507_), .B(_1301__bF_buf4), .C(_514_), .Y(_2__7_) );
OAI21X1 OAI21X1_374 ( .A(_996__bF_buf0), .B(_1002__bF_buf0), .C(PC_STACK_11__8_), .Y(_515_) );
OAI21X1 OAI21X1_375 ( .A(_1084__bF_buf4), .B(_1345_), .C(_515_), .Y(_518_) );
OAI21X1 OAI21X1_376 ( .A(_1084__bF_buf4), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_519_) );
OAI21X1 OAI21X1_377 ( .A(_517_), .B(_1301__bF_buf3), .C(_521_), .Y(_2__8_) );
OAI21X1 OAI21X1_378 ( .A(_1369_), .B(_1084__bF_buf4), .C(_522_), .Y(_523_) );
OAI21X1 OAI21X1_379 ( .A(_1344_), .B(_1301__bF_buf5), .C(_1348_), .Y(_12__8_) );
OAI21X1 OAI21X1_380 ( .A(_996__bF_buf4), .B(_1002__bF_buf1), .C(PC_STACK_11__9_), .Y(_524_) );
OAI21X1 OAI21X1_381 ( .A(_1084__bF_buf4), .B(_1373_), .C(_524_), .Y(_525_) );
OAI21X1 OAI21X1_382 ( .A(_523_), .B(_1301__bF_buf3), .C(_526_), .Y(_2__9_) );
OAI21X1 OAI21X1_383 ( .A(_986__bF_buf2), .B(_982__bF_buf6), .C(PC_STACK_5__0_), .Y(_528_) );
OAI21X1 OAI21X1_384 ( .A(_1032_), .B(_527__bF_buf0), .C(_528_), .Y(_529_) );
OAI21X1 OAI21X1_385 ( .A(_527__bF_buf0), .B(_1035_), .C(_528_), .Y(_531_) );
OAI21X1 OAI21X1_386 ( .A(_527__bF_buf0), .B(_1043_), .C(_528_), .Y(_533_) );
OAI21X1 OAI21X1_387 ( .A(_986__bF_buf2), .B(_982__bF_buf6), .C(PC_STACK_5__1_), .Y(_535_) );
OAI21X1 OAI21X1_388 ( .A(_1067_), .B(_527__bF_buf3), .C(_535_), .Y(_536_) );
OAI21X1 OAI21X1_389 ( .A(_527__bF_buf3), .B(_1070_), .C(_535_), .Y(_538_) );
OAI21X1 OAI21X1_390 ( .A(_1020__bF_buf2), .B(_1353_), .C(_1099__bF_buf4), .Y(_1354_) );
OAI21X1 OAI21X1_391 ( .A(_527__bF_buf3), .B(_1073_), .C(_535_), .Y(_540_) );
OAI21X1 OAI21X1_392 ( .A(_986__bF_buf2), .B(_982__bF_buf6), .C(PC_STACK_5__2_), .Y(_542_) );
OAI21X1 OAI21X1_393 ( .A(_1142_), .B(_527__bF_buf0), .C(_542_), .Y(_543_) );
OAI21X1 OAI21X1_394 ( .A(_527__bF_buf0), .B(_1145_), .C(_542_), .Y(_545_) );
OAI21X1 OAI21X1_395 ( .A(_527__bF_buf0), .B(_1148_), .C(_542_), .Y(_547_) );
OAI21X1 OAI21X1_396 ( .A(_986__bF_buf2), .B(_982__bF_buf6), .C(PC_STACK_5__3_), .Y(_549_) );
OAI21X1 OAI21X1_397 ( .A(_1182_), .B(_527__bF_buf3), .C(_549_), .Y(_550_) );
OAI21X1 OAI21X1_398 ( .A(_527__bF_buf3), .B(_1185_), .C(_549_), .Y(_552_) );
OAI21X1 OAI21X1_399 ( .A(_527__bF_buf3), .B(_1188_), .C(_549_), .Y(_554_) );
OAI21X1 OAI21X1_400 ( .A(_986__bF_buf1), .B(_982__bF_buf4), .C(PC_STACK_5__4_), .Y(_556_) );
OAI21X1 OAI21X1_401 ( .A(_1302_), .B(_1338_), .C(_1543__9_), .Y(_1368_) );
OAI21X1 OAI21X1_402 ( .A(_1214_), .B(_527__bF_buf2), .C(_556_), .Y(_557_) );
OAI21X1 OAI21X1_403 ( .A(_527__bF_buf2), .B(_1217_), .C(_556_), .Y(_559_) );
OAI21X1 OAI21X1_404 ( .A(_527__bF_buf2), .B(_1220_), .C(_556_), .Y(_561_) );
OAI21X1 OAI21X1_405 ( .A(_986__bF_buf1), .B(_982__bF_buf4), .C(PC_STACK_5__5_), .Y(_563_) );
OAI21X1 OAI21X1_406 ( .A(_1239_), .B(_527__bF_buf2), .C(_563_), .Y(_564_) );
OAI21X1 OAI21X1_407 ( .A(_527__bF_buf2), .B(_1242_), .C(_563_), .Y(_566_) );
OAI21X1 OAI21X1_408 ( .A(_527__bF_buf2), .B(_1245_), .C(_563_), .Y(_568_) );
OAI21X1 OAI21X1_409 ( .A(_986__bF_buf1), .B(_982__bF_buf4), .C(PC_STACK_5__6_), .Y(_570_) );
OAI21X1 OAI21X1_410 ( .A(_572_), .B(_571_), .C(_1030__bF_buf5), .Y(_573_) );
OAI21X1 OAI21X1_411 ( .A(_527__bF_buf1), .B(_1497_), .C(_570_), .Y(_575_) );
OAI21X1 OAI21X1_412 ( .A(_1369_), .B(_1019__bF_buf3), .C(_1370_), .Y(_1371_) );
OAI21X1 OAI21X1_413 ( .A(_1304_), .B(rst_bF_buf3), .C(_987__bF_buf0), .Y(_579_) );
OAI21X1 OAI21X1_414 ( .A(PC_STACK_5__7_), .B(_987__bF_buf0), .C(_579_), .Y(_580_) );
OAI21X1 OAI21X1_415 ( .A(_986__bF_buf1), .B(_982__bF_buf2), .C(PC_STACK_5__7_), .Y(_581_) );
OAI21X1 OAI21X1_416 ( .A(_527__bF_buf1), .B(_1504_), .C(_581_), .Y(_582_) );
OAI21X1 OAI21X1_417 ( .A(_585_), .B(_1311__bF_buf2), .C(_583_), .Y(_586_) );
OAI21X1 OAI21X1_418 ( .A(_580_), .B(_1301__bF_buf6), .C(_587_), .Y(_11__7_) );
OAI21X1 OAI21X1_419 ( .A(_986__bF_buf1), .B(_982__bF_buf2), .C(PC_STACK_5__8_), .Y(_588_) );
OAI21X1 OAI21X1_420 ( .A(_527__bF_buf1), .B(_1345_), .C(_588_), .Y(_591_) );
OAI21X1 OAI21X1_421 ( .A(_527__bF_buf1), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_592_) );
OAI21X1 OAI21X1_422 ( .A(_590_), .B(_1301__bF_buf6), .C(_594_), .Y(_11__8_) );
OAI21X1 OAI21X1_423 ( .A(_999__bF_buf5), .B(_982__bF_buf3), .C(PC_STACK_6__9_), .Y(_1372_) );
OAI21X1 OAI21X1_424 ( .A(_986__bF_buf1), .B(_982__bF_buf4), .C(_595_), .Y(_596_) );
OAI21X1 OAI21X1_425 ( .A(_1369_), .B(_527__bF_buf1), .C(_596_), .Y(_597_) );
OAI21X1 OAI21X1_426 ( .A(_986__bF_buf1), .B(_982__bF_buf4), .C(PC_STACK_5__9_), .Y(_598_) );
OAI21X1 OAI21X1_427 ( .A(_527__bF_buf1), .B(_1373_), .C(_598_), .Y(_599_) );
OAI21X1 OAI21X1_428 ( .A(_597_), .B(_1301__bF_buf6), .C(_600_), .Y(_11__9_) );
OAI21X1 OAI21X1_429 ( .A(_982__bF_buf5), .B(_983__bF_buf4), .C(PC_STACK_4__0_), .Y(_601_) );
OAI21X1 OAI21X1_430 ( .A(_1032_), .B(_1250__bF_buf2), .C(_601_), .Y(_602_) );
OAI21X1 OAI21X1_431 ( .A(_1250__bF_buf2), .B(_1035_), .C(_601_), .Y(_604_) );
OAI21X1 OAI21X1_432 ( .A(_1250__bF_buf2), .B(_1043_), .C(_601_), .Y(_606_) );
OAI21X1 OAI21X1_433 ( .A(_982__bF_buf6), .B(_983__bF_buf6), .C(PC_STACK_4__1_), .Y(_608_) );
OAI21X1 OAI21X1_434 ( .A(_1019__bF_buf3), .B(_1373_), .C(_1372_), .Y(_1374_) );
OAI21X1 OAI21X1_435 ( .A(_1067_), .B(_1250__bF_buf2), .C(_608_), .Y(_609_) );
OAI21X1 OAI21X1_436 ( .A(_1250__bF_buf2), .B(_1070_), .C(_608_), .Y(_611_) );
OAI21X1 OAI21X1_437 ( .A(_1250__bF_buf1), .B(_1073_), .C(_608_), .Y(_613_) );
OAI21X1 OAI21X1_438 ( .A(_982__bF_buf5), .B(_983__bF_buf4), .C(PC_STACK_4__2_), .Y(_615_) );
OAI21X1 OAI21X1_439 ( .A(_1142_), .B(_1250__bF_buf3), .C(_615_), .Y(_616_) );
OAI21X1 OAI21X1_440 ( .A(_1250__bF_buf3), .B(_1145_), .C(_615_), .Y(_618_) );
OAI21X1 OAI21X1_441 ( .A(_1250__bF_buf3), .B(_1148_), .C(_615_), .Y(_620_) );
OAI21X1 OAI21X1_442 ( .A(_982__bF_buf6), .B(_983__bF_buf3), .C(PC_STACK_4__3_), .Y(_622_) );
OAI21X1 OAI21X1_443 ( .A(_1182_), .B(_1250__bF_buf1), .C(_622_), .Y(_623_) );
OAI21X1 OAI21X1_444 ( .A(_1250__bF_buf1), .B(_1185_), .C(_622_), .Y(_625_) );
OAI21X1 OAI21X1_445 ( .A(_999__bF_buf5), .B(_982__bF_buf0), .C(PC_STACK_6__1_), .Y(_1064_) );
OAI21X1 OAI21X1_446 ( .A(_1371_), .B(_1301__bF_buf5), .C(_1375_), .Y(_12__9_) );
OAI21X1 OAI21X1_447 ( .A(_1250__bF_buf1), .B(_1188_), .C(_622_), .Y(_627_) );
OAI21X1 OAI21X1_448 ( .A(_982__bF_buf5), .B(_983__bF_buf4), .C(PC_STACK_4__4_), .Y(_629_) );
OAI21X1 OAI21X1_449 ( .A(_1214_), .B(_1250__bF_buf3), .C(_629_), .Y(_630_) );
OAI21X1 OAI21X1_450 ( .A(_1250__bF_buf3), .B(_1217_), .C(_629_), .Y(_632_) );
OAI21X1 OAI21X1_451 ( .A(_1250__bF_buf3), .B(_1220_), .C(_629_), .Y(_634_) );
OAI21X1 OAI21X1_452 ( .A(_982__bF_buf1), .B(_983__bF_buf5), .C(PC_STACK_4__5_), .Y(_636_) );
OAI21X1 OAI21X1_453 ( .A(_1239_), .B(_1250__bF_buf2), .C(_636_), .Y(_637_) );
OAI21X1 OAI21X1_454 ( .A(_1250__bF_buf4), .B(_1242_), .C(_636_), .Y(_639_) );
OAI21X1 OAI21X1_455 ( .A(_1250__bF_buf4), .B(_1245_), .C(_636_), .Y(_641_) );
OAI21X1 OAI21X1_456 ( .A(_982__bF_buf4), .B(_983__bF_buf0), .C(PC_STACK_4__6_), .Y(_643_) );
OAI21X1 OAI21X1_457 ( .A(_983__bF_buf4), .B(_991__bF_buf1), .C(PC_STACK_12__0_), .Y(_1376_) );
OAI21X1 OAI21X1_458 ( .A(_645_), .B(_644_), .C(_1030__bF_buf5), .Y(_646_) );
OAI21X1 OAI21X1_459 ( .A(_1250__bF_buf0), .B(_1497_), .C(_643_), .Y(_648_) );
OAI21X1 OAI21X1_460 ( .A(_1249_), .B(_984_), .C(_649_), .Y(_650_) );
OAI21X1 OAI21X1_461 ( .A(_1304_), .B(rst_bF_buf3), .C(_984_), .Y(_652_) );
OAI21X1 OAI21X1_462 ( .A(PC_STACK_4__7_), .B(_984_), .C(_652_), .Y(_653_) );
OAI21X1 OAI21X1_463 ( .A(_982__bF_buf2), .B(_983__bF_buf0), .C(PC_STACK_4__7_), .Y(_654_) );
OAI21X1 OAI21X1_464 ( .A(_1250__bF_buf0), .B(_1504_), .C(_654_), .Y(_655_) );
OAI21X1 OAI21X1_465 ( .A(_658_), .B(_1311__bF_buf1), .C(_656_), .Y(_659_) );
OAI21X1 OAI21X1_466 ( .A(_653_), .B(_1301__bF_buf2), .C(_660_), .Y(_10__7_) );
OAI21X1 OAI21X1_467 ( .A(_982__bF_buf1), .B(_983__bF_buf5), .C(_1332_), .Y(_661_) );
OAI21X1 OAI21X1_468 ( .A(_1032_), .B(_1117__bF_buf2), .C(_1376_), .Y(_1377_) );
OAI21X1 OAI21X1_469 ( .A(_1343_), .B(_1250__bF_buf4), .C(_661_), .Y(_662_) );
OAI21X1 OAI21X1_470 ( .A(_982__bF_buf1), .B(_983__bF_buf5), .C(PC_STACK_4__8_), .Y(_663_) );
OAI21X1 OAI21X1_471 ( .A(_1250__bF_buf4), .B(_1345_), .C(_663_), .Y(_664_) );
OAI21X1 OAI21X1_472 ( .A(_1250__bF_buf0), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_665_) );
OAI21X1 OAI21X1_473 ( .A(_662_), .B(_1301__bF_buf0), .C(_667_), .Y(_10__8_) );
OAI21X1 OAI21X1_474 ( .A(_982__bF_buf1), .B(_983__bF_buf5), .C(_1356_), .Y(_668_) );
OAI21X1 OAI21X1_475 ( .A(_1369_), .B(_1250__bF_buf0), .C(_668_), .Y(_669_) );
OAI21X1 OAI21X1_476 ( .A(_982__bF_buf1), .B(_983__bF_buf5), .C(PC_STACK_4__9_), .Y(_670_) );
OAI21X1 OAI21X1_477 ( .A(_1250__bF_buf4), .B(_1373_), .C(_670_), .Y(_671_) );
OAI21X1 OAI21X1_478 ( .A(_669_), .B(_1301__bF_buf0), .C(_672_), .Y(_10__9_) );
OAI21X1 OAI21X1_479 ( .A(_1035_), .B(_1117__bF_buf2), .C(_1376_), .Y(_1379_) );
OAI21X1 OAI21X1_480 ( .A(_989__bF_buf0), .B(_1002__bF_buf4), .C(PC_STACK_3__0_), .Y(_673_) );
OAI21X1 OAI21X1_481 ( .A(_1032_), .B(_1013__bF_buf4), .C(_673_), .Y(_674_) );
OAI21X1 OAI21X1_482 ( .A(_1035_), .B(_1013__bF_buf4), .C(_673_), .Y(_676_) );
OAI21X1 OAI21X1_483 ( .A(_1013__bF_buf4), .B(_1043_), .C(_673_), .Y(_678_) );
OAI21X1 OAI21X1_484 ( .A(_989__bF_buf0), .B(_1002__bF_buf4), .C(PC_STACK_3__1_), .Y(_680_) );
OAI21X1 OAI21X1_485 ( .A(_1067_), .B(_1013__bF_buf1), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_486 ( .A(_1013__bF_buf1), .B(_1070_), .C(_680_), .Y(_683_) );
OAI21X1 OAI21X1_487 ( .A(_1073_), .B(_1013__bF_buf1), .C(_680_), .Y(_685_) );
OAI21X1 OAI21X1_488 ( .A(_989__bF_buf2), .B(_1002__bF_buf2), .C(PC_STACK_3__2_), .Y(_687_) );
OAI21X1 OAI21X1_489 ( .A(_1142_), .B(_1013__bF_buf0), .C(_687_), .Y(_688_) );
OAI21X1 OAI21X1_490 ( .A(_1117__bF_buf2), .B(_1043_), .C(_1376_), .Y(_1381_) );
OAI21X1 OAI21X1_491 ( .A(_1013__bF_buf0), .B(_1145_), .C(_687_), .Y(_690_) );
OAI21X1 OAI21X1_492 ( .A(_1148_), .B(_1013__bF_buf0), .C(_687_), .Y(_692_) );
OAI21X1 OAI21X1_493 ( .A(_989__bF_buf0), .B(_1002__bF_buf4), .C(PC_STACK_3__3_), .Y(_694_) );
OAI21X1 OAI21X1_494 ( .A(_1182_), .B(_1013__bF_buf1), .C(_694_), .Y(_695_) );
OAI21X1 OAI21X1_495 ( .A(_1185_), .B(_1013__bF_buf1), .C(_694_), .Y(_697_) );
OAI21X1 OAI21X1_496 ( .A(_1013__bF_buf2), .B(_1188_), .C(_694_), .Y(_699_) );
OAI21X1 OAI21X1_497 ( .A(_989__bF_buf5), .B(_1002__bF_buf4), .C(PC_STACK_3__4_), .Y(_701_) );
OAI21X1 OAI21X1_498 ( .A(_1214_), .B(_1013__bF_buf2), .C(_701_), .Y(_702_) );
OAI21X1 OAI21X1_499 ( .A(_1217_), .B(_1013__bF_buf2), .C(_701_), .Y(_704_) );
OAI21X1 OAI21X1_500 ( .A(_1013__bF_buf2), .B(_1220_), .C(_701_), .Y(_706_) );
OAI21X1 OAI21X1_501 ( .A(_983__bF_buf6), .B(_991__bF_buf5), .C(PC_STACK_12__1_), .Y(_1383_) );
OAI21X1 OAI21X1_502 ( .A(_989__bF_buf0), .B(_1002__bF_buf4), .C(PC_STACK_3__5_), .Y(_708_) );
OAI21X1 OAI21X1_503 ( .A(_1239_), .B(_1013__bF_buf1), .C(_708_), .Y(_709_) );
OAI21X1 OAI21X1_504 ( .A(_1242_), .B(_1013__bF_buf4), .C(_708_), .Y(_711_) );
OAI21X1 OAI21X1_505 ( .A(_1013__bF_buf4), .B(_1245_), .C(_708_), .Y(_713_) );
OAI21X1 OAI21X1_506 ( .A(_989__bF_buf3), .B(_1002__bF_buf3), .C(PC_STACK_3__6_), .Y(_715_) );
OAI21X1 OAI21X1_507 ( .A(_717_), .B(_716_), .C(_1030__bF_buf5), .Y(_718_) );
OAI21X1 OAI21X1_508 ( .A(_1497_), .B(_1013__bF_buf3), .C(_715_), .Y(_720_) );
OAI21X1 OAI21X1_509 ( .A(_1304_), .B(rst_bF_buf0), .C(_1196_), .Y(_724_) );
OAI21X1 OAI21X1_510 ( .A(PC_STACK_3__7_), .B(_1196_), .C(_724_), .Y(_725_) );
OAI21X1 OAI21X1_511 ( .A(_989__bF_buf3), .B(_1002__bF_buf3), .C(PC_STACK_3__7_), .Y(_726_) );
OAI21X1 OAI21X1_512 ( .A(_1067_), .B(_1117__bF_buf1), .C(_1383_), .Y(_1384_) );
OAI21X1 OAI21X1_513 ( .A(_1504_), .B(_1013__bF_buf3), .C(_726_), .Y(_727_) );
OAI21X1 OAI21X1_514 ( .A(_730_), .B(_1311__bF_buf1), .C(_728_), .Y(_731_) );
OAI21X1 OAI21X1_515 ( .A(_725_), .B(_1301__bF_buf6), .C(_732_), .Y(_9__7_) );
OAI21X1 OAI21X1_516 ( .A(_989__bF_buf4), .B(_1002__bF_buf3), .C(PC_STACK_3__8_), .Y(_733_) );
OAI21X1 OAI21X1_517 ( .A(_1013__bF_buf3), .B(_1345_), .C(_733_), .Y(_736_) );
OAI21X1 OAI21X1_518 ( .A(_1013__bF_buf3), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_737_) );
OAI21X1 OAI21X1_519 ( .A(_735_), .B(_1301__bF_buf0), .C(_739_), .Y(_9__8_) );
OAI21X1 OAI21X1_520 ( .A(_1369_), .B(_1013__bF_buf2), .C(_740_), .Y(_741_) );
OAI21X1 OAI21X1_521 ( .A(_989__bF_buf5), .B(_1002__bF_buf5), .C(PC_STACK_3__9_), .Y(_742_) );
OAI21X1 OAI21X1_522 ( .A(_1013__bF_buf3), .B(_1373_), .C(_742_), .Y(_743_) );
OAI21X1 OAI21X1_523 ( .A(_1117__bF_buf1), .B(_1070_), .C(_1383_), .Y(_1386_) );
OAI21X1 OAI21X1_524 ( .A(_741_), .B(_1301__bF_buf5), .C(_744_), .Y(_9__9_) );
OAI21X1 OAI21X1_525 ( .A(_999__bF_buf3), .B(_989__bF_buf0), .C(PC_STACK_2__0_), .Y(_745_) );
OAI21X1 OAI21X1_526 ( .A(_1032_), .B(_1011__bF_buf4), .C(_745_), .Y(_746_) );
OAI21X1 OAI21X1_527 ( .A(_1035_), .B(_1011__bF_buf4), .C(_745_), .Y(_748_) );
OAI21X1 OAI21X1_528 ( .A(_1011__bF_buf2), .B(_1043_), .C(_745_), .Y(_750_) );
OAI21X1 OAI21X1_529 ( .A(_999__bF_buf3), .B(_989__bF_buf1), .C(PC_STACK_2__1_), .Y(_752_) );
OAI21X1 OAI21X1_530 ( .A(_1067_), .B(_1011__bF_buf3), .C(_752_), .Y(_753_) );
OAI21X1 OAI21X1_531 ( .A(_1011__bF_buf3), .B(_1070_), .C(_752_), .Y(_755_) );
OAI21X1 OAI21X1_532 ( .A(_1073_), .B(_1011__bF_buf3), .C(_752_), .Y(_757_) );
OAI21X1 OAI21X1_533 ( .A(_999__bF_buf3), .B(_989__bF_buf2), .C(PC_STACK_2__2_), .Y(_759_) );
OAI21X1 OAI21X1_534 ( .A(_1073_), .B(_1117__bF_buf1), .C(_1383_), .Y(_1388_) );
OAI21X1 OAI21X1_535 ( .A(_1142_), .B(_1011__bF_buf0), .C(_759_), .Y(_760_) );
OAI21X1 OAI21X1_536 ( .A(_1011__bF_buf0), .B(_1145_), .C(_759_), .Y(_762_) );
OAI21X1 OAI21X1_537 ( .A(_1148_), .B(_1011__bF_buf0), .C(_759_), .Y(_764_) );
OAI21X1 OAI21X1_538 ( .A(_999__bF_buf3), .B(_989__bF_buf1), .C(PC_STACK_2__3_), .Y(_766_) );
OAI21X1 OAI21X1_539 ( .A(_1182_), .B(_1011__bF_buf3), .C(_766_), .Y(_767_) );
OAI21X1 OAI21X1_540 ( .A(_1185_), .B(_1011__bF_buf3), .C(_766_), .Y(_769_) );
OAI21X1 OAI21X1_541 ( .A(_1011__bF_buf3), .B(_1188_), .C(_766_), .Y(_771_) );
OAI21X1 OAI21X1_542 ( .A(_999__bF_buf3), .B(_989__bF_buf1), .C(PC_STACK_2__4_), .Y(_773_) );
OAI21X1 OAI21X1_543 ( .A(_1214_), .B(_1011__bF_buf4), .C(_773_), .Y(_774_) );
OAI21X1 OAI21X1_544 ( .A(_1217_), .B(_1011__bF_buf4), .C(_773_), .Y(_776_) );
OAI21X1 OAI21X1_545 ( .A(_983__bF_buf6), .B(_991__bF_buf5), .C(PC_STACK_12__2_), .Y(_1390_) );
OAI21X1 OAI21X1_546 ( .A(_1011__bF_buf4), .B(_1220_), .C(_773_), .Y(_778_) );
OAI21X1 OAI21X1_547 ( .A(PC_STACK_2__5_), .B(_1191_), .C(_780_), .Y(_781_) );
OAI21X1 OAI21X1_548 ( .A(_999__bF_buf5), .B(_989__bF_buf5), .C(PC_STACK_2__5_), .Y(_782_) );
OAI21X1 OAI21X1_549 ( .A(_1242_), .B(_1011__bF_buf2), .C(_782_), .Y(_783_) );
OAI21X1 OAI21X1_550 ( .A(_1011__bF_buf2), .B(_1245_), .C(_782_), .Y(_785_) );
OAI21X1 OAI21X1_551 ( .A(_781_), .B(_1301__bF_buf5), .C(_788_), .Y(_8__5_) );
OAI21X1 OAI21X1_552 ( .A(_999__bF_buf2), .B(_989__bF_buf3), .C(PC_STACK_2__6_), .Y(_789_) );
OAI21X1 OAI21X1_553 ( .A(_791_), .B(_790_), .C(_1030__bF_buf7), .Y(_792_) );
OAI21X1 OAI21X1_554 ( .A(_1497_), .B(_1011__bF_buf1), .C(_789_), .Y(_794_) );
OAI21X1 OAI21X1_555 ( .A(_1248_), .B(_1191_), .C(_795_), .Y(_796_) );
OAI21X1 OAI21X1_556 ( .A(_1543__0_), .B(_1543__1_), .C(_1042_), .Y(_1066_) );
OAI21X1 OAI21X1_557 ( .A(_1142_), .B(_1117__bF_buf0), .C(_1390_), .Y(_1391_) );
OAI21X1 OAI21X1_558 ( .A(_1304_), .B(rst_bF_buf3), .C(_1191_), .Y(_798_) );
OAI21X1 OAI21X1_559 ( .A(PC_STACK_2__7_), .B(_1191_), .C(_798_), .Y(_799_) );
OAI21X1 OAI21X1_560 ( .A(_999__bF_buf2), .B(_989__bF_buf4), .C(PC_STACK_2__7_), .Y(_800_) );
OAI21X1 OAI21X1_561 ( .A(_1504_), .B(_1011__bF_buf1), .C(_800_), .Y(_801_) );
OAI21X1 OAI21X1_562 ( .A(_804_), .B(_1311__bF_buf2), .C(_802_), .Y(_805_) );
OAI21X1 OAI21X1_563 ( .A(_799_), .B(_1301__bF_buf2), .C(_806_), .Y(_8__7_) );
OAI21X1 OAI21X1_564 ( .A(_999__bF_buf2), .B(_989__bF_buf4), .C(_1328_), .Y(_807_) );
OAI21X1 OAI21X1_565 ( .A(_1343_), .B(_1011__bF_buf1), .C(_807_), .Y(_808_) );
OAI21X1 OAI21X1_566 ( .A(_999__bF_buf2), .B(_989__bF_buf4), .C(PC_STACK_2__8_), .Y(_809_) );
OAI21X1 OAI21X1_567 ( .A(_1011__bF_buf1), .B(_1345_), .C(_809_), .Y(_810_) );
OAI21X1 OAI21X1_568 ( .A(_1117__bF_buf0), .B(_1145_), .C(_1390_), .Y(_1393_) );
OAI21X1 OAI21X1_569 ( .A(_808_), .B(_1301__bF_buf0), .C(_812_), .Y(_8__8_) );
OAI21X1 OAI21X1_570 ( .A(_1369_), .B(_1011__bF_buf2), .C(_813_), .Y(_814_) );
OAI21X1 OAI21X1_571 ( .A(_999__bF_buf5), .B(_989__bF_buf5), .C(PC_STACK_2__9_), .Y(_815_) );
OAI21X1 OAI21X1_572 ( .A(_1011__bF_buf2), .B(_1373_), .C(_815_), .Y(_816_) );
OAI21X1 OAI21X1_573 ( .A(_814_), .B(_1301__bF_buf5), .C(_817_), .Y(_8__9_) );
OAI21X1 OAI21X1_574 ( .A(_986__bF_buf2), .B(_989__bF_buf0), .C(PC_STACK_1__0_), .Y(_818_) );
OAI21X1 OAI21X1_575 ( .A(_1032_), .B(_1116__bF_buf2), .C(_818_), .Y(_819_) );
OAI21X1 OAI21X1_576 ( .A(_1035_), .B(_1116__bF_buf2), .C(_818_), .Y(_821_) );
OAI21X1 OAI21X1_577 ( .A(_1116__bF_buf2), .B(_1043_), .C(_818_), .Y(_823_) );
OAI21X1 OAI21X1_578 ( .A(_986__bF_buf2), .B(_989__bF_buf3), .C(PC_STACK_1__1_), .Y(_825_) );
OAI21X1 OAI21X1_579 ( .A(_1148_), .B(_1117__bF_buf4), .C(_1390_), .Y(_1395_) );
OAI21X1 OAI21X1_580 ( .A(_1067_), .B(_1116__bF_buf0), .C(_825_), .Y(_826_) );
OAI21X1 OAI21X1_581 ( .A(_1116__bF_buf2), .B(_1070_), .C(_825_), .Y(_828_) );
OAI21X1 OAI21X1_582 ( .A(_1073_), .B(_1116__bF_buf2), .C(_825_), .Y(_830_) );
OAI21X1 OAI21X1_583 ( .A(_986__bF_buf2), .B(_989__bF_buf0), .C(PC_STACK_1__2_), .Y(_832_) );
OAI21X1 OAI21X1_584 ( .A(_1142_), .B(_1116__bF_buf4), .C(_832_), .Y(_833_) );
OAI21X1 OAI21X1_585 ( .A(_1116__bF_buf4), .B(_1145_), .C(_832_), .Y(_835_) );
OAI21X1 OAI21X1_586 ( .A(_1148_), .B(_1116__bF_buf4), .C(_832_), .Y(_837_) );
OAI21X1 OAI21X1_587 ( .A(_986__bF_buf3), .B(_989__bF_buf5), .C(PC_STACK_1__3_), .Y(_839_) );
OAI21X1 OAI21X1_588 ( .A(_1182_), .B(_1116__bF_buf0), .C(_839_), .Y(_840_) );
OAI21X1 OAI21X1_589 ( .A(_1185_), .B(_1116__bF_buf0), .C(_839_), .Y(_842_) );
OAI21X1 OAI21X1_590 ( .A(_983__bF_buf4), .B(_991__bF_buf1), .C(PC_STACK_12__3_), .Y(_1397_) );
OAI21X1 OAI21X1_591 ( .A(_1116__bF_buf0), .B(_1188_), .C(_839_), .Y(_844_) );
OAI21X1 OAI21X1_592 ( .A(_986__bF_buf3), .B(_989__bF_buf5), .C(PC_STACK_1__4_), .Y(_846_) );
OAI21X1 OAI21X1_593 ( .A(_1214_), .B(_1116__bF_buf3), .C(_846_), .Y(_847_) );
OAI21X1 OAI21X1_594 ( .A(_1217_), .B(_1116__bF_buf3), .C(_846_), .Y(_849_) );
OAI21X1 OAI21X1_595 ( .A(_1116__bF_buf3), .B(_1220_), .C(_846_), .Y(_851_) );
OAI21X1 OAI21X1_596 ( .A(PC_STACK_1__5_), .B(_990__bF_buf0), .C(_853_), .Y(_854_) );
OAI21X1 OAI21X1_597 ( .A(_986__bF_buf3), .B(_989__bF_buf5), .C(PC_STACK_1__5_), .Y(_855_) );
OAI21X1 OAI21X1_598 ( .A(_1242_), .B(_1116__bF_buf0), .C(_855_), .Y(_856_) );
OAI21X1 OAI21X1_599 ( .A(_1116__bF_buf3), .B(_1245_), .C(_855_), .Y(_858_) );
OAI21X1 OAI21X1_600 ( .A(_854_), .B(_1301__bF_buf5), .C(_861_), .Y(_7__5_) );
OAI21X1 OAI21X1_601 ( .A(_1182_), .B(_1117__bF_buf0), .C(_1397_), .Y(_1398_) );
OAI21X1 OAI21X1_602 ( .A(_986__bF_buf2), .B(_989__bF_buf3), .C(PC_STACK_1__6_), .Y(_862_) );
OAI21X1 OAI21X1_603 ( .A(_864_), .B(_863_), .C(_1030__bF_buf5), .Y(_865_) );
OAI21X1 OAI21X1_604 ( .A(_1497_), .B(_1116__bF_buf1), .C(_862_), .Y(_867_) );
OAI21X1 OAI21X1_605 ( .A(_1304_), .B(rst_bF_buf3), .C(_990__bF_buf2), .Y(_871_) );
OAI21X1 OAI21X1_606 ( .A(PC_STACK_1__7_), .B(_990__bF_buf2), .C(_871_), .Y(_872_) );
OAI21X1 OAI21X1_607 ( .A(_986__bF_buf3), .B(_989__bF_buf4), .C(PC_STACK_1__7_), .Y(_873_) );
OAI21X1 OAI21X1_608 ( .A(_1504_), .B(_1116__bF_buf1), .C(_873_), .Y(_874_) );
OAI21X1 OAI21X1_609 ( .A(_877_), .B(_1311__bF_buf2), .C(_875_), .Y(_878_) );
OAI21X1 OAI21X1_610 ( .A(_872_), .B(_1301__bF_buf2), .C(_879_), .Y(_7__7_) );
OAI21X1 OAI21X1_611 ( .A(_986__bF_buf3), .B(_989__bF_buf4), .C(PC_STACK_1__8_), .Y(_880_) );
OAI21X1 OAI21X1_612 ( .A(_1185_), .B(_1117__bF_buf0), .C(_1397_), .Y(_1400_) );
OAI21X1 OAI21X1_613 ( .A(_1116__bF_buf1), .B(_1345_), .C(_880_), .Y(_883_) );
OAI21X1 OAI21X1_614 ( .A(_882_), .B(_1301__bF_buf0), .C(_885_), .Y(_7__8_) );
OAI21X1 OAI21X1_615 ( .A(_1369_), .B(_1116__bF_buf1), .C(_886_), .Y(_887_) );
OAI21X1 OAI21X1_616 ( .A(_986__bF_buf3), .B(_989__bF_buf4), .C(PC_STACK_1__9_), .Y(_888_) );
OAI21X1 OAI21X1_617 ( .A(_1116__bF_buf1), .B(_1373_), .C(_888_), .Y(_889_) );
OAI21X1 OAI21X1_618 ( .A(_887_), .B(_1301__bF_buf0), .C(_890_), .Y(_7__9_) );
OAI21X1 OAI21X1_619 ( .A(_989__bF_buf2), .B(_983__bF_buf1), .C(PC_STACK_0__0_), .Y(_891_) );
OAI21X1 OAI21X1_620 ( .A(_1032_), .B(_1099__bF_buf3), .C(_891_), .Y(_892_) );
OAI21X1 OAI21X1_621 ( .A(_1035_), .B(_1099__bF_buf3), .C(_891_), .Y(_894_) );
OAI21X1 OAI21X1_622 ( .A(_1099__bF_buf0), .B(_1043_), .C(_891_), .Y(_896_) );
OAI21X1 OAI21X1_623 ( .A(_1117__bF_buf0), .B(_1188_), .C(_1397_), .Y(_1402_) );
OAI21X1 OAI21X1_624 ( .A(_989__bF_buf2), .B(_983__bF_buf1), .C(PC_STACK_0__1_), .Y(_898_) );
OAI21X1 OAI21X1_625 ( .A(_1067_), .B(_1099__bF_buf3), .C(_898_), .Y(_899_) );
OAI21X1 OAI21X1_626 ( .A(_1099__bF_buf0), .B(_1070_), .C(_898_), .Y(_901_) );
OAI21X1 OAI21X1_627 ( .A(_1073_), .B(_1099__bF_buf0), .C(_898_), .Y(_903_) );
OAI21X1 OAI21X1_628 ( .A(_989__bF_buf2), .B(_983__bF_buf1), .C(PC_STACK_0__2_), .Y(_905_) );
OAI21X1 OAI21X1_629 ( .A(_1142_), .B(_1099__bF_buf2), .C(_905_), .Y(_906_) );
OAI21X1 OAI21X1_630 ( .A(_1099__bF_buf2), .B(_1145_), .C(_905_), .Y(_908_) );
OAI21X1 OAI21X1_631 ( .A(_1148_), .B(_1099__bF_buf2), .C(_905_), .Y(_910_) );
OAI21X1 OAI21X1_632 ( .A(_989__bF_buf2), .B(_983__bF_buf1), .C(PC_STACK_0__3_), .Y(_912_) );
OAI21X1 OAI21X1_633 ( .A(_1182_), .B(_1099__bF_buf1), .C(_912_), .Y(_913_) );
OAI21X1 OAI21X1_634 ( .A(_983__bF_buf5), .B(_991__bF_buf6), .C(PC_STACK_12__4_), .Y(_1404_) );
OAI21X1 OAI21X1_635 ( .A(_1185_), .B(_1099__bF_buf1), .C(_912_), .Y(_915_) );
OAI21X1 OAI21X1_636 ( .A(_1099__bF_buf1), .B(_1188_), .C(_912_), .Y(_917_) );
OAI21X1 OAI21X1_637 ( .A(_989__bF_buf2), .B(_983__bF_buf1), .C(PC_STACK_0__4_), .Y(_919_) );
OAI21X1 OAI21X1_638 ( .A(_1214_), .B(_1099__bF_buf1), .C(_919_), .Y(_920_) );
OAI21X1 OAI21X1_639 ( .A(_1217_), .B(_1099__bF_buf1), .C(_919_), .Y(_922_) );
OAI21X1 OAI21X1_640 ( .A(_1099__bF_buf0), .B(_1220_), .C(_919_), .Y(_924_) );
OAI21X1 OAI21X1_641 ( .A(_989__bF_buf2), .B(_983__bF_buf1), .C(PC_STACK_0__5_), .Y(_926_) );
OAI21X1 OAI21X1_642 ( .A(_1239_), .B(_1099__bF_buf3), .C(_926_), .Y(_927_) );
OAI21X1 OAI21X1_643 ( .A(_1242_), .B(_1099__bF_buf3), .C(_926_), .Y(_929_) );
OAI21X1 OAI21X1_644 ( .A(_1099__bF_buf3), .B(_1245_), .C(_926_), .Y(_931_) );
OAI21X1 OAI21X1_645 ( .A(_1214_), .B(_1117__bF_buf3), .C(_1404_), .Y(_1405_) );
OAI21X1 OAI21X1_646 ( .A(_989__bF_buf3), .B(_983__bF_buf6), .C(PC_STACK_0__6_), .Y(_933_) );
OAI21X1 OAI21X1_647 ( .A(_935_), .B(_934_), .C(_1030__bF_buf5), .Y(_936_) );
OAI21X1 OAI21X1_648 ( .A(_1497_), .B(_1099__bF_buf4), .C(_933_), .Y(_938_) );
OAI21X1 OAI21X1_649 ( .A(_1304_), .B(rst_bF_buf2), .C(_1025_), .Y(_942_) );
OAI21X1 OAI21X1_650 ( .A(PC_STACK_0__7_), .B(_1025_), .C(_942_), .Y(_943_) );
OAI21X1 OAI21X1_651 ( .A(_989__bF_buf3), .B(_983__bF_buf0), .C(PC_STACK_0__7_), .Y(_944_) );
OAI21X1 OAI21X1_652 ( .A(_1504_), .B(_1099__bF_buf4), .C(_944_), .Y(_945_) );
OAI21X1 OAI21X1_653 ( .A(_948_), .B(_1311__bF_buf1), .C(_946_), .Y(_949_) );
OAI21X1 OAI21X1_654 ( .A(_943_), .B(_1301__bF_buf2), .C(_950_), .Y(_0__7_) );
OAI21X1 OAI21X1_655 ( .A(_989__bF_buf1), .B(_983__bF_buf3), .C(_1333_), .Y(_951_) );
OAI21X1 OAI21X1_656 ( .A(_1217_), .B(_1117__bF_buf3), .C(_1404_), .Y(_1407_) );
OAI21X1 OAI21X1_657 ( .A(_1343_), .B(_1099__bF_buf2), .C(_951_), .Y(_952_) );
OAI21X1 OAI21X1_658 ( .A(_989__bF_buf1), .B(_983__bF_buf3), .C(PC_STACK_0__8_), .Y(_953_) );
OAI21X1 OAI21X1_659 ( .A(_1099__bF_buf2), .B(_1345_), .C(_953_), .Y(_954_) );
OAI21X1 OAI21X1_660 ( .A(_952_), .B(_1301__bF_buf1), .C(_956_), .Y(_0__8_) );
OAI21X1 OAI21X1_661 ( .A(_989__bF_buf1), .B(_983__bF_buf4), .C(_1349_), .Y(_957_) );
OAI21X1 OAI21X1_662 ( .A(_1369_), .B(_1099__bF_buf4), .C(_957_), .Y(_958_) );
OAI21X1 OAI21X1_663 ( .A(_989__bF_buf1), .B(_983__bF_buf3), .C(PC_STACK_0__9_), .Y(_959_) );
OAI21X1 OAI21X1_664 ( .A(_1099__bF_buf2), .B(_1373_), .C(_959_), .Y(_960_) );
OAI21X1 OAI21X1_665 ( .A(_958_), .B(_1301__bF_buf1), .C(_961_), .Y(_0__9_) );
OAI21X1 OAI21X1_666 ( .A(_1067_), .B(_1019__bF_buf1), .C(_1064_), .Y(_1068_) );
OAI21X1 OAI21X1_667 ( .A(_1117__bF_buf3), .B(_1220_), .C(_1404_), .Y(_1409_) );
OAI21X1 OAI21X1_668 ( .A(_983__bF_buf5), .B(_991__bF_buf6), .C(PC_STACK_12__5_), .Y(_1411_) );
OAI21X1 OAI21X1_669 ( .A(_1239_), .B(_1117__bF_buf1), .C(_1411_), .Y(_1412_) );
OAI21X1 OAI21X1_670 ( .A(_1242_), .B(_1117__bF_buf3), .C(_1411_), .Y(_1414_) );
OAI21X1 OAI21X1_671 ( .A(_1117__bF_buf1), .B(_1245_), .C(_1411_), .Y(_1416_) );
OAI21X1 OAI21X1_672 ( .A(_983__bF_buf0), .B(_991__bF_buf6), .C(PC_STACK_12__6_), .Y(_1418_) );
OAI21X1 OAI21X1_673 ( .A(_1420_), .B(_1419_), .C(_1030__bF_buf7), .Y(_1421_) );
OAI21X1 OAI21X1_674 ( .A(_1304_), .B(rst_bF_buf3), .C(_992__bF_buf3), .Y(_1428_) );
OAI21X1 OAI21X1_675 ( .A(PC_STACK_12__7_), .B(_992__bF_buf3), .C(_1428_), .Y(_1429_) );
OAI21X1 OAI21X1_676 ( .A(_983__bF_buf0), .B(_991__bF_buf6), .C(PC_STACK_12__7_), .Y(_1430_) );
OAI21X1 OAI21X1_677 ( .A(_1019__bF_buf1), .B(_1070_), .C(_1064_), .Y(_1071_) );
OAI21X1 OAI21X1_678 ( .A(_1435_), .B(_1311__bF_buf2), .C(_1433_), .Y(_1436_) );
OAI21X1 OAI21X1_679 ( .A(_1429_), .B(_1301__bF_buf2), .C(_1437_), .Y(_3__7_) );
OAI21X1 OAI21X1_680 ( .A(_983__bF_buf6), .B(_991__bF_buf0), .C(_1321_), .Y(_1438_) );
OAI21X1 OAI21X1_681 ( .A(_1343_), .B(_1117__bF_buf4), .C(_1438_), .Y(_1439_) );
OAI21X1 OAI21X1_682 ( .A(_983__bF_buf6), .B(_991__bF_buf0), .C(PC_STACK_12__8_), .Y(_1440_) );
OAI21X1 OAI21X1_683 ( .A(_1117__bF_buf4), .B(_1345_), .C(_1440_), .Y(_1441_) );
OAI21X1 OAI21X1_684 ( .A(_1117__bF_buf4), .B(CORE_PC_ctrl[0]), .C(INTERRUPT_flag), .Y(_1442_) );
OAI21X1 OAI21X1_685 ( .A(_1439_), .B(_1301__bF_buf6), .C(_1444_), .Y(_3__8_) );
OAI21X1 OAI21X1_686 ( .A(_1369_), .B(_1117__bF_buf3), .C(_1445_), .Y(_1446_) );
OAI21X1 OAI21X1_687 ( .A(_983__bF_buf6), .B(_991__bF_buf6), .C(PC_STACK_12__9_), .Y(_1447_) );
OAI21X1 OAI21X1_688 ( .A(_1019__bF_buf1), .B(_1073_), .C(_1064_), .Y(_1074_) );
OAI21X1 OAI21X1_689 ( .A(_1117__bF_buf4), .B(_1373_), .C(_1447_), .Y(_1448_) );
OAI21X1 OAI21X1_690 ( .A(_1446_), .B(_1301__bF_buf2), .C(_1449_), .Y(_3__9_) );
OAI21X1 OAI21X1_691 ( .A(_986__bF_buf4), .B(_991__bF_buf5), .C(PC_STACK_13__0_), .Y(_1450_) );
OAI21X1 OAI21X1_692 ( .A(_1032_), .B(_1080__bF_buf3), .C(_1450_), .Y(_1451_) );
OAI21X1 OAI21X1_693 ( .A(_1035_), .B(_1080__bF_buf2), .C(_1450_), .Y(_1453_) );
OAI21X1 OAI21X1_694 ( .A(_1080__bF_buf2), .B(_1043_), .C(_1450_), .Y(_1455_) );
OAI21X1 OAI21X1_695 ( .A(_986__bF_buf5), .B(_991__bF_buf2), .C(PC_STACK_13__1_), .Y(_1457_) );
OAI21X1 OAI21X1_696 ( .A(_1067_), .B(_1080__bF_buf1), .C(_1457_), .Y(_1458_) );
OAI21X1 OAI21X1_697 ( .A(_1080__bF_buf1), .B(_1070_), .C(_1457_), .Y(_1460_) );
OAI21X1 OAI21X1_698 ( .A(_1073_), .B(_1080__bF_buf1), .C(_1457_), .Y(_1462_) );
OAI22X1 OAI22X1_1 ( .A(_1013__bF_buf4), .B(_1009_), .C(_1011__bF_buf4), .D(_1008_), .Y(_1014_) );
OAI22X1 OAI22X1_2 ( .A(_1085__bF_buf0), .B(_1120_), .C(_1119_), .D(_1095__bF_buf1), .Y(_1121_) );
OAI22X1 OAI22X1_3 ( .A(_1080__bF_buf2), .B(_1125_), .C(_1124_), .D(_1109__bF_buf3), .Y(_1126_) );
OAI22X1 OAI22X1_4 ( .A(_1117__bF_buf2), .B(_1130_), .C(_1116__bF_buf4), .D(_1131_), .Y(_1132_) );
OAI22X1 OAI22X1_5 ( .A(_1085__bF_buf4), .B(_1134_), .C(_1133_), .D(_1095__bF_buf1), .Y(_1135_) );
OAI22X1 OAI22X1_6 ( .A(_1112_), .B(_1123_), .C(_1128_), .D(_1137_), .Y(_1138_) );
OAI22X1 OAI22X1_7 ( .A(_1152_), .B(_1011__bF_buf0), .C(_1080__bF_buf2), .D(_1151_), .Y(_1153_) );
OAI22X1 OAI22X1_8 ( .A(_1155_), .B(_1095__bF_buf0), .C(_1084__bF_buf2), .D(_1154_), .Y(_1156_) );
OAI22X1 OAI22X1_9 ( .A(_1161_), .B(_1085__bF_buf4), .C(_1109__bF_buf1), .D(_1162_), .Y(_1163_) );
OAI22X1 OAI22X1_10 ( .A(_1173_), .B(_1116__bF_buf3), .C(_1020__bF_buf0), .D(_1174_), .Y(_1175_) );
OAI22X1 OAI22X1_11 ( .A(_1200_), .B(_1085__bF_buf0), .C(_1201__bF_buf0), .D(_1199_), .Y(_1202_) );
OAI22X1 OAI22X1_12 ( .A(_1016_), .B(_1020__bF_buf2), .C(_1019__bF_buf1), .D(_1015_), .Y(_1021_) );
OAI22X1 OAI22X1_13 ( .A(_1203_), .B(_1095__bF_buf3), .C(_1080__bF_buf0), .D(_1204_), .Y(_1205_) );
OAI22X1 OAI22X1_14 ( .A(_1248_), .B(_1011__bF_buf1), .C(_1250__bF_buf0), .D(_1249_), .Y(_1251_) );
OAI22X1 OAI22X1_15 ( .A(_1109__bF_buf4), .B(_1253_), .C(_1252_), .D(_1084__bF_buf4), .Y(_1254_) );
OAI22X1 OAI22X1_16 ( .A(_1260_), .B(_1095__bF_buf4), .C(_1201__bF_buf2), .D(_1259_), .Y(_1261_) );
OAI22X1 OAI22X1_17 ( .A(_1262_), .B(_1085__bF_buf4), .C(_1080__bF_buf3), .D(_1263_), .Y(_1264_) );
OAI22X1 OAI22X1_18 ( .A(_1287_), .B(_1013__bF_buf3), .C(_1020__bF_buf4), .D(_1288_), .Y(_1289_) );
OAI22X1 OAI22X1_19 ( .A(_1321_), .B(_1117__bF_buf4), .C(_1080__bF_buf4), .D(_1320_), .Y(_1322_) );
OAI22X1 OAI22X1_20 ( .A(_1323_), .B(_1085__bF_buf3), .C(_1109__bF_buf4), .D(_1324_), .Y(_1325_) );
OAI22X1 OAI22X1_21 ( .A(_1328_), .B(_1011__bF_buf1), .C(_1020__bF_buf4), .D(_1329_), .Y(_1330_) );
OAI22X1 OAI22X1_22 ( .A(_1333_), .B(_1099__bF_buf4), .C(_1250__bF_buf4), .D(_1332_), .Y(_1334_) );
OAI22X1 OAI22X1_23 ( .A(_1013__bF_buf0), .B(_1055_), .C(_1011__bF_buf0), .D(_1054_), .Y(_1056_) );
OAI22X1 OAI22X1_24 ( .A(_1355_), .B(_1080__bF_buf2), .C(_1250__bF_buf1), .D(_1356_), .Y(_1357_) );
OAI22X1 OAI22X1_25 ( .A(_1058_), .B(_1020__bF_buf2), .C(_1019__bF_buf1), .D(_1057_), .Y(_1059_) );
OAI22X1 OAI22X1_26 ( .A(_1078_), .B(_1011__bF_buf0), .C(_1080__bF_buf3), .D(_1077_), .Y(_1081_) );
OAI22X1 OAI22X1_27 ( .A(_1083_), .B(_1085__bF_buf0), .C(_1084__bF_buf3), .D(_1082_), .Y(_1086_) );
OAI22X1 OAI22X1_28 ( .A(_1097_), .B(_1099__bF_buf0), .C(_1013__bF_buf0), .D(_1098_), .Y(_1100_) );
OAI22X1 OAI22X1_29 ( .A(_1080__bF_buf2), .B(_1108_), .C(_1107_), .D(_1109__bF_buf3), .Y(_1110_) );
OAI22X1 OAI22X1_30 ( .A(_1117__bF_buf2), .B(_1114_), .C(_1116__bF_buf4), .D(_1115_), .Y(_1118_) );
OR2X2 OR2X2_1 ( .A(PC_pointer_0_), .B(PC_pointer_1_), .Y(_983_) );
OR2X2 OR2X2_2 ( .A(_992__bF_buf2), .B(PC_STACK_12__9_), .Y(_1445_) );
OR2X2 OR2X2_3 ( .A(_1023_), .B(PC_STACK_14__9_), .Y(_65_) );
OR2X2 OR2X2_4 ( .A(_1003_), .B(PC_STACK_15__9_), .Y(_233_) );
OR2X2 OR2X2_5 ( .A(_997__bF_buf0), .B(PC_STACK_9__9_), .Y(_305_) );
OR2X2 OR2X2_6 ( .A(_1000__bF_buf2), .B(PC_STACK_10__9_), .Y(_377_) );
OR2X2 OR2X2_7 ( .A(_1004__bF_buf3), .B(PC_STACK_8__9_), .Y(_450_) );
OR2X2 OR2X2_8 ( .A(_1026_), .B(PC_STACK_11__9_), .Y(_522_) );
OR2X2 OR2X2_9 ( .A(_1196_), .B(PC_STACK_3__9_), .Y(_740_) );
OR2X2 OR2X2_10 ( .A(_1191_), .B(PC_STACK_2__9_), .Y(_813_) );
OR2X2 OR2X2_11 ( .A(_990__bF_buf3), .B(PC_STACK_1__9_), .Y(_886_) );
OR2X2 OR2X2_12 ( .A(PC_pointer_2_), .B(PC_pointer_3_), .Y(_989_) );
OR2X2 OR2X2_13 ( .A(_1543__0_), .B(rst_bF_buf2), .Y(_1032_) );
OR2X2 OR2X2_14 ( .A(_1066_), .B(_1065_), .Y(_1067_) );
OR2X2 OR2X2_15 ( .A(_1106_), .B(_1090_), .Y(_1543__2_) );
OR2X2 OR2X2_16 ( .A(_1177_), .B(_1160_), .Y(_1543__3_) );
OR2X2 OR2X2_17 ( .A(_1181_), .B(_1180_), .Y(_1182_) );
OR2X2 OR2X2_18 ( .A(_1209_), .B(_1198_), .Y(_1543__4_) );
OR2X2 OR2X2_19 ( .A(_1102__bF_buf0), .B(PC_STACK_6__9_), .Y(_1370_) );
XNOR2X1 XNOR2X1_1 ( .A(_76_), .B(PC_pointer_0_), .Y(_16__0_) );
BUFX2 BUFX2_38 ( .A(_0__6_), .Y(CORE_InstructionIN[6]) );
BUFX2 BUFX2_39 ( .A(_0__7_), .Y(CORE_InstructionIN[7]) );
BUFX2 BUFX2_40 ( .A(_0__8_), .Y(CORE_InstructionIN[8]) );
BUFX2 BUFX2_41 ( .A(_0__9_), .Y(CORE_InstructionIN[9]) );
BUFX2 BUFX2_42 ( .A(_0__10_), .Y(CORE_InstructionIN[10]) );
BUFX2 BUFX2_43 ( .A(_0__13_), .Y(CORE_InstructionIN[13]) );
BUFX2 BUFX2_44 ( .A(_0__14_), .Y(CORE_InstructionIN[14]) );
BUFX2 BUFX2_45 ( .A(_0__15_), .Y(CORE_InstructionIN[15]) );
BUFX2 BUFX2_46 ( .A(_1__0_), .Y(IDATA_CORE_addr[0]) );
BUFX2 BUFX2_47 ( .A(_1__1_), .Y(IDATA_CORE_addr[1]) );
BUFX2 BUFX2_48 ( .A(_1__2_), .Y(IDATA_CORE_addr[2]) );
BUFX2 BUFX2_49 ( .A(_1__3_), .Y(IDATA_CORE_addr[3]) );
BUFX2 BUFX2_50 ( .A(_1__4_), .Y(IDATA_CORE_addr[4]) );
BUFX2 BUFX2_51 ( .A(_1__5_), .Y(IDATA_CORE_addr[5]) );
BUFX2 BUFX2_52 ( .A(_1__6_), .Y(IDATA_CORE_addr[6]) );
BUFX2 BUFX2_53 ( .A(_1__7_), .Y(IDATA_CORE_addr[7]) );
BUFX2 BUFX2_54 ( .A(_1__8_), .Y(IDATA_CORE_addr[8]) );
BUFX2 BUFX2_55 ( .A(_1__9_), .Y(IDATA_CORE_addr[9]) );
BUFX2 BUFX2_56 ( .A(_2_), .Y(IDATA_clk) );
BUFX2 BUFX2_57 ( .A(_3__0_), .Y(REG_R0[0]) );
BUFX2 BUFX2_58 ( .A(_3__1_), .Y(REG_R0[1]) );
BUFX2 BUFX2_59 ( .A(_3__2_), .Y(REG_R0[2]) );
BUFX2 BUFX2_60 ( .A(_3__3_), .Y(REG_R0[3]) );
BUFX2 BUFX2_61 ( .A(_3__4_), .Y(REG_R0[4]) );
BUFX2 BUFX2_62 ( .A(_3__5_), .Y(REG_R0[5]) );
BUFX2 BUFX2_63 ( .A(_3__6_), .Y(REG_R0[6]) );
BUFX2 BUFX2_64 ( .A(_3__7_), .Y(REG_R0[7]) );
BUFX2 BUFX2_65 ( .A(_3__8_), .Y(REG_R0[8]) );
BUFX2 BUFX2_66 ( .A(_3__9_), .Y(REG_R0[9]) );
BUFX2 BUFX2_67 ( .A(_0__11_), .Y(CORE_InstructionIN[11]) );
BUFX2 BUFX2_68 ( .A(_0__12_), .Y(CORE_InstructionIN[12]) );
BUFX2 BUFX2_69 ( .A(_0__0_), .Y(CORE_InstructionIN[0]) );
BUFX2 BUFX2_70 ( .A(_0__1_), .Y(CORE_InstructionIN[1]) );
BUFX2 BUFX2_71 ( .A(_0__2_), .Y(CORE_InstructionIN[2]) );
BUFX2 BUFX2_72 ( .A(_0__3_), .Y(CORE_InstructionIN[3]) );
BUFX2 BUFX2_73 ( .A(_0__4_), .Y(CORE_InstructionIN[4]) );
BUFX2 BUFX2_74 ( .A(_0__5_), .Y(CORE_InstructionIN[5]) );
endmodule
