magic
tech scmos
magscale 1 4
timestamp 1515870181
<< metal1 >>
rect 4237 5377 4259 5383
rect 4253 5363 4259 5377
rect 6200 5377 6211 5383
rect 3661 5357 3684 5363
rect 4253 5357 4291 5363
rect 3676 5354 3684 5357
rect 616 5337 627 5343
rect 904 5337 915 5343
rect 1336 5337 1347 5343
rect 1752 5337 1780 5343
rect 2349 5337 2360 5343
rect 2397 5337 2408 5343
rect 3405 5337 3427 5343
rect 3608 5337 3619 5343
rect 5036 5343 5044 5348
rect 5036 5337 5059 5343
rect 5420 5343 5428 5348
rect 5420 5337 5443 5343
rect 5724 5343 5732 5348
rect 5677 5337 5699 5343
rect 5709 5337 5732 5343
rect 6157 5337 6184 5343
rect 6428 5343 6436 5348
rect 6413 5337 6436 5343
rect 6925 5343 6931 5363
rect 6925 5337 6963 5343
rect 45 5317 72 5323
rect 300 5317 339 5323
rect 300 5314 308 5317
rect 477 5317 504 5323
rect 877 5317 915 5323
rect 36 5296 40 5304
rect 909 5297 915 5317
rect 1037 5317 1048 5323
rect 1261 5317 1272 5323
rect 1309 5317 1347 5323
rect 1341 5297 1347 5317
rect 1421 5317 1459 5323
rect 1453 5297 1459 5317
rect 2013 5317 2051 5323
rect 1476 5296 1480 5304
rect 2013 5297 2019 5317
rect 2216 5317 2227 5323
rect 2349 5317 2387 5323
rect 2349 5297 2355 5317
rect 2925 5317 2936 5323
rect 3469 5317 3507 5323
rect 3565 5317 3592 5323
rect 3469 5297 3475 5317
rect 4621 5317 4648 5323
rect 4685 5323 4691 5332
rect 4685 5317 4696 5323
rect 4765 5317 4803 5323
rect 3556 5296 3560 5304
rect 4733 5297 4744 5303
rect 4797 5297 4803 5317
rect 5181 5317 5192 5323
rect 5549 5317 5560 5323
rect 5597 5317 5635 5323
rect 5172 5296 5176 5304
rect 5565 5297 5576 5303
rect 5629 5297 5635 5317
rect 5933 5317 5971 5323
rect 5965 5297 5971 5317
rect 6045 5317 6083 5323
rect 6109 5317 6120 5323
rect 6077 5297 6083 5317
rect 6100 5296 6104 5304
rect 262 5276 264 5284
rect 1910 5276 1912 5284
rect 5768 5276 5770 5284
rect 1293 5137 1304 5143
rect 5896 5136 5898 5144
rect 6216 5137 6227 5143
rect 269 5097 280 5103
rect 445 5103 451 5123
rect 445 5097 483 5103
rect 557 5103 563 5123
rect 557 5097 595 5103
rect 765 5103 771 5123
rect 765 5097 803 5103
rect 893 5097 904 5103
rect 1357 5103 1363 5123
rect 1325 5097 1363 5103
rect 1725 5103 1731 5123
rect 1693 5097 1731 5103
rect 1837 5103 1843 5123
rect 1837 5097 1875 5103
rect 2125 5097 2168 5103
rect 2493 5103 2499 5123
rect 2605 5103 2611 5123
rect 3149 5117 3204 5123
rect 3196 5112 3204 5117
rect 2493 5097 2531 5103
rect 2573 5097 2611 5103
rect 4232 5097 4259 5103
rect 4312 5097 4323 5103
rect 188 5077 212 5083
rect 765 5077 776 5083
rect 1837 5077 1848 5083
rect 2493 5077 2504 5083
rect 3773 5077 3784 5083
rect 4205 5077 4232 5083
rect 4285 5077 4296 5083
rect 4317 5077 4323 5097
rect 4429 5103 4435 5123
rect 4488 5117 4499 5123
rect 4376 5097 4403 5103
rect 4429 5097 4467 5103
rect 4941 5103 4947 5123
rect 4964 5116 4968 5124
rect 4909 5097 4947 5103
rect 5208 5097 5219 5103
rect 6093 5103 6099 5123
rect 6061 5097 6099 5103
rect 4477 5077 4488 5083
rect 4716 5077 4728 5083
rect 4744 5077 4755 5083
rect 5180 5077 5203 5083
rect 5180 5072 5188 5077
rect 5496 5077 5523 5083
rect 5613 5077 5635 5083
rect 6141 5077 6163 5083
rect 6173 5077 6200 5083
rect 7320 5077 7347 5083
rect 4172 5063 4180 5066
rect 4172 5057 4195 5063
rect 5469 5057 5507 5063
rect 6429 5057 6467 5063
rect 7117 5057 7155 5063
rect 7229 5057 7267 5063
rect 7373 5057 7411 5063
rect 7405 4977 7416 4983
rect 5741 4957 5779 4963
rect 5853 4957 5891 4963
rect 6157 4957 6195 4963
rect 6525 4957 6563 4963
rect 152 4937 163 4943
rect 1368 4937 1379 4943
rect 1416 4937 1427 4943
rect 1629 4937 1640 4943
rect 1933 4937 1944 4943
rect 1981 4937 1992 4943
rect 2300 4937 2312 4943
rect 2504 4937 2515 4943
rect 24 4917 35 4923
rect 125 4917 163 4923
rect 157 4897 163 4917
rect 429 4917 467 4923
rect 493 4917 504 4923
rect 461 4897 467 4917
rect 653 4917 680 4923
rect 1021 4917 1032 4923
rect 1357 4923 1363 4932
rect 1341 4917 1363 4923
rect 1389 4917 1427 4923
rect 1453 4917 1480 4923
rect 829 4897 867 4903
rect 1421 4897 1427 4917
rect 1613 4917 1640 4923
rect 1896 4917 1907 4923
rect 1933 4917 1971 4923
rect 1604 4896 1608 4904
rect 1933 4897 1939 4917
rect 2509 4923 2515 4937
rect 3165 4937 3192 4943
rect 3388 4943 3396 4948
rect 3388 4937 3411 4943
rect 3448 4937 3459 4943
rect 4216 4937 4259 4943
rect 4349 4937 4360 4943
rect 4477 4937 4499 4943
rect 4520 4937 4531 4943
rect 5100 4943 5108 4948
rect 4936 4937 4963 4943
rect 5053 4937 5075 4943
rect 5085 4937 5108 4943
rect 5612 4943 5620 4948
rect 5612 4937 5635 4943
rect 7212 4937 7236 4943
rect 2509 4917 2531 4923
rect 2696 4917 2723 4923
rect 3000 4917 3011 4923
rect 3117 4917 3155 4923
rect 3117 4897 3123 4917
rect 3421 4917 3459 4923
rect 3453 4897 3459 4917
rect 3581 4917 3619 4923
rect 3613 4897 3619 4917
rect 3773 4917 3811 4923
rect 3773 4897 3779 4917
rect 4189 4917 4259 4923
rect 4253 4897 4259 4917
rect 4397 4917 4435 4923
rect 4429 4897 4435 4917
rect 5341 4917 5379 4923
rect 5028 4896 5032 4904
rect 5373 4897 5379 4917
rect 6040 4917 6067 4923
rect 5396 4896 5400 4904
rect 397 4877 408 4883
rect 4904 4877 4915 4883
rect 6605 4877 6659 4883
rect 6925 4877 6952 4883
rect 3308 4737 3336 4743
rect 3308 4732 3316 4737
rect 5309 4743 5315 4763
rect 5244 4737 5315 4743
rect 5837 4743 5843 4763
rect 6429 4743 6435 4763
rect 5837 4737 5876 4743
rect 6396 4737 6435 4743
rect 6712 4737 6739 4743
rect 6888 4737 6899 4743
rect 253 4703 259 4723
rect 221 4697 259 4703
rect 605 4697 632 4703
rect 925 4703 931 4723
rect 1076 4716 1080 4724
rect 925 4697 963 4703
rect 1085 4697 1096 4703
rect 1549 4703 1555 4723
rect 2546 4716 2552 4724
rect 2804 4716 2808 4724
rect 5224 4716 5228 4724
rect 5272 4717 5299 4723
rect 5736 4717 5747 4723
rect 6525 4717 6552 4723
rect 7101 4717 7128 4723
rect 1517 4697 1555 4703
rect 1917 4697 1928 4703
rect 1917 4688 1923 4697
rect 3896 4697 3923 4703
rect 4648 4697 4659 4703
rect 4877 4697 4888 4703
rect 5165 4697 5192 4703
rect 5208 4697 5219 4703
rect 5624 4697 5635 4703
rect 6072 4697 6083 4703
rect 7293 4697 7304 4703
rect 520 4677 531 4683
rect 1101 4677 1144 4683
rect 1245 4677 1299 4683
rect 1245 4657 1251 4677
rect 1320 4677 1347 4683
rect 2172 4677 2184 4683
rect 2216 4677 2227 4683
rect 2365 4677 2435 4683
rect 2504 4677 2515 4683
rect 2733 4677 2744 4683
rect 2861 4677 2872 4683
rect 3101 4677 3123 4683
rect 3469 4677 3491 4683
rect 3980 4677 4004 4683
rect 4376 4677 4387 4683
rect 4925 4677 4948 4683
rect 4940 4672 4948 4677
rect 5528 4677 5555 4683
rect 5917 4677 5928 4683
rect 6056 4677 6067 4683
rect 7016 4677 7032 4683
rect 3068 4663 3076 4666
rect 3068 4657 3091 4663
rect 3804 4663 3812 4666
rect 3789 4657 3812 4663
rect 5432 4657 5443 4663
rect 6173 4657 6211 4663
rect 6824 4657 6835 4663
rect 3165 4637 3192 4643
rect 6888 4637 6899 4643
rect 1618 4577 1656 4583
rect 3736 4577 3747 4583
rect 5656 4577 5726 4583
rect 61 4537 72 4543
rect 1048 4537 1059 4543
rect 1517 4537 1587 4543
rect 1869 4537 1908 4543
rect 2253 4537 2275 4543
rect 61 4517 99 4523
rect 61 4497 67 4517
rect 381 4517 392 4523
rect 653 4517 691 4523
rect 653 4497 659 4517
rect 824 4517 835 4523
rect 1021 4517 1048 4523
rect 1069 4517 1107 4523
rect 1101 4497 1107 4517
rect 2253 4523 2259 4537
rect 2600 4537 2616 4543
rect 2701 4543 2707 4563
rect 3948 4557 3971 4563
rect 3948 4554 3956 4557
rect 3420 4548 3428 4554
rect 4989 4557 5027 4563
rect 5917 4557 5955 4563
rect 6760 4557 6771 4563
rect 6909 4557 6947 4563
rect 6968 4557 6980 4563
rect 6972 4554 6980 4557
rect 2701 4537 2755 4543
rect 2776 4537 2803 4543
rect 2989 4537 3000 4543
rect 3388 4543 3396 4548
rect 3373 4537 3396 4543
rect 3613 4537 3640 4543
rect 4136 4537 4147 4543
rect 4157 4537 4168 4543
rect 4237 4537 4248 4543
rect 5032 4537 5043 4543
rect 2248 4517 2259 4523
rect 2285 4517 2323 4523
rect 1124 4496 1128 4504
rect 2125 4497 2136 4503
rect 2317 4497 2323 4517
rect 2573 4517 2600 4523
rect 2877 4517 2915 4523
rect 2564 4496 2568 4504
rect 2877 4497 2883 4517
rect 2989 4517 3027 4523
rect 2989 4497 2995 4517
rect 3325 4517 3363 4523
rect 3325 4497 3331 4517
rect 4072 4517 4083 4523
rect 4424 4517 4435 4523
rect 4605 4517 4643 4523
rect 4088 4496 4092 4504
rect 4637 4497 4643 4517
rect 4888 4517 4899 4523
rect 4920 4517 4963 4523
rect 5453 4517 5480 4523
rect 5517 4517 5544 4523
rect 5880 4517 5891 4523
rect 5181 4497 5192 4503
rect 6109 4497 6131 4503
rect 6717 4488 6723 4503
rect 3910 4476 3912 4484
rect 6365 4477 6419 4483
rect 6520 4477 6547 4483
rect 6557 4477 6568 4483
rect 6648 4477 6675 4483
rect 6808 4477 6835 4483
rect 3021 4337 3032 4343
rect 3848 4337 3859 4343
rect 3896 4336 3898 4344
rect 5517 4343 5523 4363
rect 5484 4337 5523 4343
rect 6141 4343 6147 4363
rect 6136 4337 6147 4343
rect 6909 4337 6936 4343
rect 6989 4343 6995 4363
rect 6989 4337 7027 4343
rect 61 4303 67 4323
rect 24 4297 35 4303
rect 61 4297 99 4303
rect 653 4303 659 4323
rect 653 4297 691 4303
rect 957 4303 963 4323
rect 980 4316 984 4324
rect 1517 4317 1528 4323
rect 1693 4317 1704 4323
rect 2616 4316 2620 4324
rect 925 4297 963 4303
rect 1213 4297 1224 4303
rect 1405 4297 1416 4303
rect 2157 4297 2184 4303
rect 3085 4303 3091 4323
rect 3496 4316 3500 4324
rect 3053 4297 3091 4303
rect 3224 4297 3235 4303
rect 3517 4303 3523 4323
rect 3517 4297 3555 4303
rect 3789 4303 3795 4323
rect 3789 4297 3827 4303
rect 4157 4303 4163 4323
rect 4472 4316 4476 4324
rect 4157 4297 4195 4303
rect 4493 4303 4499 4323
rect 4781 4317 4819 4323
rect 5076 4316 5080 4324
rect 5912 4317 5923 4323
rect 6280 4317 6291 4323
rect 6813 4317 6835 4323
rect 7021 4317 7027 4337
rect 7128 4337 7155 4343
rect 4456 4297 4467 4303
rect 4493 4297 4531 4303
rect 6093 4297 6104 4303
rect 61 4277 72 4283
rect 317 4277 355 4283
rect 1005 4277 1016 4283
rect 1213 4277 1240 4283
rect 1416 4277 1459 4283
rect 1645 4277 1672 4283
rect 1709 4277 1732 4283
rect 1724 4272 1732 4277
rect 2200 4277 2211 4283
rect 2280 4277 2291 4283
rect 1341 4257 1352 4263
rect 1756 4263 1764 4272
rect 1389 4257 1443 4263
rect 1756 4257 1784 4263
rect 2285 4257 2291 4277
rect 3080 4277 3091 4283
rect 3165 4277 3219 4283
rect 3576 4277 3587 4283
rect 3581 4257 3587 4277
rect 4157 4277 4168 4283
rect 4813 4277 4835 4283
rect 5292 4277 5347 4283
rect 5292 4272 5300 4277
rect 6397 4277 6435 4283
rect 4952 4256 4956 4264
rect 6397 4257 6403 4277
rect 6664 4277 6675 4283
rect 1101 4237 1128 4243
rect 5432 4177 5470 4183
rect 317 4143 323 4163
rect 1528 4157 1556 4163
rect 1548 4148 1556 4157
rect 2413 4157 2467 4163
rect 5693 4157 5731 4163
rect 7277 4157 7315 4163
rect 312 4137 323 4143
rect 333 4137 355 4143
rect 636 4137 675 4143
rect 861 4137 883 4143
rect 925 4137 947 4143
rect 1580 4143 1588 4148
rect 1388 4137 1412 4143
rect 1580 4137 1603 4143
rect 1640 4137 1651 4143
rect 1709 4137 1731 4143
rect 77 4117 88 4123
rect 253 4117 291 4123
rect 253 4097 259 4117
rect 360 4117 371 4123
rect 701 4117 712 4123
rect 1064 4117 1075 4123
rect 1085 4117 1144 4123
rect 1304 4117 1331 4123
rect 1613 4117 1651 4123
rect 1144 4097 1155 4103
rect 1645 4097 1651 4117
rect 1709 4123 1715 4137
rect 1784 4137 1795 4143
rect 1869 4137 1896 4143
rect 2008 4137 2019 4143
rect 2589 4143 2595 4152
rect 2472 4137 2483 4143
rect 2589 4137 2611 4143
rect 2648 4137 2659 4143
rect 3085 4137 3128 4143
rect 3448 4137 3475 4143
rect 4632 4137 4643 4143
rect 4920 4137 4931 4143
rect 5048 4137 5059 4143
rect 5544 4137 5555 4143
rect 5768 4137 5811 4143
rect 6072 4137 6083 4143
rect 6221 4137 6243 4143
rect 1688 4117 1715 4123
rect 2077 4117 2115 4123
rect 2109 4097 2115 4117
rect 2829 4117 2867 4123
rect 2690 4096 2696 4104
rect 2829 4097 2835 4117
rect 4013 4117 4024 4123
rect 4077 4117 4115 4123
rect 4296 4117 4323 4123
rect 4525 4117 4552 4123
rect 4893 4117 4931 4123
rect 3368 4096 3372 4104
rect 3389 4097 3427 4103
rect 3917 4097 3928 4103
rect 4269 4097 4307 4103
rect 4925 4097 4931 4117
rect 5512 4117 5571 4123
rect 5837 4117 5848 4123
rect 6029 4117 6056 4123
rect 6088 4117 6099 4123
rect 6205 4117 6216 4123
rect 6237 4123 6243 4137
rect 6424 4137 6435 4143
rect 6748 4143 6756 4148
rect 6733 4137 6756 4143
rect 6237 4117 6280 4123
rect 6856 4117 6867 4123
rect 5341 4097 5363 4103
rect 5613 4097 5624 4103
rect 6989 4097 7016 4103
rect 2573 4077 2584 4083
rect 3286 4076 3288 4084
rect 3533 4077 3572 4083
rect 3533 4057 3539 4077
rect 3900 4077 3939 4083
rect 3933 4057 3939 4077
rect 4461 4077 4500 4083
rect 4461 4057 4467 4077
rect 5596 4077 5635 4083
rect 5629 4057 5635 4077
rect 6316 4077 6355 4083
rect 6349 4057 6355 4077
rect 6572 4077 6611 4083
rect 6605 4057 6611 4077
rect 1286 3936 1288 3944
rect 3469 3937 3492 3943
rect 3484 3932 3492 3937
rect 5357 3943 5363 3963
rect 5324 3937 5363 3943
rect 6941 3943 6947 3963
rect 6941 3937 6979 3943
rect 77 3897 88 3903
rect 269 3903 275 3923
rect 248 3897 275 3903
rect 461 3903 467 3923
rect 429 3897 467 3903
rect 573 3903 579 3923
rect 573 3897 611 3903
rect 632 3897 659 3903
rect 941 3903 947 3923
rect 909 3897 947 3903
rect 1053 3903 1059 3923
rect 1053 3897 1091 3903
rect 1324 3903 1332 3906
rect 1324 3897 1363 3903
rect 1485 3903 1491 3923
rect 1453 3897 1491 3903
rect 1656 3897 1667 3903
rect 1928 3897 1939 3903
rect 2397 3903 2403 3923
rect 2365 3897 2403 3903
rect 2509 3903 2515 3923
rect 3128 3916 3132 3924
rect 2477 3897 2515 3903
rect 3149 3903 3155 3923
rect 3501 3917 3539 3923
rect 3556 3916 3560 3924
rect 3149 3897 3187 3903
rect 3357 3897 3368 3903
rect 3629 3897 3667 3903
rect 3741 3897 3779 3903
rect 4045 3903 4051 3923
rect 4360 3916 4364 3924
rect 4045 3897 4083 3903
rect 4312 3897 4328 3903
rect 4381 3903 4387 3923
rect 4701 3917 4712 3923
rect 4820 3916 4824 3924
rect 6829 3917 6851 3923
rect 6973 3917 6979 3937
rect 4381 3897 4392 3903
rect 4717 3897 4744 3903
rect 312 3877 323 3883
rect 333 3877 355 3883
rect 317 3857 323 3877
rect 573 3877 584 3883
rect 1053 3877 1064 3883
rect 1101 3877 1128 3883
rect 1773 3877 1800 3883
rect 2445 3877 2451 3892
rect 2637 3877 2691 3883
rect 2685 3857 2691 3877
rect 2792 3877 2803 3883
rect 4045 3877 4056 3883
rect 4477 3877 4488 3883
rect 4589 3877 4600 3883
rect 4717 3877 4723 3897
rect 5628 3906 5636 3912
rect 6189 3883 6195 3903
rect 6253 3897 6280 3903
rect 6141 3877 6179 3883
rect 6189 3877 6216 3883
rect 3436 3868 3444 3872
rect 5528 3857 5539 3863
rect 5837 3857 5875 3863
rect 6141 3857 6147 3877
rect 6573 3877 6584 3883
rect 7160 3877 7171 3883
rect 6253 3857 6323 3863
rect 7117 3857 7155 3863
rect 1693 3757 1747 3763
rect 604 3737 628 3743
rect 1037 3737 1048 3743
rect 1256 3737 1267 3743
rect 1544 3737 1555 3743
rect 1832 3737 1859 3743
rect 2477 3737 2488 3743
rect 3165 3743 3171 3763
rect 3517 3757 3528 3763
rect 3629 3757 3640 3763
rect 3741 3757 3752 3763
rect 3812 3757 3843 3763
rect 4776 3757 4787 3763
rect 3160 3737 3171 3743
rect 3181 3737 3235 3743
rect 3277 3737 3288 3743
rect 5053 3737 5092 3743
rect 5357 3743 5363 3763
rect 5661 3757 5699 3763
rect 5357 3737 5395 3743
rect 5853 3743 5859 3763
rect 5853 3737 5891 3743
rect 6476 3743 6484 3748
rect 6909 3743 6915 3763
rect 6312 3737 6339 3743
rect 6429 3737 6451 3743
rect 6461 3737 6484 3743
rect 6877 3737 6915 3743
rect 216 3717 227 3723
rect 824 3717 835 3723
rect 856 3717 883 3723
rect 877 3697 883 3717
rect 968 3717 979 3723
rect 1128 3717 1171 3723
rect 1197 3717 1235 3723
rect 1277 3717 1315 3723
rect 1197 3697 1203 3717
rect 1309 3697 1315 3717
rect 1421 3717 1432 3723
rect 1560 3717 1571 3723
rect 1768 3717 1779 3723
rect 1848 3717 1875 3723
rect 2429 3717 2467 3723
rect 1576 3696 1580 3704
rect 2429 3697 2435 3717
rect 3096 3717 3112 3723
rect 3373 3717 3411 3723
rect 2509 3697 2547 3703
rect 2824 3696 2828 3704
rect 3117 3697 3123 3712
rect 3373 3697 3379 3717
rect 4573 3717 4584 3723
rect 4733 3717 4771 3723
rect 4941 3717 4952 3723
rect 5608 3717 5635 3723
rect 5784 3717 5811 3723
rect 6440 3717 6451 3723
rect 7064 3717 7091 3723
rect 4184 3696 4188 3704
rect 4413 3697 4424 3703
rect 4616 3696 4620 3704
rect 5469 3697 5491 3703
rect 472 3676 474 3684
rect 2742 3676 2744 3684
rect 3629 3677 3672 3683
rect 5222 3676 5224 3684
rect 6054 3676 6056 3684
rect 2870 3536 2872 3544
rect 3368 3537 3395 3543
rect 3912 3537 3923 3543
rect 4344 3537 4392 3543
rect 4877 3543 4883 3563
rect 4844 3537 4883 3543
rect 5677 3537 5731 3543
rect 6333 3543 6339 3563
rect 6573 3543 6579 3563
rect 6333 3537 6372 3543
rect 6540 3537 6579 3543
rect 6893 3543 6899 3563
rect 6893 3537 6931 3543
rect 285 3517 296 3523
rect 829 3508 835 3523
rect 109 3497 136 3503
rect 925 3497 936 3503
rect 1117 3497 1128 3503
rect 1405 3503 1411 3523
rect 1373 3497 1411 3503
rect 1437 3497 1448 3503
rect 1533 3497 1544 3503
rect 1613 3503 1619 3523
rect 1636 3516 1640 3524
rect 2088 3516 2092 3524
rect 1581 3497 1619 3503
rect 2109 3503 2115 3523
rect 2908 3517 2931 3523
rect 2908 3512 2916 3517
rect 2109 3497 2147 3503
rect 2344 3497 2371 3503
rect 2957 3497 2984 3503
rect 525 3477 547 3483
rect 989 3477 1011 3483
rect 1400 3477 1411 3483
rect 1852 3477 1876 3483
rect 2285 3477 2296 3483
rect 2653 3477 2664 3483
rect 2957 3477 2963 3497
rect 3005 3497 3016 3503
rect 3469 3503 3475 3523
rect 4824 3516 4828 3524
rect 5612 3517 5635 3523
rect 5612 3512 5620 3517
rect 5869 3517 5880 3523
rect 6925 3517 6931 3537
rect 7112 3537 7123 3543
rect 3469 3497 3507 3503
rect 3629 3497 3640 3503
rect 4760 3497 4771 3503
rect 4781 3497 4792 3503
rect 5277 3497 5315 3503
rect 5373 3497 5395 3503
rect 6056 3497 6067 3503
rect 3212 3477 3224 3483
rect 3357 3477 3368 3483
rect 3469 3477 3480 3483
rect 3517 3477 3528 3483
rect 6648 3477 6659 3483
rect 6728 3477 6755 3483
rect 492 3463 500 3466
rect 492 3457 515 3463
rect 3533 3457 3539 3472
rect 5352 3457 5363 3463
rect 6296 3377 6318 3383
rect 2157 3357 2184 3363
rect 5272 3357 5308 3363
rect 5485 3357 5523 3363
rect 6013 3357 6051 3363
rect 7229 3357 7267 3363
rect 1052 3343 1060 3348
rect 1052 3337 1075 3343
rect 1112 3337 1155 3343
rect 1437 3337 1448 3343
rect 1644 3343 1652 3348
rect 1644 3337 1667 3343
rect 1704 3337 1715 3343
rect 2301 3337 2339 3343
rect 2429 3337 2440 3343
rect 2568 3337 2579 3343
rect 3181 3343 3187 3352
rect 2861 3337 2883 3343
rect 3149 3337 3171 3343
rect 3181 3337 3235 3343
rect 3928 3337 3944 3343
rect 120 3317 131 3323
rect 312 3317 323 3323
rect 445 3317 483 3323
rect 573 3317 584 3323
rect 445 3297 451 3317
rect 712 3317 723 3323
rect 1085 3317 1155 3323
rect 1149 3297 1155 3317
rect 1533 3317 1560 3323
rect 1677 3317 1715 3323
rect 1709 3297 1715 3317
rect 1976 3317 1987 3323
rect 2008 3317 2035 3323
rect 2029 3297 2035 3317
rect 3245 3317 3283 3323
rect 2509 3297 2547 3303
rect 3277 3297 3283 3317
rect 3741 3317 3779 3323
rect 3741 3297 3747 3317
rect 4061 3323 4067 3343
rect 4440 3337 4451 3343
rect 4653 3337 4664 3343
rect 4904 3337 4915 3343
rect 5128 3337 5139 3343
rect 5341 3343 5347 3352
rect 5325 3337 5347 3343
rect 5368 3337 5395 3343
rect 6077 3337 6104 3343
rect 6205 3337 6280 3343
rect 6760 3337 6771 3343
rect 6893 3337 6904 3343
rect 7021 3337 7032 3343
rect 7192 3337 7203 3343
rect 7288 3337 7315 3343
rect 4061 3317 4088 3323
rect 4200 3317 4243 3323
rect 4376 3317 4387 3323
rect 4728 3317 4739 3323
rect 6749 3317 6771 3323
rect 6792 3317 6803 3323
rect 7352 3317 7363 3323
rect 4744 3296 4748 3304
rect 5848 3297 5859 3303
rect 5917 3297 5928 3303
rect 6445 3297 6467 3303
rect 4045 3277 4056 3283
rect 5565 3277 5635 3283
rect 5629 3257 5635 3277
rect 5928 3277 5971 3283
rect 6557 3277 6596 3283
rect 6557 3257 6563 3277
rect 1128 3137 1139 3143
rect 1176 3136 1178 3144
rect 1526 3136 1528 3144
rect 3741 3137 3768 3143
rect 4632 3137 4643 3143
rect 4989 3143 4995 3163
rect 4956 3137 4995 3143
rect 520 3116 524 3124
rect 541 3103 547 3123
rect 541 3097 579 3103
rect 600 3097 643 3103
rect 733 3103 739 3123
rect 733 3097 771 3103
rect 1037 3103 1043 3123
rect 1037 3097 1075 3103
rect 1629 3103 1635 3123
rect 1597 3097 1635 3103
rect 1960 3097 1971 3103
rect 2845 3103 2851 3123
rect 3133 3117 3171 3123
rect 3277 3117 3288 3123
rect 2813 3097 2851 3103
rect 3032 3097 3043 3103
rect 3053 3097 3064 3103
rect 3293 3097 3320 3103
rect 605 3077 616 3083
rect 733 3077 744 3083
rect 1037 3077 1048 3083
rect 1085 3077 1112 3083
rect 1564 3077 1587 3083
rect 1564 3072 1572 3077
rect 1688 3077 1699 3083
rect 2077 3077 2099 3083
rect 2141 3077 2184 3083
rect 2221 3077 2232 3083
rect 2840 3077 2851 3083
rect 3016 3077 3027 3083
rect 3293 3077 3299 3097
rect 3341 3097 3368 3103
rect 3421 3103 3427 3123
rect 3660 3117 3683 3123
rect 3660 3112 3668 3117
rect 3789 3117 3800 3123
rect 3421 3097 3459 3103
rect 3965 3103 3971 3123
rect 4413 3117 4424 3123
rect 4477 3117 4488 3123
rect 4936 3116 4940 3124
rect 3965 3097 4003 3103
rect 5160 3097 5176 3103
rect 7389 3097 7400 3103
rect 3965 3077 3976 3083
rect 4013 3077 4035 3083
rect 4029 3068 4035 3077
rect 5048 3077 5059 3083
rect 5112 3077 5123 3083
rect 5917 3077 5944 3083
rect 6205 3077 6248 3083
rect 6301 3077 6312 3083
rect 5437 3057 5475 3063
rect 5933 3057 5971 3063
rect 5996 3063 6004 3066
rect 5992 3057 6004 3063
rect 6232 3057 6248 3063
rect 6829 3057 6867 3063
rect 2168 3037 2195 3043
rect 4685 2957 4696 2963
rect 4925 2957 4936 2963
rect 4996 2957 5027 2963
rect 5533 2957 5571 2963
rect 88 2937 99 2943
rect 253 2937 264 2943
rect 525 2937 547 2943
rect 637 2937 675 2943
rect 1565 2937 1576 2943
rect 1997 2937 2008 2943
rect 2861 2937 2872 2943
rect 3000 2937 3012 2943
rect 3613 2937 3635 2943
rect 3933 2937 3944 2943
rect 4269 2937 4280 2943
rect 4589 2937 4611 2943
rect 4860 2943 4868 2944
rect 4860 2937 4872 2943
rect 5592 2937 5619 2943
rect 6093 2943 6099 2963
rect 6093 2937 6131 2943
rect 6556 2937 6568 2943
rect 6621 2943 6627 2963
rect 6829 2957 6867 2963
rect 7325 2957 7363 2963
rect 6621 2937 6659 2943
rect 7256 2937 7267 2943
rect 61 2917 72 2923
rect 253 2917 291 2923
rect 253 2897 259 2917
rect 701 2917 739 2923
rect 733 2897 739 2917
rect 1053 2917 1091 2923
rect 1085 2897 1091 2917
rect 1421 2917 1459 2923
rect 1108 2896 1112 2904
rect 1421 2897 1427 2917
rect 1645 2917 1683 2923
rect 1645 2897 1651 2917
rect 2061 2917 2072 2923
rect 2109 2917 2152 2923
rect 2461 2917 2472 2923
rect 2936 2917 2947 2923
rect 3581 2917 3592 2923
rect 3896 2917 3907 2923
rect 3933 2917 3971 2923
rect 2125 2897 2136 2903
rect 3224 2897 3235 2903
rect 3245 2897 3283 2903
rect 3300 2896 3304 2904
rect 3933 2897 3939 2917
rect 4269 2917 4307 2923
rect 4269 2897 4275 2917
rect 5053 2917 5064 2923
rect 6093 2917 6104 2923
rect 4541 2897 4568 2903
rect 5096 2896 5100 2904
rect 5720 2897 5731 2903
rect 5901 2897 5912 2903
rect 1318 2876 1320 2884
rect 2310 2876 2312 2884
rect 2780 2883 2788 2888
rect 2776 2877 2788 2883
rect 3142 2876 3144 2884
rect 4764 2883 4772 2888
rect 4764 2877 4803 2883
rect 4797 2857 4803 2877
rect 5116 2877 5155 2883
rect 5149 2857 5155 2877
rect 5704 2877 5747 2883
rect 5741 2857 5747 2877
rect 445 2737 456 2743
rect 2461 2737 2472 2743
rect 3309 2737 3320 2743
rect 4669 2743 4675 2763
rect 4669 2737 4708 2743
rect 5517 2743 5523 2763
rect 5517 2737 5555 2743
rect 253 2703 259 2723
rect 413 2717 424 2723
rect 776 2717 787 2723
rect 221 2697 259 2703
rect 701 2697 712 2703
rect 1325 2697 1336 2703
rect 1805 2703 1811 2723
rect 1805 2697 1843 2703
rect 2525 2703 2531 2723
rect 2893 2717 2931 2723
rect 2493 2697 2531 2703
rect 349 2677 360 2683
rect 461 2677 488 2683
rect 525 2677 563 2683
rect 968 2677 995 2683
rect 1160 2677 1203 2683
rect 1912 2677 1923 2683
rect 3021 2697 3048 2703
rect 2120 2677 2131 2683
rect 2520 2677 2531 2683
rect 2621 2677 2632 2683
rect 2973 2677 2984 2683
rect 3021 2677 3027 2697
rect 3197 2697 3208 2703
rect 3373 2703 3379 2723
rect 3341 2697 3379 2703
rect 3469 2697 3496 2703
rect 3469 2677 3475 2697
rect 3661 2703 3667 2723
rect 4557 2717 4579 2723
rect 4680 2717 4691 2723
rect 4724 2716 4728 2724
rect 5320 2716 5324 2724
rect 5549 2717 5555 2737
rect 6013 2743 6019 2763
rect 5992 2737 6019 2743
rect 7112 2737 7155 2743
rect 7272 2736 7274 2744
rect 5640 2716 5644 2724
rect 5981 2717 6008 2723
rect 6157 2717 6168 2723
rect 3661 2697 3699 2703
rect 4013 2697 4040 2703
rect 4408 2697 4419 2703
rect 4760 2697 4771 2703
rect 5197 2697 5256 2703
rect 6168 2697 6211 2703
rect 6456 2697 6467 2703
rect 6733 2697 6744 2703
rect 3661 2677 3672 2683
rect 3709 2677 3731 2683
rect 3725 2668 3731 2677
rect 4157 2677 4179 2683
rect 4221 2677 4248 2683
rect 4440 2677 4467 2683
rect 5288 2677 5299 2683
rect 6616 2677 6627 2683
rect 7260 2668 7268 2672
rect 1064 2657 1075 2663
rect 4124 2663 4132 2666
rect 4124 2657 4147 2663
rect 5576 2637 5587 2643
rect 5213 2577 5240 2583
rect 1053 2557 1080 2563
rect 733 2537 760 2543
rect 925 2543 931 2552
rect 925 2537 947 2543
rect 1101 2537 1144 2543
rect 1709 2537 1720 2543
rect 1837 2537 1848 2543
rect 3165 2543 3171 2563
rect 3160 2537 3171 2543
rect 3181 2537 3224 2543
rect 45 2517 83 2523
rect 120 2517 132 2523
rect 124 2512 132 2517
rect 205 2517 243 2523
rect 317 2517 355 2523
rect 349 2497 355 2517
rect 957 2517 984 2523
rect 1080 2517 1091 2523
rect 1453 2517 1491 2523
rect 372 2496 376 2504
rect 845 2497 856 2503
rect 893 2497 915 2503
rect 1453 2497 1459 2517
rect 1837 2517 1875 2523
rect 1837 2497 1843 2517
rect 2008 2517 2019 2523
rect 2669 2517 2707 2523
rect 2136 2497 2147 2503
rect 2669 2497 2675 2517
rect 3261 2523 3267 2543
rect 3373 2537 3400 2543
rect 3597 2537 3608 2543
rect 4332 2543 4340 2544
rect 4332 2537 4344 2543
rect 4589 2537 4616 2543
rect 4680 2537 4691 2543
rect 4968 2537 4979 2543
rect 5309 2543 5315 2563
rect 5309 2537 5347 2543
rect 5741 2543 5747 2563
rect 6397 2557 6435 2563
rect 6765 2557 6803 2563
rect 5709 2537 5747 2543
rect 6685 2537 6696 2543
rect 6861 2537 6872 2543
rect 3101 2517 3139 2523
rect 3261 2517 3288 2523
rect 3080 2496 3084 2504
rect 3101 2497 3107 2517
rect 3533 2517 3544 2523
rect 3741 2517 3779 2523
rect 3245 2497 3256 2503
rect 3741 2497 3747 2517
rect 4045 2517 4083 2523
rect 4045 2497 4051 2517
rect 4941 2517 4979 2523
rect 4413 2497 4435 2503
rect 4973 2497 4979 2517
rect 5101 2517 5112 2523
rect 5613 2497 5635 2503
rect 6045 2497 6067 2503
rect 6573 2497 6595 2503
rect 6941 2497 6968 2503
rect 7133 2497 7155 2503
rect 1896 2477 1907 2483
rect 3757 2477 3763 2492
rect 4909 2477 4920 2483
rect 5405 2477 5444 2483
rect 5405 2457 5411 2477
rect 6936 2477 6984 2483
rect 7144 2477 7187 2483
rect 7341 2483 7347 2503
rect 7309 2477 7347 2483
rect 7309 2457 7315 2477
rect 6280 2437 6291 2443
rect 653 2337 664 2343
rect 1688 2337 1699 2343
rect 2573 2337 2584 2343
rect 3992 2337 4003 2343
rect 4040 2336 4042 2344
rect 4328 2337 4339 2343
rect 5798 2336 5800 2344
rect 6168 2337 6184 2343
rect 6648 2337 6675 2343
rect 6861 2343 6867 2363
rect 6861 2337 6899 2343
rect 253 2303 259 2323
rect 221 2297 259 2303
rect 717 2303 723 2323
rect 685 2297 723 2303
rect 749 2297 760 2303
rect 845 2297 856 2303
rect 925 2303 931 2323
rect 893 2297 931 2303
rect 1085 2303 1091 2323
rect 1053 2297 1091 2303
rect 1533 2303 1539 2323
rect 1501 2297 1539 2303
rect 1565 2297 1576 2303
rect 1997 2303 2003 2323
rect 2312 2316 2316 2324
rect 1965 2297 2003 2303
rect 2333 2303 2339 2323
rect 2296 2297 2307 2303
rect 2333 2297 2371 2303
rect 2637 2303 2643 2323
rect 2605 2297 2643 2303
rect 2941 2303 2947 2323
rect 2909 2297 2947 2303
rect 3053 2303 3059 2323
rect 2984 2297 3027 2303
rect 3053 2297 3091 2303
rect 3389 2303 3395 2323
rect 3357 2297 3395 2303
rect 3821 2303 3827 2323
rect 3789 2297 3827 2303
rect 3933 2303 3939 2323
rect 3933 2297 3971 2303
rect 4269 2303 4275 2323
rect 6152 2317 6163 2323
rect 6685 2317 6707 2323
rect 6893 2317 6899 2337
rect 7080 2337 7123 2343
rect 7069 2317 7080 2323
rect 4269 2297 4307 2303
rect 5101 2297 5112 2303
rect 5596 2303 5604 2308
rect 5596 2297 5608 2303
rect 5949 2288 5955 2303
rect 248 2277 259 2283
rect 397 2277 419 2283
rect 1133 2277 1160 2283
rect 1480 2277 1491 2283
rect 2264 2277 2291 2283
rect 2632 2277 2643 2283
rect 2876 2277 2899 2283
rect 2876 2272 2884 2277
rect 2936 2277 2947 2283
rect 3053 2277 3064 2283
rect 3101 2277 3156 2283
rect 3148 2272 3156 2277
rect 3768 2277 3779 2283
rect 3869 2277 3880 2283
rect 3933 2277 3944 2283
rect 4269 2277 4280 2283
rect 4813 2277 4824 2283
rect 1724 2263 1732 2272
rect 1724 2257 1752 2263
rect 4813 2257 4819 2277
rect 5309 2277 5347 2283
rect 5309 2257 5315 2277
rect 5901 2277 5939 2283
rect 5421 2257 5459 2263
rect 5901 2257 5907 2277
rect 5960 2277 5987 2283
rect 6605 2277 6616 2283
rect 7181 2277 7224 2283
rect 7261 2277 7299 2283
rect 7261 2257 7267 2277
rect 6728 2237 6739 2243
rect 1469 2157 1523 2163
rect 3436 2157 3464 2163
rect 3436 2148 3444 2157
rect 5693 2157 5731 2163
rect 6541 2157 6579 2163
rect 781 2137 803 2143
rect 797 2128 803 2137
rect 1821 2137 1832 2143
rect 2200 2137 2243 2143
rect 2285 2137 2296 2143
rect 2348 2143 2356 2148
rect 2344 2137 2356 2143
rect 3197 2137 3240 2143
rect 3341 2137 3352 2143
rect 3404 2143 3412 2148
rect 3389 2137 3412 2143
rect 3645 2137 3656 2143
rect 3965 2137 3987 2143
rect 4029 2137 4040 2143
rect 4157 2137 4179 2143
rect 4200 2137 4259 2143
rect 253 2117 291 2123
rect 253 2097 259 2117
rect 685 2117 723 2123
rect 685 2097 691 2117
rect 808 2117 819 2123
rect 1160 2117 1176 2123
rect 1357 2117 1384 2123
rect 1821 2117 1860 2123
rect 1852 2114 1860 2117
rect 2216 2117 2259 2123
rect 2285 2117 2323 2123
rect 2285 2097 2291 2117
rect 2792 2117 2819 2123
rect 3341 2117 3379 2123
rect 3341 2097 3347 2117
rect 3645 2117 3683 2123
rect 3645 2097 3651 2117
rect 4909 2117 4920 2123
rect 5261 2117 5272 2123
rect 3884 2103 3892 2108
rect 3884 2097 3907 2103
rect 5581 2097 5592 2103
rect 6717 2097 6739 2103
rect 7160 2097 7171 2103
rect 3917 2077 3944 2083
rect 4552 2077 4563 2083
rect 5965 2077 6035 2083
rect 6029 2057 6035 2077
rect 6438 2076 6440 2084
rect 7021 2077 7091 2083
rect 7021 2057 7027 2077
rect 6253 2037 6264 2043
rect 3693 1937 3704 1943
rect 7053 1943 7059 1963
rect 7053 1937 7123 1943
rect 205 1917 216 1923
rect 61 1897 72 1903
rect 312 1897 323 1903
rect 568 1897 579 1903
rect 861 1903 867 1923
rect 829 1897 867 1903
rect 973 1903 979 1923
rect 941 1897 979 1903
rect 1133 1903 1139 1923
rect 1277 1903 1283 1923
rect 1133 1897 1203 1903
rect 1245 1897 1283 1903
rect 1352 1897 1363 1903
rect 1485 1903 1491 1923
rect 1874 1916 1880 1924
rect 1453 1897 1491 1903
rect 1720 1897 1736 1903
rect 2237 1903 2243 1923
rect 2205 1897 2243 1903
rect 2605 1897 2648 1903
rect 3277 1897 3288 1903
rect 3453 1903 3459 1923
rect 4429 1917 4451 1923
rect 5000 1916 5004 1924
rect 6093 1917 6104 1923
rect 3453 1897 3491 1903
rect 4317 1897 4355 1903
rect 4717 1897 4755 1903
rect 4920 1897 4931 1903
rect 4984 1897 4995 1903
rect 5133 1897 5155 1903
rect 5192 1897 5219 1903
rect 5229 1897 5283 1903
rect 5533 1897 5576 1903
rect 6173 1897 6200 1903
rect 285 1877 307 1883
rect 1224 1877 1235 1883
rect 1693 1877 1763 1883
rect 2168 1877 2195 1883
rect 2520 1877 2531 1883
rect 1800 1857 1811 1863
rect 2525 1857 2531 1877
rect 2648 1877 2659 1883
rect 2872 1877 2883 1883
rect 3021 1877 3032 1883
rect 3453 1877 3464 1883
rect 3725 1877 3747 1883
rect 3853 1877 3875 1883
rect 3885 1877 3907 1883
rect 3885 1868 3891 1877
rect 5341 1877 5352 1883
rect 5384 1877 5416 1883
rect 5804 1877 5816 1883
rect 5901 1877 5944 1883
rect 6733 1877 6771 1883
rect 2589 1857 2643 1863
rect 5837 1857 5875 1863
rect 5981 1857 6019 1863
rect 6429 1857 6440 1863
rect 6765 1857 6771 1877
rect 7261 1877 7299 1883
rect 7261 1857 7267 1877
rect 2690 1837 2728 1843
rect 6120 1837 6158 1843
rect 7112 1837 7123 1843
rect 3165 1777 3176 1783
rect 4093 1777 4104 1783
rect 4301 1757 4312 1763
rect 6925 1757 6963 1763
rect 632 1737 643 1743
rect 776 1737 787 1743
rect 1404 1743 1412 1748
rect 1404 1737 1427 1743
rect 1464 1737 1475 1743
rect 1736 1737 1747 1743
rect 2552 1737 2563 1743
rect 2605 1737 2616 1743
rect 2669 1737 2680 1743
rect 2972 1737 2996 1743
rect 3192 1737 3219 1743
rect 3309 1737 3320 1743
rect 616 1717 659 1723
rect 669 1717 707 1723
rect 701 1697 707 1717
rect 813 1717 824 1723
rect 872 1717 899 1723
rect 1437 1717 1475 1723
rect 845 1697 856 1703
rect 1469 1697 1475 1717
rect 2029 1717 2067 1723
rect 2029 1697 2035 1717
rect 2104 1717 2115 1723
rect 2525 1717 2563 1723
rect 2557 1697 2563 1717
rect 2616 1717 2643 1723
rect 2669 1717 2707 1723
rect 2669 1697 2675 1717
rect 3229 1717 3267 1723
rect 3293 1717 3304 1723
rect 3261 1697 3267 1717
rect 3373 1717 3411 1723
rect 3373 1697 3379 1717
rect 3517 1717 3528 1723
rect 3565 1723 3571 1743
rect 4365 1737 4376 1743
rect 5341 1737 5368 1743
rect 5672 1737 5683 1743
rect 6157 1737 6168 1743
rect 6600 1737 6611 1743
rect 7400 1737 7411 1743
rect 3565 1717 3592 1723
rect 4520 1717 4531 1723
rect 4541 1717 4568 1723
rect 5133 1717 5171 1723
rect 3549 1697 3560 1703
rect 4484 1696 4488 1704
rect 4957 1697 4968 1703
rect 5133 1697 5139 1717
rect 5320 1717 5331 1723
rect 5688 1717 5699 1723
rect 5933 1717 5960 1723
rect 6536 1717 6547 1723
rect 6333 1697 6355 1703
rect 4104 1677 4136 1683
rect 4301 1677 4312 1683
rect 4429 1677 4468 1683
rect 4429 1657 4435 1677
rect 6280 1677 6323 1683
rect 360 1536 362 1544
rect 4669 1543 4675 1563
rect 4669 1537 4708 1543
rect 6061 1543 6067 1563
rect 6028 1537 6067 1543
rect 6872 1536 6874 1544
rect 253 1503 259 1523
rect 221 1497 259 1503
rect 605 1497 616 1503
rect 1069 1503 1075 1523
rect 1069 1497 1107 1503
rect 1581 1503 1587 1523
rect 1604 1516 1608 1524
rect 1549 1497 1587 1503
rect 1613 1497 1624 1503
rect 1932 1503 1940 1506
rect 1901 1497 1940 1503
rect 2205 1503 2211 1523
rect 2141 1497 2211 1503
rect 2381 1503 2387 1523
rect 2792 1516 2796 1524
rect 2381 1497 2419 1503
rect 2504 1497 2515 1503
rect 2813 1503 2819 1523
rect 2813 1497 2851 1503
rect 2920 1497 2931 1503
rect 2941 1497 2952 1503
rect 3293 1503 3299 1523
rect 3261 1497 3299 1503
rect 3405 1503 3411 1523
rect 4200 1517 4227 1523
rect 4461 1517 4472 1523
rect 3405 1497 3443 1503
rect 3885 1497 3912 1503
rect 4237 1497 4243 1512
rect 4684 1503 4692 1508
rect 4684 1497 4696 1503
rect 5128 1497 5155 1503
rect 5533 1503 5539 1523
rect 5773 1517 5795 1523
rect 6584 1517 6595 1523
rect 5501 1497 5539 1503
rect 5624 1497 5651 1503
rect 6920 1497 6947 1503
rect 7240 1497 7267 1503
rect 248 1477 259 1483
rect 1016 1477 1027 1483
rect 1069 1477 1080 1483
rect 1117 1477 1144 1483
rect 2872 1477 2883 1483
rect 2893 1477 2915 1483
rect 2877 1457 2883 1477
rect 3224 1477 3251 1483
rect 3405 1477 3416 1483
rect 3960 1477 3971 1483
rect 3981 1477 4003 1483
rect 3965 1457 3971 1477
rect 4360 1477 4371 1483
rect 4520 1477 4547 1483
rect 5016 1477 5027 1483
rect 5229 1477 5272 1483
rect 5976 1477 5987 1483
rect 6284 1477 6312 1483
rect 6733 1477 6771 1483
rect 4500 1457 4531 1463
rect 5629 1457 5640 1463
rect 6765 1457 6771 1477
rect 7053 1477 7080 1483
rect 1144 1437 1171 1443
rect 1997 1357 2008 1363
rect 2412 1357 2424 1363
rect 2412 1354 2420 1357
rect 616 1337 627 1343
rect 1933 1337 1960 1343
rect 2008 1337 2051 1343
rect 2445 1337 2467 1343
rect 2748 1337 2787 1343
rect 3000 1337 3011 1343
rect 3128 1337 3139 1343
rect 3565 1337 3587 1343
rect 4669 1337 4680 1343
rect 4732 1343 4740 1348
rect 4717 1337 4740 1343
rect 5437 1343 5443 1363
rect 5933 1357 5971 1363
rect 5405 1337 5443 1343
rect 6173 1343 6179 1363
rect 6141 1337 6179 1343
rect 6920 1337 6947 1343
rect 216 1317 227 1323
rect 253 1317 291 1323
rect 365 1317 376 1323
rect 232 1296 236 1304
rect 253 1297 259 1317
rect 397 1317 435 1323
rect 429 1297 435 1317
rect 541 1317 579 1323
rect 541 1297 547 1317
rect 829 1317 840 1323
rect 968 1317 979 1323
rect 1005 1317 1043 1323
rect 984 1296 988 1304
rect 1005 1297 1011 1317
rect 1101 1317 1144 1323
rect 1501 1317 1539 1323
rect 1117 1297 1128 1303
rect 1501 1297 1507 1317
rect 2152 1317 2179 1323
rect 2925 1317 2952 1323
rect 2973 1317 3011 1323
rect 1876 1296 1880 1304
rect 2109 1297 2152 1303
rect 2572 1303 2580 1308
rect 2509 1297 2547 1303
rect 2557 1297 2580 1303
rect 3005 1297 3011 1317
rect 3261 1317 3299 1323
rect 3261 1297 3267 1317
rect 3549 1317 3560 1323
rect 3656 1317 3667 1323
rect 4189 1317 4259 1323
rect 4568 1317 4579 1323
rect 4669 1317 4707 1323
rect 4216 1297 4243 1303
rect 4669 1297 4675 1317
rect 5725 1317 5736 1323
rect 7293 1317 7304 1323
rect 5149 1297 5176 1303
rect 5549 1297 5571 1303
rect 5624 1297 5635 1303
rect 5677 1297 5699 1303
rect 3752 1277 3768 1283
rect 4381 1277 4392 1283
rect 7117 1277 7144 1283
rect 684 1137 707 1143
rect 2829 1137 2840 1143
rect 3181 1137 3192 1143
rect 3517 1137 3540 1143
rect 3532 1132 3540 1137
rect 3885 1137 3912 1143
rect 4685 1143 4691 1163
rect 4685 1137 4724 1143
rect 4813 1143 4819 1163
rect 4813 1137 4852 1143
rect 232 1116 236 1124
rect 253 1103 259 1123
rect 973 1117 1011 1123
rect 216 1097 227 1103
rect 253 1097 291 1103
rect 669 1097 680 1103
rect 732 1106 740 1112
rect 1149 1103 1155 1123
rect 1293 1117 1304 1123
rect 1085 1097 1155 1103
rect 1661 1103 1667 1123
rect 1661 1097 1699 1103
rect 2029 1103 2035 1123
rect 1997 1097 2035 1103
rect 2173 1103 2179 1123
rect 2312 1116 2318 1124
rect 2109 1097 2179 1103
rect 2893 1103 2899 1123
rect 2861 1097 2899 1103
rect 2925 1097 2936 1103
rect 3148 1106 3156 1112
rect 3277 1103 3283 1123
rect 3677 1117 3699 1123
rect 3800 1117 3811 1123
rect 3912 1117 3923 1123
rect 4573 1117 4595 1123
rect 5245 1117 5272 1123
rect 3245 1097 3283 1103
rect 3405 1097 3416 1103
rect 3448 1097 3459 1103
rect 3804 1103 3812 1108
rect 3804 1097 3816 1103
rect 4152 1097 4163 1103
rect 4445 1097 4483 1103
rect 4728 1097 4739 1103
rect 1256 1077 1267 1083
rect 1304 1077 1315 1083
rect 1421 1077 1448 1083
rect 1496 1077 1507 1083
rect 1661 1077 1672 1083
rect 2381 1077 2424 1083
rect 2621 1077 2660 1083
rect 2888 1077 2899 1083
rect 3208 1077 3235 1083
rect 3645 1077 3651 1092
rect 5293 1103 5299 1123
rect 5229 1097 5299 1103
rect 5485 1103 5491 1123
rect 5508 1116 5512 1124
rect 6056 1116 6060 1124
rect 6077 1117 6088 1123
rect 5453 1097 5491 1103
rect 5517 1097 5528 1103
rect 6141 1103 6147 1123
rect 6484 1116 6488 1124
rect 7096 1117 7107 1123
rect 6109 1097 6147 1103
rect 6173 1097 6200 1103
rect 6493 1097 6504 1103
rect 7080 1097 7123 1103
rect 4104 1077 4120 1083
rect 4925 1077 4936 1083
rect 5256 1077 5299 1083
rect 5533 1077 5555 1083
rect 5565 1077 5588 1083
rect 5580 1072 5588 1077
rect 5912 1077 5939 1083
rect 6344 1077 6371 1083
rect 6680 1077 6691 1083
rect 6984 1077 7011 1083
rect 3484 1068 3492 1072
rect 2509 1057 2563 1063
rect 3668 1056 3672 1064
rect 3773 1057 3784 1063
rect 3956 1056 3960 1064
rect 4429 1057 4440 1063
rect 7005 1057 7016 1063
rect 4200 1037 4232 1043
rect 4312 1037 4323 1043
rect 6317 977 6328 983
rect 6456 977 6478 983
rect 1693 957 1736 963
rect 1800 957 1811 963
rect 2189 957 2275 963
rect 2285 957 2296 963
rect 3693 957 3724 963
rect 4100 956 4104 964
rect 4148 957 4179 963
rect 5629 957 5667 963
rect 413 937 424 943
rect 461 937 483 943
rect 1101 937 1144 943
rect 1805 937 1875 943
rect 1896 937 1923 943
rect 2077 937 2088 943
rect 2296 937 2323 943
rect 2808 937 2819 943
rect 2893 937 2915 943
rect 3005 937 3027 943
rect 253 917 291 923
rect 253 897 259 917
rect 376 917 387 923
rect 936 917 947 923
rect 973 917 1011 923
rect 952 896 956 904
rect 973 897 979 917
rect 1432 917 1443 923
rect 1885 917 1896 923
rect 2061 917 2104 923
rect 2248 917 2259 923
rect 2541 917 2580 923
rect 2572 914 2580 917
rect 2781 917 2819 923
rect 1624 896 1630 904
rect 2813 897 2819 917
rect 2920 917 2931 923
rect 3021 923 3027 937
rect 3133 937 3160 943
rect 3757 943 3763 948
rect 3672 937 3683 943
rect 3741 937 3768 943
rect 4509 937 4520 943
rect 4621 937 4632 943
rect 5416 937 5427 943
rect 5884 943 5892 948
rect 5869 937 5892 943
rect 6413 937 6440 943
rect 6845 937 6883 943
rect 3021 917 3048 923
rect 3085 917 3123 923
rect 3085 897 3091 917
rect 3421 917 3459 923
rect 3421 897 3427 917
rect 4264 917 4275 923
rect 4637 917 4675 923
rect 4797 917 4808 923
rect 5005 917 5016 923
rect 5389 917 5427 923
rect 4280 896 4284 904
rect 4740 896 4744 904
rect 5421 897 5427 917
rect 5480 917 5491 923
rect 5597 917 5608 923
rect 5821 917 5832 923
rect 6397 917 6408 923
rect 6621 917 6632 923
rect 6808 917 6819 923
rect 6877 917 6883 937
rect 6925 943 6931 963
rect 7085 957 7096 963
rect 6925 937 6963 943
rect 7037 937 7091 943
rect 7176 897 7187 903
rect 7204 896 7208 904
rect 4045 877 4072 883
rect 4045 857 4051 877
rect 4205 877 4232 883
rect 3848 737 3875 743
rect 3965 737 3992 743
rect 4136 737 4179 743
rect 4712 737 4723 743
rect 36 716 40 724
rect 488 716 492 724
rect 509 703 515 723
rect 472 697 483 703
rect 509 697 547 703
rect 797 697 808 703
rect 973 703 979 723
rect 973 697 1011 703
rect 1245 703 1251 723
rect 1432 716 1436 724
rect 1176 697 1219 703
rect 1245 697 1283 703
rect 1304 697 1315 703
rect 1453 703 1459 723
rect 1416 697 1427 703
rect 1453 697 1491 703
rect 1565 703 1571 723
rect 1528 697 1539 703
rect 1565 697 1603 703
rect 2349 703 2355 723
rect 2349 697 2387 703
rect 2845 703 2851 723
rect 2808 697 2819 703
rect 2845 697 2883 703
rect 3000 697 3011 703
rect 3597 703 3603 723
rect 3773 717 3811 723
rect 3837 717 3848 723
rect 4120 717 4131 723
rect 3597 697 3635 703
rect 4349 703 4355 723
rect 4372 716 4376 724
rect 4317 697 4355 703
rect 4381 697 4392 703
rect 4653 703 4659 723
rect 4653 697 4691 703
rect 5037 703 5043 723
rect 5037 697 5075 703
rect 5085 697 5096 703
rect 1032 677 1043 683
rect 1037 657 1043 677
rect 1400 677 1411 683
rect 1565 677 1576 683
rect 2109 677 2211 683
rect 2349 677 2360 683
rect 2397 677 2408 683
rect 2845 677 2856 683
rect 3244 677 3272 683
rect 3656 677 3667 683
rect 2061 657 2072 663
rect 2136 657 2195 663
rect 3661 657 3667 677
rect 4653 677 4664 683
rect 5037 677 5048 683
rect 5085 677 5091 697
rect 5149 703 5155 723
rect 5533 717 5544 723
rect 6420 716 6424 724
rect 5149 697 5187 703
rect 5965 697 6003 703
rect 5197 677 5208 683
rect 5629 677 5640 683
rect 5997 677 6003 697
rect 6584 697 6611 703
rect 6477 677 6500 683
rect 6492 672 6500 677
rect 7117 657 7155 663
rect 2152 556 2156 564
rect 5148 557 5171 563
rect 5148 554 5156 557
rect 908 543 916 548
rect 908 537 931 543
rect 1528 537 1539 543
rect 3357 537 3368 543
rect 4173 537 4195 543
rect 4621 537 4632 543
rect 5181 537 5203 543
rect 6492 543 6500 548
rect 6408 537 6419 543
rect 6477 537 6500 543
rect 6968 537 6979 543
rect 7421 537 7432 543
rect 109 517 147 523
rect 109 497 115 517
rect 429 517 467 523
rect 408 496 412 504
rect 429 497 435 517
rect 701 517 712 523
rect 968 517 995 523
rect 1389 517 1416 523
rect 1992 517 2003 523
rect 2109 517 2136 523
rect 2573 517 2616 523
rect 2909 517 2920 523
rect 3320 517 3331 523
rect 3757 517 3795 523
rect 552 497 563 503
rect 1821 497 1859 503
rect 2564 496 2568 504
rect 3757 497 3763 517
rect 3992 517 4003 523
rect 4429 517 4472 523
rect 4621 517 4659 523
rect 4093 497 4104 503
rect 4509 497 4547 503
rect 4621 497 4627 517
rect 5245 517 5315 523
rect 5245 497 5251 517
rect 6152 517 6163 523
rect 6189 517 6227 523
rect 6189 497 6195 517
rect 6328 517 6339 523
rect 6333 497 6339 517
rect 6808 517 6836 523
rect 6989 517 7016 523
rect 6828 516 6836 517
rect 6356 496 6360 504
rect 7108 496 7112 504
rect 189 337 200 343
rect 77 297 88 303
rect 253 303 259 323
rect 221 297 259 303
rect 285 297 312 303
rect 461 297 472 303
rect 781 303 787 323
rect 804 316 808 324
rect 749 297 787 303
rect 813 297 824 303
rect 1208 297 1219 303
rect 248 277 259 283
rect 349 277 371 283
rect 365 268 371 277
rect 653 277 675 283
rect 1069 277 1080 283
rect 1213 283 1219 297
rect 1517 303 1523 323
rect 1896 316 1900 324
rect 1517 297 1555 303
rect 1581 297 1603 303
rect 1213 277 1235 283
rect 1581 283 1587 297
rect 1917 303 1923 323
rect 2392 316 2396 324
rect 1880 297 1891 303
rect 1917 297 1955 303
rect 2237 297 2248 303
rect 2413 303 2419 323
rect 2792 316 2796 324
rect 2376 297 2387 303
rect 2413 297 2451 303
rect 2477 297 2499 303
rect 1576 277 1587 283
rect 2477 283 2483 297
rect 2813 303 2819 323
rect 2893 317 2904 323
rect 2813 297 2851 303
rect 2909 297 2936 303
rect 2472 277 2483 283
rect 2861 277 2872 283
rect 2909 277 2915 297
rect 3261 303 3267 323
rect 3229 297 3267 303
rect 3373 303 3379 323
rect 3336 297 3347 303
rect 3373 297 3411 303
rect 3773 303 3779 323
rect 4221 317 4291 323
rect 3544 297 3555 303
rect 3741 297 3779 303
rect 3805 297 3816 303
rect 4365 303 4371 323
rect 5661 317 5699 323
rect 4365 297 4403 303
rect 5416 297 5427 303
rect 5437 297 5448 303
rect 5501 297 5539 303
rect 5501 288 5507 297
rect 5645 297 5672 303
rect 5965 303 5971 323
rect 5965 297 6003 303
rect 6317 303 6323 323
rect 6317 297 6344 303
rect 6381 303 6387 323
rect 6692 316 6696 324
rect 7028 316 7032 324
rect 6381 297 6419 303
rect 6701 297 6712 303
rect 7341 303 7347 323
rect 7309 297 7347 303
rect 3192 277 3219 283
rect 3256 277 3267 283
rect 3309 277 3320 283
rect 3373 277 3384 283
rect 3720 277 3731 283
rect 3853 277 3875 283
rect 4248 277 4275 283
rect 4413 277 4424 283
rect 4984 277 4995 283
rect 5096 277 5107 283
rect 5149 277 5192 283
rect 5581 277 5619 283
rect 5965 277 5976 283
rect 6045 277 6068 283
rect 6060 272 6068 277
rect 6328 277 6339 283
rect 6717 277 6739 283
rect 6749 277 6772 283
rect 6764 272 6772 277
rect 7053 277 7075 283
rect 7085 277 7108 283
rect 7100 272 7108 277
rect 5165 257 5203 263
rect 5197 243 5203 257
rect 5197 237 5219 243
rect 5869 157 5892 163
rect 5884 154 5892 157
rect 6264 157 6291 163
rect 6301 157 6324 163
rect 6316 154 6324 157
rect 1628 148 1636 152
rect 696 137 707 143
rect 1352 137 1379 143
rect 1533 137 1544 143
rect 1596 143 1604 148
rect 1581 137 1604 143
rect 2476 137 2500 143
rect 2760 137 2771 143
rect 3208 137 3251 143
rect 4781 137 4792 143
rect 4844 143 4852 148
rect 4829 137 4852 143
rect 5592 137 5619 143
rect 5725 137 5736 143
rect 5848 137 5859 143
rect 6060 137 6099 143
rect 6216 137 6227 143
rect 6237 137 6264 143
rect 6716 143 6724 148
rect 6669 137 6691 143
rect 6701 137 6724 143
rect 269 117 280 123
rect 408 117 419 123
rect 669 117 707 123
rect 701 97 707 117
rect 1325 117 1352 123
rect 1533 117 1571 123
rect 1005 97 1043 103
rect 1533 97 1539 117
rect 2269 117 2280 123
rect 2733 117 2771 123
rect 2141 97 2184 103
rect 2205 97 2243 103
rect 2260 96 2264 104
rect 2765 97 2771 117
rect 3069 117 3107 123
rect 3069 97 3075 117
rect 3165 117 3224 123
rect 3581 117 3592 123
rect 4013 117 4051 123
rect 3181 97 3192 103
rect 4045 97 4051 117
rect 4413 117 4440 123
rect 4744 117 4755 123
rect 4781 117 4819 123
rect 4429 97 4467 103
rect 4781 97 4787 117
rect 5416 117 5427 123
rect 5645 117 5656 123
rect 5757 117 5795 123
rect 5789 97 5795 117
rect 6184 117 6211 123
rect 5812 96 5816 104
rect 6164 96 6168 104
rect 6205 97 6211 117
rect 6424 117 6435 123
rect 6589 117 6627 123
rect 6621 97 6627 117
rect 6644 96 6648 104
rect 5165 37 5192 43
<< m2contact >>
rect 2157 5402 2193 5418
rect 4205 5402 4241 5418
rect 6237 5402 6273 5418
rect 296 5372 312 5388
rect 664 5372 680 5388
rect 1512 5372 1528 5388
rect 1944 5372 1960 5388
rect 2888 5372 2904 5388
rect 3048 5372 3080 5388
rect 3112 5372 3128 5388
rect 3192 5372 3208 5388
rect 3640 5372 3656 5388
rect 4008 5372 4024 5388
rect 3384 5352 3400 5368
rect 4344 5372 4376 5388
rect 4568 5372 4584 5388
rect 6184 5372 6200 5388
rect 6680 5372 6696 5388
rect 6392 5352 6408 5368
rect 56 5332 72 5348
rect 104 5332 120 5348
rect 600 5332 616 5348
rect 824 5332 840 5348
rect 856 5332 872 5348
rect 888 5332 904 5348
rect 952 5332 968 5348
rect 1032 5332 1048 5348
rect 1288 5332 1304 5348
rect 1320 5332 1336 5348
rect 1384 5332 1416 5348
rect 1496 5332 1512 5348
rect 1672 5332 1688 5348
rect 1736 5332 1752 5348
rect 1960 5332 1976 5348
rect 1992 5332 2008 5348
rect 2056 5332 2072 5348
rect 2120 5332 2136 5348
rect 2296 5332 2312 5348
rect 2360 5332 2376 5348
rect 2408 5332 2424 5348
rect 2664 5332 2680 5348
rect 3000 5332 3016 5348
rect 3352 5332 3368 5348
rect 3512 5332 3528 5348
rect 3576 5332 3608 5348
rect 3624 5332 3640 5348
rect 3832 5332 3848 5348
rect 3928 5332 3944 5348
rect 3960 5332 3976 5348
rect 4072 5332 4088 5348
rect 4520 5332 4536 5348
rect 4552 5332 4568 5348
rect 4632 5332 4648 5348
rect 4680 5332 4712 5348
rect 4744 5332 4760 5348
rect 4840 5332 4856 5348
rect 5064 5332 5080 5348
rect 5192 5332 5208 5348
rect 5448 5332 5464 5348
rect 5528 5332 5544 5348
rect 5576 5332 5592 5348
rect 5880 5332 5896 5348
rect 5912 5332 5928 5348
rect 5976 5332 5992 5348
rect 6008 5332 6040 5348
rect 6120 5332 6152 5348
rect 6184 5332 6200 5348
rect 6360 5332 6376 5348
rect 6584 5332 6600 5348
rect 6648 5332 6664 5348
rect 6776 5332 6792 5348
rect 6888 5332 6920 5348
rect 6936 5352 6952 5368
rect 7208 5352 7224 5368
rect 7336 5352 7352 5368
rect 7064 5332 7080 5348
rect 7208 5332 7224 5348
rect 72 5312 88 5328
rect 184 5312 200 5328
rect 232 5312 248 5328
rect 376 5312 408 5328
rect 504 5312 536 5328
rect 648 5312 664 5328
rect 792 5314 808 5330
rect 8 5292 24 5308
rect 40 5292 56 5308
rect 72 5292 104 5308
rect 888 5292 904 5308
rect 936 5312 952 5328
rect 1048 5312 1064 5328
rect 1192 5312 1224 5328
rect 1272 5312 1288 5328
rect 1320 5292 1336 5308
rect 1368 5312 1384 5328
rect 1432 5292 1448 5308
rect 1480 5312 1496 5328
rect 1624 5312 1640 5328
rect 1704 5312 1720 5328
rect 1832 5312 1848 5328
rect 1976 5312 1992 5328
rect 1480 5292 1496 5308
rect 2168 5312 2184 5328
rect 2200 5312 2216 5328
rect 2312 5312 2328 5328
rect 2024 5292 2040 5308
rect 2424 5312 2440 5328
rect 2472 5312 2504 5328
rect 2568 5312 2584 5328
rect 2616 5312 2632 5328
rect 2744 5312 2760 5328
rect 2808 5312 2824 5328
rect 2872 5312 2888 5328
rect 2936 5312 2952 5328
rect 3016 5312 3032 5328
rect 3096 5312 3112 5328
rect 3144 5312 3160 5328
rect 3304 5312 3320 5328
rect 3432 5312 3448 5328
rect 2360 5292 2376 5308
rect 3592 5312 3608 5328
rect 3736 5312 3752 5328
rect 3784 5312 3800 5328
rect 3992 5312 4008 5328
rect 4040 5312 4056 5328
rect 4120 5312 4136 5328
rect 4312 5312 4328 5328
rect 4488 5314 4504 5330
rect 4648 5312 4680 5328
rect 4696 5312 4712 5328
rect 3480 5292 3496 5308
rect 3528 5292 3544 5308
rect 3560 5292 3576 5308
rect 3592 5292 3608 5308
rect 3880 5292 3896 5308
rect 4584 5292 4600 5308
rect 4604 5292 4620 5308
rect 4648 5292 4664 5308
rect 4744 5292 4760 5308
rect 4776 5292 4792 5308
rect 4808 5312 4840 5328
rect 4904 5314 4920 5330
rect 4968 5312 4984 5328
rect 5080 5312 5096 5328
rect 5192 5312 5208 5328
rect 5288 5314 5304 5330
rect 5352 5312 5368 5328
rect 5464 5312 5480 5328
rect 5560 5312 5576 5328
rect 5144 5292 5160 5308
rect 5176 5292 5192 5308
rect 5496 5292 5512 5308
rect 5576 5292 5592 5308
rect 5608 5292 5624 5308
rect 5640 5312 5672 5328
rect 5832 5312 5848 5328
rect 5944 5292 5960 5308
rect 5992 5312 6008 5328
rect 6056 5292 6072 5308
rect 6120 5312 6136 5328
rect 6312 5312 6328 5328
rect 6536 5312 6552 5328
rect 6616 5312 6632 5328
rect 6744 5312 6760 5328
rect 6808 5314 6824 5330
rect 6872 5312 6888 5328
rect 6968 5312 6984 5328
rect 7048 5312 7064 5328
rect 7224 5312 7240 5328
rect 7304 5312 7320 5328
rect 7352 5312 7368 5328
rect 6104 5292 6120 5308
rect 264 5272 280 5288
rect 1144 5272 1160 5288
rect 1912 5272 1928 5288
rect 2504 5272 2520 5288
rect 3432 5272 3448 5288
rect 4712 5272 4728 5288
rect 5752 5272 5768 5288
rect 360 5232 376 5248
rect 584 5232 600 5248
rect 616 5232 632 5248
rect 1240 5232 1256 5248
rect 2280 5232 2296 5248
rect 2456 5232 2472 5248
rect 2712 5232 2728 5248
rect 2776 5232 2792 5248
rect 2840 5232 2856 5248
rect 2984 5232 3000 5248
rect 3400 5232 3416 5248
rect 3912 5232 3928 5248
rect 4296 5232 4312 5248
rect 5064 5232 5080 5248
rect 5112 5232 5128 5248
rect 5448 5232 5464 5248
rect 5688 5232 5704 5248
rect 7160 5232 7176 5248
rect 7272 5232 7288 5248
rect 7320 5232 7336 5248
rect 7384 5232 7400 5248
rect 1117 5202 1153 5218
rect 3165 5202 3201 5218
rect 5213 5202 5249 5218
rect 520 5172 536 5188
rect 1032 5172 1048 5188
rect 1448 5172 1464 5188
rect 2392 5172 2408 5188
rect 3480 5172 3496 5188
rect 3720 5172 3736 5188
rect 3768 5172 3784 5188
rect 3848 5172 3864 5188
rect 3896 5172 3912 5188
rect 3976 5172 3992 5188
rect 4328 5172 4344 5188
rect 376 5132 392 5148
rect 408 5132 424 5148
rect 1304 5132 1320 5148
rect 4392 5132 4408 5148
rect 5832 5132 5848 5148
rect 5880 5132 5896 5148
rect 6200 5132 6216 5148
rect 136 5090 152 5106
rect 280 5092 296 5108
rect 408 5092 424 5108
rect 456 5112 472 5128
rect 520 5092 536 5108
rect 568 5112 584 5128
rect 616 5092 648 5108
rect 680 5092 696 5108
rect 728 5092 744 5108
rect 776 5112 792 5128
rect 1336 5112 1352 5128
rect 904 5092 920 5108
rect 1064 5092 1080 5108
rect 1176 5092 1192 5108
rect 1372 5112 1388 5128
rect 1704 5112 1720 5128
rect 1384 5092 1400 5108
rect 1416 5092 1432 5108
rect 1544 5092 1560 5108
rect 1608 5090 1624 5106
rect 1752 5092 1768 5108
rect 1800 5092 1816 5108
rect 1848 5112 1864 5128
rect 2136 5112 2152 5128
rect 2424 5112 2440 5128
rect 1960 5092 1976 5108
rect 2104 5092 2120 5108
rect 2168 5092 2184 5108
rect 2248 5092 2264 5108
rect 2392 5092 2408 5108
rect 2456 5092 2472 5108
rect 2504 5112 2520 5128
rect 2584 5112 2600 5128
rect 2904 5112 2920 5128
rect 3800 5112 3816 5128
rect 4360 5112 4376 5128
rect 2632 5092 2648 5108
rect 2728 5092 2744 5108
rect 2872 5092 2904 5108
rect 2984 5092 3000 5108
rect 3304 5092 3320 5108
rect 3384 5092 3400 5108
rect 3448 5092 3464 5108
rect 3608 5092 3624 5108
rect 3688 5092 3704 5108
rect 3736 5092 3752 5108
rect 3880 5092 3896 5108
rect 3928 5092 3960 5108
rect 4056 5092 4072 5108
rect 4216 5092 4232 5108
rect 4296 5092 4312 5108
rect 264 5072 280 5088
rect 392 5072 408 5088
rect 488 5072 520 5088
rect 600 5072 616 5088
rect 712 5072 728 5088
rect 776 5072 792 5088
rect 808 5072 824 5088
rect 840 5072 856 5088
rect 1032 5072 1048 5088
rect 1128 5072 1144 5088
rect 1304 5072 1320 5088
rect 1400 5072 1416 5088
rect 1672 5072 1688 5088
rect 1720 5072 1736 5088
rect 1768 5072 1800 5088
rect 1848 5072 1864 5088
rect 1880 5072 1896 5088
rect 1912 5072 1928 5088
rect 2088 5072 2104 5088
rect 2200 5072 2216 5088
rect 2376 5072 2392 5088
rect 2440 5072 2456 5088
rect 2504 5072 2520 5088
rect 2536 5072 2568 5088
rect 2648 5072 2664 5088
rect 2680 5072 2696 5088
rect 2760 5072 2776 5088
rect 2856 5072 2872 5088
rect 2968 5072 2984 5088
rect 3112 5072 3128 5088
rect 3352 5072 3368 5088
rect 3656 5072 3672 5088
rect 3784 5072 3800 5088
rect 3832 5072 3848 5088
rect 4072 5072 4088 5088
rect 4104 5072 4120 5088
rect 4232 5072 4248 5088
rect 4296 5072 4312 5088
rect 4328 5092 4344 5108
rect 4360 5092 4376 5108
rect 4440 5112 4456 5128
rect 4472 5112 4488 5128
rect 4504 5112 4520 5128
rect 4824 5112 4840 5128
rect 4872 5112 4888 5128
rect 4920 5112 4936 5128
rect 4648 5092 4664 5108
rect 4776 5092 4792 5108
rect 4968 5112 4984 5128
rect 5560 5112 5576 5128
rect 6072 5112 6088 5128
rect 4968 5092 4984 5108
rect 5048 5090 5064 5106
rect 5112 5092 5128 5108
rect 5192 5092 5208 5108
rect 5320 5092 5336 5108
rect 5384 5090 5400 5106
rect 5480 5092 5496 5108
rect 5544 5092 5560 5108
rect 5576 5092 5608 5108
rect 5720 5092 5736 5108
rect 5912 5092 5928 5108
rect 5960 5092 5976 5108
rect 6120 5092 6136 5108
rect 6280 5092 6296 5108
rect 6328 5092 6344 5108
rect 6440 5092 6456 5108
rect 6504 5092 6520 5108
rect 6568 5090 6584 5106
rect 6776 5092 6792 5108
rect 6824 5092 6840 5108
rect 6968 5092 6984 5108
rect 7032 5090 7048 5106
rect 7128 5092 7144 5108
rect 7192 5092 7208 5108
rect 7240 5092 7256 5108
rect 7304 5092 7336 5108
rect 7384 5092 7400 5108
rect 4376 5072 4392 5088
rect 4488 5072 4504 5088
rect 4520 5072 4536 5088
rect 4728 5072 4744 5088
rect 4792 5072 4808 5088
rect 4840 5072 4856 5088
rect 4888 5072 4904 5088
rect 4984 5072 5000 5088
rect 5416 5072 5432 5088
rect 5480 5072 5496 5088
rect 5528 5072 5544 5088
rect 5640 5072 5656 5088
rect 5672 5072 5688 5088
rect 6008 5072 6024 5088
rect 6040 5072 6056 5088
rect 6104 5072 6120 5088
rect 6200 5072 6216 5088
rect 6376 5072 6392 5088
rect 6488 5072 6504 5088
rect 6536 5072 6552 5088
rect 6872 5072 6888 5088
rect 7176 5072 7192 5088
rect 7288 5072 7320 5088
rect 5448 5052 5464 5068
rect 6408 5052 6424 5068
rect 6472 5052 6488 5068
rect 7096 5052 7112 5068
rect 7208 5052 7224 5068
rect 7416 5052 7432 5068
rect 8 5032 24 5048
rect 664 5032 680 5048
rect 1000 5032 1016 5048
rect 1288 5032 1304 5048
rect 1480 5032 1496 5048
rect 2072 5032 2088 5048
rect 2360 5032 2376 5048
rect 2600 5032 2616 5048
rect 2840 5032 2856 5048
rect 3096 5032 3112 5048
rect 3144 5032 3160 5048
rect 3192 5032 3208 5048
rect 3416 5032 3432 5048
rect 3496 5032 3512 5048
rect 3816 5032 3832 5048
rect 4536 5032 4552 5048
rect 4824 5032 4840 5048
rect 4872 5032 4888 5048
rect 5256 5032 5272 5048
rect 5624 5032 5640 5048
rect 5848 5032 5864 5048
rect 6152 5032 6168 5048
rect 6696 5032 6728 5048
rect 6904 5032 6920 5048
rect 7160 5032 7176 5048
rect 7272 5032 7288 5048
rect 7352 5032 7368 5048
rect 2157 5002 2193 5018
rect 4205 5002 4241 5018
rect 6237 5002 6273 5018
rect 760 4972 776 4988
rect 904 4972 920 4988
rect 1256 4972 1272 4988
rect 1864 4972 1880 4988
rect 2120 4972 2136 4988
rect 2328 4972 2344 4988
rect 2456 4972 2472 4988
rect 2600 4972 2616 4988
rect 2904 4972 2920 4988
rect 2952 4972 2968 4988
rect 3032 4972 3048 4988
rect 3112 4972 3128 4988
rect 3608 4972 3624 4988
rect 3704 4972 3720 4988
rect 3976 4972 3992 4988
rect 4424 4972 4440 4988
rect 4600 4972 4616 4988
rect 5688 4972 5704 4988
rect 5784 4972 5800 4988
rect 5944 4972 5960 4988
rect 6280 4972 6296 4988
rect 6504 4972 6520 4988
rect 7032 4972 7048 4988
rect 7416 4972 7432 4988
rect 264 4952 280 4968
rect 456 4952 472 4968
rect 1128 4952 1144 4968
rect 4104 4952 4120 4968
rect 4504 4952 4520 4968
rect 4728 4952 4744 4968
rect 5224 4952 5240 4968
rect 5480 4952 5496 4968
rect 5640 4952 5656 4968
rect 5720 4952 5736 4968
rect 5832 4952 5848 4968
rect 6136 4952 6152 4968
rect 6568 4952 6584 4968
rect 104 4932 120 4948
rect 136 4932 152 4948
rect 200 4932 216 4948
rect 408 4932 424 4948
rect 504 4932 552 4948
rect 648 4932 664 4948
rect 776 4932 792 4948
rect 808 4932 824 4948
rect 840 4932 856 4948
rect 1352 4932 1368 4948
rect 1400 4932 1416 4948
rect 1464 4932 1480 4948
rect 1640 4932 1656 4948
rect 1672 4932 1688 4948
rect 1704 4932 1720 4948
rect 1880 4932 1896 4948
rect 1944 4932 1960 4948
rect 1992 4932 2008 4948
rect 2312 4932 2328 4948
rect 2344 4932 2360 4948
rect 2488 4932 2504 4948
rect 8 4912 24 4928
rect 72 4912 104 4928
rect 136 4892 152 4908
rect 184 4912 200 4928
rect 280 4912 296 4928
rect 440 4892 456 4908
rect 504 4912 520 4928
rect 568 4912 584 4928
rect 680 4912 696 4928
rect 792 4912 808 4928
rect 936 4912 984 4928
rect 1032 4912 1048 4928
rect 1144 4912 1160 4928
rect 1272 4912 1304 4928
rect 872 4892 888 4908
rect 1400 4892 1416 4908
rect 1480 4912 1512 4928
rect 1544 4912 1576 4928
rect 1640 4912 1672 4928
rect 1752 4912 1768 4928
rect 1880 4912 1896 4928
rect 1576 4892 1592 4908
rect 1608 4892 1624 4908
rect 1640 4892 1656 4908
rect 2008 4912 2024 4928
rect 2056 4912 2088 4928
rect 2184 4912 2200 4928
rect 2232 4912 2248 4928
rect 2360 4912 2392 4928
rect 2424 4912 2440 4928
rect 2920 4932 2936 4948
rect 3064 4932 3080 4948
rect 3192 4932 3208 4948
rect 3224 4932 3240 4948
rect 3432 4932 3448 4948
rect 3496 4932 3512 4948
rect 3544 4932 3576 4948
rect 3656 4932 3672 4948
rect 3720 4932 3736 4948
rect 3816 4932 3832 4948
rect 3880 4932 3912 4948
rect 4168 4932 4184 4948
rect 4200 4932 4216 4948
rect 4296 4932 4312 4948
rect 4360 4932 4392 4948
rect 4504 4932 4520 4948
rect 4792 4932 4824 4948
rect 4872 4932 4904 4948
rect 4920 4932 4936 4948
rect 5320 4932 5336 4948
rect 5416 4932 5432 4948
rect 5800 4932 5816 4948
rect 5912 4932 5928 4948
rect 6008 4932 6024 4948
rect 6216 4932 6232 4948
rect 6376 4932 6392 4948
rect 6488 4932 6504 4948
rect 7144 4932 7160 4948
rect 2568 4912 2600 4928
rect 2664 4912 2696 4928
rect 2792 4912 2824 4928
rect 2856 4912 2872 4928
rect 2984 4912 3000 4928
rect 3080 4912 3096 4928
rect 1944 4892 1960 4908
rect 2312 4892 2328 4908
rect 2456 4892 2472 4908
rect 2888 4892 2904 4908
rect 3272 4912 3288 4928
rect 3128 4892 3144 4908
rect 3432 4892 3448 4908
rect 3480 4912 3496 4928
rect 3512 4892 3528 4908
rect 3592 4892 3608 4908
rect 3640 4912 3656 4928
rect 3672 4912 3688 4928
rect 3736 4912 3768 4928
rect 3864 4912 3880 4928
rect 4104 4914 4120 4930
rect 3784 4892 3800 4908
rect 3832 4892 3848 4908
rect 4200 4892 4216 4908
rect 4280 4912 4296 4928
rect 4312 4912 4328 4928
rect 4408 4892 4424 4908
rect 4456 4912 4472 4928
rect 4664 4912 4680 4928
rect 4728 4914 4744 4930
rect 4840 4912 4872 4928
rect 4984 4912 5000 4928
rect 5032 4912 5048 4928
rect 5208 4912 5224 4928
rect 4824 4892 4840 4908
rect 4920 4892 4936 4908
rect 5000 4892 5016 4908
rect 5032 4892 5048 4908
rect 5352 4892 5368 4908
rect 5400 4912 5416 4928
rect 5480 4914 5496 4930
rect 5656 4912 5672 4928
rect 5752 4912 5768 4928
rect 5816 4912 5832 4928
rect 5864 4912 5880 4928
rect 5896 4912 5912 4928
rect 5928 4912 5944 4928
rect 6024 4912 6040 4928
rect 6168 4912 6184 4928
rect 6200 4912 6216 4928
rect 6232 4912 6248 4928
rect 6392 4912 6408 4928
rect 6472 4912 6488 4928
rect 6536 4912 6552 4928
rect 6600 4912 6616 4928
rect 6680 4912 6696 4928
rect 6744 4912 6760 4928
rect 6808 4912 6824 4928
rect 6872 4912 6888 4928
rect 6936 4912 6952 4928
rect 7000 4912 7016 4928
rect 7160 4914 7176 4930
rect 7288 4912 7304 4928
rect 5400 4892 5416 4908
rect 6632 4892 6648 4908
rect 6696 4892 6712 4908
rect 6760 4892 6776 4908
rect 6824 4892 6840 4908
rect 6888 4892 6904 4908
rect 6952 4892 6968 4908
rect 7016 4892 7032 4908
rect 408 4872 424 4888
rect 3912 4872 3928 4888
rect 4888 4872 4904 4888
rect 6664 4872 6680 4888
rect 6728 4872 6744 4888
rect 6792 4872 6808 4888
rect 6856 4872 6872 4888
rect 6952 4872 6968 4888
rect 6984 4872 7000 4888
rect 56 4832 72 4848
rect 392 4832 408 4848
rect 1000 4832 1016 4848
rect 1320 4832 1336 4848
rect 1512 4832 1528 4848
rect 2024 4832 2040 4848
rect 2408 4832 2424 4848
rect 2536 4832 2552 4848
rect 2824 4832 2840 4848
rect 3032 4832 3048 4848
rect 3384 4832 3400 4848
rect 3528 4832 3544 4848
rect 3864 4832 3880 4848
rect 4488 4832 4504 4848
rect 4568 4832 4584 4848
rect 5064 4832 5080 4848
rect 6584 4832 6600 4848
rect 6744 4832 6760 4848
rect 6808 4832 6824 4848
rect 6872 4832 6888 4848
rect 6936 4832 6952 4848
rect 7000 4832 7016 4848
rect 1117 4802 1153 4818
rect 3165 4802 3201 4818
rect 5213 4802 5249 4818
rect 8 4772 24 4788
rect 1816 4772 1832 4788
rect 3224 4772 3240 4788
rect 3368 4772 3384 4788
rect 3400 4772 3416 4788
rect 3608 4772 3624 4788
rect 3720 4772 3736 4788
rect 4232 4772 4248 4788
rect 4440 4772 4456 4788
rect 4488 4772 4504 4788
rect 4760 4772 4776 4788
rect 4792 4772 4808 4788
rect 5672 4772 5688 4788
rect 6552 4772 6568 4788
rect 6600 4772 6616 4788
rect 6664 4772 6680 4788
rect 6968 4772 6984 4788
rect 1608 4752 1624 4768
rect 2680 4752 2696 4768
rect 856 4732 872 4748
rect 1464 4732 1480 4748
rect 3240 4732 3256 4748
rect 3336 4732 3368 4748
rect 3416 4732 3432 4748
rect 3624 4732 3640 4748
rect 3736 4732 3752 4748
rect 3768 4732 3784 4748
rect 4248 4732 4264 4748
rect 4456 4732 4472 4748
rect 5368 4752 5384 4768
rect 5752 4752 5768 4768
rect 5320 4732 5336 4748
rect 5384 4732 5400 4748
rect 5560 4732 5576 4748
rect 5688 4732 5704 4748
rect 5768 4732 5784 4748
rect 5816 4732 5832 4748
rect 7128 4752 7144 4768
rect 6440 4732 6456 4748
rect 6488 4732 6504 4748
rect 6568 4732 6584 4748
rect 6616 4732 6632 4748
rect 6680 4732 6712 4748
rect 6744 4732 6760 4748
rect 6824 4732 6840 4748
rect 6872 4732 6888 4748
rect 6952 4732 6968 4748
rect 7016 4732 7032 4748
rect 7064 4732 7080 4748
rect 7144 4732 7160 4748
rect 232 4712 248 4728
rect 136 4690 152 4706
rect 268 4712 284 4728
rect 568 4712 584 4728
rect 632 4712 648 4728
rect 280 4692 296 4708
rect 376 4692 392 4708
rect 552 4692 568 4708
rect 632 4692 664 4708
rect 744 4692 760 4708
rect 888 4692 920 4708
rect 936 4712 952 4728
rect 984 4712 1000 4728
rect 1048 4712 1064 4728
rect 1080 4712 1096 4728
rect 1528 4712 1544 4728
rect 1016 4692 1032 4708
rect 1096 4692 1112 4708
rect 1208 4692 1224 4708
rect 1304 4692 1320 4708
rect 1352 4692 1368 4708
rect 1384 4692 1400 4708
rect 1416 4692 1432 4708
rect 1448 4692 1464 4708
rect 1864 4712 1880 4728
rect 1928 4712 1944 4728
rect 2264 4712 2280 4728
rect 2552 4712 2568 4728
rect 2632 4712 2648 4728
rect 2808 4712 2824 4728
rect 3160 4712 3176 4728
rect 3208 4712 3224 4728
rect 3320 4712 3336 4728
rect 3384 4712 3400 4728
rect 3528 4712 3560 4728
rect 3592 4712 3608 4728
rect 3688 4712 3720 4728
rect 4216 4712 4232 4728
rect 4312 4712 4344 4728
rect 4408 4712 4440 4728
rect 4888 4712 4904 4728
rect 5128 4712 5144 4728
rect 5208 4712 5224 4728
rect 5256 4712 5272 4728
rect 5352 4712 5368 4728
rect 5592 4712 5608 4728
rect 5656 4712 5672 4728
rect 5720 4712 5736 4728
rect 5848 4712 5864 4728
rect 6104 4712 6120 4728
rect 6168 4712 6184 4728
rect 6408 4712 6424 4728
rect 6472 4712 6488 4728
rect 6552 4712 6568 4728
rect 6648 4712 6664 4728
rect 6712 4712 6728 4728
rect 6776 4712 6808 4728
rect 6856 4712 6872 4728
rect 6920 4712 6936 4728
rect 6984 4712 7000 4728
rect 7048 4712 7064 4728
rect 7128 4712 7144 4728
rect 1576 4692 1592 4708
rect 1720 4692 1736 4708
rect 1848 4692 1864 4708
rect 1896 4692 1912 4708
rect 1928 4692 1944 4708
rect 1960 4692 1976 4708
rect 2056 4692 2072 4708
rect 2104 4692 2120 4708
rect 2216 4692 2264 4708
rect 2344 4692 2360 4708
rect 2440 4692 2472 4708
rect 2520 4692 2536 4708
rect 2552 4692 2568 4708
rect 2600 4692 2616 4708
rect 2680 4692 2712 4708
rect 2776 4692 2792 4708
rect 2808 4692 2824 4708
rect 2840 4692 2856 4708
rect 2952 4692 2968 4708
rect 3128 4692 3144 4708
rect 3224 4692 3240 4708
rect 3336 4692 3352 4708
rect 3400 4692 3416 4708
rect 3496 4692 3512 4708
rect 3608 4692 3624 4708
rect 3720 4692 3736 4708
rect 3880 4692 3896 4708
rect 4040 4690 4056 4706
rect 4232 4692 4248 4708
rect 4440 4692 4456 4708
rect 4520 4692 4536 4708
rect 4632 4692 4648 4708
rect 4728 4692 4744 4708
rect 4824 4692 4840 4708
rect 4856 4692 4872 4708
rect 4888 4692 4904 4708
rect 5000 4692 5016 4708
rect 5048 4692 5064 4708
rect 5192 4692 5208 4708
rect 5304 4692 5320 4708
rect 5368 4692 5384 4708
rect 5464 4692 5480 4708
rect 5560 4692 5576 4708
rect 5608 4692 5624 4708
rect 5704 4692 5720 4708
rect 5752 4692 5768 4708
rect 5832 4692 5848 4708
rect 5896 4692 5912 4708
rect 5976 4692 5992 4708
rect 6056 4692 6072 4708
rect 6136 4692 6152 4708
rect 6232 4692 6248 4708
rect 6360 4692 6376 4708
rect 6424 4692 6440 4708
rect 6504 4692 6520 4708
rect 6552 4692 6568 4708
rect 6632 4692 6648 4708
rect 6696 4692 6712 4708
rect 6760 4692 6776 4708
rect 6808 4692 6824 4708
rect 6872 4692 6888 4708
rect 6936 4692 6952 4708
rect 7000 4692 7016 4708
rect 7080 4692 7096 4708
rect 7128 4692 7144 4708
rect 7176 4692 7192 4708
rect 7304 4692 7320 4708
rect 168 4672 184 4688
rect 200 4672 216 4688
rect 296 4672 312 4688
rect 424 4672 440 4688
rect 504 4672 520 4688
rect 568 4672 584 4688
rect 616 4672 632 4688
rect 664 4672 680 4688
rect 696 4672 712 4688
rect 872 4672 888 4688
rect 968 4672 984 4688
rect 1032 4672 1048 4688
rect 1144 4672 1160 4688
rect 1224 4672 1240 4688
rect 984 4652 1000 4668
rect 1304 4672 1320 4688
rect 1368 4672 1384 4688
rect 1432 4686 1448 4688
rect 1416 4672 1448 4686
rect 1496 4672 1512 4688
rect 1560 4672 1576 4688
rect 1592 4672 1608 4688
rect 1704 4672 1720 4688
rect 1880 4672 1896 4688
rect 1912 4672 1928 4688
rect 1976 4672 1992 4688
rect 2184 4672 2216 4688
rect 2488 4672 2504 4688
rect 2568 4672 2600 4688
rect 2744 4672 2776 4688
rect 2824 4672 2840 4688
rect 2872 4672 2888 4688
rect 2904 4672 2920 4688
rect 3000 4672 3016 4688
rect 3272 4672 3288 4688
rect 3512 4672 3528 4688
rect 3576 4672 3592 4688
rect 3656 4672 3672 4688
rect 3912 4672 3928 4688
rect 4280 4672 4296 4688
rect 4360 4672 4376 4688
rect 4664 4672 4680 4688
rect 4840 4672 4856 4688
rect 5176 4672 5208 4688
rect 5448 4672 5464 4688
rect 5512 4672 5528 4688
rect 5608 4672 5624 4688
rect 5880 4672 5896 4688
rect 5928 4672 5944 4688
rect 5960 4672 5976 4688
rect 6040 4672 6056 4688
rect 6088 4672 6104 4688
rect 6120 4672 6136 4688
rect 6216 4672 6232 4688
rect 6344 4672 6360 4688
rect 6376 4672 6392 4688
rect 7000 4672 7016 4688
rect 1416 4670 1432 4672
rect 1272 4652 1288 4668
rect 1320 4652 1336 4668
rect 1480 4652 1496 4668
rect 2376 4652 2392 4668
rect 2408 4652 2424 4668
rect 2472 4652 2504 4668
rect 2632 4652 2664 4668
rect 2872 4652 2888 4668
rect 3448 4652 3464 4668
rect 5416 4652 5432 4668
rect 5960 4652 5976 4668
rect 6808 4652 6824 4668
rect 7208 4652 7224 4668
rect 7272 4652 7288 4668
rect 8 4632 24 4648
rect 488 4632 504 4648
rect 1224 4632 1240 4648
rect 1928 4632 1944 4648
rect 1992 4632 2008 4648
rect 2360 4632 2376 4648
rect 3064 4632 3080 4648
rect 3192 4632 3208 4648
rect 3288 4632 3304 4648
rect 3560 4632 3576 4648
rect 3688 4632 3704 4648
rect 4168 4632 4184 4648
rect 4312 4632 4344 4648
rect 4392 4632 4408 4648
rect 4536 4632 4552 4648
rect 4760 4632 4776 4648
rect 4904 4632 4920 4648
rect 5128 4632 5144 4648
rect 5448 4632 5464 4648
rect 5656 4632 5672 4648
rect 5960 4632 5976 4648
rect 6216 4632 6232 4648
rect 6872 4632 6888 4648
rect 7192 4632 7208 4648
rect 7400 4632 7416 4648
rect 2157 4602 2193 4618
rect 4205 4602 4241 4618
rect 6237 4602 6273 4618
rect 296 4572 312 4588
rect 584 4572 600 4588
rect 936 4572 952 4588
rect 984 4572 1000 4588
rect 1192 4572 1208 4588
rect 1400 4572 1416 4588
rect 1656 4572 1672 4588
rect 1688 4572 1704 4588
rect 1752 4572 1768 4588
rect 1816 4572 1832 4588
rect 2072 4572 2088 4588
rect 2120 4572 2136 4588
rect 2392 4572 2408 4588
rect 2504 4572 2520 4588
rect 2680 4572 2696 4588
rect 2872 4572 2888 4588
rect 3224 4572 3240 4588
rect 3720 4572 3736 4588
rect 4040 4572 4056 4588
rect 4456 4572 4472 4588
rect 4632 4572 4648 4588
rect 5032 4572 5048 4588
rect 5416 4572 5432 4588
rect 5576 4572 5592 4588
rect 5640 4572 5656 4588
rect 5960 4572 5976 4588
rect 168 4552 184 4568
rect 856 4552 872 4568
rect 1256 4552 1272 4568
rect 1320 4552 1336 4568
rect 1384 4552 1400 4568
rect 1496 4552 1512 4568
rect 1560 4552 1576 4568
rect 8 4532 24 4548
rect 72 4532 88 4548
rect 104 4532 120 4548
rect 424 4532 440 4548
rect 600 4532 616 4548
rect 632 4532 648 4548
rect 696 4532 712 4548
rect 904 4532 920 4548
rect 952 4532 968 4548
rect 1000 4532 1016 4548
rect 1032 4532 1048 4548
rect 1144 4532 1176 4548
rect 1240 4532 1256 4548
rect 1304 4532 1320 4548
rect 1368 4532 1384 4548
rect 1704 4532 1720 4548
rect 1784 4532 1800 4548
rect 2008 4532 2024 4548
rect 2088 4532 2104 4548
rect 24 4512 40 4528
rect 168 4514 184 4530
rect 232 4512 248 4528
rect 312 4512 344 4528
rect 392 4512 408 4528
rect 472 4512 488 4528
rect 520 4512 536 4528
rect 616 4512 632 4528
rect 72 4492 88 4508
rect 712 4512 744 4528
rect 776 4512 792 4528
rect 808 4512 824 4528
rect 872 4512 904 4528
rect 1048 4512 1064 4528
rect 664 4492 680 4508
rect 936 4492 952 4508
rect 984 4492 1000 4508
rect 1032 4492 1048 4508
rect 1080 4492 1096 4508
rect 1128 4512 1144 4528
rect 1224 4512 1240 4528
rect 1272 4512 1304 4528
rect 1320 4512 1336 4528
rect 1352 4512 1368 4528
rect 1416 4512 1432 4528
rect 1480 4512 1496 4528
rect 1528 4512 1544 4528
rect 1592 4512 1608 4528
rect 1720 4512 1736 4528
rect 1832 4512 1848 4528
rect 1960 4512 1976 4528
rect 2168 4512 2200 4528
rect 2232 4512 2248 4528
rect 2360 4532 2376 4548
rect 2440 4532 2456 4548
rect 2488 4532 2504 4548
rect 2584 4532 2600 4548
rect 2616 4532 2632 4548
rect 2680 4532 2696 4548
rect 2728 4552 2744 4568
rect 2808 4552 2824 4568
rect 3976 4552 3992 4568
rect 4792 4552 4808 4568
rect 5304 4552 5320 4568
rect 5560 4552 5576 4568
rect 5768 4552 5784 4568
rect 6184 4552 6200 4568
rect 6744 4552 6760 4568
rect 6952 4552 6968 4568
rect 2760 4532 2776 4548
rect 2824 4532 2840 4548
rect 2920 4532 2952 4548
rect 3000 4532 3016 4548
rect 3032 4532 3048 4548
rect 3064 4532 3080 4548
rect 3272 4532 3288 4548
rect 3416 4532 3432 4548
rect 3544 4532 3560 4548
rect 3640 4532 3656 4548
rect 3784 4532 3800 4548
rect 3992 4532 4008 4548
rect 4056 4532 4072 4548
rect 4120 4532 4136 4548
rect 4168 4532 4184 4548
rect 4248 4532 4296 4548
rect 4344 4532 4360 4548
rect 4440 4532 4456 4548
rect 4568 4532 4600 4548
rect 4680 4532 4696 4548
rect 4776 4532 4792 4548
rect 4824 4532 4840 4548
rect 4920 4532 4952 4548
rect 5016 4532 5032 4548
rect 5464 4532 5480 4548
rect 5496 4532 5512 4548
rect 5528 4532 5544 4548
rect 5576 4532 5592 4548
rect 5752 4532 5768 4548
rect 5800 4532 5816 4548
rect 5864 4532 5880 4548
rect 5960 4532 5976 4548
rect 6056 4532 6072 4548
rect 6232 4532 6248 4548
rect 6872 4532 6888 4548
rect 7128 4532 7144 4548
rect 7176 4532 7192 4548
rect 7400 4532 7416 4548
rect 1128 4492 1144 4508
rect 1192 4492 1208 4508
rect 1672 4492 1688 4508
rect 1816 4492 1832 4508
rect 2136 4492 2152 4508
rect 2296 4492 2312 4508
rect 2344 4512 2360 4528
rect 2424 4512 2440 4528
rect 2600 4512 2616 4528
rect 2664 4512 2680 4528
rect 2760 4512 2792 4528
rect 2840 4512 2856 4528
rect 2332 4492 2348 4508
rect 2472 4492 2488 4508
rect 2520 4492 2552 4508
rect 2568 4492 2584 4508
rect 2952 4512 2968 4528
rect 2888 4492 2904 4508
rect 3096 4514 3112 4530
rect 3288 4512 3304 4528
rect 3000 4492 3016 4508
rect 3300 4492 3316 4508
rect 3496 4512 3512 4528
rect 3576 4512 3592 4528
rect 3656 4512 3672 4528
rect 3720 4512 3736 4528
rect 3832 4512 3848 4528
rect 3880 4512 3896 4528
rect 4008 4512 4024 4528
rect 4056 4512 4072 4528
rect 4296 4512 4312 4528
rect 4360 4512 4392 4528
rect 4408 4512 4424 4528
rect 4488 4512 4504 4528
rect 3336 4492 3352 4508
rect 3688 4492 3720 4508
rect 4040 4492 4056 4508
rect 4072 4492 4088 4508
rect 4104 4492 4136 4508
rect 4328 4492 4344 4508
rect 4392 4492 4424 4508
rect 4616 4492 4632 4508
rect 4664 4512 4680 4528
rect 4760 4512 4776 4528
rect 4872 4512 4888 4528
rect 4904 4512 4920 4528
rect 5048 4512 5064 4528
rect 5160 4512 5176 4528
rect 5208 4512 5224 4528
rect 5320 4512 5336 4528
rect 5384 4512 5400 4528
rect 5480 4512 5496 4528
rect 5544 4512 5560 4528
rect 5592 4512 5608 4528
rect 5736 4512 5752 4528
rect 5816 4512 5832 4528
rect 5864 4512 5880 4528
rect 5976 4512 5992 4528
rect 6072 4512 6104 4528
rect 6152 4512 6168 4528
rect 6216 4512 6232 4528
rect 6296 4512 6312 4528
rect 6376 4512 6392 4528
rect 6440 4512 6456 4528
rect 6472 4512 6488 4528
rect 6504 4512 6536 4528
rect 6568 4512 6584 4528
rect 6632 4512 6648 4528
rect 6696 4512 6712 4528
rect 6744 4512 6760 4528
rect 6808 4512 6824 4528
rect 6856 4512 6872 4528
rect 6920 4512 6936 4528
rect 7080 4512 7096 4528
rect 7240 4514 7256 4530
rect 7304 4512 7320 4528
rect 4856 4492 4888 4508
rect 4984 4492 5000 4508
rect 5192 4492 5208 4508
rect 5336 4492 5352 4508
rect 5400 4492 5432 4508
rect 5480 4492 5496 4508
rect 5848 4492 5864 4508
rect 5912 4492 5928 4508
rect 6168 4492 6200 4508
rect 6280 4492 6296 4508
rect 6392 4492 6408 4508
rect 6456 4492 6472 4508
rect 6584 4492 6600 4508
rect 6648 4492 6664 4508
rect 6728 4492 6744 4508
rect 6792 4492 6808 4508
rect 6904 4492 6920 4508
rect 3736 4472 3752 4488
rect 3912 4472 3928 4488
rect 5128 4472 5160 4488
rect 5224 4472 5240 4488
rect 5304 4472 5320 4488
rect 5368 4472 5384 4488
rect 5816 4472 5832 4488
rect 6136 4472 6152 4488
rect 6312 4472 6344 4488
rect 6424 4472 6440 4488
rect 6488 4472 6520 4488
rect 6568 4472 6584 4488
rect 6616 4472 6648 4488
rect 6680 4472 6696 4488
rect 6712 4472 6728 4488
rect 6760 4472 6776 4488
rect 6792 4472 6808 4488
rect 2392 4452 2408 4468
rect 2456 4452 2472 4468
rect 4712 4452 4728 4468
rect 5208 4452 5224 4468
rect 5384 4452 5400 4468
rect 6632 4452 6648 4468
rect 360 4432 376 4448
rect 760 4432 776 4448
rect 1448 4432 1464 4448
rect 2216 4432 2232 4448
rect 3656 4432 3672 4448
rect 3976 4432 3992 4448
rect 4184 4432 4200 4448
rect 4296 4432 4312 4448
rect 4520 4432 4536 4448
rect 4840 4432 4856 4448
rect 6344 4432 6360 4448
rect 6808 4432 6824 4448
rect 7160 4432 7176 4448
rect 7368 4432 7400 4448
rect 1117 4402 1153 4418
rect 3165 4402 3201 4418
rect 5213 4402 5249 4418
rect 792 4372 808 4388
rect 2120 4372 2136 4388
rect 2360 4372 2376 4388
rect 3624 4372 3640 4388
rect 4056 4372 4072 4388
rect 4920 4372 4936 4388
rect 5000 4372 5016 4388
rect 5896 4372 5912 4388
rect 6040 4372 6056 4388
rect 6200 4372 6216 4388
rect 6760 4372 6776 4388
rect 7032 4372 7048 4388
rect 1256 4352 1272 4368
rect 584 4332 600 4348
rect 3032 4332 3048 4348
rect 3448 4332 3464 4348
rect 3640 4332 3656 4348
rect 3832 4332 3848 4348
rect 3880 4332 3896 4348
rect 4072 4332 4088 4348
rect 4424 4332 4440 4348
rect 4840 4332 4856 4348
rect 5016 4332 5032 4348
rect 5960 4352 5976 4368
rect 5528 4332 5544 4348
rect 5880 4332 5896 4348
rect 6024 4332 6040 4348
rect 6120 4332 6136 4348
rect 6728 4352 6744 4368
rect 6152 4332 6168 4348
rect 6216 4332 6232 4348
rect 6456 4332 6472 4348
rect 6712 4332 6728 4348
rect 6776 4332 6792 4348
rect 6840 4332 6856 4348
rect 6936 4332 6952 4348
rect 6968 4332 6984 4348
rect 7080 4352 7096 4368
rect 8 4292 24 4308
rect 72 4312 88 4328
rect 372 4312 388 4328
rect 392 4312 408 4328
rect 168 4290 184 4306
rect 232 4292 248 4308
rect 360 4292 376 4308
rect 472 4292 488 4308
rect 520 4292 536 4308
rect 616 4292 648 4308
rect 664 4312 680 4328
rect 728 4312 744 4328
rect 888 4312 904 4328
rect 936 4312 952 4328
rect 760 4292 776 4308
rect 824 4292 840 4308
rect 856 4292 872 4308
rect 984 4312 1000 4328
rect 1096 4312 1112 4328
rect 1528 4312 1544 4328
rect 1576 4312 1592 4328
rect 1672 4312 1688 4328
rect 1704 4312 1720 4328
rect 1912 4312 1928 4328
rect 2600 4312 2616 4328
rect 2632 4312 2648 4328
rect 3064 4312 3080 4328
rect 984 4292 1000 4308
rect 1032 4292 1064 4308
rect 1144 4292 1176 4308
rect 1224 4292 1240 4308
rect 1256 4292 1272 4308
rect 1288 4292 1304 4308
rect 1352 4292 1368 4308
rect 1416 4292 1432 4308
rect 1464 4292 1480 4308
rect 1544 4292 1560 4308
rect 1608 4292 1624 4308
rect 1848 4290 1864 4306
rect 1944 4292 1960 4308
rect 1976 4292 1992 4308
rect 2088 4292 2104 4308
rect 2184 4292 2200 4308
rect 2216 4292 2232 4308
rect 2248 4292 2264 4308
rect 2312 4292 2344 4308
rect 2456 4292 2472 4308
rect 2600 4292 2616 4308
rect 2712 4292 2728 4308
rect 2904 4292 2920 4308
rect 3256 4312 3272 4328
rect 3480 4312 3496 4328
rect 3112 4292 3128 4308
rect 3208 4292 3224 4308
rect 3336 4292 3352 4308
rect 3480 4292 3496 4308
rect 3528 4312 3544 4328
rect 3608 4312 3624 4328
rect 3672 4312 3688 4328
rect 3624 4292 3640 4308
rect 3704 4292 3720 4308
rect 3752 4292 3768 4308
rect 3800 4312 3816 4328
rect 4040 4312 4056 4328
rect 3960 4292 3976 4308
rect 4056 4292 4072 4308
rect 4120 4292 4136 4308
rect 4168 4312 4184 4328
rect 4456 4312 4472 4328
rect 4296 4290 4312 4306
rect 4440 4292 4456 4308
rect 4504 4312 4520 4328
rect 4872 4312 4888 4328
rect 4936 4312 4952 4328
rect 4984 4312 5000 4328
rect 5048 4312 5064 4328
rect 5080 4312 5096 4328
rect 5496 4312 5512 4328
rect 5848 4312 5864 4328
rect 5896 4312 5912 4328
rect 5992 4312 6008 4328
rect 6056 4312 6072 4328
rect 6120 4312 6136 4328
rect 6184 4312 6200 4328
rect 6264 4312 6280 4328
rect 6648 4312 6664 4328
rect 6744 4312 6760 4328
rect 6872 4312 6888 4328
rect 7000 4312 7016 4328
rect 7048 4332 7064 4348
rect 7096 4332 7128 4348
rect 7160 4332 7176 4348
rect 7128 4312 7144 4328
rect 7192 4312 7208 4328
rect 4680 4290 4696 4306
rect 4840 4292 4856 4308
rect 4888 4292 4904 4308
rect 5000 4292 5016 4308
rect 5080 4292 5096 4308
rect 5160 4290 5176 4306
rect 5416 4292 5432 4308
rect 5448 4292 5464 4308
rect 5512 4292 5528 4308
rect 5560 4292 5576 4308
rect 5736 4292 5752 4308
rect 5896 4292 5912 4308
rect 5928 4292 5944 4308
rect 6008 4292 6024 4308
rect 6104 4292 6120 4308
rect 6136 4292 6152 4308
rect 6200 4292 6216 4308
rect 6312 4292 6328 4308
rect 6344 4292 6360 4308
rect 6392 4292 6408 4308
rect 6440 4292 6456 4308
rect 6568 4292 6584 4308
rect 6728 4292 6744 4308
rect 6792 4292 6808 4308
rect 6856 4292 6872 4308
rect 6888 4292 6904 4308
rect 6920 4292 6952 4308
rect 6984 4292 7000 4308
rect 7032 4292 7048 4308
rect 7112 4292 7128 4308
rect 7176 4292 7192 4308
rect 7272 4292 7288 4308
rect 7320 4292 7336 4308
rect 8 4272 24 4288
rect 72 4272 88 4288
rect 104 4272 120 4288
rect 600 4272 616 4288
rect 696 4272 712 4288
rect 840 4272 856 4288
rect 904 4272 920 4288
rect 1016 4272 1032 4288
rect 1064 4272 1080 4288
rect 1240 4272 1256 4288
rect 1304 4272 1320 4288
rect 1400 4272 1416 4288
rect 1672 4272 1688 4288
rect 1880 4272 1896 4288
rect 1960 4272 1976 4288
rect 2184 4272 2200 4288
rect 2232 4272 2248 4288
rect 2264 4272 2280 4288
rect 328 4252 344 4268
rect 1016 4252 1032 4268
rect 1320 4252 1336 4268
rect 1352 4252 1384 4268
rect 1784 4252 1800 4268
rect 1912 4252 1928 4268
rect 2408 4272 2424 4288
rect 2488 4272 2504 4288
rect 2584 4272 2600 4288
rect 2664 4272 2680 4288
rect 2856 4272 2872 4288
rect 2952 4272 2968 4288
rect 3032 4272 3048 4288
rect 3064 4272 3080 4288
rect 3128 4272 3144 4288
rect 3288 4272 3304 4288
rect 3464 4272 3480 4288
rect 3560 4272 3576 4288
rect 3144 4252 3160 4268
rect 3592 4272 3608 4288
rect 3720 4272 3752 4288
rect 3784 4272 3800 4288
rect 3832 4272 3848 4288
rect 4008 4272 4024 4288
rect 4104 4272 4120 4288
rect 4168 4272 4184 4288
rect 4200 4272 4216 4288
rect 4264 4272 4280 4288
rect 4440 4272 4456 4288
rect 4536 4272 4552 4288
rect 4712 4272 4728 4288
rect 4744 4272 4760 4288
rect 4968 4272 4984 4288
rect 5096 4272 5112 4288
rect 5128 4272 5144 4288
rect 5384 4272 5400 4288
rect 5432 4272 5448 4288
rect 5784 4272 5800 4288
rect 5816 4272 5832 4288
rect 6104 4272 6120 4288
rect 6328 4272 6344 4288
rect 6360 4272 6376 4288
rect 4792 4252 4808 4268
rect 4936 4252 4952 4268
rect 6616 4272 6632 4288
rect 6648 4272 6664 4288
rect 6680 4272 6696 4288
rect 6408 4252 6424 4268
rect 296 4232 312 4248
rect 888 4232 904 4248
rect 1128 4232 1144 4248
rect 2008 4232 2024 4248
rect 2056 4232 2072 4248
rect 2120 4232 2136 4248
rect 2296 4232 2312 4248
rect 2568 4232 2584 4248
rect 2824 4232 2840 4248
rect 3256 4232 3272 4248
rect 3672 4232 3688 4248
rect 4552 4232 4568 4248
rect 4776 4232 4792 4248
rect 5352 4232 5368 4248
rect 5480 4232 5496 4248
rect 5592 4232 5608 4248
rect 5624 4232 5640 4248
rect 5848 4232 5864 4248
rect 6056 4232 6072 4248
rect 6280 4232 6296 4248
rect 7208 4232 7224 4248
rect 2157 4202 2193 4218
rect 4205 4202 4241 4218
rect 6237 4202 6273 4218
rect 184 4172 200 4188
rect 392 4172 424 4188
rect 808 4172 824 4188
rect 952 4172 968 4188
rect 1016 4172 1032 4188
rect 1208 4172 1224 4188
rect 2200 4172 2216 4188
rect 2632 4172 2648 4188
rect 2744 4172 2760 4188
rect 3320 4172 3336 4188
rect 3704 4172 3720 4188
rect 3816 4172 3832 4188
rect 4056 4172 4072 4188
rect 4680 4172 4696 4188
rect 5144 4172 5160 4188
rect 5416 4172 5432 4188
rect 5736 4172 5752 4188
rect 5800 4172 5816 4188
rect 5864 4172 5880 4188
rect 5944 4172 5960 4188
rect 5992 4172 6008 4188
rect 6072 4172 6088 4188
rect 6424 4172 6440 4188
rect 7080 4172 7096 4188
rect 7160 4172 7176 4188
rect 7224 4172 7240 4188
rect 7320 4172 7336 4188
rect 7400 4172 7416 4188
rect 72 4132 88 4148
rect 200 4132 216 4148
rect 232 4132 248 4148
rect 296 4132 312 4148
rect 840 4152 856 4168
rect 1512 4152 1528 4168
rect 2392 4152 2408 4168
rect 2584 4152 2600 4168
rect 2760 4152 2776 4168
rect 2952 4152 2968 4168
rect 3000 4152 3016 4168
rect 3480 4152 3496 4168
rect 3688 4152 3704 4168
rect 3800 4152 3816 4168
rect 3976 4152 3992 4168
rect 4040 4152 4056 4168
rect 4808 4152 4824 4168
rect 5512 4152 5528 4168
rect 5672 4152 5688 4168
rect 6072 4152 6088 4168
rect 6424 4152 6440 4168
rect 6712 4152 6728 4168
rect 7256 4152 7272 4168
rect 440 4132 456 4148
rect 904 4132 920 4148
rect 1032 4132 1064 4148
rect 1192 4132 1208 4148
rect 1624 4132 1640 4148
rect 1688 4132 1704 4148
rect 88 4112 104 4128
rect 216 4112 232 4128
rect 344 4112 360 4128
rect 568 4112 584 4128
rect 712 4112 728 4128
rect 760 4112 792 4128
rect 888 4112 904 4128
rect 984 4112 1000 4128
rect 1048 4112 1064 4128
rect 1144 4112 1192 4128
rect 1272 4112 1304 4128
rect 1464 4112 1480 4128
rect 264 4092 280 4108
rect 392 4092 424 4108
rect 920 4092 936 4108
rect 968 4092 984 4108
rect 1096 4092 1112 4108
rect 1128 4092 1144 4108
rect 1624 4092 1640 4108
rect 1672 4112 1688 4128
rect 1768 4132 1784 4148
rect 1896 4132 1912 4148
rect 1992 4132 2008 4148
rect 2056 4132 2072 4148
rect 2152 4132 2168 4148
rect 2456 4132 2472 4148
rect 2632 4132 2648 4148
rect 2712 4132 2728 4148
rect 2776 4132 2792 4148
rect 2808 4132 2824 4148
rect 2872 4132 2888 4148
rect 3128 4132 3144 4148
rect 3160 4132 3176 4148
rect 3336 4132 3352 4148
rect 3400 4132 3416 4148
rect 3432 4132 3448 4148
rect 3560 4132 3576 4148
rect 3608 4132 3624 4148
rect 3848 4132 3864 4148
rect 3880 4132 3896 4148
rect 4024 4132 4040 4148
rect 4136 4132 4152 4148
rect 4280 4132 4296 4148
rect 4344 4132 4360 4148
rect 4536 4132 4552 4148
rect 4600 4132 4632 4148
rect 4872 4132 4888 4148
rect 4904 4132 4920 4148
rect 4968 4132 4984 4148
rect 5016 4132 5048 4148
rect 5192 4132 5208 4148
rect 5272 4132 5304 4148
rect 5480 4132 5496 4148
rect 5528 4132 5544 4148
rect 5576 4132 5592 4148
rect 5752 4132 5768 4148
rect 6056 4132 6072 4148
rect 1752 4112 1768 4128
rect 1816 4112 1848 4128
rect 1912 4112 1928 4128
rect 1960 4112 1992 4128
rect 2040 4112 2056 4128
rect 2088 4092 2104 4108
rect 2136 4112 2152 4128
rect 2264 4112 2280 4128
rect 2312 4112 2328 4128
rect 2424 4112 2440 4128
rect 2488 4112 2504 4128
rect 2664 4112 2680 4128
rect 2696 4112 2712 4128
rect 2728 4112 2744 4128
rect 2792 4112 2808 4128
rect 2632 4092 2648 4108
rect 2696 4092 2712 4108
rect 2888 4112 2904 4128
rect 3032 4112 3064 4128
rect 3208 4112 3224 4128
rect 3352 4112 3368 4128
rect 3448 4112 3464 4128
rect 3512 4112 3528 4128
rect 3592 4112 3608 4128
rect 3640 4112 3656 4128
rect 3720 4112 3736 4128
rect 3768 4112 3784 4128
rect 3832 4112 3848 4128
rect 3864 4112 3880 4128
rect 3928 4112 3944 4128
rect 4024 4112 4040 4128
rect 4120 4112 4136 4128
rect 4200 4112 4216 4128
rect 4280 4112 4296 4128
rect 4328 4112 4344 4128
rect 4392 4112 4408 4128
rect 4456 4112 4472 4128
rect 4552 4112 4568 4128
rect 4584 4112 4600 4128
rect 4664 4112 4680 4128
rect 4808 4114 4824 4130
rect 2840 4092 2856 4108
rect 2920 4092 2936 4108
rect 3352 4092 3368 4108
rect 3432 4092 3448 4108
rect 3544 4092 3560 4108
rect 3624 4092 3640 4108
rect 3784 4092 3800 4108
rect 3928 4092 3944 4108
rect 3976 4092 3992 4108
rect 4088 4092 4104 4108
rect 4248 4092 4264 4108
rect 4408 4092 4424 4108
rect 4472 4092 4488 4108
rect 4552 4092 4568 4108
rect 4904 4092 4920 4108
rect 4952 4112 4968 4128
rect 4984 4112 5000 4128
rect 5176 4112 5192 4128
rect 5208 4112 5224 4128
rect 5304 4112 5320 4128
rect 5384 4112 5400 4128
rect 5480 4112 5512 4128
rect 5624 4112 5640 4128
rect 5704 4112 5720 4128
rect 5768 4112 5784 4128
rect 5848 4112 5864 4128
rect 5896 4112 5928 4128
rect 6056 4112 6088 4128
rect 6216 4112 6232 4128
rect 6264 4132 6280 4148
rect 6296 4132 6312 4148
rect 6408 4132 6424 4148
rect 6520 4132 6536 4148
rect 6552 4132 6568 4148
rect 6680 4132 6696 4148
rect 6904 4132 6920 4148
rect 7336 4132 7352 4148
rect 6280 4112 6296 4128
rect 6344 4112 6360 4128
rect 6440 4112 6456 4128
rect 6536 4112 6552 4128
rect 6600 4112 6616 4128
rect 6648 4112 6664 4128
rect 6840 4112 6856 4128
rect 6968 4112 6984 4128
rect 7016 4112 7032 4128
rect 7112 4112 7144 4128
rect 7192 4112 7208 4128
rect 7288 4112 7304 4128
rect 7352 4112 7384 4128
rect 5240 4092 5256 4108
rect 5400 4092 5416 4108
rect 5624 4092 5640 4108
rect 6168 4092 6184 4108
rect 6328 4092 6344 4108
rect 6584 4092 6600 4108
rect 7016 4092 7032 4108
rect 2136 4072 2152 4088
rect 2584 4072 2600 4088
rect 3288 4072 3304 4088
rect 3512 4072 3528 4088
rect 3656 4072 3672 4088
rect 3752 4072 3768 4088
rect 3944 4072 3960 4088
rect 4376 4072 4392 4088
rect 4440 4072 4456 4088
rect 4392 4052 4408 4068
rect 5368 4072 5384 4088
rect 5640 4072 5656 4088
rect 6200 4072 6216 4088
rect 6360 4072 6376 4088
rect 6616 4072 6632 4088
rect 6952 4072 6968 4088
rect 7032 4072 7048 4088
rect 456 4032 472 4048
rect 664 4032 680 4048
rect 728 4032 744 4048
rect 808 4032 824 4048
rect 1016 4032 1032 4048
rect 1944 4032 1960 4048
rect 2536 4032 2552 4048
rect 2968 4032 2984 4048
rect 3000 4032 3016 4048
rect 3080 4032 3096 4048
rect 3320 4032 3336 4048
rect 3640 4032 3656 4048
rect 3768 4032 3784 4048
rect 4168 4032 4184 4048
rect 4520 4032 4536 4048
rect 4584 4032 4600 4048
rect 5064 4032 5080 4048
rect 5208 4032 5224 4048
rect 5304 4032 5320 4048
rect 5800 4032 5816 4048
rect 6936 4032 6952 4048
rect 7016 4032 7032 4048
rect 7224 4032 7240 4048
rect 1117 4002 1153 4018
rect 3165 4002 3201 4018
rect 5213 4002 5249 4018
rect 488 3972 504 3988
rect 2424 3972 2440 3988
rect 3608 3972 3624 3988
rect 3720 3972 3736 3988
rect 3848 3972 3864 3988
rect 3912 3972 3928 3988
rect 3960 3972 3976 3988
rect 4520 3972 4536 3988
rect 4632 3972 4648 3988
rect 4904 3972 4920 3988
rect 5128 3972 5144 3988
rect 5400 3972 5416 3988
rect 6520 3972 6536 3988
rect 6776 3972 6792 3988
rect 7016 3972 7032 3988
rect 2296 3952 2312 3968
rect 264 3932 280 3948
rect 1288 3932 1304 3948
rect 1320 3932 1336 3948
rect 1544 3932 1560 3948
rect 2216 3932 2232 3948
rect 2760 3932 2776 3948
rect 3832 3932 3848 3948
rect 3896 3932 3912 3948
rect 4280 3932 4296 3948
rect 4424 3932 4440 3948
rect 4536 3932 4552 3948
rect 4648 3932 4664 3948
rect 4888 3932 4904 3948
rect 4920 3932 4936 3948
rect 6744 3952 6760 3968
rect 5368 3932 5384 3948
rect 5416 3932 5432 3948
rect 6072 3932 6088 3948
rect 6728 3932 6744 3948
rect 6792 3932 6808 3948
rect 6856 3932 6872 3948
rect 6920 3932 6936 3948
rect 7048 3952 7064 3968
rect 200 3912 216 3928
rect 88 3892 104 3908
rect 232 3892 248 3908
rect 392 3912 408 3928
rect 440 3912 456 3928
rect 280 3892 296 3908
rect 344 3892 392 3908
rect 488 3892 504 3908
rect 536 3892 552 3908
rect 584 3912 600 3928
rect 680 3912 696 3928
rect 920 3912 936 3928
rect 616 3892 632 3908
rect 744 3890 760 3906
rect 968 3892 984 3908
rect 1016 3892 1032 3908
rect 1064 3912 1080 3928
rect 1464 3912 1480 3928
rect 1192 3890 1208 3906
rect 1400 3892 1432 3908
rect 1864 3912 1880 3928
rect 1960 3912 1976 3928
rect 2376 3912 2392 3928
rect 1512 3892 1528 3908
rect 1640 3892 1656 3908
rect 1736 3892 1752 3908
rect 1848 3892 1864 3908
rect 1912 3892 1928 3908
rect 2024 3890 2040 3906
rect 2232 3892 2280 3908
rect 2312 3892 2328 3908
rect 2488 3912 2504 3928
rect 2424 3892 2456 3908
rect 2824 3912 2840 3928
rect 3112 3912 3128 3928
rect 2520 3892 2552 3908
rect 2568 3892 2584 3908
rect 2616 3892 2632 3908
rect 2712 3892 2728 3908
rect 2888 3892 2904 3908
rect 2968 3892 2984 3908
rect 3112 3892 3128 3908
rect 3160 3912 3176 3928
rect 3272 3912 3288 3928
rect 3560 3912 3576 3928
rect 3640 3912 3656 3928
rect 3752 3912 3768 3928
rect 3864 3912 3880 3928
rect 3928 3912 3944 3928
rect 3368 3892 3384 3908
rect 3560 3892 3576 3908
rect 3672 3892 3688 3908
rect 3784 3892 3800 3908
rect 3848 3892 3864 3908
rect 3912 3892 3928 3908
rect 3976 3892 3992 3908
rect 4008 3892 4024 3908
rect 4056 3912 4072 3928
rect 4344 3912 4360 3928
rect 4168 3892 4184 3908
rect 4216 3892 4232 3908
rect 4296 3892 4312 3908
rect 4328 3892 4360 3908
rect 4392 3912 4408 3928
rect 4504 3912 4520 3928
rect 4616 3912 4632 3928
rect 4680 3912 4696 3928
rect 4712 3912 4728 3928
rect 4776 3912 4808 3928
rect 4824 3912 4840 3928
rect 4856 3912 4872 3928
rect 5336 3912 5352 3928
rect 5448 3912 5464 3928
rect 5624 3912 5640 3928
rect 6632 3912 6648 3928
rect 6664 3912 6680 3928
rect 6760 3912 6776 3928
rect 6888 3912 6904 3928
rect 6952 3912 6968 3928
rect 7000 3932 7016 3948
rect 7064 3932 7080 3948
rect 7032 3912 7048 3928
rect 4392 3892 4408 3908
rect 4424 3892 4440 3908
rect 4488 3892 4504 3908
rect 4520 3892 4536 3908
rect 4600 3892 4616 3908
rect 4632 3892 4648 3908
rect 72 3872 88 3888
rect 200 3872 216 3888
rect 248 3872 264 3888
rect 296 3872 312 3888
rect 408 3872 424 3888
rect 504 3872 536 3888
rect 584 3872 600 3888
rect 616 3872 648 3888
rect 760 3872 776 3888
rect 888 3872 904 3888
rect 952 3872 968 3888
rect 984 3872 1016 3888
rect 1064 3872 1080 3888
rect 1128 3872 1144 3888
rect 1224 3872 1240 3888
rect 1432 3872 1448 3888
rect 1496 3872 1512 3888
rect 1528 3872 1544 3888
rect 1704 3872 1720 3888
rect 1800 3872 1816 3888
rect 1896 3872 1928 3888
rect 1960 3872 1976 3888
rect 2344 3872 2360 3888
rect 2456 3872 2472 3888
rect 2552 3872 2568 3888
rect 1384 3852 1400 3868
rect 2024 3852 2040 3868
rect 2200 3852 2216 3868
rect 2584 3852 2616 3868
rect 2648 3852 2664 3868
rect 2696 3872 2712 3888
rect 2776 3872 2792 3888
rect 3096 3872 3112 3888
rect 3192 3872 3208 3888
rect 3240 3872 3256 3888
rect 3304 3872 3320 3888
rect 3512 3872 3528 3888
rect 3576 3872 3592 3888
rect 3688 3872 3704 3888
rect 3800 3872 3816 3888
rect 3992 3872 4008 3888
rect 4056 3872 4072 3888
rect 4088 3872 4104 3888
rect 4328 3872 4344 3888
rect 4440 3872 4456 3888
rect 4488 3872 4504 3888
rect 4600 3872 4616 3888
rect 4744 3892 4760 3908
rect 4824 3892 4840 3908
rect 4872 3892 4888 3908
rect 5032 3892 5048 3908
rect 5176 3892 5192 3908
rect 5288 3892 5304 3908
rect 5352 3892 5368 3908
rect 5432 3892 5448 3908
rect 5512 3892 5528 3908
rect 5720 3890 5736 3906
rect 5784 3892 5800 3908
rect 5848 3892 5864 3908
rect 5960 3892 5976 3908
rect 6088 3892 6104 3908
rect 6120 3892 6136 3908
rect 4728 3872 4744 3888
rect 4840 3872 4856 3888
rect 5192 3872 5208 3888
rect 5272 3872 5288 3888
rect 5320 3872 5336 3888
rect 5496 3872 5512 3888
rect 5688 3872 5704 3888
rect 5800 3872 5816 3888
rect 5912 3872 5928 3888
rect 5960 3872 5976 3888
rect 6104 3872 6120 3888
rect 6200 3892 6216 3908
rect 6280 3892 6312 3908
rect 6392 3890 6408 3906
rect 6456 3892 6472 3908
rect 6536 3892 6552 3908
rect 6696 3892 6712 3908
rect 6744 3892 6760 3908
rect 6808 3892 6824 3908
rect 6872 3892 6888 3908
rect 6936 3892 6952 3908
rect 6984 3892 7000 3908
rect 7048 3892 7064 3908
rect 7128 3892 7144 3908
rect 7192 3892 7208 3908
rect 7336 3890 7352 3906
rect 2952 3852 2968 3868
rect 3432 3852 3448 3868
rect 3592 3852 3608 3868
rect 3704 3852 3720 3868
rect 3944 3852 3960 3868
rect 4456 3852 4472 3868
rect 4568 3852 4584 3868
rect 5048 3852 5064 3868
rect 5208 3852 5224 3868
rect 5496 3852 5528 3868
rect 5880 3852 5896 3868
rect 6216 3872 6232 3888
rect 6584 3872 6616 3888
rect 7144 3872 7160 3888
rect 7176 3872 7192 3888
rect 7320 3872 7336 3888
rect 6152 3852 6168 3868
rect 6328 3852 6344 3868
rect 7096 3852 7112 3868
rect 184 3832 200 3848
rect 680 3832 696 3848
rect 872 3832 888 3848
rect 1816 3832 1832 3848
rect 1880 3832 1896 3848
rect 2152 3832 2168 3848
rect 2824 3832 2840 3848
rect 2856 3832 2872 3848
rect 3080 3832 3096 3848
rect 3272 3832 3288 3848
rect 4776 3832 4792 3848
rect 5592 3832 5608 3848
rect 5816 3832 5832 3848
rect 6616 3832 6632 3848
rect 7208 3832 7224 3848
rect 2157 3802 2193 3818
rect 4205 3802 4241 3818
rect 6237 3802 6273 3818
rect 344 3772 360 3788
rect 392 3772 408 3788
rect 424 3772 440 3788
rect 792 3772 808 3788
rect 888 3772 904 3788
rect 920 3772 936 3788
rect 1096 3772 1112 3788
rect 1448 3772 1464 3788
rect 2088 3772 2120 3788
rect 2776 3772 2792 3788
rect 3032 3772 3048 3788
rect 3368 3772 3384 3788
rect 3464 3772 3480 3788
rect 3592 3772 3608 3788
rect 3704 3772 3720 3788
rect 3848 3772 3864 3788
rect 3960 3772 3976 3788
rect 3992 3772 4008 3788
rect 4056 3772 4072 3788
rect 4104 3772 4120 3788
rect 4408 3772 4424 3788
rect 4456 3772 4472 3788
rect 4488 3772 4504 3788
rect 4552 3772 4568 3788
rect 4680 3772 4696 3788
rect 4968 3772 4984 3788
rect 5048 3772 5064 3788
rect 5256 3772 5272 3788
rect 5704 3772 5720 3788
rect 5832 3772 5848 3788
rect 6088 3772 6104 3788
rect 6120 3772 6136 3788
rect 6680 3772 6696 3788
rect 6760 3772 6776 3788
rect 6808 3772 6824 3788
rect 6968 3772 6984 3788
rect 7160 3772 7176 3788
rect 7384 3772 7400 3788
rect 664 3752 680 3768
rect 1192 3752 1208 3768
rect 1496 3752 1512 3768
rect 1624 3752 1640 3768
rect 1672 3752 1688 3768
rect 72 3732 88 3748
rect 104 3732 120 3748
rect 168 3732 184 3748
rect 248 3732 264 3748
rect 312 3732 328 3748
rect 360 3732 376 3748
rect 408 3732 424 3748
rect 856 3732 872 3748
rect 904 3732 920 3748
rect 952 3732 968 3748
rect 1048 3732 1080 3748
rect 1144 3732 1160 3748
rect 1240 3732 1256 3748
rect 1352 3732 1384 3748
rect 1528 3732 1544 3748
rect 1608 3732 1624 3748
rect 1640 3732 1656 3748
rect 1752 3732 1768 3748
rect 1816 3732 1832 3748
rect 1896 3732 1912 3748
rect 1976 3732 1992 3748
rect 2024 3732 2040 3748
rect 2136 3732 2152 3748
rect 2200 3732 2216 3748
rect 2376 3732 2392 3748
rect 2488 3732 2504 3748
rect 2520 3732 2536 3748
rect 2552 3732 2568 3748
rect 2584 3732 2600 3748
rect 2648 3732 2664 3748
rect 2792 3732 2808 3748
rect 2872 3732 2888 3748
rect 2952 3732 2968 3748
rect 3048 3732 3064 3748
rect 3096 3732 3112 3748
rect 3144 3732 3160 3748
rect 3288 3752 3304 3768
rect 3528 3752 3544 3768
rect 3640 3752 3656 3768
rect 3752 3752 3768 3768
rect 4536 3752 4552 3768
rect 4760 3752 4776 3768
rect 4792 3752 4808 3768
rect 3288 3732 3304 3748
rect 3320 3732 3336 3748
rect 3416 3732 3432 3748
rect 3560 3732 3576 3748
rect 3672 3732 3688 3748
rect 3784 3732 3800 3748
rect 3896 3732 3912 3748
rect 3944 3732 3960 3748
rect 4024 3732 4056 3748
rect 4152 3732 4168 3748
rect 4328 3732 4344 3748
rect 4376 3732 4392 3748
rect 4424 3732 4440 3748
rect 4584 3732 4600 3748
rect 4696 3732 4712 3748
rect 4872 3732 4888 3748
rect 5320 3732 5336 3748
rect 5368 3752 5384 3768
rect 5480 3752 5496 3768
rect 5528 3732 5560 3748
rect 5576 3732 5592 3748
rect 5608 3732 5624 3748
rect 5704 3732 5720 3748
rect 5816 3732 5832 3748
rect 5864 3752 5880 3768
rect 5960 3752 5976 3768
rect 6888 3752 6904 3768
rect 6232 3732 6248 3748
rect 6296 3732 6312 3748
rect 7400 3752 7416 3768
rect 6936 3732 6952 3748
rect 7128 3732 7144 3748
rect 7320 3732 7336 3748
rect 7368 3732 7384 3748
rect 136 3714 152 3730
rect 200 3712 216 3728
rect 232 3712 248 3728
rect 280 3712 312 3728
rect 536 3712 552 3728
rect 680 3712 696 3728
rect 808 3712 824 3728
rect 840 3712 856 3728
rect 200 3692 216 3708
rect 264 3692 280 3708
rect 328 3692 344 3708
rect 376 3692 392 3708
rect 808 3692 824 3708
rect 952 3712 968 3728
rect 984 3712 1000 3728
rect 1032 3712 1048 3728
rect 1112 3712 1128 3728
rect 920 3692 936 3708
rect 1096 3692 1112 3708
rect 1208 3692 1224 3708
rect 1288 3692 1304 3708
rect 1336 3712 1352 3728
rect 1432 3712 1448 3728
rect 1480 3712 1496 3728
rect 1528 3712 1560 3728
rect 1592 3712 1608 3728
rect 1656 3712 1672 3728
rect 1704 3712 1720 3728
rect 1752 3712 1768 3728
rect 1832 3712 1848 3728
rect 1960 3714 1976 3730
rect 2248 3712 2264 3728
rect 2392 3712 2424 3728
rect 1560 3692 1576 3708
rect 1896 3692 1912 3708
rect 2104 3692 2120 3708
rect 2568 3712 2584 3728
rect 2664 3712 2680 3728
rect 2808 3712 2824 3728
rect 2920 3712 2936 3728
rect 3080 3712 3096 3728
rect 3112 3712 3128 3728
rect 3240 3712 3256 3728
rect 3336 3712 3352 3728
rect 2440 3692 2456 3708
rect 2488 3692 2504 3708
rect 2808 3692 2824 3708
rect 2840 3692 2856 3708
rect 3048 3692 3064 3708
rect 3128 3692 3144 3708
rect 3272 3692 3288 3708
rect 3432 3712 3448 3728
rect 3528 3712 3544 3728
rect 3640 3712 3656 3728
rect 3752 3712 3768 3728
rect 3864 3712 3880 3728
rect 3912 3712 3928 3728
rect 4136 3712 4152 3728
rect 4168 3712 4184 3728
rect 4280 3712 4296 3728
rect 4344 3712 4360 3728
rect 4520 3712 4536 3728
rect 4584 3712 4616 3728
rect 4648 3712 4664 3728
rect 4712 3712 4728 3728
rect 4952 3712 4968 3728
rect 5000 3712 5032 3728
rect 5144 3712 5160 3728
rect 5304 3712 5320 3728
rect 5352 3712 5368 3728
rect 5400 3712 5416 3728
rect 5432 3712 5448 3728
rect 5512 3712 5528 3728
rect 5560 3712 5576 3728
rect 5592 3712 5608 3728
rect 5720 3712 5736 3728
rect 5768 3712 5784 3728
rect 5896 3712 5912 3728
rect 5976 3712 5992 3728
rect 6152 3712 6184 3728
rect 6360 3712 6376 3728
rect 6408 3712 6440 3728
rect 6536 3712 6552 3728
rect 6584 3712 6600 3728
rect 6712 3712 6744 3728
rect 6840 3712 6872 3728
rect 6920 3712 6936 3728
rect 6952 3712 6968 3728
rect 7048 3712 7064 3728
rect 7224 3712 7240 3728
rect 7272 3712 7288 3728
rect 7352 3712 7368 3728
rect 3384 3692 3400 3708
rect 3544 3692 3560 3708
rect 3592 3692 3608 3708
rect 3656 3692 3672 3708
rect 3704 3692 3720 3708
rect 3768 3692 3784 3708
rect 3816 3692 3832 3708
rect 3928 3692 3944 3708
rect 3976 3692 4008 3708
rect 4072 3692 4088 3708
rect 4168 3692 4184 3708
rect 4200 3692 4216 3708
rect 4296 3692 4312 3708
rect 4360 3692 4376 3708
rect 4424 3692 4440 3708
rect 4456 3692 4472 3708
rect 4600 3692 4616 3708
rect 4632 3692 4648 3708
rect 4744 3692 4760 3708
rect 5416 3692 5432 3708
rect 5592 3692 5608 3708
rect 5656 3692 5672 3708
rect 6264 3692 6280 3708
rect 6376 3692 6392 3708
rect 456 3672 472 3688
rect 2360 3672 2376 3688
rect 2744 3672 2760 3688
rect 3512 3672 3528 3688
rect 3672 3672 3688 3688
rect 3736 3672 3752 3688
rect 3896 3672 3912 3688
rect 4264 3672 4280 3688
rect 4328 3672 4344 3688
rect 5224 3672 5240 3688
rect 5448 3672 5464 3688
rect 6056 3672 6072 3688
rect 6248 3672 6264 3688
rect 6408 3672 6424 3688
rect 1336 3652 1352 3668
rect 4280 3652 4296 3668
rect 8 3632 24 3648
rect 424 3632 440 3648
rect 1384 3632 1400 3648
rect 1448 3632 1464 3648
rect 1528 3632 1544 3648
rect 1816 3632 1832 3648
rect 2776 3632 2792 3648
rect 3304 3632 3320 3648
rect 3464 3632 3480 3648
rect 4824 3632 4840 3648
rect 4904 3632 4920 3648
rect 6200 3632 6216 3648
rect 6760 3632 6776 3648
rect 1117 3602 1153 3618
rect 3165 3602 3201 3618
rect 5213 3602 5249 3618
rect 24 3572 40 3588
rect 552 3572 568 3588
rect 808 3572 824 3588
rect 888 3572 904 3588
rect 968 3572 984 3588
rect 1080 3572 1096 3588
rect 1512 3572 1528 3588
rect 3336 3572 3352 3588
rect 3544 3572 3560 3588
rect 3768 3572 3784 3588
rect 3832 3572 3848 3588
rect 3896 3572 3912 3588
rect 3960 3572 3976 3588
rect 4040 3572 4056 3588
rect 4088 3572 4104 3588
rect 4152 3572 4168 3588
rect 4248 3572 4264 3588
rect 4296 3572 4312 3588
rect 4408 3572 4424 3588
rect 4440 3572 4456 3588
rect 4504 3572 4520 3588
rect 4632 3572 4648 3588
rect 4696 3572 4712 3588
rect 4936 3572 4952 3588
rect 5000 3572 5016 3588
rect 5128 3572 5144 3588
rect 5208 3572 5224 3588
rect 5384 3572 5400 3588
rect 5704 3572 5720 3588
rect 5816 3572 5832 3588
rect 5896 3572 5912 3588
rect 6440 3572 6456 3588
rect 6936 3572 6952 3588
rect 6984 3572 7000 3588
rect 7384 3572 7400 3588
rect 56 3532 72 3548
rect 120 3532 136 3548
rect 184 3532 200 3548
rect 600 3532 616 3548
rect 1160 3532 1176 3548
rect 1672 3532 1688 3548
rect 2040 3532 2056 3548
rect 2872 3532 2888 3548
rect 2936 3532 2952 3548
rect 3272 3532 3288 3548
rect 3352 3532 3368 3548
rect 3784 3532 3800 3548
rect 3848 3532 3864 3548
rect 3896 3532 3912 3548
rect 3976 3532 3992 3548
rect 4024 3532 4040 3548
rect 4104 3532 4120 3548
rect 4168 3532 4184 3548
rect 4264 3532 4280 3548
rect 4312 3532 4344 3548
rect 4392 3532 4408 3548
rect 4456 3532 4472 3548
rect 4520 3532 4536 3548
rect 4648 3532 4664 3548
rect 4712 3532 4728 3548
rect 5768 3552 5784 3568
rect 6232 3552 6248 3568
rect 4888 3532 4904 3548
rect 4952 3532 4968 3548
rect 5016 3532 5032 3548
rect 5656 3532 5672 3548
rect 5784 3532 5800 3548
rect 5832 3532 5848 3548
rect 5912 3532 5928 3548
rect 6152 3532 6168 3548
rect 6312 3532 6328 3548
rect 6584 3532 6600 3548
rect 6872 3532 6888 3548
rect 7048 3552 7064 3568
rect 164 3512 180 3528
rect 200 3512 216 3528
rect 264 3512 280 3528
rect 296 3512 312 3528
rect 584 3512 600 3528
rect 936 3512 952 3528
rect 1384 3512 1400 3528
rect 24 3492 40 3508
rect 88 3492 104 3508
rect 136 3492 168 3508
rect 232 3492 248 3508
rect 376 3492 392 3508
rect 424 3492 440 3508
rect 552 3492 568 3508
rect 712 3492 728 3508
rect 824 3492 840 3508
rect 856 3492 872 3508
rect 904 3492 920 3508
rect 936 3492 952 3508
rect 968 3492 984 3508
rect 1048 3492 1064 3508
rect 1096 3492 1112 3508
rect 1128 3492 1144 3508
rect 1224 3492 1240 3508
rect 1288 3490 1304 3506
rect 1592 3512 1608 3528
rect 1448 3492 1496 3508
rect 1544 3492 1560 3508
rect 1640 3512 1656 3528
rect 2072 3512 2088 3528
rect 1640 3492 1656 3508
rect 1784 3492 1800 3508
rect 1928 3492 1944 3508
rect 1976 3492 1992 3508
rect 2072 3492 2088 3508
rect 2120 3512 2136 3528
rect 2296 3512 2312 3528
rect 2392 3512 2408 3528
rect 2600 3512 2616 3528
rect 2712 3512 2728 3528
rect 3016 3512 3032 3528
rect 3304 3512 3336 3528
rect 3400 3512 3416 3528
rect 2248 3492 2264 3508
rect 2312 3492 2344 3508
rect 2376 3492 2392 3508
rect 2472 3492 2488 3508
rect 2616 3492 2648 3508
rect 2680 3492 2712 3508
rect 2792 3492 2808 3508
rect 8 3472 24 3488
rect 72 3472 88 3488
rect 136 3472 152 3488
rect 248 3472 264 3488
rect 296 3472 312 3488
rect 760 3472 776 3488
rect 792 3472 808 3488
rect 1320 3472 1336 3488
rect 1352 3472 1368 3488
rect 1384 3472 1400 3488
rect 1448 3472 1464 3488
rect 1560 3472 1576 3488
rect 1656 3472 1672 3488
rect 2056 3472 2072 3488
rect 2152 3472 2168 3488
rect 2296 3472 2312 3488
rect 2328 3472 2360 3488
rect 2424 3472 2440 3488
rect 2664 3472 2680 3488
rect 2744 3472 2760 3488
rect 2984 3492 3000 3508
rect 3016 3492 3032 3508
rect 3096 3492 3112 3508
rect 3160 3490 3176 3506
rect 3272 3492 3288 3508
rect 3432 3492 3448 3508
rect 3480 3512 3496 3528
rect 3752 3512 3768 3528
rect 3816 3512 3832 3528
rect 3880 3512 3896 3528
rect 3944 3512 3960 3528
rect 4056 3512 4088 3528
rect 4136 3512 4152 3528
rect 4232 3512 4248 3528
rect 4344 3512 4376 3528
rect 4424 3512 4440 3528
rect 4488 3512 4504 3528
rect 4584 3512 4600 3528
rect 4616 3512 4632 3528
rect 4680 3512 4696 3528
rect 4808 3512 4824 3528
rect 4856 3512 4872 3528
rect 4920 3512 4936 3528
rect 4984 3512 5000 3528
rect 5064 3512 5080 3528
rect 5688 3512 5704 3528
rect 5752 3512 5768 3528
rect 5880 3512 5896 3528
rect 6344 3512 6360 3528
rect 6552 3512 6568 3528
rect 6776 3512 6792 3528
rect 6824 3512 6840 3528
rect 6904 3512 6920 3528
rect 6952 3532 6968 3548
rect 7000 3532 7016 3548
rect 7064 3532 7080 3548
rect 7096 3532 7112 3548
rect 7032 3512 7048 3528
rect 3640 3492 3656 3508
rect 3768 3492 3784 3508
rect 3832 3492 3848 3508
rect 3912 3492 3928 3508
rect 3960 3492 3976 3508
rect 4040 3492 4056 3508
rect 4088 3492 4104 3508
rect 4152 3492 4168 3508
rect 4248 3492 4264 3508
rect 4328 3492 4344 3508
rect 4376 3492 4392 3508
rect 4440 3492 4456 3508
rect 4504 3492 4520 3508
rect 4552 3492 4568 3508
rect 4632 3492 4648 3508
rect 4712 3492 4728 3508
rect 4744 3492 4760 3508
rect 4792 3492 4824 3508
rect 4872 3492 4888 3508
rect 4936 3492 4952 3508
rect 5000 3492 5016 3508
rect 5096 3492 5112 3508
rect 5160 3492 5192 3508
rect 5480 3490 5496 3506
rect 5640 3492 5656 3508
rect 5704 3492 5720 3508
rect 5768 3492 5784 3508
rect 5848 3492 5864 3508
rect 5896 3492 5912 3508
rect 6040 3492 6056 3508
rect 6184 3492 6216 3508
rect 6328 3492 6344 3508
rect 6392 3492 6408 3508
rect 6472 3492 6488 3508
rect 6504 3492 6520 3508
rect 6568 3492 6584 3508
rect 6664 3492 6680 3508
rect 6792 3492 6808 3508
rect 6888 3492 6904 3508
rect 6936 3492 6952 3508
rect 7016 3492 7032 3508
rect 7080 3492 7128 3508
rect 7208 3490 7224 3506
rect 7352 3492 7368 3508
rect 2968 3472 2984 3488
rect 3224 3472 3240 3488
rect 3256 3472 3272 3488
rect 3368 3472 3384 3488
rect 3416 3472 3432 3488
rect 3480 3472 3496 3488
rect 3528 3472 3544 3488
rect 3576 3472 3592 3488
rect 4776 3472 4808 3488
rect 5320 3472 5336 3488
rect 5448 3472 5464 3488
rect 6056 3472 6072 3488
rect 6408 3472 6424 3488
rect 6488 3472 6504 3488
rect 6536 3472 6552 3488
rect 6632 3472 6648 3488
rect 6712 3472 6728 3488
rect 7224 3472 7240 3488
rect 1016 3452 1032 3468
rect 2264 3452 2280 3468
rect 4744 3452 4760 3468
rect 5288 3452 5304 3468
rect 5336 3452 5352 3468
rect 5416 3452 5432 3468
rect 6232 3452 6248 3468
rect 6632 3452 6648 3468
rect 7144 3452 7160 3468
rect 200 3432 216 3448
rect 488 3432 504 3448
rect 2216 3432 2232 3448
rect 2584 3432 2600 3448
rect 2904 3432 2920 3448
rect 3032 3432 3048 3448
rect 3736 3432 3752 3448
rect 5128 3432 5144 3448
rect 5400 3432 5416 3448
rect 5608 3432 5624 3448
rect 5944 3432 5960 3448
rect 6360 3432 6376 3448
rect 6648 3432 6664 3448
rect 6760 3432 6776 3448
rect 7128 3432 7144 3448
rect 7336 3432 7352 3448
rect 2157 3402 2193 3418
rect 4205 3402 4241 3418
rect 6237 3402 6273 3418
rect 200 3372 216 3388
rect 440 3372 456 3388
rect 680 3372 696 3388
rect 808 3372 824 3388
rect 840 3372 856 3388
rect 1048 3372 1064 3388
rect 1224 3372 1240 3388
rect 1352 3372 1368 3388
rect 1640 3372 1656 3388
rect 1944 3372 1960 3388
rect 2104 3372 2120 3388
rect 2216 3372 2232 3388
rect 2296 3372 2312 3388
rect 2504 3372 2520 3388
rect 2600 3372 2616 3388
rect 2648 3372 2664 3388
rect 2728 3372 2744 3388
rect 2808 3372 2824 3388
rect 3080 3372 3112 3388
rect 3352 3372 3368 3388
rect 3448 3372 3464 3388
rect 3672 3372 3688 3388
rect 3800 3372 3816 3388
rect 3848 3372 3864 3388
rect 4168 3372 4184 3388
rect 4280 3372 4296 3388
rect 4360 3372 4376 3388
rect 4408 3372 4424 3388
rect 4472 3372 4488 3388
rect 4504 3372 4520 3388
rect 4568 3372 4584 3388
rect 4616 3372 4632 3388
rect 4680 3372 4696 3388
rect 4808 3372 4824 3388
rect 5080 3372 5096 3388
rect 5416 3372 5432 3388
rect 5464 3372 5480 3388
rect 5560 3372 5576 3388
rect 5736 3372 5752 3388
rect 5800 3372 5816 3388
rect 6056 3372 6072 3388
rect 6120 3372 6136 3388
rect 6280 3372 6296 3388
rect 6584 3372 6600 3388
rect 6728 3372 6744 3388
rect 6824 3372 6840 3388
rect 7016 3372 7032 3388
rect 7208 3372 7224 3388
rect 7384 3372 7400 3388
rect 920 3352 936 3368
rect 2136 3352 2152 3368
rect 2184 3352 2200 3368
rect 2776 3352 2792 3368
rect 2888 3352 2904 3368
rect 2952 3352 2968 3368
rect 3176 3352 3192 3368
rect 3272 3352 3288 3368
rect 4120 3352 4136 3368
rect 4248 3352 4264 3368
rect 4664 3352 4680 3368
rect 5096 3352 5112 3368
rect 5256 3352 5272 3368
rect 5336 3352 5352 3368
rect 5528 3352 5544 3368
rect 5992 3352 6008 3368
rect 6360 3352 6376 3368
rect 6712 3352 6728 3368
rect 6776 3352 6792 3368
rect 7272 3352 7288 3368
rect 312 3332 328 3348
rect 392 3332 408 3348
rect 488 3332 504 3348
rect 744 3332 776 3348
rect 856 3332 872 3348
rect 1096 3332 1112 3348
rect 1192 3332 1208 3348
rect 1448 3332 1464 3348
rect 1528 3332 1544 3348
rect 1688 3332 1704 3348
rect 1752 3332 1768 3348
rect 1816 3332 1832 3348
rect 2008 3332 2024 3348
rect 2056 3332 2072 3348
rect 2440 3332 2472 3348
rect 2520 3332 2536 3348
rect 2552 3332 2568 3348
rect 2680 3332 2696 3348
rect 2760 3332 2776 3348
rect 3320 3332 3352 3348
rect 3384 3332 3400 3348
rect 3480 3332 3496 3348
rect 3544 3332 3560 3348
rect 3688 3332 3704 3348
rect 3784 3332 3800 3348
rect 3832 3332 3848 3348
rect 3880 3332 3896 3348
rect 3912 3332 3928 3348
rect 56 3314 72 3330
rect 104 3312 120 3328
rect 296 3312 312 3328
rect 408 3312 424 3328
rect 584 3312 600 3328
rect 616 3312 632 3328
rect 696 3312 712 3328
rect 728 3312 744 3328
rect 776 3312 792 3328
rect 936 3312 952 3328
rect 456 3292 472 3308
rect 696 3292 712 3308
rect 808 3292 840 3308
rect 1096 3292 1112 3308
rect 1176 3312 1192 3328
rect 1256 3312 1272 3328
rect 1320 3312 1336 3328
rect 1384 3312 1416 3328
rect 1560 3312 1576 3328
rect 1688 3292 1704 3308
rect 1736 3312 1752 3328
rect 1832 3312 1848 3328
rect 1960 3312 1976 3328
rect 1992 3312 2008 3328
rect 1960 3292 1976 3308
rect 2072 3312 2088 3328
rect 2248 3312 2280 3328
rect 2344 3312 2360 3328
rect 2392 3312 2408 3328
rect 2472 3312 2488 3328
rect 2616 3312 2632 3328
rect 2840 3312 2856 3328
rect 2968 3312 2984 3328
rect 3128 3312 3144 3328
rect 2040 3292 2056 3308
rect 2376 3292 2392 3308
rect 2552 3292 2568 3308
rect 2600 3292 2616 3308
rect 2696 3292 2744 3308
rect 2808 3292 2824 3308
rect 3096 3292 3112 3308
rect 3256 3292 3272 3308
rect 3304 3312 3320 3328
rect 3400 3312 3432 3328
rect 3560 3312 3576 3328
rect 3704 3312 3720 3328
rect 3368 3292 3384 3308
rect 3432 3292 3464 3308
rect 3912 3312 3928 3328
rect 3976 3312 3992 3328
rect 4072 3332 4088 3348
rect 4328 3332 4344 3348
rect 4424 3332 4440 3348
rect 4664 3332 4680 3348
rect 4712 3332 4728 3348
rect 4776 3332 4792 3348
rect 4888 3332 4904 3348
rect 4920 3332 4936 3348
rect 5112 3332 5128 3348
rect 5176 3332 5192 3348
rect 5352 3332 5368 3348
rect 5448 3332 5464 3348
rect 6104 3332 6120 3348
rect 6280 3332 6296 3348
rect 6344 3332 6360 3348
rect 6392 3332 6408 3348
rect 6424 3332 6440 3348
rect 6632 3332 6648 3348
rect 6696 3332 6712 3348
rect 6744 3332 6760 3348
rect 6904 3332 6920 3348
rect 7032 3332 7048 3348
rect 7176 3332 7192 3348
rect 7272 3332 7288 3348
rect 4088 3312 4104 3328
rect 4136 3312 4152 3328
rect 4184 3312 4200 3328
rect 4312 3312 4328 3328
rect 4360 3312 4376 3328
rect 4536 3312 4552 3328
rect 4600 3312 4616 3328
rect 4696 3312 4728 3328
rect 4840 3312 4856 3328
rect 4936 3312 4952 3328
rect 5000 3312 5016 3328
rect 5064 3312 5080 3328
rect 5160 3312 5176 3328
rect 5368 3312 5384 3328
rect 5432 3312 5448 3328
rect 5496 3312 5512 3328
rect 5576 3312 5592 3328
rect 5624 3312 5640 3328
rect 5704 3312 5736 3328
rect 5768 3312 5784 3328
rect 5832 3312 5848 3328
rect 5896 3312 5912 3328
rect 5944 3312 5960 3328
rect 6024 3312 6040 3328
rect 6088 3312 6104 3328
rect 6152 3312 6184 3328
rect 6328 3312 6344 3328
rect 6408 3312 6424 3328
rect 6488 3312 6504 3328
rect 6552 3312 6568 3328
rect 6616 3312 6632 3328
rect 6680 3312 6696 3328
rect 6776 3312 6792 3328
rect 6856 3312 6872 3328
rect 6952 3312 6968 3328
rect 6984 3312 7000 3328
rect 7064 3312 7080 3328
rect 7144 3312 7160 3328
rect 7176 3312 7192 3328
rect 7240 3312 7256 3328
rect 7336 3312 7352 3328
rect 3752 3292 3768 3308
rect 3800 3292 3816 3308
rect 3848 3292 3864 3308
rect 3896 3292 3912 3308
rect 3960 3292 3976 3308
rect 4024 3292 4040 3308
rect 4120 3292 4136 3308
rect 4360 3292 4376 3308
rect 4472 3292 4488 3308
rect 4616 3292 4632 3308
rect 4728 3292 4744 3308
rect 4760 3292 4776 3308
rect 4808 3292 4840 3308
rect 4888 3292 4904 3308
rect 4968 3292 4984 3308
rect 5288 3292 5304 3308
rect 5416 3292 5432 3308
rect 5592 3292 5624 3308
rect 5784 3292 5800 3308
rect 5832 3292 5848 3308
rect 5864 3292 5880 3308
rect 5928 3292 5944 3308
rect 6504 3292 6520 3308
rect 6568 3292 6584 3308
rect 6968 3292 6984 3308
rect 7048 3292 7064 3308
rect 7112 3292 7128 3308
rect 7160 3292 7176 3308
rect 3704 3272 3720 3288
rect 3928 3272 3944 3288
rect 3992 3272 4008 3288
rect 4056 3272 4072 3288
rect 4856 3272 4872 3288
rect 3976 3252 3992 3268
rect 4840 3252 4856 3268
rect 5640 3272 5656 3288
rect 5672 3272 5704 3288
rect 5752 3272 5768 3288
rect 5816 3272 5832 3288
rect 5880 3272 5896 3288
rect 5912 3272 5928 3288
rect 6472 3272 6488 3288
rect 6536 3272 6552 3288
rect 5944 3252 5960 3268
rect 6936 3272 6952 3288
rect 7080 3272 7096 3288
rect 7128 3272 7144 3288
rect 6952 3252 6968 3268
rect 7064 3252 7080 3268
rect 184 3232 200 3248
rect 680 3232 696 3248
rect 1288 3232 1304 3248
rect 2216 3232 2232 3248
rect 2344 3232 2360 3248
rect 2792 3232 2808 3248
rect 4568 3232 4584 3248
rect 4904 3232 4920 3248
rect 5032 3232 5048 3248
rect 5192 3232 5208 3248
rect 5224 3232 5240 3248
rect 6648 3232 6664 3248
rect 6744 3232 6760 3248
rect 1117 3202 1153 3218
rect 3165 3202 3201 3218
rect 5213 3202 5249 3218
rect 24 3172 40 3188
rect 152 3172 168 3188
rect 216 3172 232 3188
rect 264 3172 280 3188
rect 632 3172 648 3188
rect 2008 3172 2024 3188
rect 2504 3172 2520 3188
rect 2712 3172 2728 3188
rect 3752 3172 3768 3188
rect 3832 3172 3848 3188
rect 4040 3172 4056 3188
rect 4328 3172 4344 3188
rect 4376 3172 4392 3188
rect 4424 3172 4440 3188
rect 4520 3172 4536 3188
rect 4616 3172 4632 3188
rect 4680 3172 4696 3188
rect 4776 3172 4792 3188
rect 4808 3172 4824 3188
rect 4872 3172 4888 3188
rect 5528 3172 5544 3188
rect 5592 3172 5608 3188
rect 5672 3172 5688 3188
rect 5704 3172 5720 3188
rect 5784 3172 5800 3188
rect 5816 3172 5832 3188
rect 6424 3172 6440 3188
rect 6680 3172 6696 3188
rect 6728 3172 6744 3188
rect 7096 3172 7112 3188
rect 120 3132 136 3148
rect 472 3132 488 3148
rect 552 3132 568 3148
rect 664 3132 680 3148
rect 968 3132 984 3148
rect 1112 3132 1128 3148
rect 1160 3132 1176 3148
rect 1528 3132 1544 3148
rect 2472 3132 2488 3148
rect 3768 3132 3784 3148
rect 3816 3132 3832 3148
rect 4312 3132 4328 3148
rect 4360 3132 4376 3148
rect 4440 3132 4456 3148
rect 4504 3132 4520 3148
rect 4616 3132 4632 3148
rect 4696 3132 4712 3148
rect 4760 3132 4776 3148
rect 4824 3132 4840 3148
rect 5000 3132 5016 3148
rect 5368 3132 5384 3148
rect 5512 3132 5528 3148
rect 5576 3132 5592 3148
rect 5656 3132 5672 3148
rect 5720 3132 5736 3148
rect 5768 3132 5784 3148
rect 5832 3132 5848 3148
rect 7064 3132 7080 3148
rect 7112 3132 7128 3148
rect 56 3112 72 3128
rect 504 3112 520 3128
rect 24 3092 40 3108
rect 88 3092 120 3108
rect 184 3092 200 3108
rect 232 3092 248 3108
rect 360 3092 376 3108
rect 408 3092 424 3108
rect 504 3092 520 3108
rect 584 3092 600 3108
rect 696 3092 712 3108
rect 744 3112 760 3128
rect 840 3090 856 3106
rect 904 3092 920 3108
rect 1000 3092 1016 3108
rect 1048 3112 1064 3128
rect 1608 3112 1624 3128
rect 1240 3092 1256 3108
rect 1368 3092 1384 3108
rect 1448 3092 1464 3108
rect 1644 3112 1660 3128
rect 1736 3112 1752 3128
rect 1944 3112 1960 3128
rect 2040 3112 2056 3128
rect 2136 3112 2152 3128
rect 2184 3112 2200 3128
rect 2488 3112 2504 3128
rect 2728 3112 2744 3128
rect 2824 3112 2840 3128
rect 1656 3092 1672 3108
rect 1704 3092 1720 3108
rect 1800 3090 1816 3106
rect 1944 3092 1960 3108
rect 2008 3092 2024 3108
rect 2104 3092 2120 3108
rect 2280 3092 2296 3108
rect 2344 3090 2360 3106
rect 2600 3092 2616 3108
rect 2760 3092 2776 3108
rect 2904 3112 2920 3128
rect 3064 3112 3080 3128
rect 3176 3112 3192 3128
rect 3256 3112 3272 3128
rect 3288 3112 3304 3128
rect 3352 3112 3368 3128
rect 2872 3092 2888 3108
rect 2952 3092 2968 3108
rect 3016 3092 3032 3108
rect 3064 3092 3080 3108
rect 3096 3092 3112 3108
rect 8 3072 24 3088
rect 72 3072 88 3088
rect 312 3072 328 3088
rect 360 3072 376 3088
rect 488 3072 504 3088
rect 616 3072 632 3088
rect 680 3072 696 3088
rect 744 3072 760 3088
rect 776 3072 792 3088
rect 984 3072 1000 3088
rect 1048 3072 1064 3088
rect 1112 3072 1128 3088
rect 1288 3072 1304 3088
rect 1336 3072 1352 3088
rect 1400 3072 1416 3088
rect 1544 3072 1560 3088
rect 1672 3072 1688 3088
rect 1736 3072 1752 3088
rect 1768 3072 1784 3088
rect 1976 3072 2008 3088
rect 2184 3072 2200 3088
rect 2232 3072 2248 3088
rect 2312 3072 2328 3088
rect 2408 3072 2424 3088
rect 2520 3072 2536 3088
rect 2552 3072 2568 3088
rect 2744 3072 2760 3088
rect 2776 3072 2808 3088
rect 2824 3072 2840 3088
rect 2888 3072 2904 3088
rect 2936 3072 2952 3088
rect 3000 3072 3016 3088
rect 3080 3072 3096 3088
rect 3144 3072 3160 3088
rect 3320 3092 3336 3108
rect 3368 3092 3400 3108
rect 3432 3112 3448 3128
rect 3768 3112 3784 3128
rect 3800 3112 3816 3128
rect 3528 3090 3544 3106
rect 3752 3092 3768 3108
rect 3800 3092 3816 3108
rect 3848 3092 3864 3108
rect 3928 3092 3944 3108
rect 3976 3112 3992 3128
rect 4280 3112 4296 3128
rect 4392 3112 4408 3128
rect 4424 3112 4440 3128
rect 4488 3112 4504 3128
rect 4552 3112 4568 3128
rect 4600 3112 4616 3128
rect 4664 3112 4680 3128
rect 4728 3112 4744 3128
rect 4792 3112 4808 3128
rect 4920 3112 4936 3128
rect 4968 3112 4984 3128
rect 5544 3112 5560 3128
rect 5608 3112 5640 3128
rect 5688 3112 5704 3128
rect 5800 3112 5816 3128
rect 5864 3112 5880 3128
rect 6824 3112 6840 3128
rect 7080 3112 7096 3128
rect 4168 3092 4184 3108
rect 4296 3092 4312 3108
rect 4376 3092 4392 3108
rect 4424 3092 4440 3108
rect 4488 3092 4504 3108
rect 4584 3092 4600 3108
rect 4616 3092 4632 3108
rect 4680 3092 4696 3108
rect 4744 3092 4760 3108
rect 4808 3092 4824 3108
rect 4888 3092 4904 3108
rect 4920 3092 4936 3108
rect 4984 3092 5000 3108
rect 5080 3092 5096 3108
rect 5144 3092 5160 3108
rect 5176 3092 5192 3108
rect 5256 3092 5272 3108
rect 5384 3092 5400 3108
rect 5448 3092 5464 3108
rect 5528 3092 5544 3108
rect 5592 3092 5608 3108
rect 5640 3092 5656 3108
rect 5704 3092 5720 3108
rect 5784 3092 5800 3108
rect 5848 3092 5864 3108
rect 5880 3092 5896 3108
rect 5944 3092 5960 3108
rect 6104 3092 6120 3108
rect 6184 3092 6200 3108
rect 6264 3092 6280 3108
rect 6376 3092 6408 3108
rect 6584 3090 6600 3106
rect 6648 3092 6664 3108
rect 6760 3092 6792 3108
rect 6840 3092 6856 3108
rect 6936 3090 6952 3106
rect 7096 3092 7112 3108
rect 7208 3092 7224 3108
rect 7336 3092 7352 3108
rect 7400 3092 7416 3108
rect 3304 3072 3320 3088
rect 3368 3072 3384 3088
rect 3416 3072 3432 3088
rect 3464 3072 3480 3088
rect 3544 3072 3560 3088
rect 3704 3072 3720 3088
rect 3912 3072 3928 3088
rect 3976 3072 3992 3088
rect 4904 3072 4920 3088
rect 5032 3072 5048 3088
rect 5096 3072 5112 3088
rect 5400 3072 5416 3088
rect 5896 3072 5912 3088
rect 5944 3072 5960 3088
rect 6152 3072 6168 3088
rect 6248 3072 6264 3088
rect 6312 3072 6328 3088
rect 6360 3072 6376 3088
rect 6568 3072 6584 3088
rect 6792 3072 6808 3088
rect 7160 3072 7176 3088
rect 7368 3072 7384 3088
rect 200 3052 216 3068
rect 2056 3052 2072 3068
rect 3224 3052 3256 3068
rect 3528 3052 3544 3068
rect 4024 3052 4040 3068
rect 4184 3052 4200 3068
rect 4856 3052 4872 3068
rect 5240 3052 5256 3068
rect 5416 3052 5432 3068
rect 5480 3052 5496 3068
rect 5976 3052 5992 3068
rect 6216 3052 6232 3068
rect 6248 3052 6264 3068
rect 6328 3052 6344 3068
rect 6424 3052 6440 3068
rect 6872 3052 6888 3068
rect 6936 3052 6952 3068
rect 7336 3052 7352 3068
rect 1928 3032 1944 3048
rect 2152 3032 2168 3048
rect 2248 3032 2264 3048
rect 2712 3032 2728 3048
rect 2920 3032 2936 3048
rect 2984 3032 3000 3048
rect 3128 3032 3144 3048
rect 3656 3032 3672 3048
rect 3688 3032 3704 3048
rect 3880 3032 3896 3048
rect 4056 3032 4072 3048
rect 6344 3032 6360 3048
rect 6456 3032 6472 3048
rect 7320 3032 7336 3048
rect 2157 3002 2193 3018
rect 4205 3002 4241 3018
rect 6237 3002 6273 3018
rect 24 2972 40 2988
rect 488 2972 504 2988
rect 584 2972 600 2988
rect 632 2972 648 2988
rect 808 2972 824 2988
rect 1352 2972 1368 2988
rect 1496 2972 1512 2988
rect 1880 2972 1896 2988
rect 1912 2972 1928 2988
rect 1960 2972 1976 2988
rect 2344 2972 2360 2988
rect 2376 2972 2392 2988
rect 2424 2972 2440 2988
rect 2488 2972 2504 2988
rect 2712 2972 2744 2988
rect 2792 2972 2808 2988
rect 2904 2972 2920 2988
rect 2968 2972 2984 2988
rect 3176 2972 3192 2988
rect 3512 2972 3528 2988
rect 3544 2972 3560 2988
rect 3784 2972 3800 2988
rect 3832 2972 3848 2988
rect 4504 2972 4520 2988
rect 4648 2972 4664 2988
rect 4744 2972 4760 2988
rect 5032 2972 5048 2988
rect 5400 2972 5416 2988
rect 6152 2972 6168 2988
rect 6376 2972 6392 2988
rect 6600 2972 6616 2988
rect 6776 2972 6792 2988
rect 7096 2972 7112 2988
rect 360 2952 376 2968
rect 504 2952 520 2968
rect 968 2952 984 2968
rect 3592 2952 3608 2968
rect 3672 2952 3688 2968
rect 4568 2952 4584 2968
rect 4696 2952 4712 2968
rect 4936 2952 4952 2968
rect 5576 2952 5592 2968
rect 72 2932 88 2948
rect 152 2932 168 2948
rect 200 2932 216 2948
rect 264 2932 280 2948
rect 296 2932 312 2948
rect 776 2932 792 2948
rect 824 2932 840 2948
rect 1032 2932 1048 2948
rect 1128 2932 1144 2948
rect 1256 2932 1272 2948
rect 1368 2932 1384 2948
rect 1464 2932 1480 2948
rect 1512 2932 1528 2948
rect 1576 2932 1608 2948
rect 1640 2932 1656 2948
rect 1688 2932 1704 2948
rect 1768 2932 1784 2948
rect 2008 2932 2040 2948
rect 2072 2932 2088 2948
rect 2248 2932 2264 2948
rect 2392 2932 2408 2948
rect 2552 2932 2568 2948
rect 2760 2932 2776 2948
rect 2808 2932 2824 2948
rect 2872 2932 2888 2948
rect 2920 2932 2936 2948
rect 2984 2932 3000 2948
rect 3256 2932 3272 2948
rect 3320 2932 3336 2948
rect 3352 2932 3368 2948
rect 3704 2932 3720 2948
rect 3736 2932 3752 2948
rect 3880 2932 3896 2948
rect 3944 2932 3960 2948
rect 3976 2932 3992 2948
rect 4216 2932 4232 2948
rect 4280 2932 4296 2948
rect 4312 2932 4328 2948
rect 4552 2932 4568 2948
rect 4728 2932 4744 2948
rect 4872 2932 4888 2948
rect 4968 2932 4984 2948
rect 5064 2932 5080 2948
rect 5240 2932 5256 2948
rect 5496 2932 5512 2948
rect 5576 2932 5592 2948
rect 6056 2932 6072 2948
rect 6104 2952 6120 2968
rect 6312 2932 6328 2948
rect 6568 2932 6600 2948
rect 6632 2952 6648 2968
rect 6808 2952 6824 2968
rect 7304 2952 7320 2968
rect 6712 2932 6728 2948
rect 6888 2932 6904 2948
rect 6936 2932 6952 2948
rect 7240 2932 7256 2948
rect 7384 2932 7400 2948
rect 72 2912 88 2928
rect 120 2912 136 2928
rect 184 2912 200 2928
rect 216 2912 232 2928
rect 360 2914 376 2930
rect 552 2912 568 2928
rect 600 2912 616 2928
rect 680 2912 696 2928
rect 264 2892 280 2908
rect 584 2892 600 2908
rect 712 2892 728 2908
rect 760 2912 776 2928
rect 952 2912 968 2928
rect 792 2892 808 2908
rect 1064 2892 1080 2908
rect 1112 2912 1128 2928
rect 1224 2914 1240 2930
rect 1384 2912 1400 2928
rect 1112 2892 1128 2908
rect 1528 2912 1544 2928
rect 1608 2912 1624 2928
rect 1432 2892 1448 2908
rect 1480 2892 1496 2908
rect 1752 2914 1768 2930
rect 1944 2912 1960 2928
rect 2072 2912 2104 2928
rect 2152 2912 2168 2928
rect 2216 2914 2232 2930
rect 2472 2912 2488 2928
rect 2520 2912 2536 2928
rect 2600 2912 2616 2928
rect 2824 2912 2840 2928
rect 2920 2912 2936 2928
rect 3064 2912 3080 2928
rect 3304 2912 3320 2928
rect 3384 2914 3400 2930
rect 3592 2912 3608 2928
rect 3640 2912 3656 2928
rect 3720 2912 3736 2928
rect 3752 2912 3768 2928
rect 3864 2912 3896 2928
rect 1656 2892 1672 2908
rect 1960 2892 1976 2908
rect 2136 2892 2152 2908
rect 2360 2892 2376 2908
rect 2728 2892 2744 2908
rect 2888 2892 2904 2908
rect 3208 2892 3224 2908
rect 3304 2892 3320 2908
rect 3672 2892 3704 2908
rect 4040 2914 4056 2930
rect 4104 2912 4120 2928
rect 4232 2912 4248 2928
rect 3944 2892 3960 2908
rect 4376 2914 4392 2930
rect 4440 2912 4456 2928
rect 4616 2912 4632 2928
rect 4696 2912 4712 2928
rect 4808 2912 4824 2928
rect 4872 2912 4888 2928
rect 4936 2912 4952 2928
rect 5064 2912 5096 2928
rect 5144 2912 5160 2928
rect 5288 2912 5304 2928
rect 5432 2912 5448 2928
rect 5480 2912 5496 2928
rect 5544 2912 5560 2928
rect 5640 2912 5656 2928
rect 5688 2912 5704 2928
rect 5736 2912 5752 2928
rect 5800 2912 5816 2928
rect 5880 2912 5896 2928
rect 5928 2912 5944 2928
rect 6024 2912 6056 2928
rect 6104 2912 6120 2928
rect 6136 2912 6152 2928
rect 6264 2912 6280 2928
rect 6440 2912 6456 2928
rect 6488 2912 6504 2928
rect 6568 2912 6584 2928
rect 6664 2912 6696 2928
rect 6744 2912 6760 2928
rect 6840 2912 6856 2928
rect 6872 2912 6888 2928
rect 6904 2912 6920 2928
rect 6968 2914 6984 2930
rect 7128 2912 7144 2928
rect 7208 2912 7224 2928
rect 7288 2912 7304 2928
rect 7336 2912 7352 2928
rect 7400 2912 7416 2928
rect 4280 2892 4296 2908
rect 4568 2892 4584 2908
rect 4648 2892 4664 2908
rect 4712 2892 4728 2908
rect 4776 2892 4808 2908
rect 4888 2892 4904 2908
rect 4952 2892 4968 2908
rect 5000 2892 5016 2908
rect 5080 2892 5096 2908
rect 5128 2892 5144 2908
rect 5416 2892 5432 2908
rect 5704 2892 5720 2908
rect 5784 2892 5800 2908
rect 5912 2892 5928 2908
rect 5992 2892 6008 2908
rect 7112 2892 7128 2908
rect 7224 2892 7240 2908
rect 760 2872 776 2888
rect 840 2872 856 2888
rect 1320 2872 1336 2888
rect 2312 2872 2328 2888
rect 2760 2872 2776 2888
rect 3144 2872 3160 2888
rect 4168 2872 4184 2888
rect 4520 2872 4536 2888
rect 4680 2872 4696 2888
rect 4808 2872 4824 2888
rect 4856 2872 4872 2888
rect 4920 2872 4936 2888
rect 5160 2872 5176 2888
rect 5448 2872 5464 2888
rect 5672 2872 5704 2888
rect 5528 2852 5544 2868
rect 5752 2872 5768 2888
rect 5816 2872 5832 2888
rect 5864 2872 5880 2888
rect 5944 2872 5960 2888
rect 7144 2872 7160 2888
rect 7176 2872 7208 2888
rect 632 2832 648 2848
rect 1384 2832 1400 2848
rect 5432 2832 5448 2848
rect 5688 2832 5704 2848
rect 5800 2832 5816 2848
rect 5848 2832 5864 2848
rect 5928 2832 5944 2848
rect 7160 2832 7176 2848
rect 7352 2832 7368 2848
rect 1117 2802 1153 2818
rect 3165 2802 3201 2818
rect 5213 2802 5249 2818
rect 392 2772 408 2788
rect 600 2772 632 2788
rect 744 2772 760 2788
rect 792 2772 808 2788
rect 1128 2772 1144 2788
rect 1432 2772 1448 2788
rect 1464 2772 1480 2788
rect 1704 2772 1720 2788
rect 1960 2772 1976 2788
rect 1992 2772 2008 2788
rect 2168 2772 2184 2788
rect 3496 2772 3512 2788
rect 3576 2772 3592 2788
rect 3736 2772 3752 2788
rect 4344 2772 4360 2788
rect 4840 2772 4856 2788
rect 4968 2772 4984 2788
rect 5016 2772 5032 2788
rect 5704 2772 5720 2788
rect 5736 2772 5752 2788
rect 6200 2772 6216 2788
rect 7080 2772 7096 2788
rect 7128 2772 7144 2788
rect 7208 2772 7240 2788
rect 1672 2752 1688 2768
rect 2056 2752 2072 2768
rect 2232 2752 2248 2768
rect 2856 2752 2872 2768
rect 3048 2752 3064 2768
rect 8 2732 24 2748
rect 456 2732 472 2748
rect 1768 2732 1784 2748
rect 2088 2732 2104 2748
rect 2472 2732 2488 2748
rect 3320 2732 3336 2748
rect 4360 2732 4376 2748
rect 4584 2732 4600 2748
rect 4648 2732 4664 2748
rect 4904 2732 4920 2748
rect 5368 2732 5384 2748
rect 5496 2732 5512 2748
rect 232 2712 248 2728
rect 136 2690 152 2706
rect 268 2712 284 2728
rect 424 2712 440 2728
rect 520 2712 536 2728
rect 728 2712 744 2728
rect 760 2712 776 2728
rect 872 2712 888 2728
rect 952 2712 968 2728
rect 1032 2712 1048 2728
rect 1144 2712 1160 2728
rect 1480 2712 1496 2728
rect 280 2692 296 2708
rect 312 2692 328 2708
rect 568 2692 584 2708
rect 680 2692 696 2708
rect 712 2692 728 2708
rect 840 2692 856 2708
rect 968 2692 984 2708
rect 1016 2692 1032 2708
rect 1080 2692 1112 2708
rect 1240 2692 1256 2708
rect 1336 2692 1352 2708
rect 1560 2692 1576 2708
rect 1736 2692 1752 2708
rect 1768 2692 1784 2708
rect 1816 2712 1832 2728
rect 1896 2712 1912 2728
rect 2104 2712 2120 2728
rect 2504 2712 2520 2728
rect 2024 2692 2040 2708
rect 2136 2692 2152 2708
rect 2264 2692 2280 2708
rect 2344 2692 2360 2708
rect 2936 2712 2952 2728
rect 2984 2712 3000 2728
rect 3080 2712 3096 2728
rect 3352 2712 3368 2728
rect 2552 2692 2568 2708
rect 2584 2692 2600 2708
rect 168 2672 184 2688
rect 200 2672 216 2688
rect 296 2672 312 2688
rect 360 2672 392 2688
rect 488 2672 520 2688
rect 648 2672 664 2688
rect 760 2672 776 2688
rect 808 2672 840 2688
rect 888 2672 904 2688
rect 920 2672 936 2688
rect 952 2672 968 2688
rect 1112 2672 1128 2688
rect 1144 2672 1160 2688
rect 1208 2676 1224 2692
rect 1320 2672 1336 2688
rect 1448 2672 1464 2688
rect 1544 2672 1560 2688
rect 1752 2672 1768 2688
rect 1848 2672 1912 2688
rect 1928 2676 1944 2692
rect 2776 2690 2792 2706
rect 2856 2692 2872 2708
rect 3000 2692 3016 2708
rect 2008 2672 2024 2688
rect 2072 2672 2088 2688
rect 2104 2672 2120 2688
rect 2296 2672 2312 2688
rect 2392 2672 2408 2688
rect 2472 2672 2488 2688
rect 2504 2672 2520 2688
rect 2568 2672 2584 2688
rect 2632 2672 2648 2688
rect 2808 2672 2824 2688
rect 2840 2672 2856 2688
rect 2904 2672 2920 2688
rect 2984 2672 3000 2688
rect 3048 2692 3064 2708
rect 3208 2692 3224 2708
rect 3388 2712 3404 2728
rect 3432 2712 3448 2728
rect 3528 2712 3544 2728
rect 3400 2692 3416 2708
rect 3448 2692 3464 2708
rect 3032 2672 3048 2688
rect 3144 2672 3160 2688
rect 3320 2672 3336 2688
rect 3416 2672 3432 2688
rect 3496 2692 3512 2708
rect 3544 2692 3560 2708
rect 3624 2692 3640 2708
rect 3672 2712 3688 2728
rect 4216 2712 4232 2728
rect 4328 2712 4344 2728
rect 4616 2712 4632 2728
rect 4664 2712 4680 2728
rect 4728 2712 4744 2728
rect 4776 2712 4792 2728
rect 4872 2712 4888 2728
rect 5144 2712 5160 2728
rect 5304 2712 5320 2728
rect 5336 2712 5352 2728
rect 5528 2712 5544 2728
rect 5576 2732 5592 2748
rect 5752 2732 5768 2748
rect 5944 2732 5960 2748
rect 5976 2732 5992 2748
rect 6024 2732 6040 2748
rect 7064 2732 7080 2748
rect 7096 2732 7112 2748
rect 7256 2732 7272 2748
rect 5624 2712 5640 2728
rect 5656 2712 5672 2728
rect 5784 2712 5800 2728
rect 5912 2712 5944 2728
rect 6008 2712 6024 2728
rect 6168 2712 6184 2728
rect 7096 2712 7128 2728
rect 3864 2692 3880 2708
rect 4040 2692 4072 2708
rect 4184 2692 4200 2708
rect 4264 2692 4280 2708
rect 4344 2692 4360 2708
rect 4392 2692 4408 2708
rect 4424 2692 4440 2708
rect 4488 2692 4504 2708
rect 4520 2692 4552 2708
rect 4600 2692 4616 2708
rect 4664 2692 4680 2708
rect 4728 2692 4760 2708
rect 4808 2692 4824 2708
rect 4888 2692 4904 2708
rect 4936 2692 4952 2708
rect 5048 2692 5080 2708
rect 5256 2692 5272 2708
rect 5304 2692 5320 2708
rect 5416 2692 5432 2708
rect 5512 2692 5528 2708
rect 5560 2692 5576 2708
rect 5624 2692 5640 2708
rect 5672 2692 5688 2708
rect 5768 2692 5784 2708
rect 5800 2692 5816 2708
rect 5880 2692 5896 2708
rect 5960 2692 5976 2708
rect 6008 2692 6024 2708
rect 6088 2692 6104 2708
rect 6152 2692 6168 2708
rect 6328 2692 6344 2708
rect 6392 2690 6408 2706
rect 6440 2692 6456 2708
rect 6536 2692 6552 2708
rect 6648 2692 6664 2708
rect 6744 2692 6760 2708
rect 6904 2692 6936 2708
rect 6984 2692 7000 2708
rect 7080 2692 7096 2708
rect 7128 2692 7144 2708
rect 7208 2692 7224 2708
rect 7288 2692 7304 2708
rect 7352 2690 7368 2706
rect 3480 2672 3496 2688
rect 3608 2672 3624 2688
rect 3672 2672 3688 2688
rect 3912 2672 3928 2688
rect 4248 2672 4264 2688
rect 4424 2672 4440 2688
rect 4504 2672 4520 2688
rect 4744 2672 4760 2688
rect 5208 2672 5224 2688
rect 5272 2672 5288 2688
rect 5432 2672 5448 2688
rect 5608 2672 5624 2688
rect 5864 2672 5880 2688
rect 5896 2672 5912 2688
rect 6104 2672 6136 2688
rect 6600 2672 6616 2688
rect 6680 2672 6696 2688
rect 392 2652 408 2668
rect 536 2652 552 2668
rect 664 2652 696 2668
rect 712 2652 728 2668
rect 1000 2652 1016 2668
rect 1048 2652 1064 2668
rect 1976 2652 1992 2668
rect 2952 2652 2968 2668
rect 3720 2652 3736 2668
rect 4296 2652 4312 2668
rect 4392 2652 4408 2668
rect 4792 2652 4808 2668
rect 5224 2652 5240 2668
rect 5448 2652 5464 2668
rect 6168 2652 6184 2668
rect 6232 2652 6248 2668
rect 7176 2652 7192 2668
rect 7256 2652 7272 2668
rect 424 2632 440 2648
rect 616 2632 632 2648
rect 744 2632 760 2648
rect 792 2632 808 2648
rect 904 2632 920 2648
rect 952 2632 968 2648
rect 1704 2632 1720 2648
rect 2648 2632 2664 2648
rect 3752 2632 3768 2648
rect 4120 2632 4136 2648
rect 4920 2632 4936 2648
rect 4968 2632 4984 2648
rect 5096 2632 5112 2648
rect 5560 2632 5576 2648
rect 5704 2632 5720 2648
rect 5832 2632 5848 2648
rect 6056 2632 6072 2648
rect 6136 2632 6152 2648
rect 6296 2632 6312 2648
rect 6520 2632 6536 2648
rect 6568 2632 6584 2648
rect 6840 2632 6856 2648
rect 6872 2632 6888 2648
rect 6952 2632 6968 2648
rect 7016 2632 7032 2648
rect 2157 2602 2193 2618
rect 4205 2602 4241 2618
rect 6237 2602 6273 2618
rect 88 2572 104 2588
rect 248 2572 264 2588
rect 584 2572 616 2588
rect 664 2572 680 2588
rect 776 2572 792 2588
rect 872 2572 888 2588
rect 1016 2572 1032 2588
rect 1384 2572 1400 2588
rect 2120 2572 2152 2588
rect 2264 2572 2296 2588
rect 2408 2572 2424 2588
rect 2600 2572 2616 2588
rect 3032 2572 3048 2588
rect 3416 2572 3432 2588
rect 3480 2572 3496 2588
rect 3640 2572 3656 2588
rect 3976 2572 3992 2588
rect 4040 2572 4056 2588
rect 4168 2572 4184 2588
rect 4392 2572 4408 2588
rect 4568 2572 4584 2588
rect 5240 2572 5256 2588
rect 5432 2572 5448 2588
rect 5976 2572 5992 2588
rect 6376 2572 6392 2588
rect 6744 2572 6760 2588
rect 104 2552 120 2568
rect 264 2552 280 2568
rect 824 2552 840 2568
rect 920 2552 936 2568
rect 1032 2552 1048 2568
rect 1080 2552 1096 2568
rect 1112 2552 1128 2568
rect 1192 2552 1208 2568
rect 2152 2552 2168 2568
rect 2904 2552 2920 2568
rect 8 2532 24 2548
rect 184 2532 200 2548
rect 280 2532 296 2548
rect 392 2532 408 2548
rect 632 2532 664 2548
rect 760 2532 776 2548
rect 856 2532 872 2548
rect 904 2532 920 2548
rect 984 2532 1000 2548
rect 1144 2532 1160 2548
rect 1400 2532 1416 2548
rect 1432 2532 1448 2548
rect 1496 2532 1512 2548
rect 1720 2532 1752 2548
rect 1784 2532 1800 2548
rect 1848 2532 1864 2548
rect 1880 2532 1896 2548
rect 2056 2532 2072 2548
rect 2088 2532 2104 2548
rect 2168 2532 2184 2548
rect 2216 2532 2232 2548
rect 2312 2532 2344 2548
rect 2376 2532 2392 2548
rect 2440 2532 2456 2548
rect 2616 2532 2632 2548
rect 2648 2532 2664 2548
rect 2712 2532 2728 2548
rect 3048 2532 3064 2548
rect 3144 2532 3160 2548
rect 3464 2552 3480 2568
rect 3224 2532 3240 2548
rect 24 2512 40 2528
rect 104 2512 120 2528
rect 136 2512 152 2528
rect 296 2512 312 2528
rect 56 2492 72 2508
rect 216 2492 232 2508
rect 328 2492 344 2508
rect 376 2512 392 2528
rect 456 2514 472 2530
rect 520 2512 536 2528
rect 696 2512 712 2528
rect 808 2512 824 2528
rect 984 2512 1000 2528
rect 1064 2512 1080 2528
rect 1160 2512 1176 2528
rect 1272 2512 1288 2528
rect 1320 2512 1336 2528
rect 1416 2512 1432 2528
rect 376 2492 392 2508
rect 600 2492 616 2508
rect 680 2492 696 2508
rect 856 2492 872 2508
rect 968 2492 984 2508
rect 1016 2492 1032 2508
rect 1512 2512 1544 2528
rect 1576 2512 1592 2528
rect 1608 2512 1624 2528
rect 1672 2512 1688 2528
rect 1800 2512 1816 2528
rect 1464 2492 1480 2508
rect 1640 2492 1656 2508
rect 1768 2492 1784 2508
rect 1992 2512 2008 2528
rect 2232 2512 2248 2528
rect 2488 2512 2504 2528
rect 2632 2512 2648 2528
rect 1848 2492 1864 2508
rect 2120 2492 2136 2508
rect 2280 2492 2296 2508
rect 2360 2492 2376 2508
rect 2408 2492 2424 2508
rect 2776 2512 2808 2528
rect 2920 2512 2936 2528
rect 3064 2512 3080 2528
rect 3272 2532 3288 2548
rect 3320 2532 3336 2548
rect 3400 2532 3416 2548
rect 3496 2532 3512 2548
rect 3608 2532 3624 2548
rect 3688 2532 3704 2548
rect 3736 2532 3752 2548
rect 3784 2532 3800 2548
rect 3992 2532 4008 2548
rect 4088 2532 4104 2548
rect 4200 2532 4216 2548
rect 4344 2532 4360 2548
rect 4376 2532 4392 2548
rect 4664 2532 4680 2548
rect 4808 2532 4824 2548
rect 4920 2532 4936 2548
rect 4952 2532 4968 2548
rect 5016 2532 5032 2548
rect 5096 2532 5112 2548
rect 5272 2532 5288 2548
rect 5320 2552 5336 2568
rect 5720 2552 5736 2568
rect 5480 2532 5496 2548
rect 6440 2552 6456 2568
rect 6808 2552 6824 2568
rect 5768 2532 5784 2548
rect 5848 2532 5864 2548
rect 6360 2532 6376 2548
rect 6696 2532 6712 2548
rect 6728 2532 6744 2548
rect 6872 2532 6888 2548
rect 7096 2532 7112 2548
rect 2680 2492 2696 2508
rect 2824 2492 2840 2508
rect 3064 2492 3080 2508
rect 3288 2512 3304 2528
rect 3336 2512 3352 2528
rect 3448 2512 3464 2528
rect 3512 2512 3528 2528
rect 3544 2512 3576 2528
rect 3672 2512 3688 2528
rect 3704 2512 3720 2528
rect 3112 2492 3128 2508
rect 3224 2492 3240 2508
rect 3256 2492 3272 2508
rect 3320 2492 3336 2508
rect 3544 2492 3560 2508
rect 3848 2514 3864 2530
rect 3912 2512 3928 2528
rect 4008 2512 4024 2528
rect 3752 2492 3768 2508
rect 4104 2512 4120 2528
rect 4248 2512 4264 2528
rect 4344 2512 4360 2528
rect 4456 2512 4472 2528
rect 4520 2512 4536 2528
rect 4632 2512 4648 2528
rect 4712 2512 4728 2528
rect 4792 2512 4808 2528
rect 4056 2492 4072 2508
rect 4136 2492 4152 2508
rect 4168 2492 4184 2508
rect 4360 2492 4376 2508
rect 4472 2492 4488 2508
rect 4536 2492 4568 2508
rect 4648 2492 4664 2508
rect 4952 2492 4968 2508
rect 5000 2512 5016 2528
rect 5112 2512 5128 2528
rect 5256 2512 5272 2528
rect 5288 2512 5304 2528
rect 5352 2512 5368 2528
rect 5400 2512 5416 2528
rect 5464 2512 5480 2528
rect 5528 2512 5544 2528
rect 5592 2512 5608 2528
rect 5656 2512 5672 2528
rect 5688 2512 5704 2528
rect 5784 2512 5800 2528
rect 5864 2512 5880 2528
rect 6008 2512 6024 2528
rect 6072 2512 6088 2528
rect 6136 2512 6152 2528
rect 6184 2512 6216 2528
rect 6296 2512 6312 2528
rect 6344 2512 6360 2528
rect 6408 2512 6424 2528
rect 6472 2512 6488 2528
rect 6552 2512 6568 2528
rect 6584 2512 6616 2528
rect 6648 2512 6664 2528
rect 6712 2512 6728 2528
rect 6776 2512 6792 2528
rect 6824 2512 6840 2528
rect 6920 2512 6936 2528
rect 6968 2512 6984 2528
rect 7032 2512 7048 2528
rect 7112 2512 7128 2528
rect 7144 2512 7176 2528
rect 7240 2512 7256 2528
rect 7304 2512 7320 2528
rect 7352 2512 7368 2528
rect 5416 2492 5432 2508
rect 5544 2492 5560 2508
rect 5672 2492 5688 2508
rect 5992 2492 6008 2508
rect 6120 2492 6136 2508
rect 6328 2492 6344 2508
rect 6456 2492 6472 2508
rect 6968 2492 6984 2508
rect 7016 2492 7032 2508
rect 7256 2492 7272 2508
rect 7320 2492 7336 2508
rect 152 2472 168 2488
rect 1176 2472 1192 2488
rect 1880 2472 1896 2488
rect 4280 2472 4296 2488
rect 4328 2472 4344 2488
rect 4440 2472 4456 2488
rect 4504 2472 4520 2488
rect 4616 2472 4632 2488
rect 4920 2472 4936 2488
rect 5384 2472 5400 2488
rect 2344 2452 2360 2468
rect 4520 2452 4536 2468
rect 5512 2472 5528 2488
rect 5576 2472 5592 2488
rect 5640 2472 5656 2488
rect 6024 2472 6040 2488
rect 6088 2472 6104 2488
rect 6152 2472 6168 2488
rect 6216 2472 6232 2488
rect 6296 2472 6312 2488
rect 6488 2472 6504 2488
rect 6536 2472 6552 2488
rect 6616 2472 6632 2488
rect 6904 2472 6936 2488
rect 6984 2472 7000 2488
rect 7048 2472 7064 2488
rect 7096 2472 7112 2488
rect 7128 2472 7144 2488
rect 7224 2472 7240 2488
rect 7288 2472 7304 2488
rect 5528 2452 5544 2468
rect 5736 2452 5752 2468
rect 6136 2452 6152 2468
rect 6200 2452 6216 2468
rect 7240 2452 7256 2468
rect 7368 2472 7384 2488
rect 136 2432 152 2448
rect 776 2432 792 2448
rect 1544 2432 1560 2448
rect 1752 2432 1768 2448
rect 1896 2432 1912 2448
rect 2744 2432 2760 2448
rect 3368 2432 3384 2448
rect 4904 2432 4920 2448
rect 5592 2432 5608 2448
rect 6072 2432 6088 2448
rect 6264 2432 6280 2448
rect 6472 2432 6488 2448
rect 6520 2432 6536 2448
rect 6600 2432 6616 2448
rect 6888 2432 6904 2448
rect 6968 2432 6984 2448
rect 7032 2432 7048 2448
rect 7160 2432 7176 2448
rect 7384 2432 7400 2448
rect 1117 2402 1153 2418
rect 3165 2402 3201 2418
rect 5213 2402 5249 2418
rect 344 2372 360 2388
rect 1624 2372 1640 2388
rect 3464 2372 3480 2388
rect 4600 2372 4616 2388
rect 4664 2372 4680 2388
rect 4744 2372 4760 2388
rect 4776 2372 4792 2388
rect 4872 2372 4888 2388
rect 5576 2372 5592 2388
rect 6040 2372 6056 2388
rect 6120 2372 6136 2388
rect 7000 2372 7016 2388
rect 7048 2372 7064 2388
rect 7096 2372 7112 2388
rect 7256 2372 7272 2388
rect 7336 2372 7352 2388
rect 7384 2372 7400 2388
rect 1656 2352 1672 2368
rect 6536 2352 6552 2368
rect 8 2332 24 2348
rect 664 2332 680 2348
rect 1000 2332 1016 2348
rect 1416 2332 1432 2348
rect 1672 2332 1688 2348
rect 2232 2332 2248 2348
rect 2584 2332 2600 2348
rect 2872 2332 2888 2348
rect 3704 2332 3720 2348
rect 3976 2332 3992 2348
rect 4024 2332 4040 2348
rect 4312 2332 4328 2348
rect 5000 2332 5016 2348
rect 5208 2332 5224 2348
rect 5496 2332 5528 2348
rect 5560 2332 5576 2348
rect 5800 2332 5816 2348
rect 5832 2332 5848 2348
rect 6104 2332 6120 2348
rect 6152 2332 6168 2348
rect 6184 2332 6200 2348
rect 6232 2332 6248 2348
rect 6392 2332 6408 2348
rect 6632 2332 6648 2348
rect 6728 2332 6744 2348
rect 6776 2332 6792 2348
rect 6840 2332 6856 2348
rect 232 2312 248 2328
rect 136 2290 152 2306
rect 456 2312 472 2328
rect 696 2312 712 2328
rect 280 2292 296 2308
rect 312 2292 328 2308
rect 424 2292 440 2308
rect 536 2292 552 2308
rect 904 2312 920 2328
rect 760 2292 808 2308
rect 856 2292 872 2308
rect 1016 2312 1032 2328
rect 1064 2312 1080 2328
rect 952 2292 968 2308
rect 1176 2312 1192 2328
rect 1512 2312 1528 2328
rect 1112 2292 1128 2308
rect 1208 2292 1224 2308
rect 1304 2292 1320 2308
rect 1432 2292 1448 2308
rect 1640 2312 1656 2328
rect 1880 2312 1896 2328
rect 1976 2312 1992 2328
rect 1576 2292 1592 2308
rect 1624 2292 1640 2308
rect 1816 2290 1832 2306
rect 1912 2292 1928 2308
rect 2296 2312 2312 2328
rect 2024 2292 2040 2308
rect 2120 2292 2136 2308
rect 2280 2292 2296 2308
rect 2344 2312 2360 2328
rect 2616 2312 2632 2328
rect 2456 2292 2472 2308
rect 2920 2312 2936 2328
rect 2664 2292 2680 2308
rect 2760 2292 2776 2308
rect 2968 2292 2984 2308
rect 3064 2312 3080 2328
rect 3368 2312 3384 2328
rect 3256 2292 3272 2308
rect 3480 2312 3496 2328
rect 3752 2312 3768 2328
rect 3800 2312 3816 2328
rect 3416 2292 3432 2308
rect 3592 2292 3608 2308
rect 3640 2292 3656 2308
rect 3848 2292 3864 2308
rect 3896 2292 3912 2308
rect 3944 2312 3960 2328
rect 4104 2292 4120 2308
rect 4232 2292 4248 2308
rect 4280 2312 4296 2328
rect 5480 2312 5496 2328
rect 5592 2312 5608 2328
rect 6136 2312 6152 2328
rect 6200 2312 6216 2328
rect 6264 2312 6280 2328
rect 6424 2312 6440 2328
rect 6632 2312 6648 2328
rect 6760 2312 6776 2328
rect 6808 2312 6824 2328
rect 6872 2312 6888 2328
rect 6920 2332 6936 2348
rect 6984 2332 7000 2348
rect 7032 2332 7048 2348
rect 7064 2332 7080 2348
rect 6952 2312 6968 2328
rect 7080 2312 7096 2328
rect 4440 2292 4456 2308
rect 4568 2292 4584 2308
rect 4632 2292 4648 2308
rect 4696 2292 4728 2308
rect 4776 2292 4792 2308
rect 4952 2292 4984 2308
rect 5112 2292 5128 2308
rect 5256 2292 5272 2308
rect 5352 2292 5384 2308
rect 5432 2292 5448 2308
rect 5496 2292 5512 2308
rect 5576 2292 5592 2308
rect 5608 2292 5624 2308
rect 5640 2292 5656 2308
rect 5720 2292 5736 2308
rect 5848 2292 5864 2308
rect 5880 2292 5896 2308
rect 6008 2292 6024 2308
rect 6072 2292 6088 2308
rect 6120 2292 6136 2308
rect 6168 2292 6184 2308
rect 6248 2292 6264 2308
rect 6360 2292 6376 2308
rect 6408 2292 6424 2308
rect 6488 2292 6520 2308
rect 6568 2292 6584 2308
rect 6648 2292 6664 2308
rect 6712 2292 6728 2308
rect 6792 2292 6808 2308
rect 6856 2292 6872 2308
rect 6904 2292 6920 2308
rect 6968 2292 6984 2308
rect 7048 2292 7064 2308
rect 7096 2292 7128 2308
rect 7144 2292 7160 2308
rect 7208 2292 7224 2308
rect 7304 2292 7320 2308
rect 7352 2292 7368 2308
rect 7416 2292 7432 2308
rect 168 2272 184 2288
rect 200 2272 216 2288
rect 232 2272 248 2288
rect 296 2272 312 2288
rect 456 2272 472 2288
rect 664 2272 680 2288
rect 760 2272 776 2288
rect 840 2272 856 2288
rect 872 2272 888 2288
rect 968 2272 1000 2288
rect 1032 2272 1048 2288
rect 1096 2272 1112 2288
rect 1160 2272 1176 2288
rect 1224 2272 1240 2288
rect 1304 2272 1336 2288
rect 1464 2272 1480 2288
rect 1528 2272 1544 2288
rect 1576 2272 1592 2288
rect 1672 2272 1688 2288
rect 1880 2272 1896 2288
rect 1928 2272 1960 2288
rect 2040 2272 2056 2288
rect 2136 2272 2152 2288
rect 2248 2272 2264 2288
rect 2376 2272 2392 2288
rect 2584 2272 2600 2288
rect 2616 2272 2632 2288
rect 2680 2272 2696 2288
rect 2808 2272 2824 2288
rect 2920 2272 2936 2288
rect 2984 2272 3016 2288
rect 3064 2272 3080 2288
rect 3240 2272 3256 2288
rect 3336 2272 3352 2288
rect 3432 2272 3448 2288
rect 3512 2272 3528 2288
rect 3544 2272 3560 2288
rect 3720 2272 3736 2288
rect 3752 2272 3768 2288
rect 3816 2272 3832 2288
rect 3880 2272 3896 2288
rect 3944 2272 3960 2288
rect 3976 2272 3992 2288
rect 4152 2272 4168 2288
rect 4216 2272 4232 2288
rect 4280 2272 4296 2288
rect 4312 2272 4328 2288
rect 4424 2272 4440 2288
rect 376 2252 392 2268
rect 520 2252 536 2268
rect 712 2252 728 2268
rect 1464 2252 1480 2268
rect 1592 2252 1608 2268
rect 1752 2252 1768 2268
rect 1816 2252 1832 2268
rect 2440 2252 2456 2268
rect 3448 2252 3464 2268
rect 4824 2272 4840 2288
rect 5096 2272 5112 2288
rect 5272 2272 5288 2288
rect 5384 2272 5400 2288
rect 5672 2272 5688 2288
rect 5864 2272 5880 2288
rect 5320 2252 5336 2268
rect 5464 2252 5480 2268
rect 5608 2252 5624 2268
rect 5944 2272 5960 2288
rect 6616 2272 6632 2288
rect 7224 2272 7240 2288
rect 5912 2252 5928 2268
rect 6328 2252 6344 2268
rect 7272 2252 7288 2268
rect 7320 2252 7336 2268
rect 344 2232 360 2248
rect 920 2232 936 2248
rect 1176 2232 1192 2248
rect 1448 2232 1464 2248
rect 1992 2232 2008 2248
rect 2568 2232 2584 2248
rect 3144 2232 3160 2248
rect 3384 2232 3400 2248
rect 3496 2232 3512 2248
rect 3752 2232 3768 2248
rect 4536 2232 4552 2248
rect 4600 2232 4616 2248
rect 4664 2232 4680 2248
rect 4920 2232 4936 2248
rect 5000 2232 5016 2248
rect 5288 2232 5304 2248
rect 5400 2232 5416 2248
rect 5512 2232 5528 2248
rect 5624 2232 5640 2248
rect 6216 2232 6232 2248
rect 6376 2232 6392 2248
rect 6456 2232 6472 2248
rect 6712 2232 6728 2248
rect 6920 2232 6936 2248
rect 2157 2202 2193 2218
rect 4205 2202 4241 2218
rect 6237 2202 6273 2218
rect 408 2172 424 2188
rect 616 2172 632 2188
rect 888 2172 904 2188
rect 1256 2172 1272 2188
rect 1320 2172 1336 2188
rect 1416 2172 1432 2188
rect 1592 2172 1608 2188
rect 1720 2172 1736 2188
rect 1848 2172 1864 2188
rect 2056 2172 2072 2188
rect 2536 2172 2552 2188
rect 3144 2172 3160 2188
rect 3272 2172 3288 2188
rect 3880 2172 3896 2188
rect 4056 2172 4072 2188
rect 5016 2172 5032 2188
rect 5064 2172 5080 2188
rect 5128 2172 5144 2188
rect 5368 2172 5384 2188
rect 5928 2172 5944 2188
rect 6472 2172 6488 2188
rect 6632 2172 6648 2188
rect 7096 2172 7112 2188
rect 7400 2172 7416 2188
rect 1528 2152 1544 2168
rect 2920 2152 2936 2168
rect 3464 2152 3480 2168
rect 3528 2152 3544 2168
rect 3752 2152 3768 2168
rect 3944 2152 3960 2168
rect 4184 2152 4200 2168
rect 4568 2152 4584 2168
rect 5496 2152 5512 2168
rect 5736 2152 5752 2168
rect 6584 2152 6600 2168
rect 7416 2152 7432 2168
rect 168 2132 184 2148
rect 200 2132 216 2148
rect 312 2132 328 2148
rect 424 2132 440 2148
rect 456 2132 472 2148
rect 520 2132 536 2148
rect 632 2132 648 2148
rect 728 2132 744 2148
rect 136 2114 152 2130
rect 1048 2132 1064 2148
rect 1448 2132 1464 2148
rect 1544 2132 1560 2148
rect 1608 2132 1624 2148
rect 1832 2132 1848 2148
rect 2008 2132 2024 2148
rect 2184 2132 2200 2148
rect 2296 2132 2312 2148
rect 2328 2132 2344 2148
rect 2440 2132 2456 2148
rect 2504 2132 2520 2148
rect 2696 2132 2712 2148
rect 2776 2132 2808 2148
rect 3016 2132 3032 2148
rect 3240 2132 3256 2148
rect 3288 2132 3304 2148
rect 3352 2132 3368 2148
rect 3592 2132 3608 2148
rect 3656 2132 3672 2148
rect 3688 2132 3704 2148
rect 3928 2132 3944 2148
rect 4040 2132 4056 2148
rect 4184 2132 4200 2148
rect 4584 2132 4600 2148
rect 4632 2132 4648 2148
rect 5208 2132 5224 2148
rect 5304 2132 5320 2148
rect 5464 2132 5496 2148
rect 5528 2132 5544 2148
rect 5656 2132 5672 2148
rect 5816 2132 5832 2148
rect 6312 2132 6328 2148
rect 6504 2132 6536 2148
rect 7384 2132 7400 2148
rect 216 2112 248 2128
rect 296 2112 312 2128
rect 328 2112 344 2128
rect 504 2112 520 2128
rect 648 2112 680 2128
rect 360 2092 376 2108
rect 392 2092 408 2108
rect 792 2112 808 2128
rect 856 2112 888 2128
rect 1000 2112 1016 2128
rect 1128 2112 1160 2128
rect 1176 2112 1192 2128
rect 1288 2112 1304 2128
rect 1384 2112 1400 2128
rect 1432 2112 1448 2128
rect 1496 2112 1512 2128
rect 1560 2112 1576 2128
rect 1592 2112 1608 2128
rect 1624 2112 1640 2128
rect 1688 2112 1704 2128
rect 1752 2112 1784 2128
rect 1960 2112 1976 2128
rect 2088 2112 2136 2128
rect 2168 2112 2184 2128
rect 2200 2112 2216 2128
rect 696 2092 712 2108
rect 744 2092 760 2108
rect 2456 2112 2472 2128
rect 2648 2112 2664 2128
rect 2744 2112 2792 2128
rect 2840 2112 2856 2128
rect 2952 2112 2968 2128
rect 3032 2112 3048 2128
rect 3304 2112 3320 2128
rect 2296 2092 2312 2108
rect 2728 2092 2744 2108
rect 2824 2092 2840 2108
rect 3160 2092 3176 2108
rect 3272 2092 3288 2108
rect 3512 2112 3528 2128
rect 3608 2112 3624 2128
rect 3352 2092 3368 2108
rect 3752 2114 3768 2130
rect 3992 2112 4008 2128
rect 4088 2112 4104 2128
rect 4136 2112 4152 2128
rect 4280 2112 4296 2128
rect 4328 2112 4344 2128
rect 4392 2112 4408 2128
rect 4456 2112 4472 2128
rect 4520 2112 4536 2128
rect 4600 2112 4616 2128
rect 4696 2114 4712 2130
rect 4760 2112 4776 2128
rect 4920 2112 4936 2128
rect 4952 2112 4968 2128
rect 5032 2112 5048 2128
rect 5096 2112 5112 2128
rect 5272 2112 5288 2128
rect 5384 2112 5400 2128
rect 5448 2112 5464 2128
rect 5560 2112 5576 2128
rect 5592 2112 5608 2128
rect 5640 2112 5656 2128
rect 5688 2112 5720 2128
rect 5800 2114 5816 2130
rect 5976 2112 5992 2128
rect 6024 2112 6040 2128
rect 6104 2112 6120 2128
rect 6152 2112 6168 2128
rect 6216 2112 6232 2128
rect 6360 2112 6376 2128
rect 6488 2112 6504 2128
rect 6552 2112 6568 2128
rect 6600 2112 6616 2128
rect 6680 2112 6696 2128
rect 6744 2112 6760 2128
rect 6808 2112 6824 2128
rect 6888 2112 6904 2128
rect 6952 2112 6968 2128
rect 7016 2112 7032 2128
rect 7064 2112 7080 2128
rect 7144 2112 7160 2128
rect 7240 2112 7256 2128
rect 7304 2114 7320 2130
rect 7368 2112 7384 2128
rect 3656 2092 3672 2108
rect 4024 2092 4040 2108
rect 4104 2092 4120 2108
rect 4124 2092 4140 2108
rect 4344 2092 4360 2108
rect 4408 2092 4424 2108
rect 4472 2092 4488 2108
rect 4536 2092 4552 2108
rect 4632 2092 4648 2108
rect 5592 2092 5608 2108
rect 5992 2092 6024 2108
rect 6120 2092 6152 2108
rect 6200 2092 6216 2108
rect 6664 2092 6680 2108
rect 6792 2092 6808 2108
rect 6904 2092 6920 2108
rect 6968 2092 6984 2108
rect 7032 2092 7064 2108
rect 7112 2092 7128 2108
rect 7144 2092 7160 2108
rect 8 2072 24 2088
rect 264 2072 280 2088
rect 3944 2072 3960 2088
rect 4312 2072 4328 2088
rect 4376 2072 4392 2088
rect 4440 2072 4456 2088
rect 4504 2072 4520 2088
rect 4536 2072 4552 2088
rect 5608 2072 5624 2088
rect 3176 2052 3192 2068
rect 6040 2072 6056 2088
rect 6088 2072 6104 2088
rect 6168 2072 6184 2088
rect 6232 2072 6248 2088
rect 6440 2072 6456 2088
rect 6696 2072 6712 2088
rect 6760 2072 6776 2088
rect 6824 2072 6840 2088
rect 6872 2072 6888 2088
rect 6936 2072 6952 2088
rect 7000 2072 7016 2088
rect 6072 2052 6088 2068
rect 6808 2052 6824 2068
rect 6952 2052 6968 2068
rect 7128 2072 7144 2088
rect 760 2032 776 2048
rect 840 2032 856 2048
rect 1096 2032 1112 2048
rect 1208 2032 1224 2048
rect 1656 2032 1672 2048
rect 1720 2032 1736 2048
rect 2152 2032 2168 2048
rect 2872 2032 2888 2048
rect 4328 2032 4344 2048
rect 4392 2032 4408 2048
rect 4424 2032 4440 2048
rect 4520 2032 4536 2048
rect 4824 2032 4840 2048
rect 5416 2032 5432 2048
rect 5592 2032 5608 2048
rect 5944 2032 5960 2048
rect 6184 2032 6200 2048
rect 6264 2032 6280 2048
rect 6744 2032 6760 2048
rect 6888 2032 6904 2048
rect 7176 2032 7192 2048
rect 1117 2002 1153 2018
rect 3165 2002 3201 2018
rect 5213 2002 5249 2018
rect 792 1972 808 1988
rect 1096 1972 1112 1988
rect 2328 1972 2344 1988
rect 2808 1972 2824 1988
rect 2952 1972 2968 1988
rect 3016 1972 3032 1988
rect 3080 1972 3096 1988
rect 3128 1972 3144 1988
rect 4808 1972 4824 1988
rect 5048 1972 5064 1988
rect 5144 1972 5160 1988
rect 6040 1972 6056 1988
rect 7160 1972 7176 1988
rect 7336 1972 7352 1988
rect 7400 1972 7416 1988
rect 1000 1952 1016 1968
rect 4248 1952 4264 1968
rect 4600 1952 4616 1968
rect 6344 1952 6360 1968
rect 3704 1932 3720 1948
rect 4072 1932 4088 1948
rect 4232 1932 4248 1948
rect 4456 1932 4472 1948
rect 4584 1932 4600 1948
rect 6056 1932 6072 1948
rect 6296 1932 6312 1948
rect 6360 1932 6376 1948
rect 7032 1932 7048 1948
rect 7176 1932 7192 1948
rect 7352 1932 7368 1948
rect 216 1912 232 1928
rect 248 1912 264 1928
rect 324 1912 340 1928
rect 344 1912 360 1928
rect 600 1912 616 1928
rect 840 1912 856 1928
rect 72 1892 104 1908
rect 136 1892 168 1908
rect 296 1892 312 1908
rect 424 1892 440 1908
rect 456 1892 488 1908
rect 552 1892 568 1908
rect 664 1890 680 1906
rect 952 1912 968 1928
rect 888 1892 904 1908
rect 1032 1912 1048 1928
rect 1000 1892 1016 1908
rect 1096 1892 1112 1908
rect 1176 1912 1192 1928
rect 1256 1912 1272 1928
rect 1464 1912 1480 1928
rect 1304 1892 1320 1908
rect 1336 1892 1352 1908
rect 1400 1892 1432 1908
rect 1880 1912 1896 1928
rect 2216 1912 2232 1928
rect 1512 1892 1528 1908
rect 1592 1892 1608 1908
rect 1672 1892 1688 1908
rect 1704 1892 1720 1908
rect 1736 1892 1752 1908
rect 1784 1892 1800 1908
rect 1848 1892 1864 1908
rect 1880 1892 1896 1908
rect 1944 1892 1960 1908
rect 2024 1892 2040 1908
rect 2744 1912 2760 1928
rect 2264 1892 2280 1908
rect 2312 1892 2328 1908
rect 2360 1892 2392 1908
rect 2424 1892 2440 1908
rect 2456 1892 2472 1908
rect 2488 1892 2504 1908
rect 2536 1892 2568 1908
rect 2648 1892 2680 1908
rect 2840 1892 2856 1908
rect 2904 1892 2936 1908
rect 2984 1892 3000 1908
rect 3048 1892 3064 1908
rect 3160 1892 3176 1908
rect 3288 1892 3304 1908
rect 3416 1892 3432 1908
rect 3464 1912 3480 1928
rect 3784 1912 3816 1928
rect 3928 1912 3960 1928
rect 4136 1912 4152 1928
rect 4264 1912 4280 1928
rect 4328 1912 4344 1928
rect 4488 1912 4504 1928
rect 4520 1912 4536 1928
rect 4616 1912 4632 1928
rect 4664 1912 4680 1928
rect 4728 1912 4744 1928
rect 4824 1912 4856 1928
rect 4952 1912 4968 1928
rect 4984 1912 5000 1928
rect 5016 1912 5032 1928
rect 5496 1912 5512 1928
rect 5608 1912 5624 1928
rect 6104 1912 6120 1928
rect 6264 1912 6280 1928
rect 6328 1912 6344 1928
rect 7064 1912 7096 1928
rect 7144 1912 7160 1928
rect 7320 1912 7336 1928
rect 3576 1892 3592 1908
rect 3752 1892 3768 1908
rect 3832 1892 3848 1908
rect 3992 1892 4008 1908
rect 4104 1892 4120 1908
rect 4168 1892 4184 1908
rect 4248 1892 4264 1908
rect 4360 1892 4376 1908
rect 4472 1892 4488 1908
rect 4552 1892 4568 1908
rect 4600 1892 4616 1908
rect 4760 1892 4776 1908
rect 4872 1892 4888 1908
rect 4904 1892 4920 1908
rect 4968 1892 4984 1908
rect 5176 1892 5192 1908
rect 5304 1892 5320 1908
rect 5432 1892 5448 1908
rect 5576 1892 5592 1908
rect 5752 1890 5768 1906
rect 5848 1892 5880 1908
rect 5912 1892 5944 1908
rect 5992 1892 6008 1908
rect 6072 1892 6088 1908
rect 6200 1892 6216 1908
rect 6280 1892 6296 1908
rect 6344 1892 6360 1908
rect 6440 1892 6456 1908
rect 6568 1892 6584 1908
rect 6632 1892 6664 1908
rect 6712 1892 6728 1908
rect 6776 1892 6792 1908
rect 6808 1892 6824 1908
rect 6872 1890 6888 1906
rect 7048 1892 7064 1908
rect 7096 1892 7112 1908
rect 7160 1892 7176 1908
rect 7208 1892 7224 1908
rect 7304 1892 7320 1908
rect 7336 1892 7352 1908
rect 7384 1892 7400 1908
rect 168 1872 184 1888
rect 216 1872 232 1888
rect 552 1872 568 1888
rect 600 1872 616 1888
rect 632 1872 648 1888
rect 808 1872 824 1888
rect 872 1872 888 1888
rect 904 1872 936 1888
rect 1016 1872 1032 1888
rect 1064 1872 1096 1888
rect 1208 1872 1224 1888
rect 1320 1872 1336 1888
rect 1432 1872 1448 1888
rect 1528 1872 1544 1888
rect 1832 1872 1848 1888
rect 1896 1872 1912 1888
rect 2008 1872 2024 1888
rect 2152 1872 2168 1888
rect 2280 1872 2296 1888
rect 2440 1872 2456 1888
rect 2472 1872 2488 1888
rect 2504 1872 2520 1888
rect 120 1852 136 1868
rect 264 1852 280 1868
rect 1384 1852 1400 1868
rect 1704 1852 1720 1868
rect 1768 1852 1800 1868
rect 1816 1852 1832 1868
rect 1912 1852 1928 1868
rect 2232 1852 2248 1868
rect 2392 1852 2408 1868
rect 2632 1872 2648 1888
rect 2776 1872 2792 1888
rect 2856 1872 2872 1888
rect 3032 1872 3048 1888
rect 3128 1872 3144 1888
rect 3224 1872 3240 1888
rect 3320 1872 3336 1888
rect 3400 1872 3416 1888
rect 3464 1872 3480 1888
rect 3496 1872 3512 1888
rect 3528 1872 3544 1888
rect 3784 1872 3800 1888
rect 3976 1872 3992 1888
rect 4376 1872 4408 1888
rect 4632 1872 4648 1888
rect 4776 1872 4808 1888
rect 4888 1872 4920 1888
rect 4968 1872 4984 1888
rect 5096 1872 5112 1888
rect 5352 1872 5384 1888
rect 5448 1872 5464 1888
rect 5544 1872 5576 1888
rect 5592 1872 5608 1888
rect 5816 1872 5832 1888
rect 5944 1872 5960 1888
rect 6184 1872 6200 1888
rect 6424 1872 6440 1888
rect 6616 1872 6632 1888
rect 2568 1852 2584 1868
rect 3704 1852 3720 1868
rect 3880 1852 3896 1868
rect 4024 1852 4040 1868
rect 4280 1852 4296 1868
rect 4680 1852 4696 1868
rect 5112 1852 5128 1868
rect 5176 1852 5208 1868
rect 5288 1852 5304 1868
rect 5464 1852 5480 1868
rect 5816 1852 5832 1868
rect 6024 1852 6040 1868
rect 6200 1852 6216 1868
rect 6440 1852 6456 1868
rect 6584 1852 6600 1868
rect 6744 1852 6760 1868
rect 6792 1872 6808 1888
rect 6840 1872 6856 1888
rect 7224 1872 7240 1888
rect 7272 1852 7288 1868
rect 7416 1852 7432 1868
rect 24 1832 40 1848
rect 200 1832 216 1848
rect 248 1832 264 1848
rect 536 1832 552 1848
rect 1048 1832 1064 1848
rect 1272 1832 1288 1848
rect 1480 1832 1496 1848
rect 1560 1832 1576 1848
rect 1688 1832 1704 1848
rect 1928 1832 1944 1848
rect 2136 1832 2168 1848
rect 2408 1832 2424 1848
rect 2728 1832 2744 1848
rect 2760 1832 2776 1848
rect 3080 1832 3096 1848
rect 3384 1832 3400 1848
rect 3800 1832 3816 1848
rect 3912 1832 3928 1848
rect 3960 1832 3976 1848
rect 4072 1832 4088 1848
rect 4296 1832 4312 1848
rect 4424 1832 4440 1848
rect 4664 1832 4680 1848
rect 4696 1832 4712 1848
rect 4840 1832 4856 1848
rect 4952 1832 4968 1848
rect 5496 1832 5512 1848
rect 5624 1832 5640 1848
rect 5960 1832 5976 1848
rect 6104 1832 6120 1848
rect 6296 1832 6312 1848
rect 6424 1832 6440 1848
rect 6536 1832 6552 1848
rect 6600 1832 6616 1848
rect 6680 1832 6696 1848
rect 7000 1832 7016 1848
rect 7096 1832 7112 1848
rect 7240 1832 7256 1848
rect 2157 1802 2193 1818
rect 4205 1802 4241 1818
rect 6237 1802 6273 1818
rect 8 1772 24 1788
rect 344 1772 360 1788
rect 376 1772 392 1788
rect 696 1772 712 1788
rect 920 1772 936 1788
rect 1176 1772 1192 1788
rect 1400 1772 1416 1788
rect 1704 1772 1720 1788
rect 2120 1772 2136 1788
rect 2456 1772 2472 1788
rect 2792 1772 2808 1788
rect 3176 1772 3192 1788
rect 3880 1772 3896 1788
rect 3976 1772 3992 1788
rect 4040 1772 4056 1788
rect 4104 1772 4120 1788
rect 4168 1772 4184 1788
rect 4936 1772 4952 1788
rect 4984 1772 5000 1788
rect 5192 1772 5208 1788
rect 5272 1772 5288 1788
rect 5384 1772 5400 1788
rect 5464 1772 5480 1788
rect 5528 1772 5544 1788
rect 5576 1772 5592 1788
rect 6040 1772 6056 1788
rect 6184 1772 6200 1788
rect 6344 1772 6360 1788
rect 6552 1772 6568 1788
rect 6872 1772 6888 1788
rect 7064 1772 7080 1788
rect 7288 1772 7304 1788
rect 2472 1752 2504 1768
rect 3032 1752 3048 1768
rect 3256 1752 3272 1768
rect 3496 1752 3512 1768
rect 4312 1752 4328 1768
rect 4552 1752 4568 1768
rect 4808 1752 4824 1768
rect 5352 1752 5368 1768
rect 5560 1752 5576 1768
rect 6568 1752 6584 1768
rect 6904 1752 6920 1768
rect 7048 1752 7064 1768
rect 7304 1752 7320 1768
rect 7416 1752 7432 1768
rect 168 1732 184 1748
rect 248 1732 264 1748
rect 312 1732 328 1748
rect 360 1732 376 1748
rect 472 1732 488 1748
rect 616 1732 632 1748
rect 744 1732 776 1748
rect 856 1732 888 1748
rect 936 1732 952 1748
rect 984 1732 1000 1748
rect 1016 1732 1032 1748
rect 1288 1732 1304 1748
rect 1448 1732 1464 1748
rect 1512 1732 1528 1748
rect 1544 1732 1560 1748
rect 1720 1732 1736 1748
rect 1944 1732 1960 1748
rect 1976 1732 1992 1748
rect 2008 1732 2024 1748
rect 2072 1732 2088 1748
rect 2296 1732 2312 1748
rect 2504 1732 2520 1748
rect 2536 1732 2552 1748
rect 2616 1732 2632 1748
rect 2680 1732 2696 1748
rect 2712 1732 2744 1748
rect 2776 1732 2792 1748
rect 3176 1732 3192 1748
rect 3320 1732 3336 1748
rect 3352 1732 3368 1748
rect 3416 1732 3432 1748
rect 120 1712 136 1728
rect 216 1712 248 1728
rect 280 1712 312 1728
rect 488 1712 504 1728
rect 600 1712 616 1728
rect 200 1692 216 1708
rect 264 1692 280 1708
rect 328 1692 344 1708
rect 568 1692 584 1708
rect 680 1692 696 1708
rect 728 1712 744 1728
rect 824 1712 840 1728
rect 856 1712 872 1728
rect 952 1712 968 1728
rect 1064 1712 1080 1728
rect 1288 1712 1304 1728
rect 1336 1712 1352 1728
rect 824 1692 840 1708
rect 856 1692 872 1708
rect 920 1692 936 1708
rect 984 1692 1000 1708
rect 1448 1692 1464 1708
rect 1496 1712 1512 1728
rect 1576 1714 1592 1730
rect 1768 1712 1784 1728
rect 1896 1712 1912 1728
rect 1992 1712 2008 1728
rect 2088 1712 2104 1728
rect 2152 1712 2184 1728
rect 2264 1712 2280 1728
rect 2344 1712 2360 1728
rect 2040 1692 2056 1708
rect 2536 1692 2552 1708
rect 2584 1712 2616 1728
rect 2744 1712 2760 1728
rect 2904 1712 2920 1728
rect 3048 1712 3064 1728
rect 2680 1692 2696 1708
rect 2776 1692 2792 1708
rect 3240 1692 3256 1708
rect 3304 1712 3320 1728
rect 3336 1712 3352 1728
rect 3432 1712 3448 1728
rect 3528 1712 3544 1728
rect 3576 1732 3592 1748
rect 3640 1732 3656 1748
rect 3720 1732 3736 1748
rect 4024 1732 4040 1748
rect 4136 1732 4152 1748
rect 4344 1732 4360 1748
rect 4376 1732 4392 1748
rect 4504 1732 4520 1748
rect 4600 1732 4616 1748
rect 4920 1732 4936 1748
rect 4968 1732 4984 1748
rect 5080 1732 5096 1748
rect 5176 1732 5192 1748
rect 5224 1732 5240 1748
rect 5304 1732 5320 1748
rect 5368 1732 5384 1748
rect 5432 1732 5448 1748
rect 5480 1732 5496 1748
rect 5576 1732 5592 1748
rect 5656 1732 5672 1748
rect 5704 1732 5720 1748
rect 6168 1732 6184 1748
rect 6232 1732 6248 1748
rect 6392 1732 6424 1748
rect 6440 1732 6456 1748
rect 6472 1732 6488 1748
rect 6504 1732 6520 1748
rect 6584 1732 6600 1748
rect 6808 1732 6824 1748
rect 6984 1732 7000 1748
rect 7272 1732 7288 1748
rect 7384 1732 7400 1748
rect 3592 1712 3608 1728
rect 3656 1712 3688 1728
rect 3752 1714 3768 1730
rect 3944 1712 3960 1728
rect 4008 1712 4024 1728
rect 4104 1712 4120 1728
rect 4232 1712 4248 1728
rect 4312 1712 4328 1728
rect 4424 1712 4440 1728
rect 4488 1712 4520 1728
rect 4568 1712 4584 1728
rect 4632 1712 4648 1728
rect 4696 1712 4712 1728
rect 4760 1712 4776 1728
rect 4840 1712 4856 1728
rect 4904 1712 4920 1728
rect 5032 1712 5048 1728
rect 5096 1712 5112 1728
rect 3384 1692 3400 1708
rect 3464 1692 3480 1708
rect 3528 1692 3544 1708
rect 3560 1692 3576 1708
rect 3624 1692 3640 1708
rect 3688 1692 3704 1708
rect 4056 1692 4072 1708
rect 4120 1692 4136 1708
rect 4168 1692 4184 1708
rect 4216 1692 4232 1708
rect 4328 1692 4344 1708
rect 4376 1692 4392 1708
rect 4440 1692 4456 1708
rect 4488 1692 4504 1708
rect 4568 1692 4584 1708
rect 4616 1692 4632 1708
rect 4680 1692 4696 1708
rect 4744 1692 4760 1708
rect 4968 1692 4984 1708
rect 5000 1692 5032 1708
rect 5304 1712 5320 1728
rect 5416 1712 5432 1728
rect 5496 1712 5512 1728
rect 5592 1712 5608 1728
rect 5672 1712 5688 1728
rect 5752 1712 5768 1728
rect 5816 1712 5832 1728
rect 5960 1712 5992 1728
rect 6088 1712 6104 1728
rect 6120 1712 6136 1728
rect 6216 1712 6232 1728
rect 6296 1712 6312 1728
rect 6376 1712 6392 1728
rect 6424 1712 6440 1728
rect 6488 1712 6504 1728
rect 6520 1712 6536 1728
rect 6632 1712 6648 1728
rect 6760 1712 6776 1728
rect 6840 1712 6856 1728
rect 6936 1712 6952 1728
rect 6968 1712 6984 1728
rect 7000 1712 7032 1728
rect 7128 1712 7144 1728
rect 7176 1712 7192 1728
rect 7256 1712 7272 1728
rect 7352 1712 7368 1728
rect 7384 1712 7400 1728
rect 5144 1692 5160 1708
rect 5192 1692 5208 1708
rect 5272 1692 5288 1708
rect 5464 1692 5480 1708
rect 5528 1692 5544 1708
rect 5720 1692 5752 1708
rect 5800 1692 5816 1708
rect 6104 1692 6120 1708
rect 6184 1692 6200 1708
rect 6280 1692 6296 1708
rect 6456 1692 6472 1708
rect 6520 1692 6536 1708
rect 7368 1692 7384 1708
rect 1784 1672 1800 1688
rect 3592 1672 3608 1688
rect 4088 1672 4104 1688
rect 4136 1672 4152 1688
rect 4248 1672 4264 1688
rect 4312 1672 4328 1688
rect 4408 1672 4424 1688
rect 4648 1672 4664 1688
rect 4712 1672 4728 1688
rect 4776 1672 4792 1688
rect 4840 1672 4856 1688
rect 5048 1672 5064 1688
rect 5768 1672 5784 1688
rect 5832 1672 5848 1688
rect 6072 1672 6088 1688
rect 6264 1672 6280 1688
rect 6648 1672 6664 1688
rect 7336 1672 7352 1688
rect 5752 1652 5768 1668
rect 5816 1652 5832 1668
rect 6088 1652 6104 1668
rect 600 1632 616 1648
rect 2232 1632 2248 1648
rect 3912 1632 3928 1648
rect 4264 1632 4280 1648
rect 4584 1632 4600 1648
rect 4664 1632 4680 1648
rect 4728 1632 4744 1648
rect 4792 1632 4808 1648
rect 4872 1632 4888 1648
rect 5064 1632 5080 1648
rect 5096 1632 5112 1648
rect 5384 1632 5400 1648
rect 5448 1632 5464 1648
rect 6872 1632 6888 1648
rect 7032 1632 7048 1648
rect 7352 1632 7368 1648
rect 1117 1602 1153 1618
rect 3165 1602 3201 1618
rect 5213 1602 5249 1618
rect 312 1572 328 1588
rect 1496 1572 1512 1588
rect 2472 1572 2488 1588
rect 4152 1572 4168 1588
rect 4328 1572 4344 1588
rect 4984 1572 5000 1588
rect 6520 1572 6536 1588
rect 6600 1572 6616 1588
rect 7144 1572 7160 1588
rect 2536 1552 2552 1568
rect 4440 1552 4456 1568
rect 8 1532 24 1548
rect 344 1532 360 1548
rect 1928 1532 1944 1548
rect 2232 1532 2248 1548
rect 4136 1532 4152 1548
rect 4248 1532 4264 1548
rect 4312 1532 4328 1548
rect 4424 1532 4440 1548
rect 4648 1532 4664 1548
rect 5288 1532 5304 1548
rect 5800 1532 5816 1548
rect 5992 1532 6008 1548
rect 6104 1552 6120 1568
rect 6072 1532 6088 1548
rect 6536 1532 6552 1548
rect 6616 1532 6632 1548
rect 6856 1532 6872 1548
rect 232 1512 248 1528
rect 120 1492 136 1508
rect 568 1512 584 1528
rect 920 1512 936 1528
rect 280 1492 296 1508
rect 424 1492 440 1508
rect 552 1492 568 1508
rect 616 1492 632 1508
rect 680 1490 696 1506
rect 744 1492 760 1508
rect 824 1492 840 1508
rect 888 1492 904 1508
rect 952 1492 968 1508
rect 1032 1492 1048 1508
rect 1080 1512 1096 1528
rect 1160 1512 1176 1528
rect 1560 1512 1576 1528
rect 1256 1490 1272 1506
rect 1320 1492 1336 1508
rect 1400 1492 1416 1508
rect 1464 1492 1480 1508
rect 1608 1512 1624 1528
rect 2152 1512 2168 1528
rect 1624 1492 1640 1508
rect 1752 1492 1768 1508
rect 1832 1492 1864 1508
rect 1992 1492 2008 1508
rect 2056 1490 2072 1506
rect 2232 1492 2248 1508
rect 2264 1492 2280 1508
rect 2344 1492 2360 1508
rect 2392 1512 2408 1528
rect 2776 1512 2792 1528
rect 2440 1492 2456 1508
rect 2488 1492 2504 1508
rect 2696 1490 2712 1506
rect 2776 1492 2792 1508
rect 2824 1512 2840 1528
rect 2952 1512 3000 1528
rect 3272 1512 3288 1528
rect 2904 1492 2920 1508
rect 2952 1492 2968 1508
rect 3144 1490 3160 1506
rect 3308 1512 3324 1528
rect 3320 1492 3336 1508
rect 3368 1492 3384 1508
rect 3416 1512 3432 1528
rect 3848 1512 3864 1528
rect 3868 1512 3884 1528
rect 3912 1512 3944 1528
rect 4040 1512 4056 1528
rect 4168 1512 4200 1528
rect 4232 1512 4248 1528
rect 4280 1512 4296 1528
rect 4472 1512 4488 1528
rect 4504 1512 4520 1528
rect 4680 1512 4696 1528
rect 4760 1512 4776 1528
rect 5128 1512 5144 1528
rect 5512 1512 5528 1528
rect 3512 1490 3528 1506
rect 3720 1492 3736 1508
rect 3912 1492 3928 1508
rect 4008 1492 4024 1508
rect 4104 1492 4120 1508
rect 4136 1492 4168 1508
rect 4296 1492 4312 1508
rect 4392 1492 4408 1508
rect 4440 1492 4456 1508
rect 4552 1492 4568 1508
rect 4616 1492 4632 1508
rect 4664 1492 4680 1508
rect 4696 1492 4712 1508
rect 4728 1492 4744 1508
rect 4856 1492 4872 1508
rect 4904 1492 4920 1508
rect 4952 1492 4968 1508
rect 5048 1492 5080 1508
rect 5112 1492 5128 1508
rect 5160 1492 5176 1508
rect 5192 1492 5208 1508
rect 5352 1492 5368 1508
rect 5416 1490 5432 1506
rect 5548 1512 5564 1528
rect 5832 1512 5848 1528
rect 6040 1512 6056 1528
rect 6568 1512 6584 1528
rect 5560 1492 5576 1508
rect 5608 1492 5624 1508
rect 5736 1492 5752 1508
rect 5816 1492 5832 1508
rect 5896 1492 5912 1508
rect 5992 1492 6008 1508
rect 6056 1492 6072 1508
rect 6168 1492 6184 1508
rect 6216 1492 6232 1508
rect 6392 1492 6408 1508
rect 6440 1492 6456 1508
rect 6552 1492 6568 1508
rect 6600 1492 6616 1508
rect 6648 1492 6664 1508
rect 6712 1492 6728 1508
rect 6776 1492 6792 1508
rect 6808 1492 6824 1508
rect 6904 1492 6920 1508
rect 7016 1492 7032 1508
rect 7096 1492 7112 1508
rect 7128 1492 7144 1508
rect 7208 1492 7240 1508
rect 7336 1492 7352 1508
rect 168 1472 184 1488
rect 200 1472 216 1488
rect 232 1472 248 1488
rect 296 1472 312 1488
rect 472 1472 488 1488
rect 568 1472 584 1488
rect 616 1472 632 1488
rect 1000 1472 1016 1488
rect 1080 1472 1096 1488
rect 1144 1472 1160 1488
rect 1192 1472 1208 1488
rect 1224 1472 1240 1488
rect 1528 1472 1544 1488
rect 1624 1472 1640 1488
rect 1752 1472 1768 1488
rect 1896 1472 1912 1488
rect 2120 1472 2136 1488
rect 2248 1472 2264 1488
rect 2296 1472 2312 1488
rect 2328 1472 2344 1488
rect 2424 1472 2440 1488
rect 2760 1472 2776 1488
rect 2856 1472 2872 1488
rect 2536 1452 2552 1468
rect 2696 1452 2712 1468
rect 3000 1472 3016 1488
rect 3128 1472 3144 1488
rect 3208 1472 3224 1488
rect 3336 1472 3368 1488
rect 3416 1472 3432 1488
rect 3448 1472 3464 1488
rect 3480 1472 3496 1488
rect 3576 1472 3592 1488
rect 3672 1472 3688 1488
rect 3896 1472 3912 1488
rect 3944 1472 3960 1488
rect 4344 1472 4360 1488
rect 4472 1472 4488 1488
rect 4504 1472 4520 1488
rect 4712 1472 4728 1488
rect 4744 1472 4760 1488
rect 4792 1472 4808 1488
rect 5000 1472 5016 1488
rect 5176 1472 5192 1488
rect 5272 1472 5288 1488
rect 5480 1472 5496 1488
rect 5576 1472 5592 1488
rect 5624 1472 5640 1488
rect 5720 1472 5736 1488
rect 5752 1472 5768 1488
rect 5880 1472 5896 1488
rect 5960 1472 5976 1488
rect 6312 1472 6328 1488
rect 4072 1452 4088 1468
rect 4264 1452 4280 1468
rect 4584 1452 4600 1468
rect 4968 1452 4984 1468
rect 5096 1452 5112 1468
rect 5640 1452 5656 1468
rect 5864 1452 5880 1468
rect 6744 1452 6760 1468
rect 6792 1472 6808 1488
rect 6984 1472 7000 1488
rect 7080 1472 7096 1488
rect 7112 1472 7128 1488
rect 7304 1472 7320 1488
rect 7352 1472 7368 1488
rect 7080 1452 7096 1468
rect 7384 1452 7400 1468
rect 520 1432 536 1448
rect 808 1432 824 1448
rect 856 1432 872 1448
rect 984 1432 1000 1448
rect 1128 1432 1144 1448
rect 1384 1432 1400 1448
rect 1432 1432 1448 1448
rect 1640 1432 1656 1448
rect 2376 1432 2392 1448
rect 2568 1432 2584 1448
rect 3016 1432 3032 1448
rect 3640 1432 3656 1448
rect 3832 1432 3848 1448
rect 4040 1432 4056 1448
rect 4760 1432 4776 1448
rect 4824 1432 4840 1448
rect 4872 1432 4888 1448
rect 4920 1432 4936 1448
rect 5624 1432 5640 1448
rect 5880 1432 5896 1448
rect 6328 1432 6344 1448
rect 6680 1432 6696 1448
rect 6824 1432 6840 1448
rect 7368 1432 7384 1448
rect 2157 1402 2193 1418
rect 4205 1402 4241 1418
rect 6237 1402 6273 1418
rect 184 1372 200 1388
rect 536 1372 552 1388
rect 936 1372 952 1388
rect 1336 1372 1352 1388
rect 1592 1372 1608 1388
rect 1800 1372 1816 1388
rect 2568 1372 2584 1388
rect 3512 1372 3528 1388
rect 3640 1372 3656 1388
rect 4728 1372 4744 1388
rect 4920 1372 4936 1388
rect 5128 1372 5144 1388
rect 5368 1372 5384 1388
rect 5448 1372 5464 1388
rect 5544 1372 5560 1388
rect 5688 1372 5704 1388
rect 5912 1372 5928 1388
rect 6184 1372 6200 1388
rect 6936 1372 6952 1388
rect 7224 1372 7240 1388
rect 1400 1352 1416 1368
rect 1560 1352 1576 1368
rect 1816 1352 1832 1368
rect 1944 1352 1960 1368
rect 2008 1352 2040 1368
rect 2280 1352 2296 1368
rect 2424 1352 2440 1368
rect 2504 1352 2520 1368
rect 2696 1352 2712 1368
rect 3256 1352 3272 1368
rect 3592 1352 3608 1368
rect 4120 1352 4136 1368
rect 4152 1352 4168 1368
rect 5416 1352 5432 1368
rect 200 1332 216 1348
rect 296 1332 312 1348
rect 376 1332 392 1348
rect 472 1332 504 1348
rect 584 1332 616 1348
rect 824 1332 840 1348
rect 952 1332 968 1348
rect 1048 1332 1080 1348
rect 1224 1332 1240 1348
rect 1448 1332 1464 1348
rect 1544 1332 1560 1348
rect 1576 1332 1592 1348
rect 1752 1332 1768 1348
rect 1832 1332 1848 1348
rect 1896 1332 1912 1348
rect 1960 1332 1976 1348
rect 1992 1332 2008 1348
rect 2248 1332 2264 1348
rect 2520 1332 2536 1348
rect 2888 1332 2904 1348
rect 2952 1332 2968 1348
rect 2984 1332 3000 1348
rect 3048 1332 3064 1348
rect 3096 1332 3128 1348
rect 3208 1332 3224 1348
rect 3304 1332 3320 1348
rect 3336 1332 3352 1348
rect 3608 1332 3624 1348
rect 4136 1332 4152 1348
rect 4280 1332 4296 1348
rect 4600 1332 4632 1348
rect 4680 1332 4696 1348
rect 4888 1332 4904 1348
rect 5080 1332 5096 1348
rect 5112 1332 5128 1348
rect 5208 1332 5224 1348
rect 5976 1352 5992 1368
rect 6152 1352 6168 1368
rect 5464 1332 5480 1348
rect 5496 1332 5512 1348
rect 5736 1332 5752 1348
rect 5896 1332 5912 1348
rect 6920 1352 6936 1368
rect 6200 1332 6216 1348
rect 6856 1332 6872 1348
rect 6888 1332 6920 1348
rect 72 1312 88 1328
rect 120 1312 136 1328
rect 200 1312 216 1328
rect 216 1292 232 1308
rect 376 1312 392 1328
rect 264 1292 280 1308
rect 408 1292 424 1308
rect 440 1312 472 1328
rect 504 1312 520 1328
rect 648 1312 664 1328
rect 680 1312 696 1328
rect 728 1312 760 1328
rect 840 1312 856 1328
rect 952 1312 968 1328
rect 552 1292 568 1308
rect 968 1292 984 1308
rect 1080 1312 1096 1328
rect 1144 1312 1160 1328
rect 1208 1314 1224 1330
rect 1368 1312 1384 1328
rect 1416 1312 1448 1328
rect 1464 1312 1480 1328
rect 1016 1292 1032 1308
rect 1128 1292 1144 1308
rect 1476 1292 1492 1308
rect 1704 1312 1720 1328
rect 1784 1312 1800 1328
rect 1848 1312 1864 1328
rect 1880 1312 1896 1328
rect 1912 1312 1928 1328
rect 1960 1312 1976 1328
rect 2056 1312 2072 1328
rect 2136 1312 2152 1328
rect 2296 1312 2312 1328
rect 2472 1312 2488 1328
rect 2696 1314 2712 1330
rect 2808 1312 2840 1328
rect 2904 1312 2920 1328
rect 2952 1312 2968 1328
rect 1512 1292 1528 1308
rect 1880 1292 1896 1308
rect 2152 1292 2168 1308
rect 2856 1292 2872 1308
rect 2936 1292 2952 1308
rect 2984 1292 3000 1308
rect 3032 1312 3048 1328
rect 3064 1312 3080 1328
rect 3224 1312 3240 1328
rect 3160 1292 3176 1308
rect 3368 1314 3384 1330
rect 3432 1312 3448 1328
rect 3560 1312 3576 1328
rect 3640 1312 3656 1328
rect 3752 1312 3768 1328
rect 3816 1312 3832 1328
rect 3880 1312 3896 1328
rect 3944 1312 3960 1328
rect 4008 1312 4024 1328
rect 4072 1312 4088 1328
rect 4168 1312 4184 1328
rect 4264 1312 4280 1328
rect 4312 1312 4328 1328
rect 4392 1312 4408 1328
rect 4456 1312 4472 1328
rect 4504 1312 4520 1328
rect 4552 1312 4568 1328
rect 4584 1312 4600 1328
rect 4632 1312 4648 1328
rect 3272 1292 3288 1308
rect 3512 1292 3528 1308
rect 3768 1292 3784 1308
rect 3832 1292 3848 1308
rect 3896 1292 3912 1308
rect 3960 1292 3976 1308
rect 4024 1292 4040 1308
rect 4088 1292 4120 1308
rect 4200 1292 4216 1308
rect 4296 1292 4312 1308
rect 4408 1292 4424 1308
rect 4472 1292 4504 1308
rect 4552 1292 4568 1308
rect 4840 1312 4856 1328
rect 5048 1314 5064 1330
rect 5256 1312 5272 1328
rect 5384 1312 5400 1328
rect 5480 1312 5496 1328
rect 5512 1312 5528 1328
rect 5592 1312 5608 1328
rect 5640 1312 5656 1328
rect 5736 1312 5752 1328
rect 5768 1312 5784 1328
rect 5832 1312 5848 1328
rect 5880 1312 5896 1328
rect 5944 1312 5960 1328
rect 5992 1312 6008 1328
rect 6088 1312 6104 1328
rect 6120 1312 6136 1328
rect 6216 1312 6232 1328
rect 6280 1312 6296 1328
rect 6360 1312 6376 1328
rect 6424 1312 6440 1328
rect 6488 1312 6504 1328
rect 6552 1312 6568 1328
rect 6616 1312 6632 1328
rect 6680 1312 6696 1328
rect 6744 1312 6760 1328
rect 6792 1312 6808 1328
rect 6872 1312 6888 1328
rect 6952 1312 6968 1328
rect 7064 1312 7080 1328
rect 7128 1312 7144 1328
rect 7192 1312 7208 1328
rect 7304 1312 7320 1328
rect 7352 1314 7368 1330
rect 4680 1292 4696 1308
rect 5176 1292 5192 1308
rect 5608 1292 5624 1308
rect 5752 1292 5768 1308
rect 5816 1292 5832 1308
rect 6104 1292 6120 1308
rect 6264 1292 6280 1308
rect 6376 1292 6392 1308
rect 6440 1292 6456 1308
rect 6504 1292 6520 1308
rect 6568 1292 6584 1308
rect 6632 1292 6648 1308
rect 6696 1292 6712 1308
rect 6760 1292 6792 1308
rect 6840 1292 6856 1308
rect 7080 1292 7096 1308
rect 7144 1292 7160 1308
rect 7208 1292 7224 1308
rect 1976 1272 1992 1288
rect 3144 1272 3160 1288
rect 3496 1272 3512 1288
rect 3640 1272 3656 1288
rect 3736 1272 3752 1288
rect 3768 1272 3784 1288
rect 3800 1272 3816 1288
rect 3864 1272 3880 1288
rect 3928 1272 3944 1288
rect 3992 1272 4008 1288
rect 4056 1272 4072 1288
rect 4328 1272 4344 1288
rect 4392 1272 4408 1288
rect 4440 1272 4456 1288
rect 4520 1272 4536 1288
rect 5576 1272 5592 1288
rect 5656 1272 5672 1288
rect 5784 1272 5800 1288
rect 5848 1272 5864 1288
rect 6072 1272 6088 1288
rect 6296 1272 6312 1288
rect 6344 1272 6360 1288
rect 6408 1272 6424 1288
rect 6472 1272 6488 1288
rect 6536 1272 6552 1288
rect 6600 1272 6616 1288
rect 6664 1272 6680 1288
rect 6728 1272 6744 1288
rect 6808 1272 6824 1288
rect 7048 1272 7064 1288
rect 7144 1272 7160 1288
rect 7176 1272 7192 1288
rect 4008 1252 4024 1268
rect 4072 1252 4088 1268
rect 6680 1252 6696 1268
rect 328 1232 344 1248
rect 712 1232 728 1248
rect 2200 1232 2216 1248
rect 3688 1232 3704 1248
rect 3720 1232 3736 1248
rect 3816 1232 3832 1248
rect 3880 1232 3896 1248
rect 3944 1232 3960 1248
rect 4344 1232 4376 1248
rect 4456 1232 4472 1248
rect 4536 1232 4552 1248
rect 5768 1232 5784 1248
rect 5832 1232 5848 1248
rect 6024 1232 6040 1248
rect 6088 1232 6104 1248
rect 6312 1232 6328 1248
rect 6360 1232 6376 1248
rect 6424 1232 6440 1248
rect 6488 1232 6504 1248
rect 6552 1232 6568 1248
rect 6616 1232 6632 1248
rect 6744 1232 6760 1248
rect 6792 1232 6808 1248
rect 7064 1232 7080 1248
rect 7128 1232 7144 1248
rect 7192 1232 7208 1248
rect 1117 1202 1153 1218
rect 3165 1202 3201 1218
rect 5213 1202 5249 1218
rect 312 1172 328 1188
rect 616 1172 632 1188
rect 5400 1172 5416 1188
rect 5544 1172 5560 1188
rect 6936 1172 6952 1188
rect 7336 1172 7352 1188
rect 7400 1172 7416 1188
rect 1576 1152 1592 1168
rect 4376 1152 4392 1168
rect 184 1132 200 1148
rect 552 1132 568 1148
rect 1176 1132 1192 1148
rect 2200 1132 2216 1148
rect 2264 1132 2280 1148
rect 2840 1132 2856 1148
rect 3192 1132 3208 1148
rect 3704 1132 3720 1148
rect 3768 1132 3784 1148
rect 3912 1132 3928 1148
rect 4104 1132 4120 1148
rect 4232 1132 4248 1148
rect 4312 1132 4328 1148
rect 4360 1132 4376 1148
rect 4552 1132 4568 1148
rect 4664 1132 4680 1148
rect 4792 1132 4808 1148
rect 6376 1152 6392 1168
rect 7192 1152 7208 1168
rect 4984 1132 5000 1148
rect 5864 1132 5880 1148
rect 216 1112 232 1128
rect 72 1092 88 1108
rect 120 1092 136 1108
rect 200 1092 216 1108
rect 264 1112 280 1128
rect 728 1112 744 1128
rect 888 1112 904 1128
rect 952 1112 968 1128
rect 1096 1112 1112 1128
rect 440 1090 456 1106
rect 504 1092 536 1108
rect 568 1092 584 1108
rect 648 1092 664 1108
rect 680 1092 696 1108
rect 808 1092 824 1108
rect 920 1092 936 1108
rect 1032 1092 1048 1108
rect 1208 1112 1224 1128
rect 1304 1112 1320 1128
rect 1336 1112 1352 1128
rect 1384 1112 1400 1128
rect 1432 1112 1464 1128
rect 1528 1112 1560 1128
rect 1176 1092 1192 1108
rect 1576 1092 1592 1108
rect 1624 1092 1640 1108
rect 1672 1112 1688 1128
rect 2008 1112 2024 1128
rect 1784 1092 1800 1108
rect 1832 1092 1848 1108
rect 1960 1092 1976 1108
rect 2120 1112 2136 1128
rect 2056 1092 2072 1108
rect 2296 1112 2312 1128
rect 2872 1112 2888 1128
rect 2200 1092 2216 1108
rect 2264 1092 2280 1108
rect 2296 1092 2312 1108
rect 2328 1092 2344 1108
rect 2360 1092 2376 1108
rect 2472 1092 2488 1108
rect 2536 1092 2552 1108
rect 2584 1092 2600 1108
rect 2712 1092 2728 1108
rect 2952 1112 2968 1128
rect 3144 1112 3160 1128
rect 3256 1112 3272 1128
rect 2936 1092 2952 1108
rect 3064 1092 3080 1108
rect 3576 1112 3592 1128
rect 3736 1112 3752 1128
rect 3784 1112 3800 1128
rect 3848 1112 3912 1128
rect 3960 1112 3976 1128
rect 4008 1112 4024 1128
rect 4072 1112 4088 1128
rect 4264 1112 4296 1128
rect 4392 1112 4408 1128
rect 4456 1112 4472 1128
rect 4520 1112 4536 1128
rect 4696 1112 4712 1128
rect 4824 1112 4840 1128
rect 4952 1112 4968 1128
rect 5272 1112 5288 1128
rect 3304 1092 3320 1108
rect 3416 1092 3448 1108
rect 3592 1092 3624 1108
rect 3640 1092 3656 1108
rect 3720 1092 3736 1108
rect 3784 1092 3800 1108
rect 3816 1092 3832 1108
rect 3896 1092 3928 1108
rect 4056 1092 4072 1108
rect 4088 1092 4104 1108
rect 4136 1092 4152 1108
rect 4168 1092 4184 1108
rect 4248 1092 4264 1108
rect 4312 1092 4328 1108
rect 4376 1092 4392 1108
rect 4488 1092 4504 1108
rect 4536 1092 4552 1108
rect 4616 1092 4632 1108
rect 4680 1092 4696 1108
rect 4712 1092 4728 1108
rect 4744 1092 4760 1108
rect 4808 1092 4824 1108
rect 4856 1092 4888 1108
rect 4936 1092 4952 1108
rect 4968 1092 4984 1108
rect 5080 1092 5096 1108
rect 200 1072 216 1088
rect 296 1072 312 1088
rect 376 1072 392 1088
rect 472 1072 488 1088
rect 632 1072 648 1088
rect 936 1072 952 1088
rect 984 1072 1000 1088
rect 1016 1072 1032 1088
rect 1048 1072 1080 1088
rect 1192 1072 1208 1088
rect 1240 1072 1256 1088
rect 1288 1072 1304 1088
rect 1352 1072 1368 1088
rect 1400 1072 1416 1088
rect 1448 1072 1464 1088
rect 1480 1072 1496 1088
rect 1592 1072 1624 1088
rect 1672 1072 1688 1088
rect 1704 1072 1720 1088
rect 1928 1072 1944 1088
rect 1976 1072 1992 1088
rect 2024 1072 2040 1088
rect 2072 1072 2104 1088
rect 2216 1072 2232 1088
rect 2280 1072 2296 1088
rect 2344 1072 2360 1088
rect 2424 1072 2440 1088
rect 2456 1072 2472 1088
rect 2488 1072 2504 1088
rect 2840 1072 2856 1088
rect 2872 1072 2888 1088
rect 2936 1072 2952 1088
rect 2984 1072 3000 1088
rect 3016 1072 3032 1088
rect 3192 1072 3208 1088
rect 3272 1072 3288 1088
rect 3320 1072 3336 1088
rect 3560 1072 3576 1088
rect 3624 1072 3640 1088
rect 5144 1090 5160 1106
rect 5464 1112 5480 1128
rect 5320 1092 5336 1108
rect 5512 1112 5528 1128
rect 5768 1112 5784 1128
rect 5832 1112 5848 1128
rect 6040 1112 6056 1128
rect 6088 1112 6104 1128
rect 6120 1112 6136 1128
rect 5528 1092 5544 1108
rect 5688 1092 5704 1108
rect 5800 1092 5816 1108
rect 5864 1092 5880 1108
rect 5944 1092 5960 1108
rect 6040 1092 6056 1108
rect 6392 1112 6408 1128
rect 6456 1112 6472 1128
rect 6488 1112 6504 1128
rect 6520 1112 6536 1128
rect 6584 1112 6600 1128
rect 6776 1112 6792 1128
rect 6796 1112 6812 1128
rect 6840 1112 6856 1128
rect 6904 1112 6920 1128
rect 7080 1112 7096 1128
rect 7160 1112 7176 1128
rect 7224 1112 7240 1128
rect 7368 1112 7384 1128
rect 6200 1092 6216 1108
rect 6280 1092 6296 1108
rect 6424 1092 6440 1108
rect 6504 1092 6520 1108
rect 6552 1092 6568 1108
rect 6616 1092 6632 1108
rect 6696 1092 6712 1108
rect 6808 1092 6824 1108
rect 6872 1092 6888 1108
rect 6936 1092 6952 1108
rect 7016 1092 7032 1108
rect 7064 1092 7080 1108
rect 7128 1092 7144 1108
rect 7192 1092 7208 1108
rect 7256 1092 7272 1108
rect 7336 1092 7352 1108
rect 7384 1092 7400 1108
rect 3816 1072 3832 1088
rect 3928 1072 3944 1088
rect 3976 1072 4008 1088
rect 4088 1072 4104 1088
rect 4504 1072 4520 1088
rect 4632 1072 4648 1088
rect 4760 1072 4776 1088
rect 4888 1072 4904 1088
rect 4936 1072 4952 1088
rect 5208 1072 5224 1088
rect 5240 1072 5256 1088
rect 5336 1072 5368 1088
rect 5432 1072 5448 1088
rect 5736 1072 5752 1088
rect 5784 1072 5800 1088
rect 5816 1072 5832 1088
rect 5880 1072 5912 1088
rect 6024 1072 6040 1088
rect 6088 1072 6104 1088
rect 6152 1072 6168 1088
rect 6184 1072 6200 1088
rect 6264 1072 6280 1088
rect 6328 1072 6344 1088
rect 6440 1072 6456 1088
rect 6504 1072 6520 1088
rect 6568 1072 6584 1088
rect 6632 1072 6648 1088
rect 6664 1072 6680 1088
rect 6824 1072 6840 1088
rect 6856 1072 6872 1088
rect 6888 1072 6904 1088
rect 6952 1072 6984 1088
rect 7144 1072 7160 1088
rect 7208 1072 7224 1088
rect 7272 1072 7288 1088
rect 7304 1072 7336 1088
rect 600 1052 616 1068
rect 824 1052 840 1068
rect 888 1052 904 1068
rect 2232 1052 2248 1068
rect 2392 1052 2408 1068
rect 2568 1052 2584 1068
rect 2696 1052 2712 1068
rect 3480 1052 3496 1068
rect 3672 1052 3688 1068
rect 3784 1052 3800 1068
rect 3960 1052 3976 1068
rect 4136 1052 4152 1068
rect 4408 1052 4424 1068
rect 4440 1052 4456 1068
rect 4904 1052 4920 1068
rect 5912 1052 5928 1068
rect 6264 1052 6280 1068
rect 6680 1052 6696 1068
rect 7016 1052 7032 1068
rect 7416 1052 7432 1068
rect 1208 1032 1224 1048
rect 1272 1032 1288 1048
rect 1336 1032 1352 1048
rect 1384 1032 1400 1048
rect 1464 1032 1480 1048
rect 1528 1032 1544 1048
rect 1896 1032 1912 1048
rect 2952 1032 2968 1048
rect 3544 1032 3560 1048
rect 3848 1032 3864 1048
rect 4024 1032 4040 1048
rect 4184 1032 4200 1048
rect 4296 1032 4312 1048
rect 4584 1032 4600 1048
rect 5000 1032 5032 1048
rect 5928 1032 5944 1048
rect 6296 1032 6312 1048
rect 6392 1032 6408 1048
rect 6520 1032 6536 1048
rect 6584 1032 6600 1048
rect 6680 1032 6696 1048
rect 7000 1032 7016 1048
rect 7224 1032 7240 1048
rect 7288 1032 7304 1048
rect 2157 1002 2193 1018
rect 4205 1002 4241 1018
rect 6237 1002 6273 1018
rect 184 972 200 988
rect 520 972 536 988
rect 584 972 600 988
rect 904 972 920 988
rect 1400 972 1416 988
rect 1800 972 1816 988
rect 2024 972 2040 988
rect 2168 972 2184 988
rect 2568 972 2584 988
rect 3352 972 3368 988
rect 3416 972 3432 988
rect 3560 972 3576 988
rect 3592 972 3608 988
rect 4408 972 4424 988
rect 4968 972 4984 988
rect 5064 972 5080 988
rect 5176 972 5192 988
rect 5752 972 5768 988
rect 6328 972 6344 988
rect 6440 972 6456 988
rect 6728 972 6744 988
rect 6840 972 6856 988
rect 6904 972 6920 988
rect 7080 972 7096 988
rect 7240 972 7256 988
rect 440 952 456 968
rect 680 952 696 968
rect 1544 952 1560 968
rect 1672 952 1688 968
rect 1736 952 1752 968
rect 1784 952 1800 968
rect 1848 952 1864 968
rect 1960 952 1976 968
rect 2296 952 2312 968
rect 2328 952 2360 968
rect 2504 952 2520 968
rect 2696 952 2712 968
rect 2872 952 2888 968
rect 4104 952 4120 968
rect 4488 952 4504 968
rect 4600 952 4616 968
rect 4808 952 4824 968
rect 5608 952 5624 968
rect 6520 952 6536 968
rect 6776 952 6792 968
rect 200 932 216 948
rect 296 932 312 948
rect 424 932 440 948
rect 536 932 552 948
rect 616 932 632 948
rect 648 932 664 948
rect 744 932 760 948
rect 824 932 840 948
rect 920 932 936 948
rect 1016 932 1032 948
rect 1144 932 1176 948
rect 1192 932 1208 948
rect 1224 932 1240 948
rect 1256 932 1272 948
rect 1288 932 1304 948
rect 1352 932 1368 948
rect 1416 932 1432 948
rect 1448 932 1464 948
rect 1480 932 1496 948
rect 1592 932 1608 948
rect 1656 932 1672 948
rect 1880 932 1896 948
rect 2008 932 2024 948
rect 2088 932 2104 948
rect 2168 932 2184 948
rect 2280 932 2296 948
rect 2392 932 2408 948
rect 2456 932 2472 948
rect 2680 932 2696 948
rect 2760 932 2776 948
rect 2792 932 2808 948
rect 2856 932 2888 948
rect 2952 932 2968 948
rect 72 912 88 928
rect 120 912 136 928
rect 216 912 248 928
rect 360 912 376 928
rect 488 912 504 928
rect 552 912 568 928
rect 632 912 648 928
rect 712 912 728 928
rect 792 912 808 928
rect 920 912 936 928
rect 264 892 280 908
rect 328 892 344 908
rect 520 892 536 908
rect 584 892 616 908
rect 936 892 952 908
rect 1032 912 1064 928
rect 1096 912 1112 928
rect 1176 912 1192 928
rect 1240 912 1256 928
rect 1304 912 1320 928
rect 1368 912 1384 928
rect 1416 912 1432 928
rect 1496 912 1512 928
rect 1576 912 1592 928
rect 1608 912 1624 928
rect 1640 912 1656 928
rect 1704 912 1720 928
rect 1784 912 1800 928
rect 1896 912 1912 928
rect 1944 912 1960 928
rect 1992 912 2008 928
rect 2024 912 2040 928
rect 2104 912 2120 928
rect 2152 912 2168 928
rect 2232 912 2248 928
rect 2296 912 2312 928
rect 2376 912 2392 928
rect 2408 912 2456 928
rect 2472 912 2504 928
rect 2696 914 2712 930
rect 984 892 1000 908
rect 1208 892 1224 908
rect 1272 892 1288 908
rect 1316 892 1332 908
rect 1336 892 1352 908
rect 1400 892 1416 908
rect 1464 892 1480 908
rect 1528 892 1544 908
rect 1608 892 1624 908
rect 2792 892 2808 908
rect 2840 912 2856 928
rect 2904 912 2920 928
rect 2968 912 2984 928
rect 3032 932 3048 948
rect 3160 932 3176 948
rect 3192 932 3208 948
rect 3368 932 3384 948
rect 3464 932 3480 948
rect 3576 932 3592 948
rect 3640 932 3672 948
rect 3832 932 3848 948
rect 3944 932 3960 948
rect 4072 932 4088 948
rect 4120 932 4136 948
rect 4248 932 4264 948
rect 4376 932 4392 948
rect 4520 932 4536 948
rect 4632 932 4648 948
rect 4696 932 4712 948
rect 4760 932 4776 948
rect 5016 932 5032 948
rect 5080 932 5096 948
rect 5336 932 5352 948
rect 5368 932 5384 948
rect 5400 932 5416 948
rect 5464 932 5480 948
rect 5512 932 5528 948
rect 5560 932 5576 948
rect 5688 932 5704 948
rect 5784 932 5800 948
rect 5848 932 5864 948
rect 5976 932 5992 948
rect 6200 932 6216 948
rect 6440 932 6456 948
rect 6488 932 6504 948
rect 6568 932 6584 948
rect 3048 912 3064 928
rect 2952 892 2968 908
rect 3060 892 3076 908
rect 3224 914 3240 930
rect 3384 912 3400 928
rect 3096 892 3112 908
rect 3496 912 3512 928
rect 3624 912 3640 928
rect 3656 912 3672 928
rect 3784 912 3800 928
rect 3848 912 3864 928
rect 3912 912 3928 928
rect 3960 912 3976 928
rect 4040 912 4056 928
rect 4200 912 4216 928
rect 4248 912 4264 928
rect 4328 912 4344 928
rect 4440 912 4456 928
rect 4520 912 4536 928
rect 4552 912 4568 928
rect 4680 912 4696 928
rect 4744 912 4760 928
rect 4776 912 4792 928
rect 4808 912 4824 928
rect 4840 912 4856 928
rect 4904 912 4920 928
rect 5016 912 5048 928
rect 5096 912 5128 928
rect 5240 912 5256 928
rect 5304 914 5320 930
rect 3432 892 3448 908
rect 3480 892 3496 908
rect 3544 892 3560 908
rect 3592 892 3608 908
rect 3704 892 3720 908
rect 3800 892 3816 908
rect 3864 892 3880 908
rect 3928 892 3944 908
rect 3992 892 4008 908
rect 4056 892 4072 908
rect 4104 892 4120 908
rect 4152 892 4168 908
rect 4264 892 4280 908
rect 4296 892 4328 908
rect 4408 892 4440 908
rect 4536 892 4552 908
rect 4648 892 4664 908
rect 4712 892 4728 908
rect 4744 892 4760 908
rect 4824 892 4840 908
rect 4888 892 4904 908
rect 5064 892 5080 908
rect 5128 892 5144 908
rect 5400 892 5416 908
rect 5448 912 5480 928
rect 5608 912 5624 928
rect 5640 912 5656 928
rect 5704 912 5736 928
rect 5800 912 5816 928
rect 5832 912 5848 928
rect 5992 912 6008 928
rect 6072 912 6088 928
rect 6184 914 6200 930
rect 6408 912 6424 928
rect 6488 912 6504 928
rect 6632 912 6648 928
rect 6744 912 6760 928
rect 6792 912 6808 928
rect 6888 932 6904 948
rect 6936 952 6952 968
rect 7096 952 7112 968
rect 6984 932 7000 948
rect 7224 932 7240 948
rect 6968 912 6984 928
rect 7000 912 7016 928
rect 7096 912 7112 928
rect 7208 912 7224 928
rect 7304 912 7320 928
rect 7352 912 7368 928
rect 5832 892 5848 908
rect 6360 892 6376 908
rect 7032 892 7048 908
rect 7160 892 7176 908
rect 7208 892 7224 908
rect 3512 872 3528 888
rect 3768 872 3784 888
rect 3832 872 3848 888
rect 3896 872 3912 888
rect 4024 872 4040 888
rect 1576 852 1592 868
rect 1992 852 2008 868
rect 3960 852 3976 868
rect 4072 872 4088 888
rect 4232 872 4248 888
rect 4344 872 4360 888
rect 4456 872 4472 888
rect 4568 872 4584 888
rect 4856 872 4872 888
rect 4920 872 4936 888
rect 1496 832 1512 848
rect 2376 832 2392 848
rect 3496 832 3512 848
rect 3912 832 3928 848
rect 4328 832 4344 848
rect 4472 832 4488 848
rect 4584 832 4600 848
rect 4872 832 4888 848
rect 4936 832 4952 848
rect 5656 832 5672 848
rect 6104 832 6120 848
rect 6392 832 6408 848
rect 1117 802 1153 818
rect 3165 802 3201 818
rect 5213 802 5249 818
rect 600 772 616 788
rect 648 772 664 788
rect 1048 772 1064 788
rect 1112 772 1128 788
rect 1352 772 1368 788
rect 1848 772 1864 788
rect 1928 772 1944 788
rect 2264 772 2280 788
rect 2440 772 2456 788
rect 2936 772 2952 788
rect 3672 772 3704 788
rect 3848 772 3864 788
rect 3976 772 3992 788
rect 4024 772 4040 788
rect 4104 772 4120 788
rect 4152 772 4168 788
rect 4264 772 4280 788
rect 5112 772 5128 788
rect 5448 772 5464 788
rect 5560 772 5576 788
rect 5768 772 5784 788
rect 5960 772 5976 788
rect 6360 772 6376 788
rect 6456 772 6472 788
rect 7208 772 7224 788
rect 7416 772 7432 788
rect 440 732 456 748
rect 904 732 920 748
rect 936 732 952 748
rect 1800 732 1816 748
rect 2552 732 2568 748
rect 3064 732 3080 748
rect 3528 732 3544 748
rect 3560 732 3576 748
rect 3832 732 3848 748
rect 3992 732 4008 748
rect 4088 732 4104 748
rect 4120 732 4136 748
rect 4248 732 4264 748
rect 4696 732 4712 748
rect 5160 732 5176 748
rect 5240 732 5256 748
rect 6120 732 6136 748
rect 6888 732 6920 748
rect 8 712 24 728
rect 40 712 56 728
rect 472 712 488 728
rect 40 692 56 708
rect 136 692 152 708
rect 328 692 344 708
rect 456 692 472 708
rect 520 712 536 728
rect 584 712 600 728
rect 552 692 568 708
rect 712 692 728 708
rect 808 692 824 708
rect 936 692 952 708
rect 984 712 1000 728
rect 1064 692 1096 708
rect 1128 692 1144 708
rect 1160 692 1176 708
rect 1256 712 1272 728
rect 1416 712 1432 728
rect 1288 692 1304 708
rect 1320 692 1336 708
rect 1368 692 1384 708
rect 1400 692 1416 708
rect 1464 712 1480 728
rect 1512 692 1528 708
rect 1576 712 1592 728
rect 1672 690 1688 706
rect 1816 692 1848 708
rect 1880 692 1896 708
rect 1960 692 1992 708
rect 2072 692 2088 708
rect 2120 692 2136 708
rect 2216 692 2232 708
rect 2312 692 2328 708
rect 2360 712 2376 728
rect 2536 712 2552 728
rect 2744 712 2760 728
rect 2424 692 2440 708
rect 2472 692 2504 708
rect 2664 692 2680 708
rect 2792 692 2808 708
rect 2856 712 2872 728
rect 2904 692 2936 708
rect 2968 692 3000 708
rect 3128 692 3144 708
rect 3176 692 3192 708
rect 3288 692 3304 708
rect 3416 692 3432 708
rect 3560 692 3576 708
rect 3608 712 3624 728
rect 3816 712 3832 728
rect 3848 712 3864 728
rect 3896 712 3912 728
rect 3992 712 4008 728
rect 4104 712 4120 728
rect 4136 712 4152 728
rect 4280 712 4296 728
rect 4328 712 4344 728
rect 3736 692 3752 708
rect 3848 692 3864 708
rect 3976 692 3992 708
rect 4056 692 4072 708
rect 4104 692 4120 708
rect 4152 692 4168 708
rect 4264 692 4280 708
rect 4376 712 4392 728
rect 4392 692 4408 708
rect 4520 692 4536 708
rect 4616 692 4632 708
rect 4664 712 4680 728
rect 4824 692 4840 708
rect 4904 692 4920 708
rect 5000 692 5016 708
rect 5048 712 5064 728
rect 56 672 72 688
rect 120 672 136 688
rect 344 672 360 688
rect 456 672 472 688
rect 568 672 584 688
rect 616 672 632 688
rect 680 672 696 688
rect 744 672 760 688
rect 920 672 936 688
rect 1016 672 1032 688
rect 632 652 648 668
rect 1192 672 1208 688
rect 1288 672 1304 688
rect 1384 672 1400 688
rect 1496 672 1528 688
rect 1576 672 1592 688
rect 1608 672 1624 688
rect 1688 672 1704 688
rect 2296 672 2312 688
rect 2360 672 2376 688
rect 2408 672 2424 688
rect 2504 672 2520 688
rect 2680 672 2696 688
rect 2776 672 2808 688
rect 2856 672 2872 688
rect 2888 672 2904 688
rect 3272 672 3288 688
rect 3400 672 3416 688
rect 3544 672 3560 688
rect 3640 672 3656 688
rect 2040 652 2056 668
rect 2072 652 2104 668
rect 2120 652 2136 668
rect 3720 672 3736 688
rect 3784 672 3800 688
rect 3928 672 3944 688
rect 4296 672 4312 688
rect 4392 672 4408 688
rect 4600 672 4616 688
rect 4664 672 4680 688
rect 4696 672 4712 688
rect 4968 672 5000 688
rect 5048 672 5064 688
rect 5096 692 5128 708
rect 5544 712 5560 728
rect 5576 712 5592 728
rect 5656 712 5672 728
rect 6020 712 6036 728
rect 6040 712 6056 728
rect 6376 712 6408 728
rect 6424 712 6440 728
rect 7144 712 7160 728
rect 5352 692 5368 708
rect 5592 692 5608 708
rect 5704 692 5720 708
rect 5880 692 5896 708
rect 5096 672 5112 688
rect 5208 672 5224 688
rect 5336 672 5352 688
rect 5432 672 5448 688
rect 5544 672 5560 688
rect 5640 672 5672 688
rect 5688 672 5704 688
rect 5928 672 5944 688
rect 5976 672 5992 688
rect 6008 692 6024 708
rect 6056 692 6072 708
rect 6232 692 6248 708
rect 6424 692 6440 708
rect 6568 692 6584 708
rect 6680 692 6696 708
rect 6760 690 6776 706
rect 7032 690 7048 706
rect 7128 692 7144 708
rect 7192 692 7208 708
rect 7288 690 7304 706
rect 6088 672 6104 688
rect 6280 672 6296 688
rect 6328 672 6360 688
rect 6440 672 6456 688
rect 6648 672 6664 688
rect 6696 672 6712 688
rect 6776 672 6792 688
rect 7176 672 7192 688
rect 7224 672 7240 688
rect 7256 672 7272 688
rect 3704 652 3720 668
rect 4536 652 4552 668
rect 4840 652 4856 668
rect 4952 652 4968 668
rect 5512 652 5528 668
rect 7032 652 7048 668
rect 7096 652 7112 668
rect 248 632 264 648
rect 1240 632 1256 648
rect 2008 632 2024 648
rect 2536 632 2552 648
rect 2744 632 2760 648
rect 3032 632 3048 648
rect 3320 632 3336 648
rect 3768 632 3784 648
rect 3896 632 3912 648
rect 4024 632 4040 648
rect 4408 632 4424 648
rect 4936 632 4952 648
rect 5672 632 5688 648
rect 5736 632 5752 648
rect 7208 632 7224 648
rect 2157 602 2193 618
rect 4205 602 4241 618
rect 6237 602 6273 618
rect 8 572 24 588
rect 504 572 520 588
rect 568 572 584 588
rect 904 572 920 588
rect 1208 572 1224 588
rect 1272 572 1288 588
rect 1496 572 1512 588
rect 1752 572 1768 588
rect 2056 572 2072 588
rect 2296 572 2312 588
rect 2344 572 2360 588
rect 2840 572 2856 588
rect 2872 572 2888 588
rect 3000 572 3016 588
rect 3048 572 3064 588
rect 3688 572 3704 588
rect 4056 572 4072 588
rect 4120 572 4136 588
rect 4264 572 4280 588
rect 4856 572 4872 588
rect 5176 572 5192 588
rect 5352 572 5368 588
rect 5432 572 5448 588
rect 5704 572 5720 588
rect 5768 572 5784 588
rect 5832 572 5864 588
rect 6040 572 6056 588
rect 6312 572 6328 588
rect 6776 572 6792 588
rect 6904 572 6920 588
rect 7016 572 7032 588
rect 7160 572 7176 588
rect 7192 572 7208 588
rect 2072 552 2088 568
rect 2136 552 2152 568
rect 4200 552 4216 568
rect 4312 552 4328 568
rect 5784 552 5800 568
rect 6456 552 6472 568
rect 40 532 72 548
rect 168 532 184 548
rect 264 532 280 548
rect 376 532 392 548
rect 488 532 504 548
rect 536 532 552 548
rect 584 532 600 548
rect 648 532 664 548
rect 712 532 728 548
rect 968 532 984 548
rect 1080 532 1096 548
rect 1336 532 1352 548
rect 1512 532 1528 548
rect 1768 532 1784 548
rect 1800 532 1816 548
rect 1832 532 1848 548
rect 2120 532 2136 548
rect 2168 532 2184 548
rect 2504 532 2520 548
rect 2584 532 2616 548
rect 2648 532 2664 548
rect 2680 532 2696 548
rect 2984 532 3000 548
rect 3224 532 3240 548
rect 3288 532 3304 548
rect 3368 532 3384 548
rect 3528 532 3544 548
rect 3704 532 3720 548
rect 3800 532 3832 548
rect 3864 532 3880 548
rect 4104 532 4120 548
rect 4328 532 4344 548
rect 4408 532 4424 548
rect 4440 532 4472 548
rect 4488 532 4504 548
rect 4520 532 4536 548
rect 4568 532 4584 548
rect 4632 532 4648 548
rect 4664 532 4680 548
rect 4872 532 4888 548
rect 4984 532 5000 548
rect 5224 532 5240 548
rect 5320 532 5352 548
rect 5384 532 5400 548
rect 5592 532 5608 548
rect 5624 532 5640 548
rect 5688 532 5704 548
rect 5800 532 5816 548
rect 5960 532 5976 548
rect 6072 532 6104 548
rect 6136 532 6152 548
rect 6168 532 6184 548
rect 6232 532 6248 548
rect 6280 532 6296 548
rect 6376 532 6408 548
rect 6648 532 6664 548
rect 6808 532 6824 548
rect 6952 532 6968 548
rect 7064 532 7080 548
rect 7128 532 7160 548
rect 7432 532 7448 548
rect 72 512 88 528
rect 8 492 24 508
rect 152 512 168 528
rect 248 512 264 528
rect 296 512 312 528
rect 392 512 408 528
rect 392 492 408 508
rect 472 512 488 528
rect 632 512 648 528
rect 680 512 696 528
rect 712 512 728 528
rect 792 512 808 528
rect 840 512 856 528
rect 952 512 968 528
rect 1000 512 1016 528
rect 1096 512 1112 528
rect 1304 512 1320 528
rect 1416 512 1432 528
rect 1560 512 1576 528
rect 1640 512 1656 528
rect 1688 512 1704 528
rect 1784 512 1800 528
rect 1944 512 1960 528
rect 1976 512 1992 528
rect 2136 512 2152 528
rect 2264 512 2280 528
rect 2328 512 2344 528
rect 2456 512 2472 528
rect 2616 512 2632 528
rect 2728 512 2744 528
rect 2920 512 2936 528
rect 2968 512 2984 528
rect 3080 512 3096 528
rect 3144 512 3160 528
rect 3192 512 3208 528
rect 3256 512 3272 528
rect 3304 512 3320 528
rect 3432 512 3464 528
rect 3576 512 3592 528
rect 3720 512 3736 528
rect 504 492 520 508
rect 536 492 552 508
rect 664 492 680 508
rect 936 492 968 508
rect 1016 492 1032 508
rect 1864 492 1880 508
rect 2072 492 2088 508
rect 2136 492 2152 508
rect 2536 492 2552 508
rect 2568 492 2584 508
rect 2648 492 2664 508
rect 3016 492 3032 508
rect 3832 512 3848 528
rect 3944 512 3960 528
rect 3976 512 3992 528
rect 4152 512 4168 528
rect 4296 512 4312 528
rect 4344 512 4360 528
rect 4472 512 4488 528
rect 4584 512 4600 528
rect 3768 492 3784 508
rect 3864 492 3880 508
rect 4104 492 4136 508
rect 4392 492 4408 508
rect 4552 492 4568 508
rect 4728 514 4744 530
rect 4792 512 4808 528
rect 4920 512 4936 528
rect 5032 512 5048 528
rect 5208 512 5224 528
rect 4632 492 4648 508
rect 4904 492 4920 508
rect 5560 514 5576 530
rect 5624 512 5656 528
rect 5976 514 5992 530
rect 6136 512 6152 528
rect 5288 492 5304 508
rect 5368 492 5384 508
rect 5416 492 5432 508
rect 5652 492 5668 508
rect 5672 492 5688 508
rect 5832 492 5848 508
rect 6040 492 6056 508
rect 6120 492 6136 508
rect 6312 512 6328 528
rect 6200 492 6216 508
rect 6312 492 6328 508
rect 6360 512 6376 528
rect 6440 512 6456 528
rect 6600 512 6616 528
rect 6680 512 6696 528
rect 6744 512 6760 528
rect 6792 512 6808 528
rect 7016 512 7032 528
rect 7048 512 7064 528
rect 7112 512 7128 528
rect 7256 512 7272 528
rect 7304 512 7320 528
rect 7384 512 7400 528
rect 6360 492 6376 508
rect 7000 492 7032 508
rect 7080 492 7096 508
rect 7112 492 7128 508
rect 7176 492 7192 508
rect 120 472 136 488
rect 360 472 376 488
rect 440 472 456 488
rect 600 472 616 488
rect 632 472 648 488
rect 2936 472 2952 488
rect 4072 472 4088 488
rect 6104 472 6120 488
rect 72 432 88 448
rect 1272 432 1288 448
rect 2232 432 2248 448
rect 3112 432 3128 448
rect 3224 432 3240 448
rect 3400 432 3416 448
rect 3480 432 3496 448
rect 3720 432 3736 448
rect 4264 432 4280 448
rect 4376 432 4392 448
rect 4888 432 4904 448
rect 4952 432 4968 448
rect 5400 432 5416 448
rect 6712 432 6728 448
rect 6824 432 6840 448
rect 1117 402 1153 418
rect 3165 402 3201 418
rect 5213 402 5249 418
rect 376 372 392 388
rect 568 372 584 388
rect 1176 372 1192 388
rect 1624 372 1640 388
rect 1992 372 2008 388
rect 2088 372 2104 388
rect 2504 372 2520 388
rect 2936 372 2952 388
rect 4104 372 4120 388
rect 4136 372 4152 388
rect 4440 372 4456 388
rect 4744 372 4760 388
rect 4824 372 4840 388
rect 4872 372 4888 388
rect 4984 372 5000 388
rect 5528 372 5544 388
rect 5576 372 5592 388
rect 6728 372 6744 388
rect 6968 372 6984 388
rect 7064 372 7080 388
rect 3688 352 3704 368
rect 5720 352 5736 368
rect 200 332 216 348
rect 1016 332 1032 348
rect 1272 332 1288 348
rect 1480 332 1496 348
rect 1848 332 1864 348
rect 2344 332 2360 348
rect 2744 332 2760 348
rect 2984 332 3000 348
rect 3608 332 3624 348
rect 4632 332 4648 348
rect 6296 332 6312 348
rect 6648 332 6664 348
rect 232 312 248 328
rect 88 292 104 308
rect 120 292 136 308
rect 312 312 328 328
rect 600 312 632 328
rect 692 312 708 328
rect 712 312 728 328
rect 760 312 776 328
rect 312 292 328 308
rect 472 292 488 308
rect 680 292 696 308
rect 808 312 824 328
rect 1256 312 1272 328
rect 824 292 840 308
rect 888 290 904 306
rect 952 292 968 308
rect 1032 292 1048 308
rect 1128 292 1160 308
rect 1192 292 1208 308
rect 200 272 216 288
rect 232 272 248 288
rect 296 272 312 288
rect 456 272 472 288
rect 584 272 600 288
rect 728 272 744 288
rect 824 272 840 288
rect 856 272 872 288
rect 1080 272 1096 288
rect 1384 292 1400 308
rect 1480 292 1496 308
rect 1528 312 1544 328
rect 1880 312 1896 328
rect 1400 272 1416 288
rect 1464 272 1480 288
rect 1560 272 1576 288
rect 1640 292 1672 308
rect 1736 292 1752 308
rect 1864 292 1880 308
rect 1928 312 1944 328
rect 2376 312 2392 328
rect 2024 292 2040 308
rect 2056 292 2072 308
rect 2104 292 2136 308
rect 2248 292 2264 308
rect 2360 292 2376 308
rect 2424 312 2440 328
rect 2776 312 2792 328
rect 1688 272 1704 288
rect 1864 272 1880 288
rect 1960 272 1976 288
rect 2232 272 2248 288
rect 2360 272 2376 288
rect 2456 272 2472 288
rect 2536 292 2568 308
rect 2632 292 2648 308
rect 2680 292 2696 308
rect 2776 292 2792 308
rect 2824 312 2840 328
rect 2872 312 2888 328
rect 2904 312 2920 328
rect 2968 312 2984 328
rect 3240 312 3256 328
rect 2760 272 2776 288
rect 2872 272 2888 288
rect 2936 292 2952 308
rect 3096 292 3112 308
rect 3288 292 3304 308
rect 3320 292 3336 308
rect 3384 312 3400 328
rect 3624 312 3640 328
rect 3672 312 3688 328
rect 3752 312 3768 328
rect 3480 290 3496 306
rect 3528 292 3544 308
rect 3788 312 3804 328
rect 3912 312 3928 328
rect 4120 312 4136 328
rect 4296 312 4312 328
rect 3816 292 3832 308
rect 3880 292 3912 308
rect 3992 292 4008 308
rect 4184 292 4200 308
rect 4328 292 4344 308
rect 4376 312 4392 328
rect 4712 312 4728 328
rect 4904 312 4920 328
rect 5400 312 5416 328
rect 5464 312 5480 328
rect 5560 312 5576 328
rect 5704 312 5720 328
rect 4504 290 4520 306
rect 4648 292 4664 308
rect 4744 292 4760 308
rect 4776 292 4792 308
rect 4872 292 4888 308
rect 4920 292 4936 308
rect 5016 292 5048 308
rect 5128 292 5144 308
rect 5336 290 5352 306
rect 5400 292 5416 308
rect 5448 292 5464 308
rect 5624 292 5640 308
rect 5672 292 5688 308
rect 5832 292 5848 308
rect 5928 292 5944 308
rect 5976 312 5992 328
rect 6168 292 6184 308
rect 6344 292 6360 308
rect 6392 312 6408 328
rect 6664 312 6680 328
rect 6696 312 6712 328
rect 6984 312 7016 328
rect 7032 312 7048 328
rect 7320 312 7336 328
rect 6520 290 6536 306
rect 6712 292 6728 308
rect 6872 292 6888 308
rect 7032 292 7048 308
rect 7208 292 7224 308
rect 7368 292 7384 308
rect 2920 272 2936 288
rect 3112 272 3128 288
rect 3176 272 3192 288
rect 3240 272 3256 288
rect 3320 272 3336 288
rect 3384 272 3400 288
rect 3416 272 3432 288
rect 3656 272 3672 288
rect 3704 272 3720 288
rect 3816 272 3832 288
rect 3944 272 3960 288
rect 3976 272 3992 288
rect 4152 272 4184 288
rect 4200 272 4216 288
rect 4232 272 4248 288
rect 4312 272 4328 288
rect 4424 272 4440 288
rect 4536 272 4552 288
rect 4760 272 4776 288
rect 4856 272 4872 288
rect 4968 272 4984 288
rect 5080 272 5096 288
rect 5192 272 5208 288
rect 5368 272 5384 288
rect 5448 272 5464 288
rect 5496 272 5528 288
rect 5672 272 5688 288
rect 5880 272 5896 288
rect 5912 272 5928 288
rect 5976 272 5992 288
rect 6008 272 6040 288
rect 6152 272 6168 288
rect 6280 272 6296 288
rect 6312 272 6328 288
rect 6376 272 6392 288
rect 6424 272 6472 288
rect 6488 272 6504 288
rect 6872 272 6888 288
rect 6952 272 6968 288
rect 7192 272 7208 288
rect 7256 272 7272 288
rect 7288 272 7304 288
rect 7384 272 7400 288
rect 56 252 72 268
rect 360 252 376 268
rect 632 252 648 268
rect 3832 252 3848 268
rect 4360 252 4376 268
rect 4424 252 4440 268
rect 4840 252 4856 268
rect 312 232 328 248
rect 1256 232 1272 248
rect 3640 232 3656 248
rect 4680 232 4696 248
rect 4808 232 4824 248
rect 4952 232 4968 248
rect 5064 232 5080 248
rect 5592 252 5608 268
rect 5464 232 5480 248
rect 7336 232 7352 248
rect 2157 202 2193 218
rect 4205 202 4241 218
rect 6237 202 6273 218
rect 184 172 200 188
rect 376 172 392 188
rect 456 172 472 188
rect 936 172 952 188
rect 1096 172 1112 188
rect 1432 172 1448 188
rect 2088 172 2104 188
rect 2296 172 2312 188
rect 2664 172 2680 188
rect 2696 172 2712 188
rect 3000 172 3016 188
rect 3448 172 3464 188
rect 3480 172 3496 188
rect 3784 172 3800 188
rect 3976 172 3992 188
rect 4104 172 4120 188
rect 4488 172 4504 188
rect 4712 172 4728 188
rect 4840 172 4856 188
rect 5208 172 5224 188
rect 5480 172 5496 188
rect 5560 172 5576 188
rect 6088 172 6104 188
rect 6680 172 6696 188
rect 6936 172 6952 188
rect 7128 172 7144 188
rect 7160 172 7176 188
rect 7384 172 7400 188
rect 56 152 72 168
rect 1624 152 1640 168
rect 2680 152 2696 168
rect 3320 152 3336 168
rect 3464 152 3480 168
rect 3656 152 3672 168
rect 3848 152 3864 168
rect 4232 152 4248 168
rect 4616 152 4632 168
rect 4968 152 4984 168
rect 6248 152 6264 168
rect 6536 152 6552 168
rect 7144 152 7160 168
rect 264 132 280 148
rect 440 132 456 148
rect 616 132 632 148
rect 648 132 664 148
rect 680 132 696 148
rect 744 132 760 148
rect 776 132 792 148
rect 840 132 856 148
rect 952 132 968 148
rect 984 132 1000 148
rect 1016 132 1032 148
rect 1192 132 1208 148
rect 1288 132 1304 148
rect 1336 132 1352 148
rect 1480 132 1496 148
rect 1544 132 1560 148
rect 1688 132 1704 148
rect 1800 132 1816 148
rect 1848 132 1864 148
rect 1976 132 1992 148
rect 2104 132 2136 148
rect 2216 132 2232 148
rect 2280 132 2296 148
rect 2568 132 2584 148
rect 2712 132 2728 148
rect 2744 132 2760 148
rect 2808 132 2824 148
rect 2904 132 2920 148
rect 3016 132 3032 148
rect 3048 132 3064 148
rect 3112 132 3144 148
rect 3192 132 3208 148
rect 3256 132 3272 148
rect 3544 132 3560 148
rect 3992 132 4008 148
rect 4088 132 4104 148
rect 4376 132 4392 148
rect 4440 132 4456 148
rect 4680 132 4696 148
rect 4728 132 4744 148
rect 4792 132 4808 148
rect 5368 132 5384 148
rect 5448 132 5464 148
rect 5528 132 5560 148
rect 5576 132 5592 148
rect 5736 132 5752 148
rect 5832 132 5848 148
rect 6184 132 6216 148
rect 6264 132 6280 148
rect 6568 132 6584 148
rect 6808 132 6824 148
rect 6872 132 6888 148
rect 6904 132 6920 148
rect 6968 132 6984 148
rect 7176 132 7192 148
rect 7224 132 7240 148
rect 72 112 88 128
rect 280 112 296 128
rect 392 112 408 128
rect 424 112 440 128
rect 584 114 600 130
rect 392 92 408 108
rect 680 92 696 108
rect 728 112 744 128
rect 824 112 840 128
rect 968 112 984 128
rect 1224 114 1240 130
rect 1352 112 1368 128
rect 1400 112 1416 128
rect 1464 112 1480 128
rect 1496 112 1512 128
rect 1048 92 1064 108
rect 1288 92 1304 108
rect 1704 112 1720 128
rect 1832 112 1848 128
rect 1864 112 1896 128
rect 1960 114 1976 130
rect 2280 112 2296 128
rect 2408 112 2424 128
rect 2552 112 2568 128
rect 1544 92 1560 108
rect 1896 92 1912 108
rect 2184 92 2200 108
rect 2264 92 2280 108
rect 2744 92 2760 108
rect 2792 112 2808 128
rect 2888 112 2904 128
rect 3032 112 3048 128
rect 3144 112 3160 128
rect 3224 112 3240 128
rect 3320 114 3336 130
rect 3496 112 3512 128
rect 3560 112 3576 128
rect 3592 112 3608 128
rect 3656 114 3672 130
rect 3864 112 3880 128
rect 3080 92 3096 108
rect 3192 92 3208 108
rect 3224 92 3240 108
rect 3592 92 3608 108
rect 4024 92 4040 108
rect 4056 112 4088 128
rect 4216 112 4232 128
rect 4328 112 4344 128
rect 4392 112 4408 128
rect 4440 112 4456 128
rect 4600 112 4616 128
rect 4728 112 4744 128
rect 4472 92 4488 108
rect 4712 92 4728 108
rect 4952 112 4968 128
rect 5032 112 5048 128
rect 5080 112 5096 128
rect 5128 112 5144 128
rect 5336 114 5352 130
rect 5400 112 5416 128
rect 5432 112 5448 128
rect 5656 112 5688 128
rect 4792 92 4808 108
rect 5400 92 5416 108
rect 5576 92 5592 108
rect 5768 92 5784 108
rect 5816 112 5832 128
rect 5992 112 6008 128
rect 6120 112 6136 128
rect 6168 112 6184 128
rect 5816 92 5832 108
rect 6136 92 6152 108
rect 6168 92 6184 108
rect 6376 112 6392 128
rect 6408 112 6424 128
rect 6504 112 6520 128
rect 6600 92 6616 108
rect 6648 112 6664 128
rect 6824 112 6840 128
rect 7016 112 7032 128
rect 7192 112 7208 128
rect 7256 114 7272 130
rect 6648 92 6664 108
rect 6936 92 6952 108
rect 3528 32 3544 48
rect 4360 32 4376 48
rect 5064 32 5080 48
rect 5112 32 5128 48
rect 5192 32 5208 48
rect 1117 2 1153 18
rect 3165 2 3201 18
rect 5213 2 5249 18
<< metal2 >>
rect 2893 5388 2899 5463
rect 3085 5428 3091 5463
rect 3053 5388 3059 5412
rect 3069 5388 3075 5392
rect 3117 5388 3123 5412
rect 3133 5408 3139 5463
rect 3165 5428 3171 5463
rect 109 5348 115 5372
rect 381 5328 387 5372
rect 861 5348 867 5372
rect 1517 5368 1523 5372
rect 877 5337 888 5343
rect 605 5328 611 5332
rect 877 5328 883 5337
rect 45 5308 51 5312
rect 77 5308 83 5312
rect 13 4968 19 5032
rect 77 4988 83 5292
rect 77 4928 83 4952
rect 141 4948 147 5090
rect 269 5088 275 5272
rect 285 5108 291 5132
rect 109 4928 115 4932
rect 13 4788 19 4912
rect 13 4648 19 4652
rect 13 4548 19 4592
rect 29 4528 35 4892
rect 61 4808 67 4832
rect 93 4648 99 4912
rect 189 4908 195 4912
rect 237 4728 243 4972
rect 269 4968 275 5072
rect 365 5028 371 5232
rect 381 5128 387 5132
rect 397 5108 403 5312
rect 509 5303 515 5312
rect 653 5308 659 5312
rect 893 5308 899 5312
rect 509 5297 531 5303
rect 525 5188 531 5297
rect 493 5128 499 5152
rect 413 5048 419 5092
rect 461 5048 467 5112
rect 493 5088 499 5112
rect 525 5108 531 5132
rect 573 5128 579 5132
rect 589 5088 595 5232
rect 621 5128 627 5232
rect 285 4928 291 4952
rect 509 4948 515 5072
rect 621 5068 627 5092
rect 637 5088 643 5092
rect 141 4706 147 4712
rect 237 4708 243 4712
rect 301 4688 307 4932
rect 413 4888 419 4932
rect 509 4908 515 4912
rect 381 4688 387 4692
rect 109 4548 115 4572
rect 173 4568 179 4672
rect 205 4668 211 4672
rect 77 4528 83 4532
rect 317 4528 323 4632
rect 333 4528 339 4572
rect 397 4528 403 4832
rect 509 4708 515 4892
rect 509 4688 515 4692
rect 429 4668 435 4672
rect 429 4548 435 4652
rect 525 4608 531 4932
rect 573 4788 579 4912
rect 637 4728 643 5032
rect 653 4948 659 5112
rect 685 5108 691 5152
rect 733 5108 739 5132
rect 781 5128 787 5132
rect 733 5088 739 5092
rect 781 5088 787 5092
rect 845 5088 851 5112
rect 717 5048 723 5072
rect 669 4768 675 5032
rect 685 4928 691 4932
rect 573 4708 579 4712
rect 637 4708 643 4712
rect 429 4528 435 4532
rect 477 4528 483 4532
rect 29 4508 35 4512
rect 13 4308 19 4312
rect 13 4268 19 4272
rect 29 3988 35 4492
rect 77 4288 83 4292
rect 109 4248 115 4272
rect 77 3888 83 4132
rect 93 4128 99 4132
rect 205 4068 211 4132
rect 221 4128 227 4312
rect 237 4308 243 4512
rect 317 4308 323 4512
rect 365 4368 371 4432
rect 381 4328 387 4452
rect 525 4328 531 4512
rect 557 4488 563 4692
rect 605 4677 616 4683
rect 605 4548 611 4677
rect 669 4648 675 4672
rect 701 4668 707 4672
rect 701 4548 707 4572
rect 733 4548 739 5072
rect 813 5048 819 5072
rect 781 4948 787 5032
rect 845 4948 851 4972
rect 781 4848 787 4932
rect 605 4528 611 4532
rect 669 4528 675 4532
rect 701 4528 707 4532
rect 781 4528 787 4632
rect 669 4508 675 4512
rect 717 4508 723 4512
rect 301 4148 307 4172
rect 269 4108 275 4112
rect 269 3948 275 4092
rect 333 4008 339 4252
rect 365 4188 371 4292
rect 397 4243 403 4312
rect 525 4308 531 4312
rect 621 4288 627 4292
rect 669 4288 675 4312
rect 701 4288 707 4332
rect 765 4308 771 4312
rect 605 4268 611 4272
rect 397 4237 419 4243
rect 397 4188 403 4212
rect 413 4188 419 4237
rect 445 4148 451 4172
rect 205 3908 211 3912
rect 349 3908 355 4112
rect 397 4088 403 4092
rect 413 4083 419 4092
rect 413 4077 435 4083
rect 93 3888 99 3892
rect 237 3883 243 3892
rect 221 3877 243 3883
rect 77 3748 83 3872
rect 173 3748 179 3752
rect 29 3588 35 3692
rect 61 3548 67 3632
rect 29 3188 35 3312
rect 77 3088 83 3472
rect 93 3108 99 3492
rect 109 3328 115 3732
rect 173 3528 179 3672
rect 189 3548 195 3612
rect 141 3508 147 3512
rect 205 3428 211 3432
rect 205 3388 211 3392
rect 221 3328 227 3877
rect 253 3808 259 3872
rect 301 3848 307 3872
rect 237 3728 243 3792
rect 349 3788 355 3872
rect 237 3348 243 3492
rect 253 3488 259 3732
rect 301 3728 307 3772
rect 365 3748 371 3892
rect 397 3888 403 3912
rect 413 3888 419 3992
rect 397 3788 403 3852
rect 429 3788 435 4077
rect 461 4008 467 4032
rect 493 3988 499 4112
rect 445 3908 451 3912
rect 541 3908 547 3972
rect 589 3928 595 3972
rect 621 3908 627 4272
rect 717 4128 723 4292
rect 781 4128 787 4472
rect 797 4388 803 4592
rect 845 4528 851 4932
rect 893 4908 899 5292
rect 957 5268 963 5332
rect 1037 5188 1043 5332
rect 1053 5328 1059 5332
rect 1277 5328 1283 5352
rect 1405 5348 1411 5352
rect 2061 5348 2067 5372
rect 1293 5328 1299 5332
rect 1069 5148 1075 5292
rect 1149 5288 1155 5312
rect 1069 5108 1075 5132
rect 1181 5108 1187 5112
rect 909 4988 915 5072
rect 973 4928 979 5032
rect 1133 4968 1139 5072
rect 1149 4928 1155 4932
rect 1197 4928 1203 5312
rect 1373 5308 1379 5312
rect 1437 5308 1443 5312
rect 1437 5288 1443 5292
rect 1245 5188 1251 5232
rect 1453 5228 1459 5292
rect 1309 5088 1315 5132
rect 1341 5108 1347 5112
rect 1293 4928 1299 5032
rect 941 4908 947 4912
rect 893 4888 899 4892
rect 877 4688 883 4832
rect 893 4708 899 4712
rect 941 4588 947 4692
rect 957 4668 963 4912
rect 973 4688 979 4732
rect 989 4708 995 4712
rect 1005 4648 1011 4832
rect 1021 4708 1027 4792
rect 1037 4748 1043 4912
rect 1053 4628 1059 4712
rect 1085 4708 1091 4712
rect 1101 4708 1107 4792
rect 989 4588 995 4612
rect 1149 4568 1155 4672
rect 1277 4668 1283 4812
rect 1325 4668 1331 4832
rect 1229 4648 1235 4652
rect 861 4548 867 4552
rect 813 4348 819 4512
rect 893 4508 899 4512
rect 909 4468 915 4532
rect 829 4308 835 4332
rect 861 4308 867 4352
rect 941 4328 947 4472
rect 957 4468 963 4532
rect 1005 4528 1011 4532
rect 813 4188 819 4272
rect 845 4168 851 4232
rect 893 4128 899 4172
rect 909 4148 915 4272
rect 269 3688 275 3692
rect 333 3648 339 3692
rect 269 3528 275 3532
rect 253 3468 259 3472
rect 269 3408 275 3512
rect 365 3488 371 3732
rect 381 3688 387 3692
rect 461 3688 467 3752
rect 429 3628 435 3632
rect 461 3508 467 3672
rect 381 3428 387 3492
rect 493 3468 499 3892
rect 509 3888 515 3892
rect 589 3888 595 3892
rect 509 3788 515 3872
rect 301 3328 307 3412
rect 445 3388 451 3412
rect 125 3148 131 3232
rect 157 3188 163 3312
rect 221 3188 227 3292
rect 269 3188 275 3312
rect 109 3108 115 3112
rect 29 2988 35 3012
rect 77 2948 83 3072
rect 93 3028 99 3092
rect 157 2928 163 2932
rect 189 2928 195 3092
rect 317 3088 323 3332
rect 461 3328 467 3452
rect 493 3348 499 3432
rect 525 3348 531 3872
rect 621 3848 627 3872
rect 669 3768 675 4032
rect 733 3988 739 4032
rect 685 3868 691 3912
rect 685 3728 691 3832
rect 557 3588 563 3652
rect 605 3508 611 3532
rect 557 3488 563 3492
rect 557 3428 563 3472
rect 685 3388 691 3692
rect 717 3508 723 3712
rect 765 3488 771 3872
rect 781 3568 787 4112
rect 925 4088 931 4092
rect 813 3948 819 4032
rect 797 3748 803 3772
rect 861 3748 867 4032
rect 904 3877 915 3883
rect 893 3788 899 3852
rect 909 3788 915 3877
rect 925 3788 931 3892
rect 909 3728 915 3732
rect 829 3717 840 3723
rect 813 3588 819 3692
rect 797 3488 803 3492
rect 765 3468 771 3472
rect 733 3328 739 3352
rect 461 3308 467 3312
rect 461 3168 467 3292
rect 557 3148 563 3172
rect 365 3108 371 3112
rect 621 3108 627 3312
rect 701 3248 707 3292
rect 669 3237 680 3243
rect 637 3188 643 3232
rect 669 3148 675 3237
rect 749 3183 755 3332
rect 765 3308 771 3332
rect 781 3328 787 3412
rect 813 3388 819 3552
rect 829 3528 835 3717
rect 941 3708 947 4312
rect 957 4188 963 4312
rect 973 4108 979 4492
rect 989 4488 995 4492
rect 973 3928 979 4092
rect 1005 4028 1011 4512
rect 1021 4308 1027 4552
rect 1149 4548 1155 4552
rect 1165 4548 1171 4552
rect 1245 4548 1251 4592
rect 1261 4568 1267 4572
rect 1293 4557 1320 4563
rect 1037 4528 1043 4532
rect 1133 4528 1139 4532
rect 1229 4528 1235 4532
rect 1293 4528 1299 4557
rect 1197 4508 1203 4512
rect 1037 4468 1043 4492
rect 1085 4488 1091 4492
rect 1053 4308 1059 4352
rect 1021 4288 1027 4292
rect 1032 4277 1043 4283
rect 1021 4248 1027 4252
rect 1021 4188 1027 4192
rect 1037 4148 1043 4277
rect 1053 4148 1059 4152
rect 1021 3968 1027 4032
rect 1021 3908 1027 3932
rect 1053 3908 1059 4112
rect 1133 4108 1139 4232
rect 1149 4188 1155 4292
rect 1165 4288 1171 4292
rect 1181 4128 1187 4312
rect 1293 4308 1299 4372
rect 1213 4188 1219 4272
rect 1229 4248 1235 4292
rect 1261 4208 1267 4292
rect 1309 4288 1315 4532
rect 1325 4528 1331 4532
rect 1341 4328 1347 5092
rect 1405 5088 1411 5192
rect 1453 5188 1459 5212
rect 1501 5208 1507 5332
rect 1837 5328 1843 5332
rect 1965 5328 1971 5332
rect 1629 5308 1635 5312
rect 1709 5308 1715 5312
rect 1421 5068 1427 5092
rect 1357 4948 1363 4972
rect 1469 4948 1475 5192
rect 1709 5148 1715 5292
rect 1613 5106 1619 5112
rect 1709 5108 1715 5112
rect 1549 5088 1555 5092
rect 1725 5088 1731 5112
rect 1805 5108 1811 5112
rect 1549 4928 1555 5032
rect 1645 4948 1651 5052
rect 1677 5048 1683 5072
rect 1677 4948 1683 4972
rect 1709 4948 1715 5072
rect 1405 4868 1411 4892
rect 1485 4868 1491 4912
rect 1421 4708 1427 4812
rect 1485 4708 1491 4852
rect 1501 4768 1507 4912
rect 1581 4908 1587 4912
rect 1645 4908 1651 4912
rect 1357 4688 1363 4692
rect 1453 4688 1459 4692
rect 1501 4688 1507 4752
rect 1373 4668 1379 4672
rect 1357 4528 1363 4612
rect 1373 4548 1379 4572
rect 1389 4568 1395 4632
rect 1405 4588 1411 4592
rect 1389 4548 1395 4552
rect 1357 4428 1363 4512
rect 1357 4308 1363 4392
rect 1293 4263 1299 4272
rect 1373 4268 1379 4372
rect 1421 4308 1427 4512
rect 1437 4288 1443 4672
rect 1501 4568 1507 4572
rect 1517 4563 1523 4832
rect 1533 4708 1539 4712
rect 1565 4568 1571 4592
rect 1512 4557 1523 4563
rect 1485 4528 1491 4532
rect 1485 4508 1491 4512
rect 1453 4328 1459 4432
rect 1533 4408 1539 4512
rect 1581 4443 1587 4692
rect 1597 4688 1603 4832
rect 1597 4508 1603 4512
rect 1581 4437 1603 4443
rect 1469 4317 1480 4323
rect 1389 4277 1400 4283
rect 1293 4257 1320 4263
rect 1357 4243 1363 4252
rect 1389 4243 1395 4277
rect 1357 4237 1395 4243
rect 1197 4148 1203 4152
rect 1149 4108 1155 4112
rect 1277 4103 1283 4112
rect 1277 4097 1299 4103
rect 1069 3948 1075 4072
rect 1069 3928 1075 3932
rect 957 3868 963 3872
rect 957 3728 963 3732
rect 893 3588 899 3672
rect 829 3508 835 3512
rect 845 3388 851 3512
rect 861 3348 867 3412
rect 909 3408 915 3492
rect 925 3368 931 3452
rect 941 3428 947 3492
rect 957 3428 963 3712
rect 973 3688 979 3892
rect 1069 3888 1075 3892
rect 989 3728 995 3832
rect 1005 3828 1011 3872
rect 1005 3808 1011 3812
rect 1101 3788 1107 4092
rect 1293 3948 1299 4097
rect 1133 3888 1139 3932
rect 1069 3748 1075 3772
rect 1053 3728 1059 3732
rect 973 3588 979 3632
rect 973 3428 979 3492
rect 733 3177 755 3183
rect 701 3108 707 3112
rect 573 3097 584 3103
rect 205 3048 211 3052
rect 205 2948 211 2972
rect 365 2968 371 3072
rect 301 2948 307 2952
rect 461 2928 467 3072
rect 509 3048 515 3092
rect 493 2968 499 2972
rect 557 2928 563 2932
rect 13 2728 19 2732
rect 13 2548 19 2552
rect 29 2528 35 2552
rect 61 2488 67 2492
rect 77 2448 83 2912
rect 125 2888 131 2912
rect 189 2908 195 2912
rect 141 2706 147 2732
rect 237 2728 243 2912
rect 269 2908 275 2912
rect 397 2788 403 2892
rect 461 2748 467 2912
rect 269 2728 275 2732
rect 205 2688 211 2712
rect 237 2708 243 2712
rect 509 2708 515 2892
rect 93 2588 99 2652
rect 109 2568 115 2592
rect 109 2528 115 2552
rect 141 2508 147 2512
rect 141 2488 147 2492
rect 13 2268 19 2332
rect 77 1908 83 2432
rect 173 2288 179 2672
rect 189 2548 195 2592
rect 237 2328 243 2692
rect 301 2688 307 2692
rect 253 2588 259 2632
rect 269 2488 275 2552
rect 301 2508 307 2512
rect 237 2288 243 2292
rect 173 2148 179 2272
rect 205 2268 211 2272
rect 205 2148 211 2152
rect 221 2128 227 2232
rect 157 1908 163 1932
rect 253 1928 259 2312
rect 269 2308 275 2472
rect 317 2448 323 2692
rect 365 2688 371 2692
rect 509 2688 515 2692
rect 381 2648 387 2672
rect 541 2668 547 2692
rect 397 2648 403 2652
rect 381 2608 387 2632
rect 429 2548 435 2632
rect 557 2628 563 2912
rect 573 2908 579 3097
rect 632 3077 643 3083
rect 589 2988 595 3052
rect 637 2988 643 3077
rect 685 2988 691 3072
rect 616 2917 627 2923
rect 589 2763 595 2892
rect 621 2888 627 2917
rect 685 2908 691 2912
rect 605 2788 611 2792
rect 621 2788 627 2872
rect 589 2757 611 2763
rect 573 2668 579 2692
rect 573 2648 579 2652
rect 605 2588 611 2757
rect 637 2708 643 2832
rect 333 2508 339 2512
rect 285 2308 291 2312
rect 317 2308 323 2432
rect 349 2388 355 2492
rect 301 2248 307 2272
rect 349 2188 355 2232
rect 301 2128 307 2172
rect 317 2108 323 2132
rect 365 2108 371 2532
rect 381 2528 387 2532
rect 397 2503 403 2512
rect 392 2497 403 2503
rect 413 2188 419 2312
rect 429 2148 435 2292
rect 525 2268 531 2512
rect 589 2508 595 2572
rect 621 2408 627 2632
rect 653 2628 659 2672
rect 685 2668 691 2692
rect 701 2668 707 3092
rect 733 2928 739 3177
rect 765 3103 771 3112
rect 749 3097 771 3103
rect 749 3088 755 3097
rect 765 2928 771 2992
rect 813 2988 819 3292
rect 829 3188 835 3292
rect 957 3143 963 3392
rect 1021 3188 1027 3452
rect 1053 3388 1059 3492
rect 957 3137 968 3143
rect 845 3106 851 3112
rect 957 3088 963 3137
rect 1005 3128 1011 3152
rect 1005 3108 1011 3112
rect 973 2968 979 3092
rect 989 3048 995 3072
rect 1069 3068 1075 3732
rect 1213 3708 1219 3912
rect 1085 3588 1091 3672
rect 1101 3508 1107 3532
rect 1133 3428 1139 3492
rect 1197 3348 1203 3552
rect 1229 3508 1235 3872
rect 1373 3748 1379 4132
rect 1453 3948 1459 4312
rect 1469 4308 1475 4317
rect 1517 4168 1523 4232
rect 1597 4108 1603 4437
rect 1469 3928 1475 3952
rect 1245 3668 1251 3732
rect 1357 3488 1363 3532
rect 1325 3468 1331 3472
rect 1229 3388 1235 3412
rect 1357 3388 1363 3452
rect 1373 3388 1379 3732
rect 1389 3568 1395 3632
rect 1389 3488 1395 3492
rect 1421 3428 1427 3892
rect 1437 3888 1443 3892
rect 1453 3788 1459 3912
rect 1517 3908 1523 3952
rect 1549 3908 1555 3932
rect 1533 3828 1539 3872
rect 1533 3748 1539 3752
rect 1517 3737 1528 3743
rect 1437 3588 1443 3712
rect 1101 3328 1107 3332
rect 1261 3328 1267 3332
rect 1437 3328 1443 3572
rect 1453 3528 1459 3632
rect 1517 3588 1523 3737
rect 1549 3728 1555 3792
rect 1613 3748 1619 4272
rect 1629 4128 1635 4132
rect 1645 4088 1651 4892
rect 1693 4588 1699 4692
rect 1709 4688 1715 4932
rect 1757 4908 1763 4912
rect 1773 4848 1779 5072
rect 1789 5068 1795 5072
rect 1725 4688 1731 4692
rect 1805 4628 1811 5092
rect 1821 4788 1827 4832
rect 1757 4588 1763 4612
rect 1821 4588 1827 4712
rect 1677 4488 1683 4492
rect 1709 4428 1715 4532
rect 1725 4528 1731 4532
rect 1789 4428 1795 4532
rect 1837 4528 1843 5292
rect 1917 5288 1923 5292
rect 1853 5088 1859 5092
rect 1917 5088 1923 5272
rect 1965 5268 1971 5312
rect 1981 5288 1987 5312
rect 2125 5308 2131 5332
rect 2301 5328 2307 5332
rect 2413 5328 2419 5332
rect 2429 5328 2435 5372
rect 3389 5368 3395 5372
rect 2621 5328 2627 5332
rect 2029 5288 2035 5292
rect 2173 5288 2179 5312
rect 1981 5088 1987 5272
rect 1885 5048 1891 5072
rect 1981 5008 1987 5072
rect 2093 5068 2099 5072
rect 2077 4988 2083 5032
rect 1885 4948 1891 4952
rect 1997 4928 2003 4932
rect 2013 4928 2019 4972
rect 1885 4888 1891 4912
rect 2077 4908 2083 4912
rect 1949 4888 1955 4892
rect 2109 4888 2115 5092
rect 2141 5048 2147 5112
rect 2205 5088 2211 5312
rect 2285 5188 2291 5232
rect 2301 5128 2307 5312
rect 2317 5228 2323 5312
rect 2365 5228 2371 5292
rect 2397 5188 2403 5272
rect 2493 5243 2499 5312
rect 2509 5288 2515 5312
rect 2573 5308 2579 5312
rect 2477 5237 2499 5243
rect 2461 5148 2467 5232
rect 2397 5088 2403 5092
rect 2381 5068 2387 5072
rect 2349 5037 2360 5043
rect 2125 4928 2131 4972
rect 2029 4728 2035 4832
rect 1869 4708 1875 4712
rect 1965 4708 1971 4712
rect 1944 4697 1955 4703
rect 1837 4508 1843 4512
rect 1805 4468 1811 4492
rect 1853 4468 1859 4692
rect 1917 4568 1923 4672
rect 1949 4568 1955 4697
rect 1981 4668 1987 4672
rect 1965 4528 1971 4532
rect 1997 4508 2003 4632
rect 2013 4548 2019 4692
rect 2077 4588 2083 4592
rect 2125 4588 2131 4712
rect 2189 4688 2195 4912
rect 2221 4708 2227 5012
rect 2333 4988 2339 5032
rect 2317 4948 2323 4952
rect 2349 4948 2355 5037
rect 2381 5008 2387 5052
rect 2237 4928 2243 4932
rect 2381 4928 2387 4972
rect 2397 4928 2403 5072
rect 2429 4988 2435 5112
rect 2445 5088 2451 5112
rect 2461 5028 2467 5092
rect 2429 4928 2435 4932
rect 2365 4908 2371 4912
rect 2461 4908 2467 4912
rect 2477 4908 2483 5237
rect 2493 4948 2499 5172
rect 2589 5128 2595 5212
rect 2669 5143 2675 5332
rect 2749 5248 2755 5312
rect 2813 5308 2819 5312
rect 2877 5308 2883 5312
rect 2717 5208 2723 5232
rect 2669 5137 2691 5143
rect 2509 5108 2515 5112
rect 2589 5108 2595 5112
rect 2685 5088 2691 5137
rect 2541 5048 2547 5072
rect 2557 4988 2563 5072
rect 2653 5068 2659 5072
rect 2605 5028 2611 5032
rect 2557 4943 2563 4972
rect 2557 4937 2579 4943
rect 2573 4928 2579 4937
rect 2669 4928 2675 4952
rect 2685 4928 2691 5012
rect 2589 4908 2595 4912
rect 2317 4883 2323 4892
rect 2312 4877 2323 4883
rect 2141 4588 2147 4612
rect 2093 4508 2099 4532
rect 2141 4508 2147 4572
rect 1645 3888 1651 3892
rect 1533 3628 1539 3632
rect 1549 3528 1555 3712
rect 1565 3708 1571 3712
rect 1597 3688 1603 3712
rect 1613 3708 1619 3732
rect 1661 3728 1667 4392
rect 1677 4288 1683 4292
rect 1789 4168 1795 4252
rect 1693 4148 1699 4152
rect 1741 4117 1752 4123
rect 1677 4108 1683 4112
rect 1741 3908 1747 4117
rect 1709 3848 1715 3872
rect 1581 3517 1592 3523
rect 1453 3508 1459 3512
rect 1565 3508 1571 3512
rect 1453 3348 1459 3472
rect 1469 3428 1475 3492
rect 1181 3308 1187 3312
rect 1101 3228 1107 3292
rect 1325 3288 1331 3312
rect 1389 3288 1395 3312
rect 1117 3148 1123 3172
rect 1117 3088 1123 3132
rect 1165 3108 1171 3132
rect 1245 3088 1251 3092
rect 1293 3088 1299 3232
rect 1373 3108 1379 3272
rect 1533 3148 1539 3332
rect 1453 3108 1459 3112
rect 1549 3088 1555 3492
rect 1565 3488 1571 3492
rect 1037 2948 1043 2952
rect 1133 2948 1139 2972
rect 1261 2948 1267 3072
rect 1501 2988 1507 3052
rect 1357 2968 1363 2972
rect 781 2928 787 2932
rect 845 2888 851 2892
rect 957 2888 963 2912
rect 1069 2908 1075 2912
rect 1229 2908 1235 2914
rect 1437 2908 1443 2912
rect 749 2788 755 2872
rect 637 2548 643 2612
rect 669 2588 675 2652
rect 717 2588 723 2652
rect 733 2608 739 2712
rect 765 2708 771 2712
rect 765 2688 771 2692
rect 653 2548 659 2552
rect 637 2308 643 2532
rect 685 2508 691 2532
rect 749 2528 755 2632
rect 765 2548 771 2652
rect 781 2588 787 2852
rect 957 2728 963 2732
rect 1149 2728 1155 2732
rect 829 2648 835 2672
rect 669 2348 675 2352
rect 765 2348 771 2532
rect 797 2523 803 2632
rect 877 2588 883 2692
rect 957 2688 963 2712
rect 893 2668 899 2672
rect 893 2588 899 2652
rect 909 2628 915 2632
rect 925 2608 931 2672
rect 829 2548 835 2552
rect 797 2517 808 2523
rect 541 2268 547 2292
rect 669 2288 675 2332
rect 701 2328 707 2332
rect 525 2148 531 2252
rect 397 2088 403 2092
rect 429 1948 435 2132
rect 232 1917 243 1923
rect 237 1908 243 1917
rect 301 1908 307 1932
rect 13 1788 19 1892
rect 125 1868 131 1872
rect 13 1508 19 1532
rect 13 588 19 712
rect 29 528 35 1832
rect 141 1508 147 1892
rect 173 1888 179 1892
rect 221 1868 227 1872
rect 173 1548 179 1732
rect 205 1708 211 1832
rect 237 1728 243 1892
rect 253 1763 259 1832
rect 301 1768 307 1892
rect 349 1788 355 1912
rect 461 1908 467 2132
rect 429 1868 435 1892
rect 381 1788 387 1852
rect 477 1848 483 1892
rect 541 1808 547 1832
rect 557 1828 563 1872
rect 253 1757 275 1763
rect 237 1648 243 1712
rect 253 1588 259 1732
rect 269 1708 275 1757
rect 365 1748 371 1752
rect 477 1748 483 1752
rect 301 1708 307 1712
rect 125 1488 131 1492
rect 173 1488 179 1532
rect 205 1488 211 1492
rect 269 1368 275 1632
rect 317 1588 323 1692
rect 285 1508 291 1512
rect 61 688 67 1332
rect 125 1108 131 1312
rect 205 1308 211 1312
rect 221 1308 227 1312
rect 269 1308 275 1352
rect 285 1308 291 1492
rect 301 1488 307 1572
rect 477 1528 483 1732
rect 589 1723 595 2172
rect 637 2148 643 2232
rect 733 2148 739 2172
rect 653 2108 659 2112
rect 749 2108 755 2312
rect 765 2308 771 2332
rect 781 2328 787 2432
rect 797 2308 803 2352
rect 765 2248 771 2272
rect 765 1948 771 2032
rect 605 1928 611 1932
rect 669 1888 675 1890
rect 637 1768 643 1872
rect 589 1717 600 1723
rect 685 1708 691 1792
rect 701 1788 707 1852
rect 733 1768 739 1812
rect 733 1728 739 1752
rect 765 1748 771 1832
rect 781 1748 787 2292
rect 797 1988 803 2112
rect 813 1948 819 2512
rect 957 2388 963 2632
rect 1005 2628 1011 2652
rect 1037 2568 1043 2652
rect 1101 2588 1107 2692
rect 1117 2688 1123 2692
rect 1149 2688 1155 2712
rect 1245 2688 1251 2692
rect 1325 2688 1331 2872
rect 1389 2788 1395 2832
rect 1469 2808 1475 2932
rect 1485 2908 1491 2952
rect 1581 2948 1587 3517
rect 1597 3508 1603 3512
rect 1613 3128 1619 3632
rect 1661 3548 1667 3712
rect 1677 3688 1683 3752
rect 1709 3728 1715 3752
rect 1741 3688 1747 3892
rect 1757 3668 1763 3712
rect 1677 3528 1683 3532
rect 1656 3517 1667 3523
rect 1661 3503 1667 3517
rect 1661 3497 1683 3503
rect 1677 3488 1683 3497
rect 1645 3388 1651 3392
rect 1661 3143 1667 3472
rect 1773 3383 1779 4132
rect 1821 4128 1827 4132
rect 1837 4128 1843 4372
rect 1981 4308 1987 4492
rect 2173 4468 2179 4512
rect 2189 4508 2195 4512
rect 2093 4308 2099 4452
rect 2205 4448 2211 4672
rect 2237 4588 2243 4692
rect 2301 4548 2307 4872
rect 2237 4528 2243 4532
rect 2301 4508 2307 4532
rect 2301 4443 2307 4492
rect 2285 4437 2307 4443
rect 2125 4388 2131 4432
rect 2221 4348 2227 4432
rect 2221 4308 2227 4312
rect 1992 4297 2003 4303
rect 1853 4268 1859 4290
rect 1885 4228 1891 4272
rect 1901 4148 1907 4172
rect 1965 4168 1971 4272
rect 1901 4128 1907 4132
rect 1917 4128 1923 4152
rect 1869 3928 1875 3932
rect 1917 3908 1923 4092
rect 1805 3888 1811 3892
rect 1821 3828 1827 3832
rect 1821 3748 1827 3812
rect 1853 3808 1859 3892
rect 1933 3883 1939 4152
rect 1997 4148 2003 4297
rect 2093 4268 2099 4292
rect 2013 4228 2019 4232
rect 2013 4188 2019 4212
rect 2061 4208 2067 4232
rect 1965 4128 1971 4132
rect 1949 3988 1955 4032
rect 2045 4028 2051 4112
rect 2093 4108 2099 4112
rect 2093 3948 2099 4092
rect 2125 4048 2131 4232
rect 2221 4208 2227 4292
rect 2157 4148 2163 4152
rect 2205 4148 2211 4172
rect 2157 4048 2163 4132
rect 1965 3908 1971 3912
rect 2029 3888 2035 3890
rect 1928 3877 1939 3883
rect 1821 3608 1827 3632
rect 1837 3508 1843 3712
rect 1885 3703 1891 3832
rect 1901 3828 1907 3872
rect 2029 3848 2035 3852
rect 2029 3748 2035 3832
rect 2093 3828 2099 3832
rect 2093 3788 2099 3812
rect 2125 3788 2131 4032
rect 2237 3908 2243 4272
rect 2253 4248 2259 4292
rect 2269 4288 2275 4332
rect 2269 4128 2275 4172
rect 2285 4108 2291 4437
rect 2317 4408 2323 4692
rect 2349 4688 2355 4692
rect 2365 4648 2371 4672
rect 2397 4588 2403 4892
rect 2413 4728 2419 4832
rect 2413 4668 2419 4712
rect 2445 4588 2451 4692
rect 2349 4528 2355 4532
rect 2317 4308 2323 4392
rect 2365 4388 2371 4532
rect 2429 4388 2435 4512
rect 2365 4308 2371 4372
rect 2445 4368 2451 4532
rect 2461 4528 2467 4692
rect 2493 4688 2499 4712
rect 2541 4703 2547 4832
rect 2701 4808 2707 5012
rect 2717 4948 2723 5192
rect 2733 5088 2739 5092
rect 2749 5028 2755 5232
rect 2781 4988 2787 5232
rect 2845 5128 2851 5232
rect 2845 5083 2851 5112
rect 2845 5077 2856 5083
rect 2813 4928 2819 5032
rect 2797 4908 2803 4912
rect 2605 4708 2611 4752
rect 2621 4717 2632 4723
rect 2541 4697 2552 4703
rect 2509 4588 2515 4612
rect 2525 4563 2531 4692
rect 2541 4668 2547 4697
rect 2573 4668 2579 4672
rect 2589 4668 2595 4672
rect 2509 4557 2531 4563
rect 2477 4488 2483 4492
rect 2461 4308 2467 4312
rect 2301 4168 2307 4232
rect 2317 4228 2323 4292
rect 2317 4088 2323 4112
rect 2157 3848 2163 3892
rect 2141 3837 2152 3843
rect 2141 3748 2147 3837
rect 2253 3828 2259 3892
rect 2269 3848 2275 3892
rect 1901 3728 1907 3732
rect 1885 3697 1896 3703
rect 1933 3508 1939 3512
rect 1981 3508 1987 3732
rect 2109 3648 2115 3692
rect 1789 3488 1795 3492
rect 1981 3468 1987 3492
rect 1757 3377 1779 3383
rect 1757 3368 1763 3377
rect 1757 3348 1763 3352
rect 2013 3348 2019 3532
rect 2045 3488 2051 3532
rect 2061 3488 2067 3532
rect 2125 3508 2131 3512
rect 2253 3508 2259 3512
rect 2109 3388 2115 3452
rect 2061 3348 2067 3372
rect 1693 3328 1699 3332
rect 1741 3308 1747 3312
rect 1661 3137 1683 3143
rect 1613 3108 1619 3112
rect 1597 2948 1603 3072
rect 1661 3063 1667 3092
rect 1677 3088 1683 3137
rect 1693 3128 1699 3292
rect 1821 3148 1827 3332
rect 1709 3108 1715 3112
rect 1741 3108 1747 3112
rect 1773 3088 1779 3132
rect 1805 3088 1811 3090
rect 1661 3057 1683 3063
rect 1437 2788 1443 2792
rect 1341 2708 1347 2772
rect 1117 2568 1123 2612
rect 1149 2548 1155 2652
rect 1213 2648 1219 2676
rect 1165 2528 1171 2572
rect 1197 2568 1203 2612
rect 1453 2608 1459 2672
rect 1277 2528 1283 2532
rect 1389 2528 1395 2572
rect 909 2328 915 2332
rect 957 2308 963 2332
rect 845 2268 851 2272
rect 861 2188 867 2292
rect 877 2183 883 2272
rect 877 2177 888 2183
rect 877 2143 883 2177
rect 861 2137 883 2143
rect 861 2128 867 2137
rect 925 2128 931 2232
rect 973 2228 979 2272
rect 1117 2268 1123 2292
rect 1053 2148 1059 2172
rect 1149 2128 1155 2372
rect 1165 2288 1171 2492
rect 1181 2328 1187 2332
rect 1261 2308 1267 2412
rect 1309 2308 1315 2312
rect 877 2088 883 2112
rect 845 1948 851 2032
rect 861 1923 867 2032
rect 1101 2008 1107 2032
rect 1037 1928 1043 1992
rect 1101 1948 1107 1952
rect 856 1917 867 1923
rect 813 1888 819 1912
rect 925 1888 931 1912
rect 1021 1888 1027 1892
rect 925 1788 931 1852
rect 1021 1848 1027 1872
rect 1037 1808 1043 1912
rect 1101 1908 1107 1932
rect 1085 1888 1091 1892
rect 1165 1888 1171 2272
rect 1213 2268 1219 2292
rect 1229 2268 1235 2272
rect 1181 2168 1187 2232
rect 1181 2108 1187 2112
rect 1213 1948 1219 2032
rect 941 1748 947 1752
rect 749 1728 755 1732
rect 861 1728 867 1732
rect 605 1548 611 1632
rect 621 1568 627 1572
rect 573 1528 579 1532
rect 429 1488 435 1492
rect 477 1488 483 1512
rect 621 1508 627 1552
rect 749 1508 755 1512
rect 829 1508 835 1672
rect 301 1348 307 1372
rect 525 1368 531 1432
rect 541 1388 547 1432
rect 365 1337 376 1343
rect 285 1123 291 1292
rect 280 1117 291 1123
rect 205 1108 211 1112
rect 221 1108 227 1112
rect 125 1088 131 1092
rect 301 1088 307 1132
rect 333 1108 339 1232
rect 365 1188 371 1337
rect 413 1308 419 1352
rect 461 1328 467 1352
rect 125 928 131 1072
rect 205 1068 211 1072
rect 397 1068 403 1272
rect 445 1106 451 1312
rect 477 1288 483 1332
rect 493 1268 499 1332
rect 509 1308 515 1312
rect 605 1308 611 1332
rect 621 1188 627 1452
rect 685 1448 691 1490
rect 877 1468 883 1732
rect 957 1728 963 1792
rect 989 1728 995 1732
rect 893 1508 899 1712
rect 1021 1528 1027 1732
rect 1053 1708 1059 1832
rect 1069 1788 1075 1872
rect 1085 1848 1091 1872
rect 1181 1828 1187 1912
rect 1229 1908 1235 2252
rect 1261 2188 1267 2292
rect 1325 2288 1331 2512
rect 1309 2188 1315 2272
rect 1405 2268 1411 2532
rect 1501 2528 1507 2532
rect 1517 2528 1523 2932
rect 1533 2788 1539 2912
rect 1565 2708 1571 2732
rect 1581 2548 1587 2932
rect 1645 2908 1651 2932
rect 1661 2908 1667 2912
rect 1677 2888 1683 3057
rect 1693 2948 1699 2952
rect 1773 2948 1779 3072
rect 1917 2988 1923 3112
rect 1933 3048 1939 3072
rect 1965 2988 1971 3132
rect 1997 3128 2003 3312
rect 2077 3308 2083 3312
rect 2077 3288 2083 3292
rect 2125 3268 2131 3492
rect 2157 3488 2163 3492
rect 2285 3463 2291 4032
rect 2333 3528 2339 4292
rect 2397 4168 2403 4192
rect 2413 4188 2419 4272
rect 2461 4148 2467 4152
rect 2429 4088 2435 4112
rect 2429 3988 2435 4012
rect 2477 3928 2483 4472
rect 2509 4248 2515 4557
rect 2557 4548 2563 4552
rect 2541 4468 2547 4492
rect 2493 4108 2499 4112
rect 2349 3888 2355 3892
rect 2429 3888 2435 3892
rect 2445 3888 2451 3892
rect 2461 3888 2467 3892
rect 2429 3868 2435 3872
rect 2541 3868 2547 3892
rect 2557 3888 2563 4532
rect 2605 4528 2611 4692
rect 2621 4628 2627 4717
rect 2685 4708 2691 4712
rect 2701 4708 2707 4792
rect 2653 4648 2659 4652
rect 2685 4588 2691 4652
rect 2733 4568 2739 4812
rect 2781 4708 2787 4812
rect 2797 4748 2803 4892
rect 2877 4888 2883 5092
rect 2909 4988 2915 5112
rect 2893 4888 2899 4892
rect 2829 4688 2835 4832
rect 2845 4708 2851 4712
rect 2909 4688 2915 4952
rect 2925 4928 2931 4932
rect 2941 4788 2947 5312
rect 3021 5028 3027 5312
rect 3149 5183 3155 5312
rect 3309 5288 3315 5312
rect 3149 5177 3171 5183
rect 3117 5068 3123 5072
rect 3037 5008 3043 5052
rect 2957 4988 2963 4992
rect 3037 4988 3043 4992
rect 3101 4928 3107 5032
rect 3117 4988 3123 5032
rect 2989 4888 2995 4912
rect 3085 4908 3091 4912
rect 2749 4568 2755 4672
rect 2829 4583 2835 4672
rect 2877 4648 2883 4652
rect 2877 4588 2883 4612
rect 2813 4577 2835 4583
rect 2621 4548 2627 4552
rect 2781 4528 2787 4572
rect 2813 4568 2819 4577
rect 2829 4548 2835 4552
rect 2925 4548 2931 4592
rect 2941 4548 2947 4632
rect 2957 4628 2963 4692
rect 2589 4308 2595 4352
rect 2589 4288 2595 4292
rect 2584 4237 2595 4243
rect 2573 3908 2579 4212
rect 2589 4168 2595 4237
rect 2605 4108 2611 4292
rect 2621 4088 2627 4512
rect 2669 4508 2675 4512
rect 2829 4408 2835 4532
rect 2845 4448 2851 4512
rect 2957 4508 2963 4512
rect 2893 4448 2899 4492
rect 2637 4188 2643 4312
rect 2637 4128 2643 4132
rect 2669 4128 2675 4232
rect 2749 4188 2755 4192
rect 2381 3748 2387 3772
rect 2525 3748 2531 3812
rect 2557 3808 2563 3872
rect 2573 3828 2579 3892
rect 2589 3888 2595 4072
rect 2605 3868 2611 3952
rect 2621 3908 2627 4072
rect 2653 3988 2659 4112
rect 2733 4103 2739 4112
rect 2712 4097 2739 4103
rect 2765 4028 2771 4152
rect 2781 4148 2787 4152
rect 2813 4148 2819 4292
rect 2909 4288 2915 4292
rect 2829 4148 2835 4232
rect 2797 4108 2803 4112
rect 2925 4108 2931 4432
rect 2957 4188 2963 4272
rect 2957 4148 2963 4152
rect 2989 4088 2995 4872
rect 3005 4568 3011 4672
rect 3037 4648 3043 4832
rect 3133 4708 3139 4732
rect 3149 4723 3155 5032
rect 3165 4928 3171 5177
rect 3357 5128 3363 5332
rect 3469 5263 3475 5463
rect 3517 5368 3523 5463
rect 3517 5348 3523 5352
rect 3581 5348 3587 5372
rect 3629 5348 3635 5463
rect 3485 5308 3491 5312
rect 3533 5308 3539 5332
rect 3565 5308 3571 5312
rect 3597 5308 3603 5312
rect 3485 5288 3491 5292
rect 3597 5288 3603 5292
rect 3469 5257 3491 5263
rect 3309 5048 3315 5092
rect 3357 5088 3363 5112
rect 3389 5108 3395 5232
rect 3197 4948 3203 5032
rect 3229 4948 3235 4952
rect 3277 4928 3283 4932
rect 3229 4788 3235 4852
rect 3213 4728 3219 4752
rect 3341 4748 3347 4832
rect 3373 4788 3379 5012
rect 3405 4803 3411 5232
rect 3485 5188 3491 5257
rect 3421 4968 3427 5032
rect 3405 4797 3427 4803
rect 3421 4768 3427 4797
rect 3149 4717 3160 4723
rect 3069 4608 3075 4632
rect 3037 4548 3043 4572
rect 3069 4548 3075 4552
rect 3005 4528 3011 4532
rect 3005 4308 3011 4492
rect 3197 4468 3203 4632
rect 3037 4328 3043 4332
rect 3037 4288 3043 4312
rect 3069 4308 3075 4312
rect 3117 4288 3123 4292
rect 3133 4288 3139 4392
rect 3053 4228 3059 4252
rect 3133 4248 3139 4272
rect 3149 4268 3155 4312
rect 3213 4308 3219 4692
rect 3229 4628 3235 4692
rect 3277 4688 3283 4692
rect 3277 4668 3283 4672
rect 3277 4548 3283 4632
rect 3293 4548 3299 4632
rect 3261 4328 3267 4532
rect 3341 4508 3347 4512
rect 3341 4448 3347 4492
rect 3405 4428 3411 4692
rect 3421 4648 3427 4732
rect 3453 4708 3459 5092
rect 3512 5037 3523 5043
rect 3501 4968 3507 4972
rect 3501 4948 3507 4952
rect 3517 4948 3523 5037
rect 3613 4988 3619 5092
rect 3661 5088 3667 5112
rect 3693 5088 3699 5092
rect 3549 4948 3555 4952
rect 3661 4948 3667 4992
rect 3709 4988 3715 5463
rect 3725 5188 3731 5232
rect 3741 5128 3747 5312
rect 3757 5248 3763 5463
rect 3853 5457 3875 5463
rect 3773 5188 3779 5272
rect 3805 5128 3811 5372
rect 3837 5328 3843 5332
rect 3869 5283 3875 5457
rect 3933 5428 3939 5463
rect 3853 5277 3875 5283
rect 3853 5188 3859 5277
rect 3901 5188 3907 5412
rect 3965 5328 3971 5332
rect 3981 5188 3987 5463
rect 4013 5457 4035 5463
rect 4013 5388 4019 5457
rect 4349 5388 4355 5463
rect 4077 5328 4083 5332
rect 3997 5268 4003 5312
rect 3741 5068 3747 5092
rect 3485 4908 3491 4912
rect 3517 4908 3523 4932
rect 3501 4708 3507 4792
rect 3533 4728 3539 4832
rect 3549 4808 3555 4932
rect 3613 4788 3619 4912
rect 3645 4908 3651 4912
rect 3645 4788 3651 4892
rect 3677 4828 3683 4912
rect 3725 4868 3731 4932
rect 3789 4928 3795 5072
rect 3821 5008 3827 5032
rect 3837 4968 3843 5072
rect 3885 4948 3891 4952
rect 3549 4728 3555 4752
rect 3693 4748 3699 4852
rect 3725 4788 3731 4812
rect 3693 4728 3699 4732
rect 3709 4708 3715 4712
rect 3501 4668 3507 4692
rect 3613 4688 3619 4692
rect 3453 4588 3459 4652
rect 3501 4508 3507 4512
rect 3341 4308 3347 4312
rect 3037 4128 3043 4132
rect 3053 4128 3059 4212
rect 3165 4148 3171 4172
rect 3261 4168 3267 4232
rect 3213 4108 3219 4112
rect 3293 4088 3299 4272
rect 3405 4148 3411 4172
rect 3437 4148 3443 4412
rect 3469 4368 3475 4412
rect 3469 4288 3475 4352
rect 3485 4288 3491 4292
rect 3517 4228 3523 4672
rect 3581 4668 3587 4672
rect 3565 4588 3571 4632
rect 3549 4528 3555 4532
rect 3581 4408 3587 4512
rect 3629 4388 3635 4692
rect 3725 4688 3731 4692
rect 3645 4677 3656 4683
rect 3645 4548 3651 4677
rect 3645 4368 3651 4532
rect 3661 4528 3667 4532
rect 3533 4308 3539 4312
rect 3565 4288 3571 4332
rect 3629 4288 3635 4292
rect 3496 4157 3507 4163
rect 3437 4108 3443 4112
rect 2557 3748 2563 3752
rect 2397 3708 2403 3712
rect 2493 3708 2499 3732
rect 2525 3728 2531 3732
rect 2493 3688 2499 3692
rect 2301 3508 2307 3512
rect 2381 3508 2387 3512
rect 2397 3508 2403 3512
rect 2333 3488 2339 3492
rect 2285 3457 2307 3463
rect 2141 3368 2147 3392
rect 2221 3388 2227 3412
rect 2269 3388 2275 3452
rect 2301 3388 2307 3457
rect 2333 3428 2339 3472
rect 2429 3468 2435 3472
rect 2461 3348 2467 3352
rect 2253 3328 2259 3332
rect 2269 3288 2275 3312
rect 2285 3308 2291 3332
rect 2477 3328 2483 3412
rect 2509 3388 2515 3412
rect 2525 3348 2531 3712
rect 2621 3688 2627 3892
rect 2653 3868 2659 3972
rect 2813 3917 2824 3923
rect 2701 3868 2707 3872
rect 2781 3788 2787 3872
rect 2797 3748 2803 3752
rect 2557 3348 2563 3432
rect 2605 3388 2611 3512
rect 2525 3328 2531 3332
rect 2349 3308 2355 3312
rect 2557 3308 2563 3332
rect 2621 3328 2627 3332
rect 2637 3308 2643 3492
rect 2653 3388 2659 3732
rect 2813 3728 2819 3917
rect 2893 3908 2899 4072
rect 2973 3968 2979 4032
rect 2973 3908 2979 3912
rect 2669 3708 2675 3712
rect 2829 3703 2835 3832
rect 2861 3788 2867 3832
rect 2957 3748 2963 3852
rect 3005 3768 3011 4032
rect 3085 3863 3091 4032
rect 3277 3928 3283 3972
rect 3293 3943 3299 4072
rect 3325 3988 3331 4032
rect 3293 3937 3315 3943
rect 3165 3908 3171 3912
rect 3101 3888 3107 3892
rect 3085 3857 3107 3863
rect 2829 3697 2840 3703
rect 2669 3488 2675 3552
rect 2685 3488 2691 3492
rect 2717 3443 2723 3512
rect 2749 3488 2755 3672
rect 2717 3437 2739 3443
rect 2733 3388 2739 3437
rect 2765 3348 2771 3392
rect 2781 3368 2787 3632
rect 2877 3548 2883 3732
rect 2925 3728 2931 3732
rect 2957 3488 2963 3732
rect 3005 3568 3011 3752
rect 3101 3748 3107 3857
rect 3101 3648 3107 3732
rect 3117 3728 3123 3892
rect 3309 3888 3315 3937
rect 3197 3848 3203 3872
rect 3149 3748 3155 3772
rect 3245 3728 3251 3872
rect 3021 3528 3027 3532
rect 3165 3506 3171 3532
rect 2973 3488 2979 3492
rect 2813 3388 2819 3452
rect 2893 3368 2899 3432
rect 2909 3408 2915 3432
rect 2957 3368 2963 3472
rect 2685 3328 2691 3332
rect 2013 3188 2019 3212
rect 2141 3128 2147 3132
rect 2189 3128 2195 3252
rect 1885 2968 1891 2972
rect 1757 2908 1763 2914
rect 1709 2788 1715 2872
rect 1613 2528 1619 2772
rect 1853 2748 1859 2752
rect 1741 2688 1747 2692
rect 1757 2688 1763 2712
rect 1773 2708 1779 2712
rect 1421 2508 1427 2512
rect 1421 2288 1427 2332
rect 1437 2308 1443 2432
rect 1469 2288 1475 2452
rect 1517 2428 1523 2512
rect 1581 2468 1587 2512
rect 1517 2328 1523 2332
rect 1533 2288 1539 2312
rect 1549 2268 1555 2432
rect 1709 2348 1715 2632
rect 1741 2548 1747 2592
rect 1581 2308 1587 2332
rect 1325 2248 1331 2252
rect 1325 2188 1331 2232
rect 1421 2188 1427 2192
rect 1293 2128 1299 2132
rect 1309 2083 1315 2172
rect 1437 2128 1443 2152
rect 1453 2148 1459 2232
rect 1501 2128 1507 2152
rect 1533 2128 1539 2152
rect 1549 2148 1555 2252
rect 1581 2188 1587 2272
rect 1597 2268 1603 2272
rect 1629 2248 1635 2292
rect 1677 2288 1683 2332
rect 1597 2188 1603 2232
rect 1613 2128 1619 2132
rect 1293 2077 1315 2083
rect 1261 1928 1267 2032
rect 1213 1868 1219 1872
rect 1229 1848 1235 1892
rect 1085 1528 1091 1792
rect 1293 1748 1299 2077
rect 1309 1908 1315 1952
rect 1421 1908 1427 2072
rect 1533 2028 1539 2112
rect 1565 2048 1571 2112
rect 1629 2108 1635 2112
rect 1693 2068 1699 2112
rect 1517 1908 1523 1932
rect 1597 1908 1603 2052
rect 1661 2008 1667 2032
rect 1325 1868 1331 1872
rect 1165 1528 1171 1692
rect 1037 1508 1043 1512
rect 685 1328 691 1372
rect 733 1328 739 1332
rect 749 1328 755 1372
rect 813 1348 819 1432
rect 525 1108 531 1132
rect 573 1108 579 1172
rect 189 968 195 972
rect 205 948 211 1052
rect 301 948 307 952
rect 365 928 371 992
rect 125 688 131 912
rect 221 908 227 912
rect 141 708 147 712
rect 221 708 227 892
rect 45 548 51 632
rect 61 563 67 672
rect 61 557 83 563
rect 77 528 83 557
rect 173 548 179 552
rect 61 168 67 252
rect 77 128 83 432
rect 125 328 131 472
rect 205 348 211 572
rect 237 508 243 692
rect 349 608 355 672
rect 253 508 259 512
rect 125 288 131 292
rect 189 188 195 312
rect 205 288 211 332
rect 237 328 243 492
rect 237 288 243 292
rect 269 288 275 532
rect 301 528 307 592
rect 381 563 387 1052
rect 477 968 483 1072
rect 429 668 435 932
rect 509 928 515 1092
rect 637 1088 643 1092
rect 525 988 531 992
rect 589 988 595 1012
rect 637 988 643 1072
rect 653 1068 659 1092
rect 509 897 520 903
rect 445 728 451 732
rect 461 708 467 752
rect 477 708 483 712
rect 381 557 403 563
rect 397 528 403 557
rect 381 388 387 452
rect 429 388 435 652
rect 317 328 323 372
rect 317 308 323 312
rect 269 148 275 272
rect 317 108 323 232
rect 365 183 371 252
rect 365 177 376 183
rect 413 163 419 372
rect 413 157 435 163
rect 429 128 435 157
rect 445 148 451 372
rect 461 288 467 592
rect 493 568 499 692
rect 509 588 515 897
rect 541 703 547 932
rect 573 708 579 972
rect 589 883 595 892
rect 589 877 611 883
rect 605 788 611 877
rect 637 708 643 912
rect 653 788 659 932
rect 525 697 547 703
rect 493 548 499 552
rect 493 528 499 532
rect 477 508 483 512
rect 509 488 515 492
rect 525 468 531 697
rect 541 548 547 552
rect 557 508 563 692
rect 573 688 579 692
rect 573 588 579 612
rect 589 568 595 692
rect 621 688 627 692
rect 637 648 643 652
rect 685 608 691 672
rect 589 548 595 552
rect 477 308 483 332
rect 541 328 547 492
rect 589 308 595 532
rect 653 528 659 532
rect 637 508 643 512
rect 669 488 675 492
rect 605 388 611 472
rect 621 328 627 372
rect 685 348 691 512
rect 701 328 707 1152
rect 717 1048 723 1232
rect 813 1068 819 1092
rect 829 1068 835 1332
rect 717 928 723 972
rect 749 948 755 952
rect 829 948 835 1052
rect 861 1008 867 1432
rect 893 1428 899 1492
rect 957 1488 963 1492
rect 1085 1488 1091 1492
rect 941 1368 947 1372
rect 957 1308 963 1312
rect 973 1308 979 1312
rect 989 1308 995 1432
rect 893 1108 899 1112
rect 989 1108 995 1292
rect 925 1068 931 1092
rect 717 708 723 912
rect 925 908 931 912
rect 941 908 947 912
rect 813 708 819 732
rect 589 288 595 292
rect 733 288 739 332
rect 765 308 771 312
rect 829 308 835 892
rect 909 728 915 732
rect 925 688 931 832
rect 909 588 915 672
rect 941 668 947 692
rect 957 648 963 1092
rect 1005 1068 1011 1472
rect 1149 1448 1155 1472
rect 1053 1348 1059 1352
rect 1069 1288 1075 1332
rect 1085 1328 1091 1392
rect 1133 1308 1139 1432
rect 1165 1408 1171 1512
rect 1197 1408 1203 1472
rect 1229 1348 1235 1472
rect 1229 1188 1235 1292
rect 1165 1103 1171 1132
rect 1165 1097 1176 1103
rect 1037 1088 1043 1092
rect 1197 1088 1203 1092
rect 1021 1068 1027 1072
rect 973 768 979 932
rect 989 908 995 992
rect 1021 948 1027 972
rect 989 768 995 892
rect 957 528 963 632
rect 973 548 979 752
rect 1021 748 1027 932
rect 1037 928 1043 1072
rect 1053 1043 1059 1072
rect 1069 1068 1075 1072
rect 1053 1037 1075 1043
rect 989 668 995 712
rect 1021 688 1027 712
rect 1037 708 1043 912
rect 1069 903 1075 1037
rect 1165 948 1171 1072
rect 1181 948 1187 1032
rect 1197 948 1203 972
rect 1149 928 1155 932
rect 1181 928 1187 932
rect 1213 908 1219 1032
rect 1229 948 1235 1172
rect 1293 1088 1299 1152
rect 1309 1148 1315 1812
rect 1341 1788 1347 1892
rect 1341 1688 1347 1712
rect 1325 1508 1331 1672
rect 1405 1508 1411 1512
rect 1405 1488 1411 1492
rect 1341 1388 1347 1392
rect 1373 1328 1379 1432
rect 1421 1388 1427 1892
rect 1437 1888 1443 1892
rect 1437 1808 1443 1872
rect 1453 1728 1459 1732
rect 1485 1728 1491 1832
rect 1565 1828 1571 1832
rect 1517 1748 1523 1812
rect 1501 1708 1507 1712
rect 1549 1688 1555 1732
rect 1501 1588 1507 1672
rect 1437 1388 1443 1432
rect 1421 1363 1427 1372
rect 1421 1357 1443 1363
rect 1437 1328 1443 1357
rect 1453 1348 1459 1552
rect 1469 1428 1475 1492
rect 1533 1448 1539 1472
rect 1469 1328 1475 1372
rect 1517 1308 1523 1372
rect 1533 1328 1539 1432
rect 1549 1348 1555 1372
rect 1565 1368 1571 1392
rect 1597 1388 1603 1652
rect 1629 1528 1635 1932
rect 1709 1908 1715 2292
rect 1725 2248 1731 2532
rect 1773 2508 1779 2652
rect 1757 2428 1763 2432
rect 1725 2188 1731 2212
rect 1757 2143 1763 2252
rect 1789 2228 1795 2532
rect 1805 2528 1811 2532
rect 1805 2508 1811 2512
rect 1821 2448 1827 2712
rect 1853 2688 1859 2732
rect 1869 2688 1875 2692
rect 1901 2688 1907 2712
rect 1933 2648 1939 2676
rect 1949 2628 1955 2912
rect 1965 2908 1971 2952
rect 1997 2788 2003 3072
rect 2013 2948 2019 3092
rect 2045 3068 2051 3112
rect 2061 3068 2067 3072
rect 2077 3048 2083 3112
rect 2221 3108 2227 3232
rect 2285 3108 2291 3292
rect 2349 3268 2355 3292
rect 2381 3268 2387 3292
rect 2349 3106 2355 3232
rect 2141 3037 2152 3043
rect 2077 2948 2083 3032
rect 2029 2928 2035 2932
rect 2077 2908 2083 2912
rect 2141 2908 2147 3037
rect 2237 2988 2243 3072
rect 2253 2948 2259 3032
rect 2061 2768 2067 2772
rect 2077 2768 2083 2892
rect 2173 2788 2179 2832
rect 1981 2668 1987 2732
rect 2013 2668 2019 2672
rect 1853 2528 1859 2532
rect 1885 2488 1891 2532
rect 2013 2508 2019 2652
rect 2029 2648 2035 2692
rect 2061 2548 2067 2652
rect 2077 2608 2083 2672
rect 2077 2588 2083 2592
rect 2093 2548 2099 2692
rect 2109 2688 2115 2712
rect 2125 2588 2131 2752
rect 2269 2708 2275 2912
rect 2317 2888 2323 3072
rect 2381 2988 2387 3232
rect 2493 3128 2499 3292
rect 2509 3188 2515 3252
rect 2717 3188 2723 3292
rect 2733 3248 2739 3292
rect 2397 2948 2403 3092
rect 2429 2988 2435 3012
rect 2493 2988 2499 3112
rect 2525 3088 2531 3132
rect 2557 2948 2563 3072
rect 2717 3048 2723 3052
rect 2733 2988 2739 3112
rect 2765 3108 2771 3232
rect 2797 3208 2803 3232
rect 2605 2928 2611 2952
rect 2717 2948 2723 2972
rect 2749 2968 2755 3072
rect 2797 3068 2803 3072
rect 2813 3043 2819 3292
rect 2845 3168 2851 3312
rect 2829 3108 2835 3112
rect 2797 3037 2819 3043
rect 2797 2988 2803 3037
rect 2845 2968 2851 3152
rect 2909 3128 2915 3132
rect 2877 3088 2883 3092
rect 2893 3088 2899 3092
rect 2813 2948 2819 2952
rect 2877 2948 2883 3072
rect 2909 2988 2915 3092
rect 2941 3088 2947 3152
rect 2957 3108 2963 3332
rect 2973 3328 2979 3352
rect 2989 3308 2995 3492
rect 3101 3488 3107 3492
rect 3229 3488 3235 3552
rect 3101 3388 3107 3392
rect 3181 3368 3187 3372
rect 3133 3308 3139 3312
rect 3245 3308 3251 3712
rect 3277 3708 3283 3832
rect 3293 3768 3299 3832
rect 3325 3748 3331 3752
rect 3325 3728 3331 3732
rect 3341 3728 3347 3752
rect 3261 3488 3267 3632
rect 3309 3548 3315 3632
rect 3325 3528 3331 3692
rect 3341 3588 3347 3672
rect 3357 3548 3363 3792
rect 3373 3788 3379 3892
rect 3389 3708 3395 3752
rect 3437 3743 3443 3852
rect 3432 3737 3443 3743
rect 3389 3668 3395 3692
rect 3261 3348 3267 3472
rect 3277 3408 3283 3492
rect 3309 3488 3315 3512
rect 3341 3348 3347 3432
rect 3357 3388 3363 3472
rect 3405 3448 3411 3512
rect 3421 3488 3427 3712
rect 3437 3588 3443 3712
rect 3437 3408 3443 3492
rect 3261 3308 3267 3312
rect 3373 3308 3379 3392
rect 3453 3388 3459 3812
rect 3469 3788 3475 3852
rect 3469 3388 3475 3632
rect 3485 3488 3491 3492
rect 3501 3408 3507 4157
rect 3517 4128 3523 4212
rect 3645 4208 3651 4332
rect 3645 4168 3651 4172
rect 3565 4128 3571 4132
rect 3645 4128 3651 4152
rect 3661 4128 3667 4432
rect 3677 4328 3683 4572
rect 3693 4508 3699 4632
rect 3725 4588 3731 4652
rect 3741 4588 3747 4732
rect 3757 4708 3763 4912
rect 3789 4908 3795 4912
rect 3933 4888 3939 5092
rect 3981 4968 3987 4972
rect 3981 4928 3987 4952
rect 4045 4908 4051 5312
rect 4061 5108 4067 5132
rect 4077 5088 4083 5312
rect 4125 5308 4131 5312
rect 4221 5108 4227 5232
rect 4301 5108 4307 5232
rect 4333 5188 4339 5292
rect 4109 4968 4115 5072
rect 4221 5048 4227 5092
rect 4173 4948 4179 4952
rect 4301 4948 4307 5072
rect 4317 4928 4323 5052
rect 4205 4908 4211 4912
rect 3917 4868 3923 4872
rect 4205 4843 4211 4892
rect 4189 4837 4211 4843
rect 3789 4528 3795 4532
rect 3725 4508 3731 4512
rect 3709 4488 3715 4492
rect 3741 4468 3747 4472
rect 3725 4288 3731 4352
rect 3757 4308 3763 4432
rect 3661 4108 3667 4112
rect 3613 3988 3619 4052
rect 3629 3988 3635 4092
rect 3565 3888 3571 3892
rect 3517 3688 3523 3832
rect 3565 3748 3571 3752
rect 3549 3648 3555 3692
rect 3581 3628 3587 3872
rect 3597 3788 3603 3852
rect 3629 3708 3635 3972
rect 3645 3928 3651 4032
rect 3661 3848 3667 4072
rect 3677 3908 3683 4232
rect 3709 4188 3715 4272
rect 3741 4248 3747 4272
rect 3757 4248 3763 4292
rect 3805 4248 3811 4312
rect 3821 4188 3827 4612
rect 3869 4348 3875 4832
rect 3885 4348 3891 4512
rect 3917 4488 3923 4672
rect 4045 4588 4051 4690
rect 4061 4548 4067 4552
rect 4173 4548 4179 4632
rect 3837 4308 3843 4332
rect 3837 4288 3843 4292
rect 3949 4263 3955 4492
rect 3965 4288 3971 4292
rect 3949 4257 3971 4263
rect 3693 3888 3699 4132
rect 3725 4128 3731 4152
rect 3773 4128 3779 4172
rect 3816 4157 3827 4163
rect 3725 3988 3731 4052
rect 3757 4048 3763 4072
rect 3773 3923 3779 4032
rect 3789 4028 3795 4092
rect 3768 3917 3779 3923
rect 3821 3863 3827 4157
rect 3837 4157 3891 4163
rect 3837 4128 3843 4157
rect 3885 4148 3891 4157
rect 3853 4128 3859 4132
rect 3933 4128 3939 4212
rect 3869 4108 3875 4112
rect 3837 3948 3843 4032
rect 3853 3988 3859 4072
rect 3805 3857 3827 3863
rect 3709 3788 3715 3852
rect 3677 3748 3683 3752
rect 3549 3588 3555 3612
rect 3597 3608 3603 3692
rect 3661 3688 3667 3692
rect 3581 3488 3587 3552
rect 3677 3508 3683 3672
rect 3709 3628 3715 3692
rect 3741 3688 3747 3832
rect 3789 3748 3795 3752
rect 3757 3728 3763 3732
rect 3773 3648 3779 3692
rect 3773 3588 3779 3612
rect 3741 3448 3747 3472
rect 3757 3468 3763 3512
rect 3773 3508 3779 3532
rect 3789 3508 3795 3532
rect 3789 3383 3795 3492
rect 3805 3388 3811 3857
rect 3821 3588 3827 3692
rect 3837 3628 3843 3932
rect 3869 3928 3875 4012
rect 3917 3988 3923 4092
rect 3933 4028 3939 4092
rect 3949 4048 3955 4072
rect 3965 3988 3971 4257
rect 3981 4188 3987 4432
rect 3997 4428 4003 4532
rect 4013 4508 4019 4512
rect 4045 4508 4051 4532
rect 4173 4528 4179 4532
rect 4061 4508 4067 4512
rect 4077 4508 4083 4512
rect 4109 4508 4115 4512
rect 4125 4488 4131 4492
rect 4189 4488 4195 4837
rect 4237 4788 4243 4892
rect 4317 4728 4323 4732
rect 4333 4728 4339 5072
rect 4365 4948 4371 5092
rect 4429 5083 4435 5312
rect 4445 5108 4451 5112
rect 4461 5083 4467 5463
rect 4509 5428 4515 5463
rect 4541 5428 4547 5463
rect 4557 5348 4563 5372
rect 4637 5348 4643 5372
rect 4685 5348 4691 5463
rect 4733 5428 4739 5463
rect 4797 5428 4803 5463
rect 4845 5408 4851 5463
rect 4941 5428 4947 5463
rect 5325 5428 5331 5463
rect 5373 5428 5379 5463
rect 5437 5408 5443 5463
rect 5533 5348 5539 5352
rect 5581 5348 5587 5352
rect 5917 5348 5923 5463
rect 6029 5348 6035 5463
rect 6125 5348 6131 5352
rect 6189 5348 6195 5372
rect 6040 5337 6051 5343
rect 4493 5308 4499 5314
rect 4493 5148 4499 5272
rect 4525 5248 4531 5332
rect 4589 5308 4595 5312
rect 4653 5308 4659 5312
rect 4477 5108 4483 5112
rect 4493 5088 4499 5132
rect 4429 5077 4451 5083
rect 4461 5077 4483 5083
rect 4381 4948 4387 4992
rect 4429 4988 4435 5052
rect 4365 4908 4371 4932
rect 4253 4548 4259 4592
rect 4285 4548 4291 4672
rect 4061 4388 4067 4472
rect 4077 4328 4083 4332
rect 4013 4268 4019 4272
rect 3853 3908 3859 3912
rect 3901 3848 3907 3932
rect 3933 3928 3939 3972
rect 4013 3968 4019 4232
rect 4061 4188 4067 4292
rect 4109 4288 4115 4412
rect 4269 4368 4275 4532
rect 4301 4528 4307 4612
rect 4301 4388 4307 4432
rect 4173 4308 4179 4312
rect 4125 4288 4131 4292
rect 4205 4288 4211 4312
rect 4301 4288 4307 4290
rect 4269 4268 4275 4272
rect 4029 4108 4035 4112
rect 3917 3908 3923 3912
rect 3981 3908 3987 3932
rect 4013 3908 4019 3952
rect 3997 3868 4003 3872
rect 3960 3857 3971 3863
rect 3853 3788 3859 3792
rect 3901 3788 3907 3832
rect 3965 3788 3971 3857
rect 4045 3863 4051 4152
rect 4141 4128 4147 4132
rect 4125 4108 4131 4112
rect 4093 4088 4099 4092
rect 4061 3928 4067 3952
rect 4061 3888 4067 3892
rect 4093 3888 4099 3912
rect 4045 3857 4067 3863
rect 3997 3788 4003 3812
rect 4061 3788 4067 3857
rect 4157 3748 4163 4132
rect 4173 3968 4179 4032
rect 4205 4008 4211 4112
rect 4253 4108 4259 4172
rect 4221 3868 4227 3892
rect 4269 3868 4275 4252
rect 4285 4108 4291 4112
rect 4317 3948 4323 4632
rect 4333 4508 4339 4632
rect 4365 4548 4371 4672
rect 4381 4608 4387 4932
rect 4413 4728 4419 4812
rect 4445 4788 4451 5077
rect 4461 4908 4467 4912
rect 4461 4728 4467 4732
rect 4429 4708 4435 4712
rect 4477 4703 4483 5077
rect 4493 4943 4499 5072
rect 4653 5068 4659 5092
rect 4509 4968 4515 5032
rect 4701 5008 4707 5312
rect 4781 5308 4787 5312
rect 4813 5308 4819 5312
rect 4749 5128 4755 5292
rect 4781 5108 4787 5252
rect 4829 5128 4835 5312
rect 4909 5308 4915 5314
rect 4973 5268 4979 5312
rect 4973 5248 4979 5252
rect 4829 5108 4835 5112
rect 4877 5108 4883 5112
rect 4605 4968 4611 4972
rect 4733 4968 4739 5072
rect 4781 5048 4787 5092
rect 4797 5068 4803 5072
rect 4797 4948 4803 4952
rect 4493 4937 4504 4943
rect 4493 4828 4499 4832
rect 4493 4788 4499 4792
rect 4669 4728 4675 4912
rect 4829 4908 4835 5032
rect 4845 5008 4851 5072
rect 4861 4928 4867 5092
rect 4893 5088 4899 5132
rect 4925 5108 4931 5112
rect 5053 5106 5059 5112
rect 4877 4968 4883 5032
rect 4893 4948 4899 5072
rect 4925 4948 4931 5092
rect 4461 4697 4483 4703
rect 4445 4668 4451 4692
rect 4381 4388 4387 4512
rect 4397 4508 4403 4632
rect 4461 4588 4467 4697
rect 4525 4688 4531 4692
rect 4541 4628 4547 4632
rect 4589 4548 4595 4612
rect 4637 4588 4643 4692
rect 4669 4688 4675 4712
rect 4733 4708 4739 4832
rect 4797 4788 4803 4892
rect 4685 4548 4691 4572
rect 4493 4508 4499 4512
rect 4621 4508 4627 4512
rect 4749 4503 4755 4652
rect 4765 4588 4771 4632
rect 4781 4548 4787 4612
rect 4797 4528 4803 4552
rect 4749 4497 4771 4503
rect 4333 4128 4339 4172
rect 4349 4148 4355 4352
rect 4413 4308 4419 4492
rect 4621 4488 4627 4492
rect 4429 4328 4435 4332
rect 4445 4308 4451 4352
rect 4461 4148 4467 4312
rect 4525 4228 4531 4432
rect 4541 4288 4547 4352
rect 4349 3968 4355 4132
rect 4397 4128 4403 4132
rect 4461 4128 4467 4132
rect 4541 4128 4547 4132
rect 4589 4128 4595 4372
rect 4621 4148 4627 4472
rect 4413 4088 4419 4092
rect 4285 3928 4291 3932
rect 4301 3908 4307 3932
rect 4333 3917 4344 3923
rect 4333 3908 4339 3917
rect 4333 3828 4339 3872
rect 4381 3788 4387 4072
rect 4429 4063 4435 4092
rect 4408 4057 4435 4063
rect 4445 4048 4451 4072
rect 4477 4028 4483 4092
rect 4397 3928 4403 3932
rect 4429 3908 4435 3912
rect 4445 3908 4451 3952
rect 3901 3728 3907 3732
rect 3917 3728 3923 3732
rect 3949 3728 3955 3732
rect 3869 3708 3875 3712
rect 3965 3697 3976 3703
rect 3933 3688 3939 3692
rect 3837 3588 3843 3592
rect 3821 3448 3827 3512
rect 3837 3508 3843 3532
rect 3773 3377 3795 3383
rect 3677 3368 3683 3372
rect 3389 3348 3395 3352
rect 3485 3348 3491 3352
rect 3693 3348 3699 3372
rect 3405 3308 3411 3312
rect 3421 3308 3427 3312
rect 3453 3308 3459 3312
rect 3005 3088 3011 3192
rect 3021 3108 3027 3292
rect 3101 3268 3107 3292
rect 3261 3208 3267 3292
rect 3213 3128 3219 3192
rect 3373 3148 3379 3292
rect 3053 3117 3064 3123
rect 3053 3108 3059 3117
rect 2925 3028 2931 3032
rect 2973 2988 2979 3052
rect 2989 2948 2995 3032
rect 3021 2948 3027 3092
rect 3085 3088 3091 3112
rect 3101 3108 3107 3112
rect 3101 3068 3107 3092
rect 3149 3068 3155 3072
rect 3133 3008 3139 3032
rect 2525 2908 2531 2912
rect 2317 2783 2323 2872
rect 2365 2808 2371 2892
rect 2525 2788 2531 2892
rect 2301 2777 2323 2783
rect 2141 2588 2147 2612
rect 2125 2548 2131 2552
rect 2173 2548 2179 2572
rect 2125 2508 2131 2532
rect 2237 2528 2243 2632
rect 2269 2623 2275 2692
rect 2301 2688 2307 2777
rect 2349 2688 2355 2692
rect 2301 2668 2307 2672
rect 2269 2617 2291 2623
rect 2269 2588 2275 2592
rect 2285 2588 2291 2617
rect 2333 2548 2339 2572
rect 2381 2548 2387 2692
rect 2477 2688 2483 2732
rect 2509 2728 2515 2752
rect 2557 2708 2563 2752
rect 2397 2548 2403 2672
rect 2573 2668 2579 2672
rect 2413 2588 2419 2612
rect 2493 2528 2499 2532
rect 2589 2528 2595 2692
rect 2621 2548 2627 2932
rect 2893 2908 2899 2932
rect 3069 2928 3075 2992
rect 3181 2988 3187 3052
rect 2733 2768 2739 2892
rect 2637 2688 2643 2692
rect 1885 2328 1891 2352
rect 1885 2288 1891 2292
rect 1789 2168 1795 2212
rect 1821 2148 1827 2252
rect 1901 2228 1907 2432
rect 1917 2308 1923 2492
rect 2365 2488 2371 2492
rect 2413 2488 2419 2492
rect 2589 2428 2595 2512
rect 2637 2508 2643 2512
rect 1981 2328 1987 2332
rect 2029 2308 2035 2332
rect 2285 2308 2291 2312
rect 2301 2308 2307 2312
rect 2381 2288 2387 2332
rect 2589 2288 2595 2332
rect 2669 2328 2675 2752
rect 2717 2548 2723 2572
rect 2765 2548 2771 2872
rect 2781 2706 2787 2752
rect 2845 2688 2851 2852
rect 2781 2528 2787 2552
rect 2797 2528 2803 2612
rect 2813 2608 2819 2672
rect 2845 2668 2851 2672
rect 2909 2668 2915 2672
rect 2909 2648 2915 2652
rect 2909 2568 2915 2592
rect 2925 2543 2931 2912
rect 3149 2888 3155 2932
rect 3213 2928 3219 3112
rect 3261 2988 3267 3112
rect 3309 3068 3315 3072
rect 3325 3068 3331 3092
rect 3389 3088 3395 3092
rect 3373 3048 3379 3072
rect 3405 3068 3411 3292
rect 3437 3288 3443 3292
rect 3421 3088 3427 3112
rect 3437 3088 3443 3112
rect 3533 3106 3539 3112
rect 3549 3088 3555 3332
rect 3565 3288 3571 3312
rect 3693 3168 3699 3332
rect 3709 3328 3715 3332
rect 3757 3188 3763 3272
rect 3773 3148 3779 3377
rect 3789 3348 3795 3352
rect 3805 3288 3811 3292
rect 3821 3223 3827 3432
rect 3853 3388 3859 3392
rect 3837 3308 3843 3332
rect 3853 3283 3859 3292
rect 3805 3217 3827 3223
rect 3837 3277 3859 3283
rect 3789 3088 3795 3132
rect 3805 3128 3811 3217
rect 3821 3148 3827 3192
rect 3837 3188 3843 3277
rect 3869 3268 3875 3652
rect 3901 3628 3907 3672
rect 3933 3568 3939 3672
rect 3965 3588 3971 3697
rect 4045 3588 4051 3732
rect 4077 3688 4083 3692
rect 3885 3388 3891 3512
rect 3901 3448 3907 3532
rect 3949 3528 3955 3572
rect 4061 3568 4067 3592
rect 3917 3408 3923 3492
rect 3949 3468 3955 3512
rect 3997 3508 4003 3532
rect 4061 3528 4067 3552
rect 4077 3528 4083 3632
rect 4093 3588 4099 3732
rect 4125 3717 4136 3723
rect 4045 3508 4051 3512
rect 3896 3337 3912 3343
rect 3917 3308 3923 3312
rect 3869 3103 3875 3252
rect 3901 3128 3907 3292
rect 3933 3288 3939 3432
rect 3965 3408 3971 3492
rect 3981 3328 3987 3332
rect 3933 3208 3939 3272
rect 3965 3168 3971 3292
rect 3997 3288 4003 3492
rect 4029 3308 4035 3352
rect 3981 3268 3987 3272
rect 4045 3188 4051 3332
rect 4061 3308 4067 3512
rect 4077 3468 4083 3512
rect 4093 3508 4099 3512
rect 4109 3448 4115 3532
rect 4125 3443 4131 3717
rect 4157 3703 4163 3712
rect 4157 3697 4168 3703
rect 4157 3588 4163 3672
rect 4205 3588 4211 3692
rect 4253 3588 4259 3692
rect 4269 3688 4275 3772
rect 4397 3763 4403 3892
rect 4445 3888 4451 3892
rect 4413 3788 4419 3832
rect 4461 3788 4467 3852
rect 4397 3757 4419 3763
rect 4285 3728 4291 3752
rect 4333 3728 4339 3732
rect 4349 3728 4355 3752
rect 4285 3668 4291 3672
rect 4301 3648 4307 3692
rect 4333 3628 4339 3672
rect 4141 3568 4147 3572
rect 4141 3528 4147 3552
rect 4333 3548 4339 3612
rect 4173 3528 4179 3532
rect 4125 3437 4147 3443
rect 4141 3328 4147 3437
rect 4157 3428 4163 3492
rect 4237 3483 4243 3512
rect 4237 3477 4259 3483
rect 4173 3388 4179 3432
rect 4253 3428 4259 3477
rect 4269 3448 4275 3532
rect 4349 3528 4355 3632
rect 4365 3608 4371 3692
rect 4381 3688 4387 3732
rect 4413 3588 4419 3757
rect 4429 3728 4435 3732
rect 4440 3697 4451 3703
rect 4445 3588 4451 3697
rect 4477 3568 4483 4012
rect 4525 4008 4531 4032
rect 4493 3908 4499 3992
rect 4541 3988 4547 4112
rect 4605 4108 4611 4132
rect 4525 3968 4531 3972
rect 4509 3897 4520 3903
rect 4509 3883 4515 3897
rect 4504 3877 4515 3883
rect 4541 3868 4547 3932
rect 4589 3903 4595 4032
rect 4637 3988 4643 4492
rect 4685 4306 4691 4332
rect 4749 4288 4755 4352
rect 4669 4048 4675 4112
rect 4589 3897 4600 3903
rect 4637 3888 4643 3892
rect 4493 3788 4499 3852
rect 4557 3788 4563 3872
rect 4653 3868 4659 3932
rect 4573 3848 4579 3852
rect 4589 3768 4595 3812
rect 4525 3708 4531 3712
rect 4509 3588 4515 3692
rect 4365 3528 4371 3552
rect 4397 3523 4403 3532
rect 4397 3517 4419 3523
rect 4253 3388 4259 3412
rect 4285 3388 4291 3512
rect 4333 3488 4339 3492
rect 4381 3488 4387 3492
rect 3864 3097 3875 3103
rect 3917 3088 3923 3152
rect 3933 3108 3939 3132
rect 3981 3128 3987 3132
rect 3933 3088 3939 3092
rect 3981 3088 3987 3092
rect 3261 2948 3267 2952
rect 3325 2948 3331 3032
rect 3517 2968 3523 2972
rect 3533 2948 3539 3052
rect 3661 3048 3667 3072
rect 3709 3068 3715 3072
rect 3549 2988 3555 3032
rect 3325 2928 3331 2932
rect 3613 2928 3619 2932
rect 3213 2908 3219 2912
rect 3389 2908 3395 2914
rect 2989 2728 2995 2732
rect 2941 2648 2947 2712
rect 3085 2708 3091 2712
rect 3053 2568 3059 2692
rect 3149 2688 3155 2872
rect 3501 2788 3507 2832
rect 3581 2788 3587 2892
rect 3597 2868 3603 2912
rect 3213 2708 3219 2732
rect 3325 2688 3331 2732
rect 3117 2548 3123 2632
rect 3149 2608 3155 2672
rect 3149 2548 3155 2572
rect 2909 2537 2931 2543
rect 2781 2488 2787 2512
rect 2669 2308 2675 2312
rect 2621 2288 2627 2292
rect 1933 2268 1939 2272
rect 1949 2208 1955 2272
rect 2045 2268 2051 2272
rect 1997 2208 2003 2232
rect 1853 2188 1859 2192
rect 1757 2137 1779 2143
rect 1773 2128 1779 2137
rect 1757 2108 1763 2112
rect 1757 2088 1763 2092
rect 1725 1888 1731 2032
rect 1789 1908 1795 1932
rect 1693 1828 1699 1832
rect 1709 1788 1715 1792
rect 1613 1508 1619 1512
rect 1629 1508 1635 1512
rect 1645 1483 1651 1732
rect 1725 1708 1731 1732
rect 1741 1708 1747 1892
rect 1837 1888 1843 2132
rect 1965 2128 1971 2192
rect 2061 2188 2067 2232
rect 1853 1908 1859 2032
rect 1896 1917 1923 1923
rect 1917 1903 1923 1917
rect 1917 1897 1944 1903
rect 1773 1868 1779 1872
rect 1821 1848 1827 1852
rect 1773 1728 1779 1792
rect 1853 1768 1859 1892
rect 1885 1848 1891 1892
rect 2013 1888 2019 2132
rect 2125 2128 2131 2212
rect 2141 2148 2147 2272
rect 2253 2248 2259 2272
rect 2445 2268 2451 2272
rect 2189 2148 2195 2152
rect 2109 2108 2115 2112
rect 2205 2108 2211 2112
rect 2029 1868 2035 1892
rect 1933 1808 1939 1832
rect 1640 1477 1651 1483
rect 1309 1128 1315 1132
rect 1341 1128 1347 1132
rect 1357 1088 1363 1152
rect 1437 1128 1443 1132
rect 1245 968 1251 1072
rect 1405 1068 1411 1072
rect 1261 948 1267 992
rect 1229 908 1235 932
rect 1245 928 1251 932
rect 1277 908 1283 1032
rect 1341 908 1347 1032
rect 1053 897 1075 903
rect 1053 788 1059 897
rect 1389 903 1395 1032
rect 1421 948 1427 1092
rect 1453 948 1459 952
rect 1389 897 1400 903
rect 1133 708 1139 732
rect 1085 688 1091 692
rect 1165 648 1171 692
rect 845 443 851 512
rect 957 508 963 512
rect 973 488 979 532
rect 1085 508 1091 532
rect 845 437 867 443
rect 861 288 867 437
rect 893 306 899 312
rect 1037 308 1043 352
rect 1085 308 1091 492
rect 1181 388 1187 872
rect 1197 808 1203 832
rect 1197 688 1203 792
rect 1357 788 1363 832
rect 1213 588 1219 672
rect 1261 648 1267 712
rect 1245 528 1251 632
rect 1277 588 1283 692
rect 1325 688 1331 692
rect 1373 688 1379 692
rect 1389 688 1395 792
rect 1421 788 1427 912
rect 1469 908 1475 1032
rect 1485 1028 1491 1072
rect 1501 943 1507 1172
rect 1496 937 1507 943
rect 1501 768 1507 832
rect 1405 708 1411 752
rect 1469 728 1475 752
rect 1517 743 1523 1292
rect 1597 1188 1603 1192
rect 1533 1128 1539 1132
rect 1549 1088 1555 1112
rect 1581 1088 1587 1092
rect 1597 1088 1603 1172
rect 1677 1168 1683 1692
rect 1837 1508 1843 1612
rect 1853 1508 1859 1672
rect 1757 1468 1763 1472
rect 1757 1348 1763 1452
rect 1837 1348 1843 1392
rect 1709 1308 1715 1312
rect 1757 1308 1763 1332
rect 1853 1328 1859 1352
rect 1885 1328 1891 1752
rect 1901 1728 1907 1752
rect 2013 1748 2019 1752
rect 1901 1368 1907 1472
rect 1901 1348 1907 1352
rect 1917 1328 1923 1692
rect 1933 1508 1939 1532
rect 1949 1468 1955 1732
rect 2045 1708 2051 1712
rect 2077 1688 2083 1732
rect 2093 1668 2099 1712
rect 2109 1628 2115 2092
rect 2157 1968 2163 2032
rect 2157 1848 2163 1872
rect 2125 1788 2131 1832
rect 2141 1783 2147 1832
rect 2141 1777 2163 1783
rect 2061 1506 2067 1532
rect 1997 1468 2003 1492
rect 2125 1488 2131 1492
rect 1997 1368 2003 1452
rect 2029 1368 2035 1372
rect 1976 1337 1992 1343
rect 2013 1343 2019 1352
rect 2013 1337 2035 1343
rect 1629 1108 1635 1152
rect 1677 1128 1683 1152
rect 1837 1108 1843 1292
rect 1789 1088 1795 1092
rect 1837 1088 1843 1092
rect 1613 1048 1619 1072
rect 1709 1048 1715 1072
rect 1533 908 1539 1032
rect 1549 968 1555 972
rect 1752 957 1784 963
rect 1597 948 1603 952
rect 1581 908 1587 912
rect 1645 908 1651 912
rect 1661 868 1667 932
rect 1677 928 1683 952
rect 1805 948 1811 972
rect 1789 928 1795 932
rect 1677 888 1683 912
rect 1709 828 1715 912
rect 1853 868 1859 952
rect 1885 948 1891 1272
rect 1917 1023 1923 1312
rect 1965 1308 1971 1312
rect 1965 1088 1971 1092
rect 2029 1088 2035 1337
rect 2141 1328 2147 1752
rect 2157 1728 2163 1777
rect 2173 1628 2179 1712
rect 2157 1508 2163 1512
rect 2205 1508 2211 2092
rect 2269 1908 2275 1992
rect 2269 1808 2275 1892
rect 2285 1888 2291 2252
rect 2445 2148 2451 2252
rect 2333 2128 2339 2132
rect 2461 2128 2467 2132
rect 2509 2028 2515 2132
rect 2333 1988 2339 2012
rect 2317 1848 2323 1892
rect 2365 1868 2371 1892
rect 2237 1568 2243 1632
rect 2253 1488 2259 1732
rect 2301 1623 2307 1732
rect 2349 1728 2355 1732
rect 2381 1628 2387 1892
rect 2397 1828 2403 1852
rect 2413 1803 2419 1832
rect 2429 1828 2435 1892
rect 2461 1888 2467 1892
rect 2413 1797 2435 1803
rect 2429 1668 2435 1797
rect 2445 1788 2451 1872
rect 2461 1788 2467 1832
rect 2477 1828 2483 1872
rect 2493 1828 2499 1892
rect 2509 1888 2515 1952
rect 2573 1928 2579 2232
rect 2461 1748 2467 1772
rect 2557 1708 2563 1892
rect 2573 1868 2579 1872
rect 2605 1728 2611 1792
rect 2621 1748 2627 2232
rect 2685 2228 2691 2272
rect 2749 2163 2755 2432
rect 2829 2408 2835 2492
rect 2909 2488 2915 2537
rect 2925 2508 2931 2512
rect 2877 2328 2883 2332
rect 2797 2188 2803 2232
rect 2749 2157 2771 2163
rect 2701 2108 2707 2132
rect 2733 2108 2739 2132
rect 2765 2128 2771 2157
rect 2781 2148 2787 2152
rect 2797 2148 2803 2172
rect 2669 1908 2675 1972
rect 2637 1888 2643 1892
rect 2541 1648 2547 1692
rect 2589 1648 2595 1712
rect 2605 1708 2611 1712
rect 2285 1617 2307 1623
rect 2269 1508 2275 1512
rect 2253 1468 2259 1472
rect 2285 1368 2291 1617
rect 2477 1588 2483 1632
rect 2397 1508 2403 1512
rect 2301 1488 2307 1492
rect 2445 1488 2451 1492
rect 2333 1448 2339 1472
rect 2253 1348 2259 1352
rect 2381 1328 2387 1432
rect 2429 1368 2435 1472
rect 2061 1168 2067 1312
rect 2077 1108 2083 1112
rect 2109 1108 2115 1312
rect 2125 1128 2131 1132
rect 2061 1088 2067 1092
rect 2077 1088 2083 1092
rect 1981 1068 1987 1072
rect 1901 1017 1923 1023
rect 1901 928 1907 1017
rect 1965 968 1971 972
rect 1997 928 2003 972
rect 2013 948 2019 952
rect 2040 917 2051 923
rect 1949 888 1955 912
rect 1853 788 1859 852
rect 1933 788 1939 792
rect 1517 737 1539 743
rect 1309 528 1315 532
rect 1341 508 1347 532
rect 1421 528 1427 712
rect 1517 708 1523 712
rect 1501 588 1507 672
rect 1517 568 1523 672
rect 1517 548 1523 552
rect 1277 368 1283 432
rect 1133 308 1139 352
rect 1277 328 1283 332
rect 1261 308 1267 312
rect 1389 308 1395 332
rect 1085 288 1091 292
rect 1149 288 1155 292
rect 648 257 659 263
rect 653 188 659 257
rect 653 148 659 172
rect 829 168 835 272
rect 861 163 867 272
rect 1021 188 1027 272
rect 845 157 867 163
rect 749 148 755 152
rect 845 148 851 157
rect 957 148 963 152
rect 1021 148 1027 172
rect 1085 148 1091 272
rect 1197 188 1203 292
rect 685 128 691 132
rect 829 128 835 132
rect 1229 130 1235 132
rect 429 108 435 112
rect 733 108 739 112
rect 1053 108 1059 112
rect 1261 108 1267 232
rect 1341 148 1347 152
rect 1357 128 1363 292
rect 1437 188 1443 472
rect 1533 328 1539 737
rect 1581 688 1587 692
rect 1613 688 1619 732
rect 1837 708 1843 732
rect 1981 708 1987 732
rect 1565 388 1571 512
rect 1629 388 1635 632
rect 1645 528 1651 552
rect 1693 528 1699 672
rect 1789 528 1795 592
rect 1805 548 1811 552
rect 1533 308 1539 312
rect 1565 288 1571 312
rect 1661 308 1667 392
rect 1629 297 1640 303
rect 1480 277 1491 283
rect 1405 128 1411 132
rect 1469 128 1475 172
rect 1485 148 1491 277
rect 1629 168 1635 297
rect 1693 288 1699 512
rect 1821 408 1827 692
rect 1837 548 1843 572
rect 1869 508 1875 592
rect 1885 588 1891 692
rect 1949 528 1955 552
rect 1693 148 1699 272
rect 1837 188 1843 452
rect 1869 328 1875 492
rect 1869 308 1875 312
rect 1885 308 1891 312
rect 1965 308 1971 332
rect 1965 288 1971 292
rect 1549 128 1555 132
rect 1837 128 1843 172
rect 1869 148 1875 272
rect 1981 148 1987 512
rect 1997 388 2003 612
rect 2013 608 2019 632
rect 2029 308 2035 792
rect 2045 668 2051 917
rect 2061 848 2067 1072
rect 2093 1068 2099 1072
rect 2077 708 2083 812
rect 2093 668 2099 932
rect 2109 928 2115 1092
rect 2109 908 2115 912
rect 2125 708 2131 912
rect 2141 808 2147 1312
rect 2205 1168 2211 1232
rect 2205 1088 2211 1092
rect 2221 1088 2227 1192
rect 2157 928 2163 972
rect 2237 868 2243 912
rect 2237 828 2243 852
rect 2253 763 2259 1152
rect 2269 1108 2275 1112
rect 2285 968 2291 1072
rect 2301 1028 2307 1092
rect 2301 948 2307 952
rect 2269 788 2275 812
rect 2253 757 2275 763
rect 2221 708 2227 752
rect 2045 648 2051 652
rect 2077 508 2083 532
rect 2093 388 2099 652
rect 2173 548 2179 572
rect 2269 528 2275 757
rect 2317 728 2323 1212
rect 2493 1188 2499 1492
rect 2525 1348 2531 1612
rect 2573 1448 2579 1452
rect 2525 1328 2531 1332
rect 2541 1108 2547 1432
rect 2589 1108 2595 1152
rect 2349 1068 2355 1072
rect 2333 968 2339 972
rect 2349 968 2355 992
rect 2365 928 2371 1092
rect 2429 1068 2435 1072
rect 2397 948 2403 952
rect 2413 928 2419 932
rect 2445 928 2451 1092
rect 2493 1068 2499 1072
rect 2461 948 2467 972
rect 2509 948 2515 952
rect 2445 788 2451 892
rect 2317 708 2323 712
rect 2301 588 2307 672
rect 2301 568 2307 572
rect 2301 548 2307 552
rect 2141 508 2147 512
rect 2237 448 2243 512
rect 2125 308 2131 392
rect 2109 183 2115 292
rect 2237 288 2243 432
rect 2104 177 2115 183
rect 2109 148 2115 177
rect 2221 148 2227 172
rect 2285 148 2291 272
rect 1501 108 1507 112
rect 1869 108 1875 112
rect 1901 108 1907 132
rect 2269 108 2275 112
rect 2285 108 2291 112
rect 2317 108 2323 692
rect 2413 688 2419 692
rect 2349 588 2355 652
rect 2429 588 2435 692
rect 2461 683 2467 932
rect 2504 917 2515 923
rect 2477 768 2483 912
rect 2493 708 2499 752
rect 2461 677 2483 683
rect 2477 508 2483 677
rect 2493 628 2499 692
rect 2509 688 2515 917
rect 2541 868 2547 1092
rect 2584 1057 2595 1063
rect 2589 1028 2595 1057
rect 2589 888 2595 1012
rect 2605 788 2611 1692
rect 2653 1448 2659 1892
rect 2717 1808 2723 1852
rect 2717 1748 2723 1792
rect 2733 1748 2739 1752
rect 2685 1723 2691 1732
rect 2749 1728 2755 1872
rect 2765 1868 2771 2112
rect 2813 2108 2819 2272
rect 2909 2143 2915 2472
rect 2925 2328 2931 2392
rect 2973 2308 2979 2392
rect 2925 2288 2931 2292
rect 2989 2268 2995 2272
rect 3005 2228 3011 2272
rect 3053 2168 3059 2532
rect 3069 2528 3075 2532
rect 3117 2508 3123 2532
rect 3293 2528 3299 2552
rect 3229 2348 3235 2492
rect 3069 2308 3075 2312
rect 3261 2288 3267 2292
rect 3229 2277 3240 2283
rect 2909 2137 2931 2143
rect 2845 2128 2851 2132
rect 2813 1988 2819 2092
rect 2829 2008 2835 2092
rect 2685 1717 2707 1723
rect 2701 1708 2707 1717
rect 2749 1628 2755 1712
rect 2765 1703 2771 1832
rect 2797 1788 2803 1792
rect 2765 1697 2776 1703
rect 2701 1506 2707 1512
rect 2765 1488 2771 1532
rect 2701 1448 2707 1452
rect 2701 1368 2707 1432
rect 2813 1328 2819 1792
rect 2829 1528 2835 1852
rect 2845 1808 2851 1892
rect 2877 1808 2883 2032
rect 2925 1908 2931 2137
rect 2957 2088 2963 2112
rect 3021 2108 3027 2132
rect 3037 2128 3043 2132
rect 3053 2048 3059 2052
rect 2957 1988 2963 1992
rect 3021 1988 3027 2012
rect 2957 1968 2963 1972
rect 3053 1908 3059 2032
rect 3085 1988 3091 2212
rect 3133 1988 3139 2252
rect 3160 2237 3171 2243
rect 3149 2128 3155 2172
rect 3165 2108 3171 2237
rect 3229 2108 3235 2277
rect 3277 2188 3283 2472
rect 3309 2143 3315 2652
rect 3341 2528 3347 2772
rect 3389 2728 3395 2732
rect 3357 2708 3363 2712
rect 3405 2548 3411 2692
rect 3437 2688 3443 2712
rect 3533 2708 3539 2712
rect 3560 2697 3571 2703
rect 3501 2688 3507 2692
rect 3421 2668 3427 2672
rect 3421 2588 3427 2632
rect 3485 2588 3491 2672
rect 3469 2568 3475 2572
rect 3517 2568 3523 2672
rect 3565 2628 3571 2697
rect 3373 2328 3379 2432
rect 3373 2308 3379 2312
rect 3437 2288 3443 2532
rect 3501 2528 3507 2532
rect 3517 2528 3523 2552
rect 3565 2528 3571 2612
rect 3469 2388 3475 2512
rect 3517 2288 3523 2512
rect 3549 2488 3555 2492
rect 3597 2468 3603 2852
rect 3613 2688 3619 2912
rect 3645 2748 3651 2912
rect 3661 2903 3667 3012
rect 3693 2908 3699 3032
rect 3709 2988 3715 3052
rect 3789 2988 3795 3072
rect 4029 3048 4035 3052
rect 3709 2948 3715 2952
rect 3661 2897 3672 2903
rect 3741 2788 3747 2932
rect 3869 2928 3875 2992
rect 3885 2968 3891 3032
rect 4093 2988 4099 3312
rect 4125 3288 4131 3292
rect 4141 3228 4147 3312
rect 3885 2948 3891 2952
rect 3949 2928 3955 2932
rect 3757 2868 3763 2912
rect 3885 2888 3891 2912
rect 3981 2888 3987 2932
rect 3757 2788 3763 2852
rect 3629 2648 3635 2692
rect 3645 2688 3651 2732
rect 3677 2708 3683 2712
rect 3869 2688 3875 2692
rect 3613 2528 3619 2532
rect 3629 2368 3635 2632
rect 3645 2588 3651 2672
rect 3725 2648 3731 2652
rect 3677 2528 3683 2552
rect 3789 2548 3795 2552
rect 3597 2308 3603 2312
rect 3645 2308 3651 2472
rect 3304 2137 3315 2143
rect 3165 1908 3171 1972
rect 2909 1748 2915 1892
rect 2909 1708 2915 1712
rect 2829 1508 2835 1512
rect 2909 1508 2915 1612
rect 2861 1468 2867 1472
rect 2829 1328 2835 1332
rect 2909 1328 2915 1492
rect 2813 1168 2819 1312
rect 2701 1028 2707 1052
rect 2701 968 2707 1012
rect 2765 948 2771 972
rect 2541 728 2547 772
rect 2557 708 2563 732
rect 2509 668 2515 672
rect 2541 508 2547 632
rect 2509 388 2515 492
rect 2557 408 2563 612
rect 2605 568 2611 612
rect 2605 548 2611 552
rect 2573 508 2579 512
rect 2589 488 2595 532
rect 2621 528 2627 772
rect 2669 688 2675 692
rect 2685 688 2691 932
rect 2797 928 2803 932
rect 2749 728 2755 772
rect 2797 728 2803 892
rect 2797 708 2803 712
rect 2653 528 2659 532
rect 2365 308 2371 312
rect 2381 308 2387 312
rect 2461 288 2467 332
rect 2557 308 2563 392
rect 2541 188 2547 292
rect 2589 288 2595 472
rect 2637 308 2643 312
rect 2685 308 2691 532
rect 2749 508 2755 632
rect 2781 588 2787 672
rect 2797 628 2803 672
rect 2813 528 2819 1152
rect 2829 748 2835 1312
rect 2845 1128 2851 1132
rect 2845 1088 2851 1112
rect 2861 948 2867 1252
rect 2925 1228 2931 1892
rect 3037 1768 3043 1872
rect 3053 1728 3059 1752
rect 3085 1548 3091 1832
rect 3085 1528 3091 1532
rect 2973 1488 2979 1512
rect 3005 1468 3011 1472
rect 3021 1448 3027 1472
rect 2957 1348 2963 1372
rect 3101 1363 3107 1732
rect 3165 1728 3171 1892
rect 3229 1888 3235 2092
rect 3245 2028 3251 2132
rect 3341 2128 3347 2272
rect 3389 2148 3395 2232
rect 3437 2168 3443 2272
rect 3453 2248 3459 2252
rect 3469 2168 3475 2272
rect 3357 2128 3363 2132
rect 3277 2108 3283 2112
rect 3309 2108 3315 2112
rect 3501 2108 3507 2232
rect 3549 2203 3555 2272
rect 3533 2197 3555 2203
rect 3533 2168 3539 2197
rect 3597 2148 3603 2252
rect 3645 2188 3651 2292
rect 3661 2128 3667 2132
rect 3309 1968 3315 2092
rect 3613 2088 3619 2112
rect 3661 2088 3667 2092
rect 3325 1868 3331 1872
rect 3181 1748 3187 1772
rect 3181 1728 3187 1732
rect 3213 1628 3219 1812
rect 3245 1808 3251 1812
rect 3245 1708 3251 1792
rect 3357 1748 3363 1892
rect 3309 1708 3315 1712
rect 3325 1568 3331 1732
rect 3341 1708 3347 1712
rect 3149 1506 3155 1532
rect 3309 1528 3315 1532
rect 3341 1528 3347 1552
rect 3373 1528 3379 1952
rect 3421 1908 3427 1952
rect 3469 1928 3475 1952
rect 3469 1888 3475 1892
rect 3533 1868 3539 1872
rect 3389 1768 3395 1832
rect 3613 1828 3619 2072
rect 3421 1748 3427 1752
rect 3437 1728 3443 1792
rect 3677 1748 3683 2512
rect 3741 2508 3747 2532
rect 3885 2528 3891 2872
rect 4109 2868 4115 2912
rect 4061 2708 4067 2852
rect 3917 2528 3923 2672
rect 4045 2588 4051 2692
rect 3981 2568 3987 2572
rect 3981 2528 3987 2552
rect 4109 2528 4115 2772
rect 4141 2648 4147 3212
rect 4189 2868 4195 3052
rect 4221 2948 4227 2952
rect 4189 2748 4195 2812
rect 4189 2708 4195 2732
rect 4221 2708 4227 2712
rect 4269 2708 4275 3192
rect 4333 3188 4339 3332
rect 4365 3328 4371 3332
rect 4376 3297 4387 3303
rect 4285 2928 4291 2932
rect 4125 2548 4131 2632
rect 4173 2588 4179 2692
rect 4189 2543 4195 2692
rect 4189 2537 4200 2543
rect 4253 2528 4259 2632
rect 3757 2508 3763 2512
rect 3853 2508 3859 2514
rect 3917 2488 3923 2512
rect 4013 2508 4019 2512
rect 3757 2328 3763 2332
rect 3757 2288 3763 2312
rect 3805 2308 3811 2312
rect 3821 2288 3827 2312
rect 3901 2308 3907 2352
rect 3949 2328 3955 2352
rect 3949 2288 3955 2292
rect 3981 2288 3987 2332
rect 3885 2268 3891 2272
rect 3757 2208 3763 2232
rect 3757 2168 3763 2172
rect 3693 2148 3699 2152
rect 3709 1888 3715 1932
rect 3789 1928 3795 2192
rect 3885 2168 3891 2172
rect 3981 2168 3987 2272
rect 3933 2128 3939 2132
rect 3805 1928 3811 2052
rect 3933 2028 3939 2112
rect 3837 1908 3843 2012
rect 3933 1928 3939 1932
rect 3709 1868 3715 1872
rect 3757 1868 3763 1892
rect 3837 1868 3843 1892
rect 3581 1728 3587 1732
rect 3608 1717 3619 1723
rect 3277 1508 3283 1512
rect 3085 1357 3107 1363
rect 3037 1308 3043 1312
rect 2941 1288 2947 1292
rect 2877 1128 2883 1152
rect 2941 1108 2947 1152
rect 2877 1088 2883 1092
rect 2877 968 2883 1032
rect 2845 908 2851 912
rect 2861 688 2867 692
rect 2877 588 2883 932
rect 2909 928 2915 1052
rect 2957 963 2963 1032
rect 2941 957 2963 963
rect 2973 963 2979 1212
rect 2989 1068 2995 1072
rect 2989 1048 2995 1052
rect 3021 1028 3027 1072
rect 2973 957 2995 963
rect 2909 768 2915 912
rect 2941 903 2947 957
rect 2941 897 2952 903
rect 2941 788 2947 872
rect 2909 708 2915 752
rect 2989 708 2995 957
rect 2909 548 2915 692
rect 2925 588 2931 692
rect 2973 688 2979 692
rect 3005 588 3011 992
rect 3053 968 3059 1332
rect 3069 1328 3075 1332
rect 3069 1108 3075 1112
rect 3037 948 3043 952
rect 2925 508 2931 512
rect 2973 508 2979 512
rect 2973 488 2979 492
rect 2685 228 2691 292
rect 2765 288 2771 472
rect 2941 388 2947 432
rect 2989 368 2995 532
rect 2877 328 2883 332
rect 2829 308 2835 312
rect 2877 288 2883 312
rect 2941 308 2947 352
rect 3021 348 3027 492
rect 3037 408 3043 632
rect 3053 588 3059 872
rect 3069 688 3075 732
rect 3085 568 3091 1357
rect 3117 1348 3123 1452
rect 3133 1448 3139 1472
rect 3213 1348 3219 1412
rect 3277 1343 3283 1492
rect 3341 1488 3347 1512
rect 3373 1508 3379 1512
rect 3613 1508 3619 1717
rect 3645 1568 3651 1732
rect 3677 1708 3683 1712
rect 3693 1708 3699 1752
rect 3725 1748 3731 1852
rect 3885 1788 3891 1852
rect 3917 1768 3923 1832
rect 3949 1728 3955 1892
rect 3981 1888 3987 1952
rect 4013 1948 4019 2492
rect 4029 2348 4035 2472
rect 4109 2328 4115 2512
rect 4173 2508 4179 2512
rect 4237 2328 4243 2492
rect 4237 2308 4243 2312
rect 4221 2268 4227 2272
rect 4061 2188 4067 2252
rect 4029 2088 4035 2092
rect 4093 2008 4099 2112
rect 4093 1988 4099 1992
rect 3757 1708 3763 1714
rect 3917 1648 3923 1712
rect 3725 1508 3731 1532
rect 3421 1488 3427 1492
rect 3341 1348 3347 1432
rect 3357 1428 3363 1472
rect 3453 1448 3459 1472
rect 3485 1388 3491 1472
rect 3261 1337 3283 1343
rect 3101 1328 3107 1332
rect 3117 1088 3123 1332
rect 3165 1263 3171 1292
rect 3149 1257 3171 1263
rect 3149 1128 3155 1257
rect 3213 1168 3219 1332
rect 3261 1308 3267 1337
rect 3277 1308 3283 1312
rect 3197 1088 3203 1132
rect 3261 1128 3267 1292
rect 3309 1288 3315 1332
rect 3373 1330 3379 1352
rect 3437 1328 3443 1372
rect 3597 1368 3603 1392
rect 3613 1348 3619 1492
rect 3645 1408 3651 1432
rect 3661 1383 3667 1392
rect 3656 1377 3667 1383
rect 3261 1108 3267 1112
rect 3277 1088 3283 1112
rect 3325 1088 3331 1152
rect 3101 908 3107 912
rect 3085 528 3091 552
rect 3101 368 3107 892
rect 3117 888 3123 1072
rect 3133 708 3139 1012
rect 3165 948 3171 972
rect 3197 948 3203 1012
rect 3373 948 3379 952
rect 3229 908 3235 914
rect 3293 708 3299 732
rect 3373 668 3379 932
rect 3389 928 3395 1312
rect 3437 1108 3443 1312
rect 3421 988 3427 1092
rect 3565 1088 3571 1312
rect 3581 1063 3587 1112
rect 3613 1108 3619 1332
rect 3645 1328 3651 1332
rect 3741 1288 3747 1452
rect 3773 1308 3779 1552
rect 3869 1528 3875 1532
rect 3917 1528 3923 1632
rect 3965 1588 3971 1832
rect 3981 1788 3987 1852
rect 4045 1803 4051 1952
rect 4109 1908 4115 1972
rect 4173 1908 4179 2232
rect 4029 1797 4051 1803
rect 3981 1768 3987 1772
rect 4029 1748 4035 1797
rect 4013 1728 4019 1732
rect 3917 1508 3923 1512
rect 3837 1448 3843 1472
rect 3901 1448 3907 1472
rect 3821 1328 3827 1352
rect 3917 1348 3923 1492
rect 4045 1483 4051 1512
rect 4029 1477 4051 1483
rect 3949 1328 3955 1352
rect 3901 1308 3907 1312
rect 3965 1308 3971 1312
rect 3784 1297 3795 1303
rect 3693 1208 3699 1232
rect 3709 1148 3715 1212
rect 3725 1128 3731 1232
rect 3773 1228 3779 1272
rect 3741 1128 3747 1152
rect 3773 1148 3779 1212
rect 3645 1108 3651 1112
rect 3613 1088 3619 1092
rect 3565 1057 3587 1063
rect 3485 943 3491 1052
rect 3549 1008 3555 1032
rect 3565 988 3571 1057
rect 3480 937 3491 943
rect 3389 908 3395 912
rect 3549 908 3555 972
rect 3581 948 3587 1032
rect 3597 988 3603 1032
rect 3613 923 3619 1072
rect 3613 917 3624 923
rect 3421 708 3427 732
rect 3197 528 3203 552
rect 3293 528 3299 532
rect 3085 308 3091 312
rect 2573 148 2579 212
rect 2701 188 2707 192
rect 2669 168 2675 172
rect 2717 148 2723 152
rect 2765 148 2771 272
rect 2909 148 2915 212
rect 2925 208 2931 272
rect 3021 148 3027 232
rect 2749 128 2755 132
rect 2893 128 2899 132
rect 3085 128 3091 292
rect 3117 288 3123 432
rect 3229 408 3235 432
rect 3117 228 3123 272
rect 3117 148 3123 172
rect 3133 148 3139 192
rect 3149 128 3155 392
rect 3309 388 3315 512
rect 3181 288 3187 332
rect 3245 328 3251 352
rect 3293 308 3299 352
rect 3325 328 3331 632
rect 3373 548 3379 652
rect 3437 548 3443 892
rect 3453 528 3459 552
rect 3437 468 3443 512
rect 3325 308 3331 312
rect 3245 288 3251 292
rect 3341 283 3347 412
rect 3389 288 3395 292
rect 3336 277 3347 283
rect 3325 208 3331 272
rect 3405 248 3411 432
rect 3485 428 3491 432
rect 3421 288 3427 332
rect 3405 208 3411 232
rect 3485 188 3491 252
rect 3453 148 3459 172
rect 3469 148 3475 152
rect 2797 108 2803 112
rect 3085 108 3091 112
rect 3149 108 3155 112
rect 3197 108 3203 132
rect 3501 128 3507 832
rect 3533 728 3539 732
rect 3613 708 3619 712
rect 3549 668 3555 672
rect 3533 528 3539 532
rect 3581 528 3587 552
rect 3533 308 3539 512
rect 3629 508 3635 912
rect 3645 908 3651 932
rect 3677 788 3683 872
rect 3693 788 3699 892
rect 3709 788 3715 892
rect 3725 868 3731 1092
rect 3741 768 3747 1112
rect 3773 888 3779 1132
rect 3789 1128 3795 1297
rect 3805 1248 3811 1272
rect 3821 1128 3827 1232
rect 3837 1168 3843 1292
rect 3885 1168 3891 1232
rect 3901 1128 3907 1292
rect 3997 1288 4003 1432
rect 4029 1408 4035 1477
rect 4045 1388 4051 1432
rect 4061 1428 4067 1692
rect 4077 1683 4083 1832
rect 4173 1788 4179 1872
rect 4141 1748 4147 1772
rect 4109 1728 4115 1732
rect 4189 1728 4195 2132
rect 4237 1948 4243 2012
rect 4253 1988 4259 2512
rect 4285 2508 4291 2892
rect 4301 2768 4307 3092
rect 4317 2948 4323 2972
rect 4349 2788 4355 3252
rect 4365 3148 4371 3272
rect 4381 3188 4387 3297
rect 4397 3128 4403 3412
rect 4413 3388 4419 3517
rect 4429 3428 4435 3512
rect 4429 3188 4435 3332
rect 4445 3248 4451 3492
rect 4461 3288 4467 3532
rect 4477 3388 4483 3452
rect 4493 3168 4499 3512
rect 4525 3488 4531 3532
rect 4509 3388 4515 3412
rect 4541 3408 4547 3752
rect 4589 3748 4595 3752
rect 4589 3703 4595 3712
rect 4589 3697 4600 3703
rect 4637 3688 4643 3692
rect 4653 3628 4659 3712
rect 4637 3588 4643 3612
rect 4669 3608 4675 4032
rect 4685 3928 4691 3972
rect 4749 3908 4755 3932
rect 4733 3888 4739 3892
rect 4685 3788 4691 3872
rect 4765 3768 4771 4497
rect 4813 4388 4819 4712
rect 4861 4708 4867 4892
rect 4829 4668 4835 4692
rect 4861 4508 4867 4692
rect 4877 4588 4883 4932
rect 4989 4928 4995 4932
rect 5005 4908 5011 4952
rect 5069 4888 5075 5232
rect 5085 5048 5091 5312
rect 5181 5308 5187 5312
rect 5149 5288 5155 5292
rect 5197 5288 5203 5312
rect 5357 5268 5363 5312
rect 5117 5248 5123 5252
rect 5117 5108 5123 5232
rect 5453 5228 5459 5232
rect 5565 5128 5571 5312
rect 5661 5308 5667 5312
rect 5581 5288 5587 5292
rect 5581 5128 5587 5272
rect 5757 5268 5763 5272
rect 5693 5188 5699 5232
rect 5597 5108 5603 5112
rect 5197 5088 5203 5092
rect 5085 5028 5091 5032
rect 4893 4728 4899 4872
rect 5085 4848 5091 5012
rect 5005 4708 5011 4712
rect 4909 4648 4915 4672
rect 4909 4528 4915 4632
rect 4925 4528 4931 4532
rect 4813 4288 4819 4372
rect 4845 4368 4851 4432
rect 4845 4308 4851 4312
rect 4861 4308 4867 4492
rect 4877 4488 4883 4492
rect 4925 4388 4931 4492
rect 4989 4468 4995 4492
rect 5005 4388 5011 4652
rect 5021 4548 5027 4712
rect 5037 4568 5043 4572
rect 5053 4448 5059 4512
rect 5053 4328 5059 4352
rect 4797 4248 4803 4252
rect 4781 3928 4787 4232
rect 4813 4168 4819 4272
rect 4845 3968 4851 4292
rect 4877 4268 4883 4312
rect 4893 4288 4899 4292
rect 5005 4268 5011 4292
rect 4877 4148 4883 4172
rect 4893 3948 4899 4172
rect 4909 4128 4915 4132
rect 4957 4128 4963 4132
rect 4989 4128 4995 4212
rect 5037 4148 5043 4272
rect 5021 4088 5027 4132
rect 5069 4128 5075 4832
rect 5133 4728 5139 4752
rect 5197 4708 5203 5072
rect 5229 4968 5235 5092
rect 5389 5088 5395 5090
rect 5533 5088 5539 5092
rect 5213 4908 5219 4912
rect 5261 4728 5267 5032
rect 5421 4988 5427 5072
rect 5453 5048 5459 5052
rect 5485 4968 5491 4972
rect 5421 4948 5427 4952
rect 5325 4908 5331 4932
rect 5357 4908 5363 4912
rect 5485 4908 5491 4914
rect 5533 4848 5539 5072
rect 5549 4868 5555 5092
rect 5549 4788 5555 4852
rect 5389 4728 5395 4732
rect 5197 4668 5203 4672
rect 5133 4628 5139 4632
rect 5165 4528 5171 4612
rect 5197 4508 5203 4552
rect 5213 4508 5219 4512
rect 5229 4468 5235 4472
rect 5133 4288 5139 4372
rect 5165 4306 5171 4312
rect 5101 4148 5107 4272
rect 5149 4188 5155 4212
rect 4909 3988 4915 4072
rect 4861 3908 4867 3912
rect 4877 3888 4883 3892
rect 4781 3788 4787 3832
rect 4845 3828 4851 3872
rect 4749 3628 4755 3692
rect 4701 3588 4707 3612
rect 4525 3188 4531 3292
rect 4557 3208 4563 3492
rect 4573 3428 4579 3472
rect 4573 3388 4579 3412
rect 4637 3408 4643 3492
rect 4653 3488 4659 3532
rect 4728 3497 4744 3503
rect 4781 3488 4787 3752
rect 4877 3748 4883 3792
rect 4973 3788 4979 3812
rect 5005 3728 5011 4032
rect 5133 3988 5139 4052
rect 5037 3908 5043 3912
rect 5053 3788 5059 3852
rect 4957 3688 4963 3712
rect 4829 3588 4835 3632
rect 4797 3517 4808 3523
rect 4797 3508 4803 3517
rect 4621 3388 4627 3392
rect 4685 3388 4691 3392
rect 4669 3368 4675 3372
rect 4701 3357 4739 3363
rect 4680 3337 4691 3343
rect 4605 3328 4611 3332
rect 4429 3128 4435 3152
rect 4493 3128 4499 3152
rect 4573 3148 4579 3232
rect 4440 3117 4451 3123
rect 4445 3108 4451 3117
rect 4589 3108 4595 3192
rect 4621 3188 4627 3292
rect 4605 3128 4611 3152
rect 4605 3097 4616 3103
rect 4381 3088 4387 3092
rect 4493 3088 4499 3092
rect 4605 3028 4611 3097
rect 4573 2968 4579 2972
rect 4557 2928 4563 2932
rect 4445 2868 4451 2912
rect 4557 2828 4563 2912
rect 4605 2848 4611 3012
rect 4333 2708 4339 2712
rect 4397 2588 4403 2652
rect 4365 2508 4371 2572
rect 4285 2288 4291 2292
rect 4317 2288 4323 2332
rect 4285 2128 4291 2212
rect 4317 2168 4323 2272
rect 4333 2128 4339 2132
rect 4349 2108 4355 2192
rect 4397 2128 4403 2132
rect 4413 2108 4419 2572
rect 4429 2288 4435 2672
rect 4445 2488 4451 2732
rect 4493 2708 4499 2772
rect 4637 2723 4643 3232
rect 4685 3188 4691 3337
rect 4701 3328 4707 3357
rect 4717 3308 4723 3312
rect 4733 3308 4739 3357
rect 4765 3268 4771 3292
rect 4781 3188 4787 3332
rect 4797 3308 4803 3472
rect 4813 3388 4819 3472
rect 4829 3388 4835 3572
rect 4861 3528 4867 3552
rect 4877 3368 4883 3492
rect 4893 3428 4899 3532
rect 4909 3528 4915 3632
rect 4941 3588 4947 3672
rect 5005 3668 5011 3712
rect 5021 3708 5027 3712
rect 4989 3528 4995 3632
rect 5021 3628 5027 3692
rect 5005 3588 5011 3612
rect 4845 3328 4851 3352
rect 5005 3328 5011 3372
rect 4813 3188 4819 3292
rect 4829 3248 4835 3292
rect 4861 3288 4867 3292
rect 4877 3188 4883 3272
rect 4653 2988 4659 3032
rect 4669 2848 4675 3112
rect 4749 2988 4755 3052
rect 4733 2948 4739 2952
rect 4701 2928 4707 2932
rect 4632 2717 4643 2723
rect 4525 2648 4531 2692
rect 4653 2668 4659 2732
rect 4669 2728 4675 2752
rect 4685 2748 4691 2872
rect 4717 2828 4723 2892
rect 4765 2888 4771 3132
rect 4797 2908 4803 3112
rect 4813 3028 4819 3092
rect 4813 2928 4819 2932
rect 4573 2588 4579 2612
rect 4461 2528 4467 2532
rect 4525 2528 4531 2532
rect 4477 2508 4483 2512
rect 4605 2508 4611 2592
rect 4557 2488 4563 2492
rect 4509 2468 4515 2472
rect 4525 2468 4531 2472
rect 4605 2388 4611 2492
rect 4621 2488 4627 2652
rect 4717 2588 4723 2812
rect 4781 2808 4787 2892
rect 4845 2828 4851 3152
rect 4893 3108 4899 3112
rect 4909 3088 4915 3232
rect 4941 3228 4947 3312
rect 5021 3308 5027 3532
rect 5085 3388 5091 3432
rect 5069 3328 5075 3352
rect 5117 3348 5123 3612
rect 5133 3588 5139 3952
rect 5165 3528 5171 4152
rect 5293 4148 5299 4652
rect 5373 4628 5379 4692
rect 5325 4528 5331 4612
rect 5389 4528 5395 4692
rect 5309 4388 5315 4472
rect 5325 4408 5331 4512
rect 5389 4508 5395 4512
rect 5405 4508 5411 4752
rect 5453 4688 5459 4732
rect 5597 4728 5603 4772
rect 5613 4708 5619 5172
rect 5885 5148 5891 5332
rect 5917 5168 5923 5332
rect 5997 5308 6003 5312
rect 5645 5088 5651 5132
rect 5421 4588 5427 4652
rect 5453 4628 5459 4632
rect 5421 4508 5427 4552
rect 5341 4488 5347 4492
rect 5405 4488 5411 4492
rect 5373 4468 5379 4472
rect 5357 4208 5363 4232
rect 5357 4148 5363 4192
rect 5373 4168 5379 4452
rect 5389 4288 5395 4292
rect 5437 4288 5443 4412
rect 5453 4308 5459 4572
rect 5469 4528 5475 4532
rect 5485 4528 5491 4612
rect 5501 4548 5507 4552
rect 5181 4108 5187 4112
rect 5197 4108 5203 4132
rect 5213 4128 5219 4132
rect 5245 4068 5251 4092
rect 5197 4037 5208 4043
rect 5197 3903 5203 4037
rect 5197 3897 5219 3903
rect 5181 3863 5187 3892
rect 5213 3868 5219 3897
rect 5277 3888 5283 4132
rect 5293 3908 5299 4112
rect 5373 4088 5379 4132
rect 5181 3857 5203 3863
rect 5165 3508 5171 3512
rect 5181 3508 5187 3592
rect 4973 3128 4979 3232
rect 5005 3148 5011 3292
rect 5037 3108 5043 3232
rect 4925 3008 4931 3092
rect 4989 3048 4995 3092
rect 5085 3088 5091 3092
rect 5101 3088 5107 3112
rect 5037 2988 5043 3052
rect 5005 2908 5011 2952
rect 4845 2788 4851 2812
rect 4744 2717 4755 2723
rect 4749 2708 4755 2717
rect 4733 2688 4739 2692
rect 4749 2668 4755 2672
rect 4637 2528 4643 2552
rect 4669 2528 4675 2532
rect 4717 2528 4723 2532
rect 4621 2468 4627 2472
rect 4749 2468 4755 2632
rect 4669 2388 4675 2432
rect 4749 2388 4755 2452
rect 4781 2388 4787 2692
rect 4797 2628 4803 2652
rect 4861 2648 4867 2872
rect 4893 2848 4899 2892
rect 4573 2308 4579 2372
rect 4797 2303 4803 2492
rect 4877 2408 4883 2712
rect 4893 2708 4899 2712
rect 4941 2708 4947 2772
rect 4925 2568 4931 2632
rect 4957 2608 4963 2892
rect 4973 2868 4979 2872
rect 4973 2788 4979 2852
rect 5021 2788 5027 2832
rect 5053 2708 5059 3072
rect 5069 2948 5075 2972
rect 5085 2928 5091 2992
rect 5069 2903 5075 2912
rect 5069 2897 5080 2903
rect 5117 2708 5123 3332
rect 5133 2948 5139 3432
rect 5149 3108 5155 3492
rect 5165 3328 5171 3472
rect 5197 3428 5203 3857
rect 5261 3708 5267 3772
rect 5229 3648 5235 3672
rect 5181 3348 5187 3352
rect 5165 3188 5171 3312
rect 5197 3208 5203 3232
rect 5149 2928 5155 3032
rect 5133 2768 5139 2892
rect 4957 2588 4963 2592
rect 4973 2548 4979 2632
rect 4925 2488 4931 2532
rect 4957 2528 4963 2532
rect 4957 2448 4963 2492
rect 5005 2448 5011 2512
rect 4792 2297 4803 2303
rect 4637 2268 4643 2292
rect 4701 2288 4707 2292
rect 4541 2208 4547 2232
rect 4461 2108 4467 2112
rect 4477 2108 4483 2172
rect 4573 2168 4579 2192
rect 4589 2148 4595 2252
rect 4637 2248 4643 2252
rect 4605 2143 4611 2232
rect 4605 2137 4627 2143
rect 4317 2068 4323 2072
rect 4333 1988 4339 2032
rect 4253 1948 4259 1952
rect 4269 1928 4275 1932
rect 4333 1908 4339 1912
rect 4253 1848 4259 1892
rect 4285 1868 4291 1872
rect 4125 1708 4131 1712
rect 4157 1697 4168 1703
rect 4077 1677 4088 1683
rect 4125 1568 4131 1692
rect 4141 1568 4147 1672
rect 4157 1588 4163 1697
rect 4141 1548 4147 1552
rect 4189 1528 4195 1712
rect 4221 1708 4227 1772
rect 4253 1728 4259 1832
rect 4301 1808 4307 1832
rect 4349 1788 4355 2092
rect 4381 2028 4387 2072
rect 4365 1848 4371 1892
rect 4397 1888 4403 2032
rect 4429 2028 4435 2032
rect 4461 1948 4467 2072
rect 4477 1948 4483 2092
rect 4509 2088 4515 2092
rect 4525 1988 4531 2032
rect 4541 1968 4547 2072
rect 4493 1863 4499 1912
rect 4477 1857 4499 1863
rect 4429 1828 4435 1832
rect 4328 1757 4339 1763
rect 4333 1743 4339 1757
rect 4333 1737 4344 1743
rect 4317 1728 4323 1732
rect 4237 1688 4243 1712
rect 4237 1528 4243 1672
rect 4269 1588 4275 1632
rect 4317 1548 4323 1672
rect 4381 1648 4387 1692
rect 4445 1648 4451 1692
rect 4333 1588 4339 1632
rect 4285 1528 4291 1532
rect 4109 1508 4115 1512
rect 4125 1497 4136 1503
rect 4093 1483 4099 1492
rect 4125 1483 4131 1497
rect 4168 1497 4296 1503
rect 4093 1477 4131 1483
rect 4317 1468 4323 1532
rect 4397 1508 4403 1572
rect 4317 1448 4323 1452
rect 4013 1368 4019 1372
rect 4013 1328 4019 1352
rect 4029 1328 4035 1372
rect 4045 1328 4051 1372
rect 4029 1308 4035 1312
rect 4093 1308 4099 1412
rect 4253 1368 4259 1412
rect 4136 1357 4152 1363
rect 4269 1328 4275 1352
rect 4413 1308 4419 1632
rect 4429 1548 4435 1552
rect 4445 1548 4451 1552
rect 4477 1528 4483 1857
rect 4493 1728 4499 1832
rect 4509 1748 4515 1772
rect 4509 1703 4515 1712
rect 4541 1708 4547 1952
rect 4573 1903 4579 2072
rect 4589 1948 4595 2052
rect 4568 1897 4579 1903
rect 4589 1828 4595 1932
rect 4605 1928 4611 1952
rect 4621 1928 4627 2137
rect 4669 2128 4675 2232
rect 4781 2208 4787 2292
rect 4701 2130 4707 2132
rect 4765 2128 4771 2152
rect 4637 2068 4643 2092
rect 4829 2088 4835 2272
rect 4733 1928 4739 2012
rect 4813 1988 4819 2052
rect 4829 1948 4835 2032
rect 4765 1908 4771 1912
rect 4637 1888 4643 1892
rect 4797 1888 4803 1932
rect 4845 1928 4851 1972
rect 4669 1808 4675 1832
rect 4557 1748 4563 1752
rect 4653 1728 4659 1792
rect 4701 1748 4707 1832
rect 4504 1697 4515 1703
rect 4621 1668 4627 1692
rect 4717 1688 4723 1852
rect 4813 1768 4819 1792
rect 4765 1728 4771 1732
rect 4589 1628 4595 1632
rect 4669 1548 4675 1632
rect 4733 1568 4739 1632
rect 4509 1528 4515 1532
rect 4621 1508 4627 1512
rect 4445 1428 4451 1492
rect 4557 1488 4563 1492
rect 4509 1328 4515 1472
rect 4653 1428 4659 1532
rect 4685 1528 4691 1552
rect 4589 1328 4595 1392
rect 4605 1328 4611 1332
rect 3917 1148 3923 1272
rect 3933 1268 3939 1272
rect 3997 1268 4003 1272
rect 4077 1268 4083 1272
rect 3949 1123 3955 1232
rect 3949 1117 3960 1123
rect 3789 1088 3795 1092
rect 3821 1068 3827 1072
rect 3853 988 3859 1032
rect 3853 928 3859 952
rect 3789 883 3795 912
rect 3869 908 3875 1092
rect 3789 877 3811 883
rect 3645 688 3651 712
rect 3741 708 3747 712
rect 3805 688 3811 877
rect 3885 883 3891 1112
rect 3901 1088 3907 1092
rect 3917 943 3923 1092
rect 3933 1088 3939 1112
rect 3981 1088 3987 1152
rect 4093 1128 4099 1292
rect 4109 1268 4115 1292
rect 4205 1288 4211 1292
rect 4109 1148 4115 1152
rect 4237 1148 4243 1232
rect 4013 1028 4019 1112
rect 4269 1108 4275 1112
rect 4061 1088 4067 1092
rect 4253 1068 4259 1092
rect 4317 1068 4323 1092
rect 3917 937 3939 943
rect 3933 928 3939 937
rect 3933 908 3939 912
rect 3965 908 3971 912
rect 3885 877 3896 883
rect 3837 748 3843 872
rect 3981 788 3987 1012
rect 4029 1008 4035 1032
rect 4077 948 4083 952
rect 4125 928 4131 932
rect 3853 728 3859 752
rect 3901 728 3907 752
rect 3997 748 4003 872
rect 3821 708 3827 712
rect 3901 708 3907 712
rect 3997 708 4003 712
rect 4045 708 4051 912
rect 4061 908 4067 912
rect 4077 888 4083 912
rect 4189 908 4195 1032
rect 4253 948 4259 952
rect 4061 708 4067 792
rect 4109 788 4115 892
rect 4125 748 4131 872
rect 4157 788 4163 892
rect 4237 888 4243 892
rect 4253 888 4259 912
rect 4269 908 4275 912
rect 4301 908 4307 1032
rect 4317 928 4323 1052
rect 4333 908 4339 912
rect 4349 903 4355 1232
rect 4365 1228 4371 1232
rect 4397 1148 4403 1272
rect 4413 1188 4419 1292
rect 4445 1248 4451 1272
rect 4413 1123 4419 1172
rect 4461 1168 4467 1232
rect 4477 1228 4483 1292
rect 4509 1208 4515 1272
rect 4525 1268 4531 1272
rect 4621 1268 4627 1332
rect 4408 1117 4419 1123
rect 4445 1123 4451 1152
rect 4525 1128 4531 1212
rect 4541 1208 4547 1232
rect 4557 1168 4563 1232
rect 4653 1223 4659 1412
rect 4669 1388 4675 1492
rect 4685 1308 4691 1312
rect 4685 1288 4691 1292
rect 4653 1217 4675 1223
rect 4669 1168 4675 1217
rect 4557 1148 4563 1152
rect 4669 1148 4675 1152
rect 4445 1117 4456 1123
rect 4685 1123 4691 1272
rect 4701 1128 4707 1492
rect 4733 1488 4739 1492
rect 4749 1488 4755 1652
rect 4797 1528 4803 1632
rect 4733 1388 4739 1452
rect 4669 1117 4691 1123
rect 4381 1048 4387 1092
rect 4413 1068 4419 1072
rect 4413 988 4419 992
rect 4349 897 4371 903
rect 4269 788 4275 872
rect 4317 828 4323 892
rect 4349 868 4355 872
rect 4141 728 4147 752
rect 4285 728 4291 752
rect 4333 748 4339 832
rect 3789 668 3795 672
rect 3693 588 3699 652
rect 3773 568 3779 632
rect 3709 528 3715 532
rect 3725 528 3731 532
rect 3709 428 3715 512
rect 3773 508 3779 532
rect 3725 428 3731 432
rect 3533 168 3539 292
rect 3629 208 3635 312
rect 3645 228 3651 232
rect 3549 148 3555 192
rect 3565 128 3571 192
rect 3677 188 3683 312
rect 3709 288 3715 392
rect 3757 328 3763 332
rect 3789 328 3795 632
rect 3805 408 3811 532
rect 3821 528 3827 532
rect 3837 528 3843 692
rect 3853 668 3859 692
rect 3821 308 3827 492
rect 3853 448 3859 652
rect 3901 588 3907 632
rect 3933 588 3939 672
rect 3981 648 3987 692
rect 4045 688 4051 692
rect 4109 688 4115 692
rect 3869 508 3875 512
rect 3901 308 3907 552
rect 3949 528 3955 532
rect 3917 328 3923 352
rect 3981 288 3987 512
rect 3997 308 4003 412
rect 4029 368 4035 632
rect 4109 568 4115 672
rect 4125 588 4131 692
rect 4157 668 4163 692
rect 4269 688 4275 692
rect 4301 648 4307 672
rect 4269 588 4275 612
rect 4301 588 4307 632
rect 4205 568 4211 572
rect 4157 528 4163 532
rect 4365 523 4371 897
rect 4381 848 4387 932
rect 4445 928 4451 1052
rect 4461 948 4467 1072
rect 4493 1028 4499 1092
rect 4509 1088 4515 1112
rect 4525 1108 4531 1112
rect 4509 1068 4515 1072
rect 4493 968 4499 972
rect 4509 968 4515 1052
rect 4541 1048 4547 1092
rect 4557 928 4563 932
rect 4589 928 4595 1032
rect 4621 1028 4627 1092
rect 4621 923 4627 1012
rect 4621 917 4643 923
rect 4413 888 4419 892
rect 4429 888 4435 892
rect 4381 708 4387 712
rect 4397 708 4403 712
rect 4397 628 4403 672
rect 4477 668 4483 832
rect 4413 548 4419 592
rect 4493 548 4499 912
rect 4589 748 4595 832
rect 4461 523 4467 532
rect 4477 528 4483 532
rect 4360 517 4371 523
rect 4445 517 4467 523
rect 4136 497 4147 503
rect 4077 408 4083 472
rect 4109 388 4115 392
rect 4141 388 4147 497
rect 3789 188 3795 272
rect 3821 268 3827 272
rect 3837 268 3843 272
rect 3869 128 3875 252
rect 3949 168 3955 272
rect 3981 188 3987 232
rect 3997 148 4003 172
rect 4077 128 4083 332
rect 4093 148 4099 272
rect 4125 248 4131 312
rect 4157 308 4163 512
rect 4301 488 4307 512
rect 4157 288 4163 292
rect 4269 288 4275 432
rect 4381 368 4387 432
rect 4445 388 4451 517
rect 4301 308 4307 312
rect 4317 288 4323 352
rect 4333 308 4339 332
rect 4381 328 4387 332
rect 4205 268 4211 272
rect 4237 248 4243 272
rect 4381 148 4387 272
rect 3565 108 3571 112
rect 4077 108 4083 112
rect 4397 108 4403 112
rect 3533 -43 3539 32
rect 4029 -43 4035 12
rect 4365 -43 4371 32
rect 4413 -43 4419 352
rect 4429 288 4435 292
rect 4509 268 4515 290
rect 4525 288 4531 532
rect 4541 508 4547 652
rect 4573 588 4579 632
rect 4637 628 4643 917
rect 4653 908 4659 992
rect 4669 728 4675 1117
rect 4749 1123 4755 1472
rect 4765 1468 4771 1512
rect 4829 1468 4835 1912
rect 4877 1908 4883 1912
rect 4909 1908 4915 2432
rect 4957 2308 4963 2412
rect 4973 2308 4979 2312
rect 4925 2188 4931 2232
rect 4925 2128 4931 2132
rect 4957 2128 4963 2152
rect 5005 2108 5011 2232
rect 5021 2228 5027 2532
rect 5053 2388 5059 2692
rect 5101 2548 5107 2632
rect 5101 2288 5107 2532
rect 5133 2348 5139 2752
rect 5165 2648 5171 2872
rect 5181 2428 5187 3092
rect 5261 3068 5267 3092
rect 5245 2948 5251 3052
rect 5245 2888 5251 2932
rect 5213 2688 5219 2712
rect 5261 2708 5267 2792
rect 5277 2688 5283 3872
rect 5293 3748 5299 3892
rect 5309 3888 5315 4032
rect 5373 3948 5379 4072
rect 5325 3748 5331 3812
rect 5309 3588 5315 3712
rect 5341 3708 5347 3912
rect 5389 3908 5395 4112
rect 5405 4108 5411 4212
rect 5421 4188 5427 4232
rect 5405 3988 5411 4052
rect 5421 3948 5427 4152
rect 5437 3968 5443 4272
rect 5453 4128 5459 4292
rect 5469 4068 5475 4512
rect 5485 4468 5491 4492
rect 5517 4428 5523 4672
rect 5613 4668 5619 4672
rect 5629 4628 5635 5032
rect 5661 5028 5667 5032
rect 5645 4948 5651 4952
rect 5661 4928 5667 5012
rect 5677 4988 5683 5072
rect 5805 5023 5811 5092
rect 5853 5028 5859 5032
rect 5789 5017 5811 5023
rect 5725 4968 5731 5012
rect 5789 4988 5795 5017
rect 5661 4728 5667 4732
rect 5693 4728 5699 4732
rect 5725 4728 5731 4952
rect 5757 4848 5763 4912
rect 5805 4848 5811 4932
rect 5821 4928 5827 4992
rect 5917 4988 5923 5092
rect 6013 5088 6019 5092
rect 6045 5088 6051 5337
rect 6317 5328 6323 5332
rect 6749 5328 6755 5332
rect 6109 5308 6115 5312
rect 6125 5308 6131 5312
rect 5933 4988 5939 4992
rect 5837 4768 5843 4952
rect 5917 4928 5923 4932
rect 5933 4928 5939 4972
rect 5949 4968 5955 4972
rect 6013 4948 6019 5072
rect 6045 5068 6051 5072
rect 5901 4908 5907 4912
rect 6029 4908 6035 4912
rect 5757 4748 5763 4752
rect 5533 4503 5539 4532
rect 5549 4528 5555 4612
rect 5581 4548 5587 4552
rect 5597 4528 5603 4572
rect 5661 4568 5667 4632
rect 5533 4497 5555 4503
rect 5533 4328 5539 4332
rect 5485 4148 5491 4232
rect 5501 4228 5507 4312
rect 5501 4128 5507 4192
rect 5533 4068 5539 4132
rect 5549 4108 5555 4497
rect 5565 4308 5571 4332
rect 5693 4328 5699 4712
rect 5581 4148 5587 4152
rect 5421 3848 5427 3932
rect 5517 3888 5523 3892
rect 5373 3708 5379 3752
rect 5405 3728 5411 3812
rect 5501 3768 5507 3852
rect 5533 3748 5539 3952
rect 5549 3748 5555 4092
rect 5597 3988 5603 4232
rect 5629 4228 5635 4232
rect 5677 4168 5683 4212
rect 5709 4148 5715 4692
rect 5757 4548 5763 4552
rect 5741 4488 5747 4512
rect 5773 4488 5779 4552
rect 5805 4548 5811 4612
rect 5821 4588 5827 4732
rect 5853 4728 5859 4772
rect 5901 4708 5907 4872
rect 5805 4528 5811 4532
rect 5837 4508 5843 4692
rect 5933 4668 5939 4672
rect 5741 4188 5747 4292
rect 5837 4288 5843 4492
rect 5853 4468 5859 4492
rect 5853 4328 5859 4352
rect 5885 4348 5891 4572
rect 5933 4488 5939 4652
rect 5885 4317 5896 4323
rect 5629 4128 5635 4132
rect 5757 4128 5763 4132
rect 5565 3748 5571 3932
rect 5629 3928 5635 4092
rect 5773 4088 5779 4112
rect 5645 4068 5651 4072
rect 5725 3906 5731 3912
rect 5597 3848 5603 3852
rect 5581 3748 5587 3752
rect 5517 3728 5523 3732
rect 5453 3668 5459 3672
rect 5293 3308 5299 3452
rect 5309 3408 5315 3572
rect 5325 3488 5331 3492
rect 5341 3468 5347 3612
rect 5389 3588 5395 3612
rect 5453 3488 5459 3632
rect 5293 3128 5299 3212
rect 5309 3128 5315 3392
rect 5341 3368 5347 3452
rect 5405 3328 5411 3432
rect 5485 3423 5491 3490
rect 5533 3468 5539 3732
rect 5469 3417 5491 3423
rect 5469 3388 5475 3417
rect 5549 3388 5555 3732
rect 5565 3728 5571 3732
rect 5597 3728 5603 3732
rect 5597 3608 5603 3692
rect 5661 3548 5667 3652
rect 5693 3648 5699 3872
rect 5709 3788 5715 3792
rect 5757 3723 5763 4072
rect 5789 3968 5795 4272
rect 5885 4268 5891 4317
rect 5901 4288 5907 4292
rect 5933 4288 5939 4292
rect 5805 4188 5811 4232
rect 5853 4208 5859 4232
rect 5869 4188 5875 4212
rect 5805 3908 5811 4032
rect 5789 3788 5795 3892
rect 5805 3888 5811 3892
rect 5805 3828 5811 3872
rect 5821 3768 5827 3832
rect 5837 3788 5843 3912
rect 5885 3868 5891 4252
rect 5901 4228 5907 4272
rect 5949 4228 5955 4832
rect 5981 4708 5987 4752
rect 6061 4708 6067 5212
rect 6125 5108 6131 5112
rect 6205 5088 6211 5132
rect 6509 5108 6515 5112
rect 6333 5088 6339 5092
rect 6445 5088 6451 5092
rect 6541 5088 6547 5092
rect 6141 4828 6147 4952
rect 6157 4748 6163 5032
rect 6285 4968 6291 4972
rect 6381 4948 6387 5072
rect 6413 5028 6419 5052
rect 6221 4928 6227 4932
rect 6205 4908 6211 4912
rect 6237 4868 6243 4912
rect 6397 4908 6403 4912
rect 6173 4728 6179 4792
rect 6237 4708 6243 4812
rect 6365 4708 6371 4872
rect 6413 4788 6419 5012
rect 6445 4848 6451 5072
rect 6509 4988 6515 5072
rect 6573 5068 6579 5090
rect 6621 5048 6627 5312
rect 6781 5108 6787 5332
rect 6797 5068 6803 5463
rect 6941 5368 6947 5372
rect 6813 5330 6819 5332
rect 6893 5288 6899 5332
rect 7069 5328 7075 5332
rect 6973 5288 6979 5312
rect 7053 5308 7059 5312
rect 7133 5108 7139 5272
rect 7277 5208 7283 5232
rect 7325 5148 7331 5232
rect 7325 5108 7331 5112
rect 6829 5088 6835 5092
rect 6877 5088 6883 5092
rect 6909 5048 6915 5052
rect 6701 5028 6707 5032
rect 6717 4988 6723 5032
rect 6573 4968 6579 4972
rect 6541 4928 6547 4932
rect 6557 4788 6563 4792
rect 6413 4728 6419 4772
rect 6445 4748 6451 4772
rect 6573 4763 6579 4952
rect 6589 4768 6595 4832
rect 6605 4788 6611 4912
rect 6685 4908 6691 4912
rect 6701 4908 6707 4932
rect 6765 4908 6771 4932
rect 6813 4908 6819 4912
rect 6829 4908 6835 4972
rect 6877 4908 6883 4912
rect 6909 4903 6915 5032
rect 6904 4897 6915 4903
rect 6637 4848 6643 4892
rect 6557 4757 6579 4763
rect 5965 4588 5971 4592
rect 6045 4548 6051 4672
rect 6093 4668 6099 4672
rect 6125 4628 6131 4672
rect 6125 4588 6131 4612
rect 5965 4528 5971 4532
rect 5981 4408 5987 4512
rect 6061 4488 6067 4532
rect 6077 4528 6083 4532
rect 6157 4528 6163 4652
rect 6029 4328 6035 4332
rect 6061 4328 6067 4352
rect 5981 4317 5992 4323
rect 5981 4268 5987 4317
rect 5997 4297 6008 4303
rect 5949 4188 5955 4212
rect 5997 4188 6003 4297
rect 5997 4148 6003 4172
rect 6029 4123 6035 4312
rect 6093 4283 6099 4472
rect 6125 4348 6131 4452
rect 6109 4308 6115 4312
rect 6093 4277 6104 4283
rect 6061 4148 6067 4232
rect 6013 4117 6035 4123
rect 5901 4108 5907 4112
rect 5869 3768 5875 3852
rect 5885 3808 5891 3852
rect 5965 3768 5971 3872
rect 5901 3728 5907 3732
rect 5981 3728 5987 3752
rect 5757 3717 5768 3723
rect 5725 3648 5731 3712
rect 5645 3468 5651 3492
rect 5565 3388 5571 3412
rect 5373 3308 5379 3312
rect 5421 3308 5427 3352
rect 5437 3328 5443 3332
rect 5453 3328 5459 3332
rect 5432 3297 5443 3303
rect 5389 3108 5395 3112
rect 5437 3008 5443 3297
rect 5453 3108 5459 3312
rect 5533 3308 5539 3352
rect 5581 3288 5587 3312
rect 5613 3308 5619 3432
rect 5517 3148 5523 3232
rect 5533 3188 5539 3252
rect 5597 3188 5603 3292
rect 5629 3168 5635 3312
rect 5693 3303 5699 3512
rect 5709 3508 5715 3532
rect 5757 3528 5763 3572
rect 5773 3548 5779 3552
rect 5725 3328 5731 3512
rect 5741 3388 5747 3492
rect 5773 3468 5779 3492
rect 5773 3368 5779 3452
rect 5805 3388 5811 3632
rect 5821 3588 5827 3592
rect 5901 3588 5907 3692
rect 6013 3668 6019 4117
rect 6061 4108 6067 4112
rect 6061 3708 6067 4092
rect 6077 4008 6083 4112
rect 6093 4048 6099 4252
rect 6109 4068 6115 4272
rect 6093 3988 6099 4032
rect 6093 3908 6099 3972
rect 6125 3948 6131 4312
rect 6141 4308 6147 4392
rect 6157 4383 6163 4512
rect 6173 4468 6179 4492
rect 6189 4488 6195 4492
rect 6205 4388 6211 4492
rect 6237 4428 6243 4532
rect 6301 4528 6307 4692
rect 6285 4468 6291 4492
rect 6157 4377 6179 4383
rect 6173 4348 6179 4377
rect 6157 4308 6163 4332
rect 6205 4308 6211 4332
rect 6269 4328 6275 4352
rect 6285 4328 6291 4452
rect 6301 4408 6307 4512
rect 6317 4488 6323 4552
rect 6349 4463 6355 4672
rect 6445 4508 6451 4512
rect 6461 4508 6467 4532
rect 6397 4488 6403 4492
rect 6493 4488 6499 4732
rect 6557 4728 6563 4757
rect 6653 4763 6659 4892
rect 6733 4848 6739 4872
rect 6669 4788 6675 4832
rect 6637 4757 6659 4763
rect 6584 4737 6595 4743
rect 6509 4668 6515 4692
rect 6509 4508 6515 4512
rect 6520 4497 6531 4503
rect 6333 4457 6355 4463
rect 6333 4428 6339 4457
rect 6173 4108 6179 4192
rect 6205 4128 6211 4292
rect 6317 4288 6323 4292
rect 6333 4288 6339 4412
rect 6429 4348 6435 4472
rect 6461 4328 6467 4332
rect 6221 4228 6227 4252
rect 6365 4248 6371 4272
rect 6413 4268 6419 4312
rect 6445 4268 6451 4292
rect 6285 4228 6291 4232
rect 6525 4228 6531 4497
rect 6557 4408 6563 4692
rect 6573 4528 6579 4672
rect 6589 4628 6595 4737
rect 6637 4708 6643 4757
rect 6685 4748 6691 4792
rect 6701 4748 6707 4812
rect 6733 4788 6739 4832
rect 6749 4748 6755 4832
rect 6797 4808 6803 4872
rect 6941 4868 6947 4912
rect 6957 4908 6963 4972
rect 6637 4688 6643 4692
rect 6589 4508 6595 4572
rect 6621 4488 6627 4552
rect 6685 4508 6691 4732
rect 6781 4728 6787 4772
rect 6813 4728 6819 4832
rect 6877 4748 6883 4832
rect 6941 4768 6947 4832
rect 6957 4748 6963 4872
rect 6989 4848 6995 4872
rect 7005 4868 7011 4912
rect 7021 4908 7027 5052
rect 7037 5048 7043 5090
rect 7133 5088 7139 5092
rect 7149 4948 7155 5092
rect 7197 5008 7203 5092
rect 7245 5068 7251 5092
rect 7293 5068 7299 5072
rect 7213 4988 7219 5052
rect 7005 4783 7011 4832
rect 7005 4777 7027 4783
rect 6701 4688 6707 4692
rect 6717 4648 6723 4712
rect 6765 4668 6771 4692
rect 6829 4628 6835 4732
rect 6877 4708 6883 4712
rect 6925 4648 6931 4712
rect 6957 4703 6963 4732
rect 6989 4728 6995 4752
rect 7005 4708 7011 4752
rect 7021 4748 7027 4777
rect 6957 4697 6979 4703
rect 6701 4528 6707 4552
rect 6749 4528 6755 4532
rect 6637 4488 6643 4492
rect 6765 4488 6771 4612
rect 6877 4608 6883 4632
rect 6797 4568 6803 4572
rect 6797 4508 6803 4552
rect 6685 4468 6691 4472
rect 6717 4448 6723 4472
rect 6765 4468 6771 4472
rect 6653 4328 6659 4392
rect 6797 4368 6803 4472
rect 6813 4463 6819 4512
rect 6877 4488 6883 4532
rect 6925 4488 6931 4512
rect 6813 4457 6835 4463
rect 6664 4317 6675 4323
rect 6285 4128 6291 4152
rect 6413 4148 6419 4212
rect 6429 4148 6435 4152
rect 6221 3988 6227 4112
rect 6093 3788 6099 3792
rect 6109 3748 6115 3872
rect 6157 3868 6163 3932
rect 6301 3908 6307 4012
rect 6333 3988 6339 4092
rect 6125 3788 6131 3852
rect 6205 3788 6211 3892
rect 5837 3548 5843 3552
rect 5853 3428 5859 3492
rect 5885 3388 5891 3512
rect 5901 3368 5907 3492
rect 5837 3328 5843 3332
rect 5773 3308 5779 3312
rect 5693 3297 5715 3303
rect 5645 3248 5651 3272
rect 5677 3188 5683 3232
rect 5693 3228 5699 3272
rect 5709 3188 5715 3297
rect 5757 3268 5763 3272
rect 5789 3188 5795 3292
rect 5805 3277 5816 3283
rect 5805 3248 5811 3277
rect 5837 3263 5843 3292
rect 5853 3288 5859 3352
rect 5821 3257 5843 3263
rect 5821 3188 5827 3257
rect 5581 3148 5587 3152
rect 5485 3108 5491 3132
rect 5453 3088 5459 3092
rect 5405 2968 5411 2972
rect 5437 2928 5443 2992
rect 5453 2948 5459 3072
rect 5485 3068 5491 3092
rect 5293 2868 5299 2912
rect 5245 2588 5251 2612
rect 5261 2528 5267 2672
rect 5277 2608 5283 2672
rect 5277 2548 5283 2552
rect 5309 2528 5315 2692
rect 5325 2628 5331 2652
rect 5325 2568 5331 2612
rect 5389 2588 5395 2912
rect 5421 2888 5427 2892
rect 5453 2888 5459 2892
rect 5357 2528 5363 2552
rect 5213 2328 5219 2332
rect 5261 2308 5267 2512
rect 5389 2488 5395 2572
rect 5405 2528 5411 2732
rect 5437 2728 5443 2832
rect 5485 2828 5491 2912
rect 5517 2908 5523 3132
rect 5533 3108 5539 3112
rect 5549 3108 5555 3112
rect 5581 3088 5587 3132
rect 5597 3128 5603 3152
rect 5597 3108 5603 3112
rect 5613 3068 5619 3112
rect 5629 3108 5635 3112
rect 5549 2928 5555 2932
rect 5661 2928 5667 3132
rect 5693 3068 5699 3112
rect 5421 2628 5427 2692
rect 5021 2188 5027 2192
rect 5069 2188 5075 2212
rect 5101 2168 5107 2272
rect 5117 2248 5123 2292
rect 5133 2188 5139 2272
rect 5037 2048 5043 2112
rect 5149 2048 5155 2252
rect 5037 1983 5043 2032
rect 5149 1988 5155 2032
rect 5037 1977 5048 1983
rect 4941 1917 4952 1923
rect 4893 1868 4899 1872
rect 4845 1728 4851 1832
rect 4893 1788 4899 1852
rect 4909 1768 4915 1872
rect 4941 1788 4947 1917
rect 4973 1908 4979 1932
rect 4973 1768 4979 1872
rect 4989 1788 4995 1852
rect 4925 1748 4931 1752
rect 4989 1703 4995 1712
rect 5005 1708 5011 1812
rect 5021 1788 5027 1912
rect 5181 1908 5187 2292
rect 5261 2288 5267 2292
rect 5213 2148 5219 2152
rect 5101 1808 5107 1872
rect 5117 1748 5123 1852
rect 5181 1848 5187 1852
rect 5181 1748 5187 1792
rect 5229 1748 5235 1752
rect 5085 1728 5091 1732
rect 5037 1708 5043 1712
rect 5149 1708 5155 1712
rect 4984 1697 4995 1703
rect 4845 1688 4851 1692
rect 4989 1588 4995 1697
rect 4909 1508 4915 1552
rect 4957 1508 4963 1512
rect 5005 1488 5011 1692
rect 5021 1688 5027 1692
rect 5197 1688 5203 1692
rect 5229 1648 5235 1732
rect 5053 1508 5059 1572
rect 5069 1528 5075 1632
rect 5101 1488 5107 1632
rect 5117 1508 5123 1612
rect 4765 1308 4771 1432
rect 4829 1428 4835 1432
rect 4877 1408 4883 1432
rect 4925 1428 4931 1432
rect 4973 1408 4979 1452
rect 4925 1388 4931 1392
rect 4845 1328 4851 1332
rect 4797 1148 4803 1152
rect 4829 1128 4835 1172
rect 4989 1148 4995 1172
rect 5005 1168 5011 1472
rect 5053 1330 5059 1472
rect 5133 1388 5139 1512
rect 5165 1508 5171 1532
rect 5181 1488 5187 1632
rect 5261 1488 5267 2272
rect 5325 2268 5331 2312
rect 5373 2308 5379 2432
rect 5389 2368 5395 2472
rect 5405 2308 5411 2512
rect 5421 2508 5427 2592
rect 5437 2588 5443 2672
rect 5453 2668 5459 2712
rect 5485 2688 5491 2812
rect 5501 2748 5507 2832
rect 5581 2748 5587 2872
rect 5645 2788 5651 2912
rect 5693 2908 5699 2912
rect 5709 2908 5715 2952
rect 5677 2888 5683 2892
rect 5501 2568 5507 2732
rect 5517 2608 5523 2692
rect 5533 2668 5539 2712
rect 5677 2708 5683 2852
rect 5693 2728 5699 2832
rect 5709 2788 5715 2872
rect 5725 2848 5731 3132
rect 5741 2928 5747 3092
rect 5773 3088 5779 3132
rect 5789 3108 5795 3112
rect 5789 3003 5795 3092
rect 5805 3028 5811 3112
rect 5853 3108 5859 3272
rect 5885 3228 5891 3272
rect 5789 2997 5811 3003
rect 5805 2928 5811 2997
rect 5757 2888 5763 2912
rect 5805 2908 5811 2912
rect 5789 2848 5795 2892
rect 5821 2888 5827 3072
rect 5869 3028 5875 3112
rect 5885 3108 5891 3192
rect 5901 3128 5907 3312
rect 5917 3288 5923 3532
rect 6045 3463 6051 3492
rect 6061 3488 6067 3672
rect 6045 3457 6067 3463
rect 5949 3388 5955 3432
rect 6061 3388 6067 3457
rect 5997 3368 6003 3372
rect 6093 3328 6099 3392
rect 6109 3348 6115 3732
rect 6173 3728 6179 3732
rect 6157 3628 6163 3712
rect 6125 3388 6131 3412
rect 6173 3328 6179 3692
rect 6189 3628 6195 3672
rect 6221 3668 6227 3872
rect 6237 3748 6243 3752
rect 6301 3748 6307 3892
rect 6333 3868 6339 3972
rect 6349 3948 6355 4112
rect 6365 4028 6371 4072
rect 6445 4028 6451 4112
rect 6461 3968 6467 4172
rect 6525 4148 6531 4192
rect 6621 4188 6627 4272
rect 6541 4128 6547 4152
rect 6653 4128 6659 4132
rect 6669 4128 6675 4317
rect 6685 4288 6691 4352
rect 6733 4348 6739 4352
rect 6797 4348 6803 4352
rect 6717 4203 6723 4332
rect 6733 4228 6739 4292
rect 6749 4248 6755 4312
rect 6829 4288 6835 4457
rect 6845 4348 6851 4472
rect 6957 4343 6963 4512
rect 6973 4348 6979 4697
rect 6989 4548 6995 4692
rect 6952 4337 6963 4343
rect 6845 4243 6851 4332
rect 6861 4268 6867 4292
rect 6845 4237 6867 4243
rect 6717 4197 6739 4203
rect 6685 4128 6691 4132
rect 6461 3908 6467 3952
rect 6461 3768 6467 3892
rect 6493 3808 6499 4052
rect 6541 3908 6547 4052
rect 6589 3988 6595 4092
rect 6589 3888 6595 3892
rect 6621 3888 6627 4072
rect 6733 3948 6739 4197
rect 6845 4108 6851 4112
rect 6781 3988 6787 3992
rect 6749 3948 6755 3952
rect 6637 3928 6643 3932
rect 6205 3648 6211 3652
rect 6189 3508 6195 3612
rect 6205 3548 6211 3632
rect 6269 3608 6275 3692
rect 6349 3528 6355 3532
rect 6365 3528 6371 3712
rect 6413 3708 6419 3712
rect 6381 3688 6387 3692
rect 6205 3488 6211 3492
rect 5949 3288 5955 3312
rect 6029 3268 6035 3312
rect 5901 3088 5907 3092
rect 5741 2788 5747 2792
rect 5757 2728 5763 2732
rect 5805 2723 5811 2832
rect 5853 2808 5859 2832
rect 5869 2768 5875 2872
rect 5885 2748 5891 2912
rect 5901 2888 5907 3072
rect 5917 2908 5923 2952
rect 5933 2943 5939 3212
rect 5965 3083 5971 3092
rect 5960 3077 5971 3083
rect 6061 2948 6067 3252
rect 6093 3128 6099 3312
rect 6157 3248 6163 3312
rect 6173 3208 6179 3312
rect 6205 3228 6211 3472
rect 6285 3388 6291 3512
rect 6333 3428 6339 3492
rect 6333 3368 6339 3412
rect 6365 3383 6371 3432
rect 6349 3377 6371 3383
rect 6285 3348 6291 3352
rect 6349 3348 6355 3377
rect 6397 3348 6403 3392
rect 6429 3383 6435 3712
rect 6445 3588 6451 3652
rect 6413 3377 6435 3383
rect 6413 3328 6419 3377
rect 6429 3348 6435 3352
rect 6381 3108 6387 3112
rect 6397 3108 6403 3292
rect 6429 3188 6435 3252
rect 6461 3208 6467 3752
rect 6477 3508 6483 3512
rect 6477 3308 6483 3492
rect 6493 3488 6499 3792
rect 6541 3728 6547 3752
rect 6557 3508 6563 3512
rect 6573 3508 6579 3832
rect 6605 3828 6611 3872
rect 6637 3848 6643 3912
rect 6621 3808 6627 3832
rect 6685 3788 6691 3832
rect 6701 3748 6707 3892
rect 6733 3848 6739 3932
rect 6765 3868 6771 3912
rect 6813 3908 6819 3952
rect 6861 3948 6867 4237
rect 6925 4228 6931 4292
rect 6909 4148 6915 4172
rect 6957 4088 6963 4337
rect 6989 4308 6995 4532
rect 7069 4528 7075 4732
rect 7085 4668 7091 4692
rect 7085 4508 7091 4512
rect 7037 4388 7043 4412
rect 7053 4348 7059 4352
rect 7101 4348 7107 4872
rect 7245 4848 7251 5052
rect 7277 4928 7283 5032
rect 7293 4928 7299 4992
rect 7309 4903 7315 5072
rect 7293 4897 7315 4903
rect 7149 4628 7155 4732
rect 7181 4708 7187 4832
rect 7165 4697 7176 4703
rect 7133 4548 7139 4552
rect 7165 4488 7171 4697
rect 7213 4648 7219 4652
rect 7197 4588 7203 4632
rect 7277 4568 7283 4652
rect 7165 4408 7171 4432
rect 7181 4348 7187 4532
rect 6973 4128 6979 4212
rect 6989 4148 6995 4292
rect 6877 3908 6883 3992
rect 6941 3968 6947 4032
rect 6957 4028 6963 4072
rect 6973 4008 6979 4112
rect 6765 3788 6771 3832
rect 6813 3788 6819 3872
rect 6589 3688 6595 3712
rect 6669 3508 6675 3592
rect 6493 3328 6499 3412
rect 6541 3288 6547 3452
rect 6573 3323 6579 3492
rect 6589 3388 6595 3452
rect 6701 3408 6707 3732
rect 6717 3703 6723 3712
rect 6717 3697 6739 3703
rect 6717 3448 6723 3472
rect 6717 3368 6723 3432
rect 6733 3388 6739 3697
rect 6765 3548 6771 3632
rect 6845 3628 6851 3712
rect 6781 3488 6787 3512
rect 6765 3388 6771 3432
rect 6781 3368 6787 3472
rect 6717 3328 6723 3352
rect 6568 3317 6579 3323
rect 6477 3268 6483 3272
rect 6461 3108 6467 3192
rect 6653 3188 6659 3232
rect 6733 3188 6739 3252
rect 6733 3168 6739 3172
rect 6781 3148 6787 3312
rect 6797 3228 6803 3492
rect 6829 3388 6835 3492
rect 6861 3343 6867 3712
rect 6877 3583 6883 3892
rect 6893 3848 6899 3912
rect 6957 3848 6963 3912
rect 6941 3728 6947 3732
rect 6957 3728 6963 3792
rect 6973 3788 6979 3952
rect 6989 3908 6995 3992
rect 7005 3968 7011 4312
rect 7037 4308 7043 4332
rect 7037 4088 7043 4212
rect 7085 4188 7091 4252
rect 7021 4008 7027 4032
rect 7053 3948 7059 3952
rect 7069 3928 7075 3932
rect 7101 3928 7107 4332
rect 7133 4308 7139 4312
rect 7117 4288 7123 4292
rect 7133 4248 7139 4292
rect 7165 4228 7171 4332
rect 7277 4308 7283 4552
rect 7181 4288 7187 4292
rect 7213 4248 7219 4292
rect 7277 4288 7283 4292
rect 7213 4228 7219 4232
rect 7229 4188 7235 4272
rect 7261 4168 7267 4212
rect 7133 4128 7139 4152
rect 7197 4128 7203 4152
rect 7293 4128 7299 4897
rect 7117 4068 7123 4112
rect 7037 3888 7043 3912
rect 7037 3868 7043 3872
rect 7101 3868 7107 3872
rect 7117 3803 7123 4052
rect 7133 3908 7139 3912
rect 7181 3888 7187 3912
rect 7149 3808 7155 3872
rect 7101 3797 7123 3803
rect 6973 3768 6979 3772
rect 6925 3708 6931 3712
rect 7053 3708 7059 3712
rect 6941 3588 6947 3592
rect 6877 3577 6899 3583
rect 6877 3508 6883 3532
rect 6893 3508 6899 3577
rect 6909 3428 6915 3512
rect 6941 3508 6947 3552
rect 6957 3548 6963 3592
rect 6989 3588 6995 3592
rect 7101 3548 7107 3797
rect 7165 3788 7171 3872
rect 7069 3528 7075 3532
rect 6845 3337 6867 3343
rect 6157 3088 6163 3092
rect 6189 3088 6195 3092
rect 6221 3028 6227 3052
rect 6269 3048 6275 3092
rect 6157 2968 6163 2972
rect 6317 2948 6323 3072
rect 6333 3068 6339 3072
rect 6349 2948 6355 3032
rect 5933 2937 5955 2943
rect 5949 2888 5955 2937
rect 6141 2928 6147 2932
rect 6317 2928 6323 2932
rect 6029 2888 6035 2912
rect 5933 2743 5939 2832
rect 5949 2748 5955 2872
rect 6045 2828 6051 2912
rect 6333 2828 6339 2872
rect 6205 2788 6211 2792
rect 5917 2737 5939 2743
rect 5917 2728 5923 2737
rect 5800 2717 5811 2723
rect 5773 2708 5779 2712
rect 5565 2668 5571 2692
rect 5629 2688 5635 2692
rect 5869 2688 5875 2692
rect 5885 2688 5891 2692
rect 5533 2648 5539 2652
rect 5885 2648 5891 2672
rect 5565 2628 5571 2632
rect 5533 2528 5539 2592
rect 5549 2508 5555 2512
rect 5421 2328 5427 2492
rect 5517 2348 5523 2472
rect 5581 2388 5587 2472
rect 5597 2468 5603 2512
rect 5645 2488 5651 2552
rect 5661 2528 5667 2592
rect 5709 2588 5715 2632
rect 5837 2603 5843 2632
rect 5821 2597 5843 2603
rect 5709 2548 5715 2572
rect 5709 2523 5715 2532
rect 5704 2517 5715 2523
rect 5565 2348 5571 2352
rect 5357 2288 5363 2292
rect 5437 2288 5443 2292
rect 5277 2128 5283 2152
rect 5309 2148 5315 2252
rect 5277 1788 5283 2072
rect 5357 1888 5363 2272
rect 5405 2168 5411 2232
rect 5453 2128 5459 2212
rect 5469 2188 5475 2252
rect 5485 2248 5491 2312
rect 5581 2308 5587 2352
rect 5597 2348 5603 2432
rect 5485 2208 5491 2232
rect 5293 1848 5299 1852
rect 5293 1708 5299 1832
rect 5357 1788 5363 1872
rect 5389 1788 5395 2092
rect 5357 1748 5363 1752
rect 5309 1708 5315 1712
rect 5277 1488 5283 1492
rect 5181 1368 5187 1472
rect 5117 1348 5123 1352
rect 4749 1117 4771 1123
rect 4685 1048 4691 1092
rect 4701 948 4707 1072
rect 4749 1028 4755 1092
rect 4765 1088 4771 1117
rect 5085 1108 5091 1332
rect 5261 1328 5267 1392
rect 4765 948 4771 1052
rect 4813 1048 4819 1092
rect 4813 968 4819 972
rect 4845 928 4851 932
rect 4781 908 4787 912
rect 4861 888 4867 1032
rect 4877 1028 4883 1092
rect 4973 1088 4979 1092
rect 4893 1068 4899 1072
rect 4909 1068 4915 1072
rect 5021 1048 5027 1052
rect 4925 888 4931 992
rect 4669 708 4675 712
rect 4701 688 4707 732
rect 4557 508 4563 552
rect 4573 548 4579 572
rect 4669 548 4675 572
rect 4701 568 4707 672
rect 4637 508 4643 512
rect 4541 288 4547 492
rect 4749 388 4755 872
rect 4829 688 4835 692
rect 4637 308 4643 332
rect 4653 308 4659 312
rect 4429 168 4435 252
rect 4541 208 4547 272
rect 4493 168 4499 172
rect 4621 168 4627 192
rect 4445 148 4451 152
rect 4653 -43 4659 292
rect 4685 248 4691 272
rect 4685 148 4691 232
rect 4717 188 4723 312
rect 4781 308 4787 652
rect 4797 508 4803 512
rect 4845 508 4851 652
rect 4877 568 4883 832
rect 4909 708 4915 732
rect 4925 668 4931 792
rect 4941 768 4947 832
rect 5005 748 5011 1032
rect 5037 928 5043 1052
rect 5069 988 5075 1012
rect 5085 988 5091 1092
rect 5181 1043 5187 1292
rect 5277 1128 5283 1472
rect 5357 1348 5363 1492
rect 5389 1468 5395 1632
rect 5405 1188 5411 2112
rect 5469 2108 5475 2132
rect 5421 1948 5427 2032
rect 5517 1923 5523 2232
rect 5597 2188 5603 2312
rect 5613 2308 5619 2392
rect 5661 2368 5667 2512
rect 5725 2508 5731 2552
rect 5789 2448 5795 2512
rect 5805 2348 5811 2432
rect 5645 2308 5651 2312
rect 5677 2268 5683 2272
rect 5613 2248 5619 2252
rect 5533 2128 5539 2132
rect 5565 2128 5571 2132
rect 5613 2103 5619 2232
rect 5629 2168 5635 2232
rect 5709 2148 5715 2272
rect 5741 2168 5747 2172
rect 5821 2148 5827 2597
rect 5853 2448 5859 2532
rect 5965 2528 5971 2692
rect 5981 2668 5987 2732
rect 6013 2608 6019 2692
rect 6093 2688 6099 2692
rect 6109 2688 6115 2692
rect 6173 2668 6179 2712
rect 6333 2708 6339 2812
rect 6237 2668 6243 2672
rect 6013 2588 6019 2592
rect 5869 2468 5875 2512
rect 5853 2308 5859 2412
rect 5917 2328 5923 2332
rect 5853 2228 5859 2292
rect 5917 2268 5923 2312
rect 5709 2128 5715 2132
rect 5608 2097 5619 2103
rect 5512 1917 5523 1923
rect 5565 1888 5571 1952
rect 5597 1923 5603 2032
rect 5597 1917 5608 1923
rect 5469 1788 5475 1832
rect 5501 1808 5507 1832
rect 5533 1788 5539 1872
rect 5549 1848 5555 1872
rect 5597 1868 5603 1872
rect 5565 1768 5571 1792
rect 5485 1748 5491 1752
rect 5597 1728 5603 1792
rect 5533 1688 5539 1692
rect 5453 1628 5459 1632
rect 5421 1506 5427 1512
rect 5485 1488 5491 1532
rect 5517 1508 5523 1512
rect 5453 1388 5459 1392
rect 5421 1368 5427 1372
rect 5469 1328 5475 1332
rect 5469 1148 5475 1312
rect 5485 1208 5491 1312
rect 5517 1308 5523 1312
rect 5277 1108 5283 1112
rect 5245 1088 5251 1092
rect 5437 1088 5443 1112
rect 5213 1068 5219 1072
rect 5181 1037 5203 1043
rect 5181 968 5187 972
rect 5021 888 5027 912
rect 5005 708 5011 712
rect 4877 503 4883 532
rect 4925 528 4931 552
rect 4909 508 4915 512
rect 4861 497 4883 503
rect 4829 388 4835 412
rect 4861 288 4867 497
rect 4877 388 4883 432
rect 4893 323 4899 432
rect 4893 317 4904 323
rect 4717 108 4723 152
rect 4797 128 4803 132
rect 4733 108 4739 112
rect 4813 -43 4819 232
rect 4845 188 4851 252
rect 4877 188 4883 292
rect 4941 28 4947 632
rect 4957 588 4963 652
rect 4989 648 4995 672
rect 4989 508 4995 532
rect 4957 268 4963 432
rect 4989 388 4995 492
rect 5021 308 5027 872
rect 5069 848 5075 892
rect 5085 728 5091 932
rect 5101 928 5107 952
rect 5117 788 5123 852
rect 5101 708 5107 732
rect 5117 708 5123 712
rect 5053 688 5059 692
rect 5117 688 5123 692
rect 5037 528 5043 552
rect 5117 548 5123 672
rect 5133 648 5139 892
rect 5181 588 5187 932
rect 5037 308 5043 312
rect 5133 308 5139 312
rect 5085 288 5091 292
rect 5197 288 5203 1037
rect 5357 988 5363 1072
rect 5245 928 5251 972
rect 5373 948 5379 952
rect 5341 688 5347 932
rect 5405 928 5411 932
rect 5437 768 5443 1072
rect 5453 928 5459 1092
rect 5485 948 5491 1192
rect 5533 1128 5539 1452
rect 5549 1388 5555 1452
rect 5597 1388 5603 1692
rect 5613 1508 5619 1772
rect 5629 1708 5635 1832
rect 5645 1648 5651 2112
rect 5661 1748 5667 1972
rect 5821 1888 5827 2132
rect 5917 1908 5923 2212
rect 5965 2128 5971 2512
rect 5981 2508 5987 2572
rect 6061 2488 6067 2632
rect 6141 2628 6147 2632
rect 6189 2528 6195 2532
rect 6301 2528 6307 2632
rect 6365 2568 6371 3072
rect 6381 2988 6387 3052
rect 6397 2728 6403 3092
rect 6525 3003 6531 3132
rect 6509 2997 6531 3003
rect 6493 2928 6499 2932
rect 6445 2768 6451 2912
rect 6445 2708 6451 2752
rect 6397 2623 6403 2690
rect 6381 2617 6403 2623
rect 6381 2588 6387 2617
rect 6365 2548 6371 2552
rect 6413 2528 6419 2552
rect 6077 2508 6083 2512
rect 6029 2368 6035 2472
rect 6045 2388 6051 2432
rect 5981 2048 5987 2112
rect 6013 2108 6019 2172
rect 5997 2068 6003 2092
rect 6045 2088 6051 2232
rect 6061 2088 6067 2432
rect 6077 2388 6083 2432
rect 6125 2408 6131 2492
rect 6141 2468 6147 2472
rect 6077 2308 6083 2332
rect 6093 2088 6099 2352
rect 6157 2348 6163 2472
rect 6205 2468 6211 2492
rect 6221 2448 6227 2472
rect 6109 2268 6115 2332
rect 5933 1948 5939 1972
rect 5933 1908 5939 1932
rect 5949 1908 5955 2032
rect 6045 1988 6051 2032
rect 6061 1948 6067 2072
rect 6109 1968 6115 2112
rect 6141 2108 6147 2172
rect 6125 2088 6131 2092
rect 6173 2088 6179 2252
rect 6189 2248 6195 2332
rect 6237 2328 6243 2332
rect 6253 2308 6259 2392
rect 6269 2328 6275 2432
rect 6301 2368 6307 2472
rect 6349 2428 6355 2512
rect 6445 2508 6451 2552
rect 6477 2528 6483 2572
rect 6365 2308 6371 2452
rect 6397 2348 6403 2372
rect 6413 2308 6419 2372
rect 6477 2328 6483 2432
rect 6493 2428 6499 2472
rect 6493 2308 6499 2312
rect 6509 2308 6515 2997
rect 6573 2948 6579 3072
rect 6589 3023 6595 3090
rect 6589 3017 6611 3023
rect 6605 2988 6611 3017
rect 6637 2968 6643 3032
rect 6653 2988 6659 3092
rect 6589 2928 6595 2932
rect 6685 2928 6691 2952
rect 6717 2928 6723 2932
rect 6733 2928 6739 3112
rect 6765 3108 6771 3112
rect 6797 3108 6803 3212
rect 6781 3083 6787 3092
rect 6765 3077 6787 3083
rect 6573 2908 6579 2912
rect 6765 2908 6771 3077
rect 6781 2988 6787 2992
rect 6797 2963 6803 3072
rect 6813 2988 6819 3292
rect 6845 3108 6851 3337
rect 6909 3328 6915 3332
rect 6813 2968 6819 2972
rect 6781 2957 6803 2963
rect 6525 2508 6531 2632
rect 6573 2568 6579 2632
rect 6573 2548 6579 2552
rect 6589 2528 6595 2592
rect 6605 2528 6611 2672
rect 6525 2408 6531 2432
rect 6557 2308 6563 2512
rect 6621 2508 6627 2732
rect 6653 2708 6659 2772
rect 6685 2688 6691 2752
rect 6701 2548 6707 2612
rect 6749 2588 6755 2692
rect 6781 2548 6787 2957
rect 6813 2568 6819 2572
rect 6621 2488 6627 2492
rect 6605 2388 6611 2432
rect 6701 2428 6707 2532
rect 6781 2528 6787 2532
rect 6829 2528 6835 3092
rect 6845 2968 6851 3052
rect 6845 2928 6851 2952
rect 6861 2788 6867 3312
rect 6909 3288 6915 3312
rect 6941 3288 6947 3452
rect 6973 3308 6979 3412
rect 7021 3388 7027 3492
rect 7037 3408 7043 3512
rect 7117 3508 7123 3512
rect 7101 3368 7107 3492
rect 7117 3488 7123 3492
rect 7149 3468 7155 3552
rect 7149 3448 7155 3452
rect 7133 3348 7139 3432
rect 6989 3328 6995 3332
rect 6877 3068 6883 3132
rect 6893 2948 6899 2952
rect 6909 2928 6915 3232
rect 6941 3188 6947 3272
rect 6957 3268 6963 3272
rect 6973 3148 6979 3292
rect 6941 3106 6947 3112
rect 6941 2948 6947 3052
rect 6909 2908 6915 2912
rect 6989 2828 6995 3312
rect 6925 2708 6931 2812
rect 6989 2708 6995 2772
rect 6845 2588 6851 2632
rect 6957 2588 6963 2632
rect 6637 2348 6643 2352
rect 6573 2308 6579 2312
rect 6365 2288 6371 2292
rect 6221 2208 6227 2232
rect 6205 2108 6211 2172
rect 6365 2128 6371 2132
rect 6205 2088 6211 2092
rect 5853 1888 5859 1892
rect 5997 1888 6003 1892
rect 5629 1468 5635 1472
rect 5597 1328 5603 1372
rect 5581 1268 5587 1272
rect 5549 1188 5555 1212
rect 5517 1108 5523 1112
rect 5533 1108 5539 1112
rect 5533 928 5539 1092
rect 5565 948 5571 1072
rect 5613 1028 5619 1292
rect 5629 1188 5635 1432
rect 5661 1348 5667 1732
rect 5757 1728 5763 1772
rect 5821 1743 5827 1852
rect 5805 1737 5827 1743
rect 5677 1228 5683 1712
rect 5805 1708 5811 1737
rect 5725 1668 5731 1692
rect 5837 1688 5843 1832
rect 5757 1668 5763 1672
rect 5773 1648 5779 1672
rect 5725 1488 5731 1612
rect 5741 1508 5747 1512
rect 5693 1388 5699 1472
rect 5757 1468 5763 1472
rect 5741 1348 5747 1392
rect 5741 1308 5747 1312
rect 5757 1308 5763 1352
rect 5613 968 5619 1012
rect 5645 968 5651 1132
rect 5645 928 5651 952
rect 5693 948 5699 952
rect 5709 948 5715 1212
rect 5741 1108 5747 1292
rect 5789 1288 5795 1632
rect 5837 1543 5843 1672
rect 5885 1628 5891 1732
rect 5965 1728 5971 1832
rect 6029 1783 6035 1852
rect 6029 1777 6040 1783
rect 5981 1668 5987 1712
rect 6045 1708 6051 1772
rect 5965 1588 5971 1612
rect 5837 1537 5859 1543
rect 5837 1508 5843 1512
rect 5821 1388 5827 1492
rect 5821 1323 5827 1372
rect 5821 1317 5832 1323
rect 5853 1288 5859 1537
rect 5869 1468 5875 1532
rect 5901 1508 5907 1552
rect 5965 1488 5971 1572
rect 6045 1528 6051 1552
rect 6061 1543 6067 1932
rect 6077 1908 6083 1952
rect 6173 1848 6179 2072
rect 6189 1948 6195 2032
rect 6205 1908 6211 1992
rect 6269 1928 6275 2032
rect 6381 2028 6387 2232
rect 6461 2108 6467 2232
rect 6477 2108 6483 2172
rect 6589 2168 6595 2272
rect 6509 2148 6515 2152
rect 6557 2148 6563 2152
rect 6557 2128 6563 2132
rect 6445 1968 6451 2072
rect 6285 1908 6291 1952
rect 6349 1908 6355 1912
rect 6109 1828 6115 1832
rect 6093 1728 6099 1772
rect 6125 1728 6131 1792
rect 6173 1788 6179 1832
rect 6189 1788 6195 1872
rect 6205 1848 6211 1852
rect 6237 1748 6243 1752
rect 6173 1728 6179 1732
rect 6189 1688 6195 1692
rect 6221 1688 6227 1712
rect 6269 1688 6275 1772
rect 6301 1768 6307 1832
rect 6349 1788 6355 1852
rect 6077 1648 6083 1672
rect 6093 1668 6099 1672
rect 6061 1537 6072 1543
rect 5997 1508 6003 1512
rect 6045 1508 6051 1512
rect 6061 1508 6067 1512
rect 6008 1497 6019 1503
rect 5917 1388 5923 1452
rect 5901 1348 5907 1352
rect 5853 1268 5859 1272
rect 5773 1128 5779 1232
rect 5837 1128 5843 1232
rect 5869 1183 5875 1332
rect 5949 1328 5955 1352
rect 5885 1228 5891 1312
rect 5965 1188 5971 1472
rect 5981 1368 5987 1492
rect 5997 1328 6003 1472
rect 5869 1177 5891 1183
rect 5741 1043 5747 1072
rect 5741 1037 5763 1043
rect 5757 988 5763 1037
rect 5757 968 5763 972
rect 5709 928 5715 932
rect 5453 908 5459 912
rect 5357 588 5363 632
rect 5437 608 5443 672
rect 5229 548 5235 552
rect 5245 528 5251 552
rect 5325 548 5331 572
rect 5389 568 5395 592
rect 5453 583 5459 632
rect 5448 577 5459 583
rect 5389 548 5395 552
rect 5325 528 5331 532
rect 5213 508 5219 512
rect 4957 148 4963 232
rect 4973 168 4979 272
rect 4861 -43 4867 12
rect 4925 -43 4931 12
rect 4973 -43 4979 12
rect 5005 -43 5011 252
rect 5037 108 5043 112
rect 5053 -43 5059 132
rect 5069 68 5075 232
rect 5085 128 5091 132
rect 5069 28 5075 32
rect 5101 -37 5107 52
rect 5101 -43 5123 -37
rect 5165 -43 5171 32
rect 5181 -37 5187 52
rect 5325 48 5331 512
rect 5373 448 5379 492
rect 5405 328 5411 432
rect 5421 308 5427 492
rect 5469 468 5475 912
rect 5565 788 5571 812
rect 5517 648 5523 652
rect 5469 343 5475 452
rect 5469 337 5491 343
rect 5373 268 5379 272
rect 5373 148 5379 252
rect 5437 128 5443 312
rect 5469 108 5475 232
rect 5485 188 5491 337
rect 5517 288 5523 532
rect 5533 388 5539 612
rect 5549 548 5555 672
rect 5597 548 5603 672
rect 5613 608 5619 912
rect 5725 888 5731 912
rect 5661 748 5667 832
rect 5773 788 5779 1012
rect 5805 948 5811 1092
rect 5821 1088 5827 1112
rect 5869 948 5875 1092
rect 5885 1088 5891 1177
rect 5885 1068 5891 1072
rect 5917 1068 5923 1112
rect 5997 1028 6003 1312
rect 5981 948 5987 952
rect 5629 548 5635 712
rect 5661 688 5667 712
rect 5645 528 5651 672
rect 5565 508 5571 514
rect 5581 388 5587 432
rect 5501 188 5507 272
rect 5517 188 5523 272
rect 5533 148 5539 272
rect 5565 188 5571 312
rect 5597 268 5603 352
rect 5629 308 5635 512
rect 5677 508 5683 632
rect 5693 548 5699 672
rect 5709 588 5715 592
rect 5549 148 5555 172
rect 5581 148 5587 232
rect 5197 -17 5203 12
rect 5197 -23 5219 -17
rect 5213 -37 5219 -23
rect 5181 -43 5203 -37
rect 5213 -43 5251 -37
rect 5277 -43 5283 32
rect 5309 -37 5315 12
rect 5309 -43 5331 -37
rect 5357 -43 5363 12
rect 5405 -43 5411 32
rect 5533 -43 5539 132
rect 5597 103 5603 132
rect 5661 128 5667 372
rect 5693 328 5699 532
rect 5741 348 5747 632
rect 5789 568 5795 592
rect 5837 588 5843 892
rect 5965 788 5971 852
rect 6013 828 6019 1497
rect 6077 1288 6083 1532
rect 6173 1508 6179 1652
rect 6093 1328 6099 1492
rect 6125 1328 6131 1352
rect 6157 1308 6163 1352
rect 6029 1228 6035 1232
rect 6029 1088 6035 1172
rect 6045 968 6051 1092
rect 6077 928 6083 1152
rect 6093 1128 6099 1232
rect 6125 1128 6131 1212
rect 6125 1108 6131 1112
rect 6093 928 6099 1072
rect 6157 928 6163 1072
rect 6173 1048 6179 1492
rect 6189 1388 6195 1472
rect 6221 1468 6227 1492
rect 6269 1468 6275 1672
rect 6205 1348 6211 1352
rect 6221 1328 6227 1432
rect 6301 1343 6307 1712
rect 6365 1588 6371 1932
rect 6445 1908 6451 1912
rect 6429 1868 6435 1872
rect 6429 1788 6435 1832
rect 6445 1748 6451 1852
rect 6461 1748 6467 2092
rect 6493 1988 6499 2112
rect 6589 2108 6595 2152
rect 6605 2128 6611 2312
rect 6637 2288 6643 2312
rect 6605 1888 6611 2112
rect 6621 1888 6627 2272
rect 6637 2228 6643 2232
rect 6637 2188 6643 2212
rect 6701 2108 6707 2412
rect 6717 2308 6723 2372
rect 6733 2328 6739 2332
rect 6701 2088 6707 2092
rect 6717 2008 6723 2232
rect 6749 2128 6755 2412
rect 6829 2348 6835 2512
rect 6845 2348 6851 2352
rect 6781 2228 6787 2332
rect 6813 2283 6819 2312
rect 6861 2308 6867 2552
rect 6877 2528 6883 2532
rect 6925 2528 6931 2552
rect 7021 2548 7027 2632
rect 7037 2568 7043 3332
rect 7069 3308 7075 3312
rect 7165 3308 7171 3352
rect 7181 3348 7187 3872
rect 7197 3788 7203 3892
rect 7229 3748 7235 4032
rect 7229 3728 7235 3732
rect 7213 3388 7219 3490
rect 7229 3488 7235 3712
rect 7245 3328 7251 3332
rect 7053 3288 7059 3292
rect 7096 3277 7107 3283
rect 7101 3188 7107 3277
rect 7133 3168 7139 3272
rect 7181 3248 7187 3312
rect 7101 3088 7107 3092
rect 7117 3008 7123 3132
rect 7133 2948 7139 3152
rect 7165 3088 7171 3192
rect 7085 2788 7091 2892
rect 7101 2768 7107 2932
rect 7133 2788 7139 2912
rect 7197 2888 7203 2992
rect 7213 2928 7219 3072
rect 7245 2928 7251 2932
rect 7165 2808 7171 2832
rect 7101 2748 7107 2752
rect 7069 2628 7075 2732
rect 7101 2628 7107 2712
rect 6909 2488 6915 2512
rect 7037 2508 7043 2512
rect 7005 2497 7016 2503
rect 6925 2488 6931 2492
rect 6909 2468 6915 2472
rect 6893 2388 6899 2432
rect 6973 2428 6979 2432
rect 6877 2308 6883 2312
rect 6909 2308 6915 2392
rect 7005 2388 7011 2497
rect 7053 2388 7059 2472
rect 6925 2348 6931 2372
rect 6797 2277 6819 2283
rect 6797 2108 6803 2277
rect 6797 2048 6803 2092
rect 6829 2088 6835 2152
rect 6813 2068 6819 2072
rect 6637 1908 6643 1972
rect 6717 1888 6723 1892
rect 6509 1748 6515 1832
rect 6541 1743 6547 1832
rect 6557 1788 6563 1852
rect 6541 1737 6563 1743
rect 6397 1728 6403 1732
rect 6381 1708 6387 1712
rect 6429 1608 6435 1712
rect 6477 1628 6483 1732
rect 6525 1728 6531 1732
rect 6525 1588 6531 1692
rect 6317 1488 6323 1492
rect 6285 1337 6307 1343
rect 6285 1328 6291 1337
rect 6221 1208 6227 1312
rect 6301 1288 6307 1312
rect 6333 1308 6339 1432
rect 6349 1288 6355 1452
rect 6365 1328 6371 1332
rect 6413 1328 6419 1572
rect 6557 1508 6563 1737
rect 6573 1688 6579 1752
rect 6573 1528 6579 1672
rect 6589 1648 6595 1732
rect 6605 1728 6611 1832
rect 6445 1488 6451 1492
rect 6429 1328 6435 1332
rect 6189 1088 6195 1152
rect 6317 1148 6323 1232
rect 6269 1088 6275 1132
rect 6365 1128 6371 1232
rect 6381 1228 6387 1292
rect 6413 1288 6419 1312
rect 6445 1308 6451 1412
rect 6557 1408 6563 1492
rect 6557 1328 6563 1392
rect 6429 1168 6435 1232
rect 6493 1148 6499 1232
rect 6509 1228 6515 1292
rect 6573 1268 6579 1292
rect 6589 1288 6595 1632
rect 6605 1588 6611 1692
rect 6621 1608 6627 1872
rect 6637 1728 6643 1872
rect 6685 1768 6691 1832
rect 6621 1548 6627 1572
rect 6653 1508 6659 1512
rect 6685 1448 6691 1492
rect 6685 1348 6691 1432
rect 6685 1328 6691 1332
rect 6701 1328 6707 1552
rect 6717 1508 6723 1592
rect 6717 1488 6723 1492
rect 6637 1308 6643 1312
rect 6701 1308 6707 1312
rect 6669 1288 6675 1292
rect 6685 1268 6691 1272
rect 6557 1188 6563 1232
rect 6397 1128 6403 1132
rect 6525 1128 6531 1152
rect 6621 1148 6627 1232
rect 6589 1128 6595 1132
rect 6285 1108 6291 1112
rect 6269 1048 6275 1052
rect 6205 948 6211 1032
rect 6301 928 6307 1032
rect 6333 988 6339 1072
rect 6413 928 6419 1092
rect 6429 968 6435 1092
rect 6445 1088 6451 1092
rect 6429 923 6435 952
rect 6493 948 6499 1112
rect 6509 1108 6515 1112
rect 6621 1108 6627 1112
rect 6637 1108 6643 1232
rect 6509 1068 6515 1072
rect 6509 948 6515 1052
rect 6525 968 6531 1032
rect 6557 1028 6563 1092
rect 6573 1088 6579 1092
rect 6573 1068 6579 1072
rect 6573 948 6579 952
rect 6456 937 6467 943
rect 6429 917 6451 923
rect 5885 708 5891 732
rect 5981 688 5987 732
rect 5853 588 5859 592
rect 5965 548 5971 672
rect 6045 588 6051 712
rect 6077 703 6083 912
rect 6072 697 6083 703
rect 6093 688 6099 692
rect 5805 448 5811 532
rect 5981 530 5987 552
rect 5709 328 5715 332
rect 5805 288 5811 432
rect 5592 97 5603 103
rect 5741 48 5747 132
rect 5821 128 5827 332
rect 5981 328 5987 492
rect 6077 368 6083 532
rect 6093 528 6099 532
rect 6109 528 6115 832
rect 6365 788 6371 892
rect 6237 708 6243 712
rect 6125 508 6131 692
rect 6317 588 6323 712
rect 6349 688 6355 752
rect 6397 748 6403 832
rect 6381 708 6387 712
rect 6445 708 6451 917
rect 6461 908 6467 937
rect 6461 788 6467 892
rect 6573 708 6579 732
rect 6141 548 6147 572
rect 6173 548 6179 552
rect 6141 508 6147 512
rect 5981 308 5987 312
rect 5997 283 6003 292
rect 6013 288 6019 312
rect 6141 288 6147 492
rect 6237 468 6243 532
rect 6285 448 6291 532
rect 6301 517 6312 523
rect 6301 488 6307 517
rect 6317 488 6323 492
rect 6285 288 6291 312
rect 5992 277 6003 283
rect 5885 268 5891 272
rect 5773 108 5779 112
rect 5997 108 6003 112
rect 6013 -43 6019 272
rect 6157 268 6163 272
rect 6093 188 6099 252
rect 6125 128 6131 172
rect 6141 108 6147 132
rect 6173 128 6179 272
rect 6189 148 6195 152
rect 6269 28 6275 132
rect 6269 -43 6275 12
rect 6333 -37 6339 672
rect 6381 548 6387 552
rect 6397 488 6403 532
rect 6429 488 6435 692
rect 6445 688 6451 692
rect 6445 528 6451 532
rect 6397 328 6403 472
rect 6381 288 6387 312
rect 6397 308 6403 312
rect 6429 288 6435 352
rect 6461 288 6467 332
rect 6525 306 6531 312
rect 6381 128 6387 252
rect 6413 108 6419 112
rect 6333 -43 6355 -37
rect 6429 -43 6435 272
rect 6493 268 6499 272
rect 6509 148 6515 172
rect 6573 148 6579 212
rect 6589 143 6595 512
rect 6605 508 6611 512
rect 6621 508 6627 1092
rect 6637 1088 6643 1092
rect 6669 1048 6675 1072
rect 6685 1068 6691 1112
rect 6717 1103 6723 1452
rect 6733 1308 6739 1992
rect 6749 1928 6755 2032
rect 6829 2008 6835 2072
rect 6845 1968 6851 2132
rect 6877 2088 6883 2092
rect 6909 2068 6915 2092
rect 6893 2008 6899 2032
rect 6781 1908 6787 1912
rect 6845 1888 6851 1952
rect 6877 1906 6883 1912
rect 6877 1788 6883 1832
rect 6909 1788 6915 2052
rect 6909 1768 6915 1772
rect 6813 1648 6819 1732
rect 6845 1728 6851 1732
rect 6861 1548 6867 1632
rect 6877 1588 6883 1632
rect 6781 1508 6787 1512
rect 6909 1508 6915 1512
rect 6925 1468 6931 2232
rect 6941 2088 6947 2352
rect 7069 2348 7075 2432
rect 7085 2343 7091 2572
rect 7101 2508 7107 2532
rect 7117 2528 7123 2692
rect 7181 2668 7187 2672
rect 7149 2528 7155 2552
rect 7165 2528 7171 2572
rect 7133 2468 7139 2472
rect 7085 2337 7107 2343
rect 6957 2308 6963 2312
rect 6989 2108 6995 2332
rect 7053 2308 7059 2312
rect 7069 2228 7075 2332
rect 7101 2308 7107 2337
rect 6957 2068 6963 2072
rect 6973 2068 6979 2092
rect 7005 2088 7011 2212
rect 7101 2188 7107 2272
rect 7117 2128 7123 2292
rect 7069 2108 7075 2112
rect 7037 2068 7043 2092
rect 7053 2088 7059 2092
rect 7133 2088 7139 2452
rect 7165 2408 7171 2432
rect 7149 2308 7155 2352
rect 7197 2348 7203 2872
rect 7229 2788 7235 2892
rect 7245 2708 7251 2912
rect 7261 2748 7267 3812
rect 7277 3728 7283 3792
rect 7293 3628 7299 4112
rect 7309 3828 7315 4512
rect 7341 4508 7347 5352
rect 7357 5068 7363 5312
rect 7389 5123 7395 5232
rect 7373 5117 7395 5123
rect 7357 5008 7363 5032
rect 7373 4468 7379 5117
rect 7389 5088 7395 5092
rect 7405 4663 7411 5052
rect 7421 4988 7427 5052
rect 7421 4948 7427 4972
rect 7405 4657 7427 4663
rect 7325 4188 7331 4292
rect 7341 4148 7347 4452
rect 7389 4348 7395 4432
rect 7405 4188 7411 4472
rect 7341 3928 7347 4132
rect 7357 4048 7363 4112
rect 7373 4068 7379 4112
rect 7325 3748 7331 3872
rect 7341 3828 7347 3890
rect 7389 3788 7395 3812
rect 7357 3728 7363 3772
rect 7405 3748 7411 3752
rect 7384 3737 7395 3743
rect 7373 3728 7379 3732
rect 7357 3508 7363 3692
rect 7341 3408 7347 3432
rect 7277 3368 7283 3392
rect 7277 3328 7283 3332
rect 7293 2928 7299 3312
rect 7357 3228 7363 3492
rect 7373 3088 7379 3712
rect 7389 3588 7395 3737
rect 7389 3388 7395 3452
rect 7341 3068 7347 3072
rect 7293 2788 7299 2912
rect 7309 2908 7315 2952
rect 7213 2648 7219 2692
rect 7293 2688 7299 2692
rect 7245 2528 7251 2572
rect 7261 2508 7267 2652
rect 7325 2628 7331 3032
rect 7309 2528 7315 2572
rect 7229 2448 7235 2472
rect 7261 2388 7267 2472
rect 7277 2363 7283 2512
rect 7325 2508 7331 2612
rect 7293 2388 7299 2472
rect 7277 2357 7299 2363
rect 7213 2268 7219 2292
rect 7229 2288 7235 2292
rect 7277 2268 7283 2312
rect 7245 2128 7251 2132
rect 7037 1948 7043 1952
rect 7069 1928 7075 2052
rect 7085 1928 7091 1992
rect 7101 1908 7107 1992
rect 7133 1968 7139 2072
rect 7149 1928 7155 2092
rect 7181 2008 7187 2032
rect 7165 1988 7171 1992
rect 6941 1748 6947 1872
rect 7005 1848 7011 1852
rect 7181 1848 7187 1932
rect 6941 1728 6947 1732
rect 7021 1728 7027 1752
rect 7005 1708 7011 1712
rect 7021 1548 7027 1712
rect 6749 1448 6755 1452
rect 6749 1428 6755 1432
rect 6749 1348 6755 1352
rect 6749 1328 6755 1332
rect 6781 1308 6787 1432
rect 6797 1328 6803 1392
rect 6733 1288 6739 1292
rect 6765 1268 6771 1292
rect 6712 1097 6723 1103
rect 6685 1008 6691 1032
rect 6749 1028 6755 1232
rect 6765 1003 6771 1252
rect 6797 1143 6803 1232
rect 6781 1137 6803 1143
rect 6781 1128 6787 1137
rect 6845 1128 6851 1132
rect 6877 1128 6883 1312
rect 6893 1248 6899 1332
rect 6909 1128 6915 1172
rect 6925 1168 6931 1352
rect 6941 1188 6947 1332
rect 6877 1108 6883 1112
rect 6941 1108 6947 1132
rect 6813 1008 6819 1092
rect 6893 1088 6899 1092
rect 6957 1088 6963 1092
rect 6861 1063 6867 1072
rect 6973 1063 6979 1072
rect 6861 1057 6979 1063
rect 6749 997 6771 1003
rect 6749 988 6755 997
rect 6845 988 6851 1032
rect 6941 968 6947 972
rect 6637 928 6643 952
rect 6893 928 6899 932
rect 6973 928 6979 972
rect 6989 968 6995 1472
rect 7037 1468 7043 1632
rect 7053 1588 7059 1752
rect 7053 1568 7059 1572
rect 7101 1568 7107 1832
rect 7133 1648 7139 1712
rect 7101 1508 7107 1512
rect 7085 1488 7091 1492
rect 7117 1488 7123 1532
rect 7069 1328 7075 1392
rect 7085 1308 7091 1372
rect 7005 1048 7011 1192
rect 7069 1123 7075 1232
rect 7069 1117 7080 1123
rect 7021 1108 7027 1112
rect 7037 1063 7043 1092
rect 7032 1057 7043 1063
rect 7005 928 7011 932
rect 6749 888 6755 912
rect 6701 688 6707 732
rect 6653 548 6659 672
rect 6685 528 6691 532
rect 6669 308 6675 312
rect 6685 188 6691 492
rect 6717 328 6723 432
rect 6733 388 6739 812
rect 6765 706 6771 712
rect 6781 588 6787 672
rect 6749 528 6755 532
rect 6797 528 6803 912
rect 7037 908 7043 1012
rect 7037 706 7043 712
rect 6909 588 6915 652
rect 7021 588 7027 672
rect 7037 648 7043 652
rect 7069 548 7075 992
rect 7085 868 7091 972
rect 7101 968 7107 1012
rect 7117 988 7123 1472
rect 7133 1328 7139 1352
rect 7149 1308 7155 1372
rect 7165 1283 7171 1832
rect 7213 1828 7219 1892
rect 7229 1888 7235 1892
rect 7277 1868 7283 1912
rect 7245 1788 7251 1832
rect 7261 1728 7267 1812
rect 7293 1788 7299 2357
rect 7309 2208 7315 2292
rect 7325 2268 7331 2492
rect 7341 2388 7347 2892
rect 7357 2706 7363 2832
rect 7373 2788 7379 3072
rect 7389 2948 7395 3332
rect 7389 2928 7395 2932
rect 7405 2928 7411 3092
rect 7405 2888 7411 2912
rect 7357 2363 7363 2512
rect 7373 2468 7379 2472
rect 7389 2428 7395 2432
rect 7389 2388 7395 2392
rect 7421 2368 7427 4657
rect 7341 2357 7363 2363
rect 7309 2130 7315 2172
rect 7341 1988 7347 2357
rect 7357 2308 7363 2312
rect 7421 2308 7427 2352
rect 7389 2148 7395 2192
rect 7405 2157 7416 2163
rect 7373 1988 7379 2112
rect 7357 1948 7363 1952
rect 7325 1928 7331 1932
rect 7341 1908 7347 1912
rect 7309 1748 7315 1752
rect 7357 1743 7363 1932
rect 7389 1908 7395 2132
rect 7405 1988 7411 2157
rect 7421 1868 7427 1992
rect 7341 1737 7363 1743
rect 7277 1728 7283 1732
rect 7261 1708 7267 1712
rect 7181 1408 7187 1672
rect 7213 1508 7219 1632
rect 7277 1608 7283 1712
rect 7341 1688 7347 1737
rect 7357 1688 7363 1712
rect 7373 1708 7379 1752
rect 7357 1528 7363 1632
rect 7229 1508 7235 1512
rect 7357 1488 7363 1492
rect 7373 1488 7379 1692
rect 7389 1508 7395 1712
rect 7197 1328 7203 1352
rect 7213 1308 7219 1472
rect 7229 1388 7235 1392
rect 7309 1328 7315 1472
rect 7160 1277 7176 1283
rect 7133 1128 7139 1232
rect 7197 1188 7203 1232
rect 7341 1188 7347 1452
rect 7373 1403 7379 1432
rect 7357 1397 7379 1403
rect 7357 1330 7363 1397
rect 7405 1188 7411 1272
rect 7229 1128 7235 1172
rect 7101 668 7107 732
rect 7165 588 7171 892
rect 7197 883 7203 1092
rect 7213 1068 7219 1072
rect 7277 1068 7283 1072
rect 7229 1028 7235 1032
rect 7293 1008 7299 1032
rect 7309 988 7315 1072
rect 7421 1068 7427 1732
rect 7309 928 7315 952
rect 7357 908 7363 912
rect 7197 877 7219 883
rect 7213 788 7219 877
rect 7181 688 7187 692
rect 6701 308 6707 312
rect 6717 308 6723 312
rect 6749 148 6755 512
rect 6813 488 6819 532
rect 6813 468 6819 472
rect 6829 428 6835 432
rect 6957 308 6963 532
rect 7032 517 7043 523
rect 7005 508 7011 512
rect 7037 508 7043 517
rect 6989 497 7000 503
rect 6973 388 6979 492
rect 6989 328 6995 497
rect 7149 488 7155 532
rect 7069 388 7075 452
rect 6813 148 6819 152
rect 6877 148 6883 272
rect 6589 137 6611 143
rect 6509 128 6515 132
rect 6573 48 6579 132
rect 6605 128 6611 137
rect 6925 143 6931 292
rect 6941 188 6947 232
rect 6957 228 6963 272
rect 7005 248 7011 312
rect 6973 148 6979 152
rect 6920 137 6931 143
rect 6605 108 6611 112
rect 6829 108 6835 112
rect 6573 -43 6579 32
rect 6909 28 6915 132
rect 7021 128 7027 212
rect 7037 128 7043 292
rect 7133 188 7139 192
rect 7165 188 7171 552
rect 7181 508 7187 652
rect 7197 628 7203 692
rect 7293 688 7299 690
rect 7213 548 7219 632
rect 7229 588 7235 672
rect 7261 648 7267 672
rect 7261 528 7267 632
rect 7389 528 7395 792
rect 7405 783 7411 972
rect 7405 777 7416 783
rect 7437 568 7443 4692
rect 7437 528 7443 532
rect 7181 308 7187 492
rect 7213 308 7219 312
rect 7261 288 7267 512
rect 7309 508 7315 512
rect 7293 328 7299 472
rect 7325 328 7331 512
rect 7293 288 7299 312
rect 7325 308 7331 312
rect 7341 228 7347 232
rect 7149 168 7155 172
rect 7229 148 7235 152
rect 7197 128 7203 132
rect 6941 108 6947 112
<< m3contact >>
rect 2157 5402 2193 5418
rect 3048 5412 3064 5428
rect 3080 5412 3096 5428
rect 3112 5412 3128 5428
rect 3064 5392 3080 5408
rect 3160 5412 3176 5428
rect 3128 5392 3144 5408
rect 104 5372 120 5388
rect 296 5372 312 5388
rect 376 5372 392 5388
rect 664 5372 680 5388
rect 856 5372 872 5388
rect 1944 5372 1960 5388
rect 2056 5372 2072 5388
rect 2424 5372 2440 5388
rect 3192 5372 3208 5388
rect 3384 5372 3400 5388
rect 56 5332 72 5348
rect 1272 5352 1288 5368
rect 1400 5352 1416 5368
rect 1512 5352 1528 5368
rect 824 5332 840 5348
rect 1032 5332 1048 5348
rect 1048 5332 1064 5348
rect 40 5312 56 5328
rect 184 5312 200 5328
rect 232 5312 248 5328
rect 520 5312 536 5328
rect 600 5312 616 5328
rect 792 5314 808 5328
rect 792 5312 808 5314
rect 872 5312 904 5328
rect 936 5312 952 5328
rect 8 5292 24 5308
rect 88 5292 104 5308
rect 72 4972 88 4988
rect 8 4952 24 4968
rect 72 4952 88 4968
rect 280 5132 296 5148
rect 232 4972 248 4988
rect 200 4932 216 4948
rect 72 4912 88 4928
rect 104 4912 120 4928
rect 184 4912 200 4928
rect 24 4892 40 4908
rect 8 4652 24 4668
rect 8 4592 24 4608
rect 56 4792 72 4808
rect 136 4892 152 4908
rect 184 4892 200 4908
rect 376 5112 392 5128
rect 648 5292 664 5308
rect 488 5152 504 5168
rect 408 5132 424 5148
rect 520 5132 536 5148
rect 568 5132 584 5148
rect 488 5112 504 5128
rect 392 5092 408 5108
rect 392 5072 408 5088
rect 680 5152 696 5168
rect 616 5112 632 5128
rect 648 5112 664 5128
rect 616 5092 632 5108
rect 504 5072 520 5088
rect 584 5072 600 5088
rect 600 5072 616 5088
rect 408 5032 424 5048
rect 456 5032 472 5048
rect 360 5012 376 5028
rect 280 4952 296 4968
rect 456 4952 472 4968
rect 632 5072 648 5088
rect 616 5052 632 5068
rect 632 5032 648 5048
rect 296 4932 312 4948
rect 536 4932 552 4948
rect 136 4712 152 4728
rect 264 4712 268 4728
rect 268 4712 280 4728
rect 232 4692 248 4708
rect 280 4692 296 4708
rect 440 4892 456 4908
rect 504 4892 520 4908
rect 376 4672 392 4688
rect 88 4632 104 4648
rect 104 4572 120 4588
rect 200 4652 216 4668
rect 312 4632 328 4648
rect 296 4572 312 4588
rect 328 4572 344 4588
rect 504 4692 520 4708
rect 424 4652 440 4668
rect 488 4632 504 4648
rect 568 4772 584 4788
rect 728 5132 744 5148
rect 776 5132 792 5148
rect 840 5112 856 5128
rect 776 5092 792 5108
rect 728 5072 744 5088
rect 712 5032 728 5048
rect 680 4932 696 4948
rect 664 4752 680 4768
rect 632 4712 648 4728
rect 568 4692 584 4708
rect 648 4692 664 4708
rect 520 4592 536 4608
rect 472 4532 488 4548
rect 72 4512 88 4528
rect 168 4514 184 4528
rect 168 4512 184 4514
rect 232 4512 248 4528
rect 424 4512 440 4528
rect 24 4492 40 4508
rect 72 4492 88 4508
rect 8 4312 24 4328
rect 8 4252 24 4268
rect 72 4312 88 4328
rect 216 4312 232 4328
rect 72 4292 88 4308
rect 168 4306 184 4308
rect 168 4292 184 4306
rect 104 4232 120 4248
rect 184 4172 200 4188
rect 88 4132 104 4148
rect 24 3972 40 3988
rect 376 4452 392 4468
rect 360 4352 376 4368
rect 568 4672 584 4688
rect 584 4572 600 4588
rect 696 4652 712 4668
rect 664 4632 680 4648
rect 696 4572 712 4588
rect 776 5032 792 5048
rect 808 5032 824 5048
rect 760 4972 776 4988
rect 840 4972 856 4988
rect 808 4932 824 4948
rect 792 4912 808 4928
rect 776 4832 792 4848
rect 744 4692 760 4708
rect 776 4632 792 4648
rect 632 4532 648 4548
rect 664 4532 680 4548
rect 728 4532 744 4548
rect 792 4592 808 4608
rect 600 4512 616 4528
rect 616 4512 632 4528
rect 664 4512 680 4528
rect 696 4512 712 4528
rect 728 4512 744 4528
rect 712 4492 728 4508
rect 552 4472 568 4488
rect 776 4472 792 4488
rect 760 4432 776 4448
rect 584 4332 600 4348
rect 696 4332 712 4348
rect 520 4312 536 4328
rect 312 4292 328 4308
rect 360 4292 376 4308
rect 296 4232 312 4248
rect 296 4172 312 4188
rect 232 4132 248 4148
rect 216 4112 232 4128
rect 264 4112 280 4128
rect 200 4052 216 4068
rect 472 4292 488 4308
rect 632 4292 648 4308
rect 728 4312 744 4328
rect 760 4312 776 4328
rect 712 4292 728 4308
rect 616 4272 632 4288
rect 664 4272 680 4288
rect 600 4252 616 4268
rect 392 4212 408 4228
rect 360 4172 376 4188
rect 440 4172 456 4188
rect 488 4112 504 4128
rect 568 4112 584 4128
rect 328 3992 344 4008
rect 392 4072 408 4088
rect 408 3992 424 4008
rect 200 3892 216 3908
rect 280 3892 296 3908
rect 376 3892 392 3908
rect 88 3872 104 3888
rect 200 3872 216 3888
rect 184 3832 200 3848
rect 168 3752 184 3768
rect 24 3692 40 3708
rect 8 3632 24 3648
rect 56 3632 72 3648
rect 24 3492 40 3508
rect 88 3492 104 3508
rect 8 3472 24 3488
rect 72 3472 88 3488
rect 24 3312 40 3328
rect 56 3314 72 3328
rect 56 3312 72 3314
rect 56 3112 72 3128
rect 40 3092 56 3108
rect 136 3714 152 3728
rect 136 3712 152 3714
rect 200 3712 216 3728
rect 200 3692 216 3708
rect 168 3672 184 3688
rect 120 3532 136 3548
rect 184 3612 200 3628
rect 136 3512 152 3528
rect 200 3512 216 3528
rect 152 3492 168 3508
rect 136 3472 152 3488
rect 200 3412 216 3428
rect 200 3392 216 3408
rect 344 3872 360 3888
rect 296 3832 312 3848
rect 232 3792 264 3808
rect 296 3772 312 3788
rect 248 3732 264 3748
rect 392 3872 408 3888
rect 392 3852 408 3868
rect 456 3992 472 4008
rect 536 3972 552 3988
rect 584 3972 600 3988
rect 952 5252 968 5268
rect 1320 5332 1336 5348
rect 1384 5332 1400 5348
rect 1496 5332 1512 5348
rect 1672 5332 1688 5348
rect 1736 5332 1752 5348
rect 1832 5332 1848 5348
rect 1992 5332 2008 5348
rect 2360 5332 2376 5348
rect 1144 5312 1160 5328
rect 1208 5312 1224 5328
rect 1288 5312 1304 5328
rect 1432 5312 1448 5328
rect 1480 5312 1496 5328
rect 1064 5292 1080 5308
rect 1117 5202 1153 5218
rect 1064 5132 1080 5148
rect 1176 5112 1192 5128
rect 904 5092 920 5108
rect 904 5072 920 5088
rect 1032 5072 1048 5088
rect 1128 5072 1144 5088
rect 968 5032 984 5048
rect 1000 5032 1016 5048
rect 1144 4932 1160 4948
rect 1320 5292 1336 5308
rect 1368 5292 1384 5308
rect 1448 5292 1464 5308
rect 1480 5292 1496 5308
rect 1432 5272 1448 5288
rect 1448 5212 1464 5228
rect 1400 5192 1416 5208
rect 1240 5172 1256 5188
rect 1368 5112 1372 5128
rect 1372 5112 1384 5128
rect 1336 5092 1352 5108
rect 1384 5092 1400 5108
rect 1256 4972 1272 4988
rect 952 4912 968 4928
rect 1192 4912 1208 4928
rect 1272 4912 1288 4928
rect 888 4892 904 4908
rect 936 4892 952 4908
rect 888 4872 904 4888
rect 872 4832 888 4848
rect 856 4732 872 4748
rect 888 4712 904 4728
rect 936 4712 952 4728
rect 904 4692 920 4708
rect 936 4692 952 4708
rect 968 4732 984 4748
rect 984 4692 1000 4708
rect 952 4652 968 4668
rect 984 4652 1000 4668
rect 1016 4792 1032 4808
rect 1096 4792 1112 4808
rect 1117 4802 1153 4818
rect 1272 4812 1288 4828
rect 1032 4732 1048 4748
rect 1032 4672 1048 4688
rect 1000 4632 1016 4648
rect 1080 4692 1096 4708
rect 1208 4692 1224 4708
rect 1224 4672 1240 4688
rect 984 4612 1000 4628
rect 1048 4612 1064 4628
rect 1304 4692 1320 4708
rect 1304 4672 1320 4688
rect 1224 4652 1240 4668
rect 1320 4652 1336 4668
rect 1240 4592 1256 4608
rect 1192 4572 1208 4588
rect 1016 4552 1032 4568
rect 1144 4552 1176 4568
rect 856 4532 872 4548
rect 840 4512 856 4528
rect 872 4512 888 4528
rect 888 4492 904 4508
rect 936 4492 952 4508
rect 936 4472 952 4488
rect 904 4452 920 4468
rect 856 4352 872 4368
rect 808 4332 840 4348
rect 1000 4512 1016 4528
rect 968 4492 984 4508
rect 952 4452 968 4468
rect 888 4312 904 4328
rect 952 4312 968 4328
rect 856 4292 872 4308
rect 808 4272 824 4288
rect 840 4272 856 4288
rect 840 4232 856 4248
rect 888 4232 904 4248
rect 888 4172 904 4188
rect 760 4112 776 4128
rect 440 3892 456 3908
rect 488 3892 504 3908
rect 504 3892 520 3908
rect 584 3892 600 3908
rect 456 3752 472 3768
rect 312 3732 328 3748
rect 360 3732 376 3748
rect 408 3732 424 3748
rect 280 3712 296 3728
rect 264 3672 280 3688
rect 328 3632 344 3648
rect 264 3532 280 3548
rect 296 3512 312 3528
rect 248 3452 264 3468
rect 376 3672 392 3688
rect 424 3612 440 3628
rect 424 3492 440 3508
rect 456 3492 472 3508
rect 296 3472 312 3488
rect 360 3472 376 3488
rect 520 3872 536 3888
rect 632 3872 648 3888
rect 504 3772 520 3788
rect 456 3452 472 3468
rect 488 3452 504 3468
rect 296 3412 312 3428
rect 376 3412 392 3428
rect 440 3412 456 3428
rect 264 3392 280 3408
rect 232 3332 248 3348
rect 392 3332 408 3348
rect 152 3312 168 3328
rect 216 3312 232 3328
rect 264 3312 280 3328
rect 120 3232 136 3248
rect 216 3292 232 3308
rect 184 3232 200 3248
rect 104 3112 120 3128
rect 184 3092 200 3108
rect 232 3092 248 3108
rect 8 3072 24 3088
rect 24 3012 40 3028
rect 88 3012 104 3028
rect 616 3832 632 3848
rect 728 3972 744 3988
rect 744 3906 760 3908
rect 744 3892 760 3906
rect 680 3852 696 3868
rect 536 3712 552 3728
rect 712 3712 728 3728
rect 680 3692 696 3708
rect 552 3652 568 3668
rect 584 3512 600 3528
rect 600 3492 616 3508
rect 552 3472 568 3488
rect 552 3412 568 3428
rect 920 4072 936 4088
rect 856 4032 872 4048
rect 808 3932 824 3948
rect 920 3912 936 3928
rect 920 3892 936 3908
rect 888 3852 904 3868
rect 872 3832 888 3848
rect 904 3772 920 3788
rect 792 3732 808 3748
rect 904 3732 920 3748
rect 808 3712 824 3728
rect 776 3552 792 3568
rect 808 3552 824 3568
rect 792 3492 808 3508
rect 760 3452 776 3468
rect 776 3412 792 3428
rect 728 3352 744 3368
rect 520 3332 536 3348
rect 408 3312 424 3328
rect 456 3312 472 3328
rect 584 3312 600 3328
rect 696 3312 712 3328
rect 552 3172 568 3188
rect 456 3152 472 3168
rect 472 3132 488 3148
rect 552 3132 568 3148
rect 360 3112 376 3128
rect 504 3112 520 3128
rect 632 3232 648 3248
rect 696 3232 712 3248
rect 904 3712 920 3728
rect 984 4472 1000 4488
rect 984 4312 1000 4328
rect 984 4292 1000 4308
rect 984 4112 1000 4128
rect 1256 4572 1272 4588
rect 1128 4532 1144 4548
rect 1224 4532 1240 4548
rect 1320 4532 1336 4548
rect 1032 4512 1048 4528
rect 1048 4512 1064 4528
rect 1192 4512 1208 4528
rect 1272 4512 1288 4528
rect 1032 4492 1048 4508
rect 1128 4492 1144 4508
rect 1080 4472 1096 4488
rect 1032 4452 1048 4468
rect 1117 4402 1153 4418
rect 1288 4372 1304 4388
rect 1048 4352 1064 4368
rect 1256 4352 1272 4368
rect 1096 4312 1112 4328
rect 1176 4312 1192 4328
rect 1016 4292 1032 4308
rect 1032 4292 1048 4308
rect 1016 4232 1032 4248
rect 1016 4192 1032 4208
rect 1064 4272 1080 4288
rect 1048 4152 1064 4168
rect 1032 4132 1048 4148
rect 1000 4012 1016 4028
rect 1016 3952 1032 3968
rect 1016 3932 1032 3948
rect 968 3912 984 3928
rect 1160 4272 1176 4288
rect 1144 4172 1160 4188
rect 1208 4272 1224 4288
rect 1240 4272 1256 4288
rect 1224 4232 1240 4248
rect 1960 5312 1976 5328
rect 1624 5292 1640 5308
rect 1704 5292 1720 5308
rect 1832 5292 1848 5308
rect 1912 5292 1928 5308
rect 1464 5192 1480 5208
rect 1496 5192 1512 5208
rect 1416 5052 1432 5068
rect 1352 4972 1368 4988
rect 1704 5132 1720 5148
rect 1608 5112 1624 5128
rect 1720 5112 1736 5128
rect 1800 5112 1816 5128
rect 1704 5092 1720 5108
rect 1752 5092 1768 5108
rect 1544 5072 1560 5088
rect 1704 5072 1720 5088
rect 1640 5052 1656 5068
rect 1480 5032 1496 5048
rect 1544 5032 1560 5048
rect 1400 4932 1416 4948
rect 1672 5032 1688 5048
rect 1672 4972 1688 4988
rect 1560 4912 1576 4928
rect 1576 4912 1592 4928
rect 1656 4912 1672 4928
rect 1400 4852 1416 4868
rect 1480 4852 1496 4868
rect 1416 4812 1432 4828
rect 1464 4732 1480 4748
rect 1608 4892 1624 4908
rect 1592 4832 1608 4848
rect 1496 4752 1512 4768
rect 1368 4692 1384 4708
rect 1480 4692 1496 4708
rect 1352 4672 1368 4688
rect 1416 4686 1432 4688
rect 1416 4672 1432 4686
rect 1448 4672 1464 4688
rect 1368 4652 1384 4668
rect 1384 4632 1400 4648
rect 1352 4612 1368 4628
rect 1368 4572 1384 4588
rect 1400 4592 1416 4608
rect 1384 4532 1400 4548
rect 1416 4512 1432 4528
rect 1352 4412 1368 4428
rect 1352 4392 1368 4408
rect 1336 4312 1352 4328
rect 1368 4372 1384 4388
rect 1288 4272 1304 4288
rect 1304 4272 1320 4288
rect 1464 4652 1480 4668
rect 1496 4572 1512 4588
rect 1528 4692 1544 4708
rect 1576 4692 1592 4708
rect 1560 4672 1576 4688
rect 1560 4592 1576 4608
rect 1480 4532 1496 4548
rect 1480 4492 1496 4508
rect 1608 4752 1624 4768
rect 1592 4492 1608 4508
rect 1528 4392 1544 4408
rect 1448 4312 1464 4328
rect 1432 4272 1448 4288
rect 1256 4192 1272 4208
rect 1192 4152 1208 4168
rect 1368 4132 1384 4148
rect 1160 4112 1176 4128
rect 1288 4112 1304 4128
rect 1144 4092 1160 4108
rect 1064 4072 1080 4088
rect 1064 3932 1080 3948
rect 968 3892 984 3908
rect 1048 3892 1080 3908
rect 952 3852 968 3868
rect 920 3692 936 3708
rect 936 3692 952 3708
rect 888 3672 904 3688
rect 824 3512 856 3528
rect 936 3512 952 3528
rect 856 3492 872 3508
rect 856 3412 872 3428
rect 920 3452 936 3468
rect 904 3392 920 3408
rect 984 3872 1000 3888
rect 984 3832 1000 3848
rect 1000 3812 1016 3828
rect 1000 3792 1016 3808
rect 1117 4002 1153 4018
rect 1128 3932 1144 3948
rect 1320 3932 1336 3948
rect 1208 3912 1224 3928
rect 1192 3906 1208 3908
rect 1192 3892 1208 3906
rect 1064 3772 1080 3788
rect 1192 3752 1208 3768
rect 1144 3732 1160 3748
rect 1032 3712 1048 3728
rect 1048 3712 1064 3728
rect 968 3672 984 3688
rect 968 3632 984 3648
rect 936 3412 984 3428
rect 952 3392 968 3408
rect 936 3312 952 3328
rect 760 3292 776 3308
rect 696 3112 712 3128
rect 408 3092 424 3108
rect 456 3072 472 3088
rect 488 3072 504 3088
rect 200 3032 216 3048
rect 200 2972 216 2988
rect 296 2952 312 2968
rect 264 2932 280 2948
rect 504 3032 520 3048
rect 488 2952 504 2968
rect 504 2952 520 2968
rect 552 2932 568 2948
rect 152 2912 168 2928
rect 216 2912 232 2928
rect 232 2912 248 2928
rect 264 2912 280 2928
rect 360 2914 376 2928
rect 360 2912 376 2914
rect 456 2912 472 2928
rect 8 2712 24 2728
rect 8 2552 40 2568
rect 24 2512 40 2528
rect 56 2472 72 2488
rect 184 2892 200 2908
rect 120 2872 136 2888
rect 136 2732 152 2748
rect 392 2892 408 2908
rect 504 2892 520 2908
rect 264 2732 280 2748
rect 200 2712 216 2728
rect 424 2712 440 2728
rect 520 2712 536 2728
rect 232 2692 248 2708
rect 280 2692 296 2708
rect 296 2692 312 2708
rect 360 2692 376 2708
rect 504 2692 520 2708
rect 536 2692 552 2708
rect 88 2652 104 2668
rect 104 2592 120 2608
rect 136 2492 152 2508
rect 136 2472 152 2488
rect 152 2472 168 2488
rect 72 2432 88 2448
rect 136 2432 152 2448
rect 8 2252 24 2268
rect 8 2072 24 2088
rect 136 2306 152 2308
rect 136 2292 152 2306
rect 184 2592 200 2608
rect 216 2492 232 2508
rect 248 2632 264 2648
rect 280 2532 296 2548
rect 296 2492 312 2508
rect 264 2472 280 2488
rect 232 2312 248 2328
rect 248 2312 264 2328
rect 232 2292 248 2308
rect 200 2252 216 2268
rect 216 2232 232 2248
rect 200 2152 216 2168
rect 168 2132 184 2148
rect 136 2114 152 2128
rect 136 2112 152 2114
rect 232 2112 248 2128
rect 152 1932 168 1948
rect 488 2672 504 2688
rect 376 2632 408 2648
rect 376 2592 392 2608
rect 616 3092 632 3108
rect 584 3052 600 3068
rect 680 2972 696 2988
rect 568 2892 584 2908
rect 680 2892 696 2908
rect 616 2872 632 2888
rect 600 2792 616 2808
rect 568 2652 584 2668
rect 568 2632 584 2648
rect 552 2612 568 2628
rect 632 2692 648 2708
rect 360 2532 392 2548
rect 392 2532 408 2548
rect 424 2532 440 2548
rect 328 2512 344 2528
rect 344 2492 360 2508
rect 312 2432 328 2448
rect 280 2312 296 2328
rect 264 2292 280 2308
rect 296 2232 312 2248
rect 296 2172 312 2188
rect 344 2172 360 2188
rect 344 2112 360 2128
rect 392 2512 408 2528
rect 456 2514 472 2528
rect 456 2512 472 2514
rect 408 2312 424 2328
rect 456 2312 472 2328
rect 376 2252 392 2268
rect 424 2292 440 2308
rect 456 2272 472 2288
rect 584 2492 600 2508
rect 600 2492 616 2508
rect 744 3112 760 3128
rect 760 3112 776 3128
rect 776 3072 792 3088
rect 760 2992 776 3008
rect 824 3172 840 3188
rect 1016 3172 1032 3188
rect 1000 3152 1016 3168
rect 840 3112 856 3128
rect 904 3092 920 3108
rect 1000 3112 1016 3128
rect 1048 3112 1064 3128
rect 968 3092 984 3108
rect 952 3072 968 3088
rect 1048 3072 1064 3088
rect 1112 3712 1128 3728
rect 1096 3692 1112 3708
rect 1080 3672 1096 3688
rect 1117 3602 1153 3618
rect 1192 3552 1208 3568
rect 1096 3532 1112 3548
rect 1160 3532 1176 3548
rect 1128 3412 1144 3428
rect 1480 4312 1496 4328
rect 1528 4312 1544 4328
rect 1576 4312 1592 4328
rect 1544 4292 1560 4308
rect 1512 4232 1528 4248
rect 1464 4112 1480 4128
rect 1608 4292 1624 4308
rect 1608 4272 1624 4288
rect 1592 4092 1608 4108
rect 1464 3952 1480 3968
rect 1512 3952 1528 3968
rect 1448 3932 1464 3948
rect 1448 3912 1464 3928
rect 1400 3892 1416 3908
rect 1432 3892 1448 3908
rect 1384 3852 1400 3868
rect 1336 3712 1352 3728
rect 1288 3692 1304 3708
rect 1240 3652 1256 3668
rect 1336 3652 1352 3668
rect 1352 3532 1368 3548
rect 1288 3506 1304 3508
rect 1288 3492 1304 3506
rect 1320 3452 1336 3468
rect 1352 3452 1368 3468
rect 1224 3412 1240 3428
rect 1384 3552 1400 3568
rect 1384 3512 1400 3528
rect 1384 3492 1400 3508
rect 1544 3892 1560 3908
rect 1496 3872 1512 3888
rect 1528 3812 1544 3828
rect 1544 3792 1560 3808
rect 1496 3752 1512 3768
rect 1528 3752 1544 3768
rect 1480 3712 1496 3728
rect 1432 3572 1448 3588
rect 1416 3412 1432 3428
rect 1368 3372 1384 3388
rect 1192 3332 1208 3348
rect 1256 3332 1272 3348
rect 1624 4112 1640 4128
rect 1624 4092 1640 4108
rect 1688 4692 1704 4708
rect 1752 4892 1768 4908
rect 1784 5052 1800 5068
rect 1768 4832 1784 4848
rect 1720 4672 1736 4688
rect 1816 4832 1832 4848
rect 1816 4712 1832 4728
rect 1752 4612 1768 4628
rect 1800 4612 1816 4628
rect 1656 4572 1672 4588
rect 1720 4532 1736 4548
rect 1672 4472 1688 4488
rect 1848 5112 1864 5128
rect 1848 5092 1864 5108
rect 2616 5332 2632 5348
rect 3000 5332 3016 5348
rect 2296 5312 2312 5328
rect 2408 5312 2424 5328
rect 2472 5312 2488 5328
rect 2504 5312 2520 5328
rect 2120 5292 2136 5308
rect 1976 5272 1992 5288
rect 2024 5272 2040 5288
rect 2168 5272 2184 5288
rect 1960 5252 1976 5268
rect 1960 5092 1976 5108
rect 1976 5072 1992 5088
rect 1880 5032 1896 5048
rect 2088 5052 2104 5068
rect 2072 5032 2088 5048
rect 1976 4992 1992 5008
rect 1864 4972 1880 4988
rect 2008 4972 2024 4988
rect 2072 4972 2088 4988
rect 1880 4952 1896 4968
rect 1944 4932 1960 4948
rect 1992 4912 2008 4928
rect 2056 4912 2072 4928
rect 2072 4892 2088 4908
rect 2168 5092 2184 5108
rect 2280 5172 2296 5188
rect 2392 5272 2408 5288
rect 2312 5212 2328 5228
rect 2360 5212 2376 5228
rect 2568 5292 2584 5308
rect 2456 5132 2472 5148
rect 2296 5112 2312 5128
rect 2440 5112 2456 5128
rect 2248 5092 2264 5108
rect 2392 5072 2408 5088
rect 2376 5052 2392 5068
rect 2136 5032 2152 5048
rect 2328 5032 2344 5048
rect 2157 5002 2193 5018
rect 2216 5012 2232 5028
rect 2120 4912 2136 4928
rect 1880 4872 1896 4888
rect 1944 4872 1960 4888
rect 2104 4872 2120 4888
rect 1928 4712 1944 4728
rect 1960 4712 1976 4728
rect 2024 4712 2040 4728
rect 2120 4712 2136 4728
rect 1864 4692 1880 4708
rect 1896 4692 1912 4708
rect 1800 4492 1816 4508
rect 1832 4492 1848 4508
rect 1880 4672 1896 4688
rect 1928 4632 1944 4648
rect 1960 4692 1976 4708
rect 2008 4692 2024 4708
rect 2056 4692 2072 4708
rect 2104 4692 2120 4708
rect 1976 4652 1992 4668
rect 1912 4552 1928 4568
rect 1944 4552 1960 4568
rect 1960 4532 1976 4548
rect 2072 4592 2088 4608
rect 2312 4952 2328 4968
rect 2376 4992 2392 5008
rect 2376 4972 2392 4988
rect 2232 4932 2248 4948
rect 2344 4932 2360 4948
rect 2456 5092 2472 5108
rect 2456 5012 2472 5028
rect 2424 4972 2440 4988
rect 2456 4972 2472 4988
rect 2424 4932 2440 4948
rect 2392 4912 2408 4928
rect 2456 4912 2472 4928
rect 2584 5212 2600 5228
rect 2488 5172 2504 5188
rect 3112 5312 3128 5328
rect 2808 5292 2824 5308
rect 2872 5292 2888 5308
rect 2744 5232 2760 5248
rect 2712 5192 2728 5208
rect 2504 5092 2520 5108
rect 2584 5092 2600 5108
rect 2632 5092 2648 5108
rect 2504 5072 2520 5088
rect 2536 5032 2552 5048
rect 2648 5052 2664 5068
rect 2600 5012 2616 5028
rect 2680 5012 2712 5028
rect 2552 4972 2568 4988
rect 2600 4972 2616 4988
rect 2664 4952 2680 4968
rect 2360 4892 2376 4908
rect 2392 4892 2408 4908
rect 2472 4892 2488 4908
rect 2584 4892 2600 4908
rect 2296 4872 2312 4888
rect 2264 4712 2280 4728
rect 2248 4692 2264 4708
rect 2136 4612 2152 4628
rect 2157 4602 2193 4618
rect 2136 4572 2152 4588
rect 1976 4492 2008 4508
rect 2088 4492 2104 4508
rect 1800 4452 1816 4468
rect 1848 4452 1864 4468
rect 1704 4412 1720 4428
rect 1784 4412 1800 4428
rect 1656 4392 1672 4408
rect 1640 4072 1656 4088
rect 1640 3872 1656 3888
rect 1624 3752 1640 3768
rect 1640 3732 1656 3748
rect 1528 3712 1544 3728
rect 1560 3712 1576 3728
rect 1528 3612 1544 3628
rect 1832 4372 1848 4388
rect 1672 4312 1688 4328
rect 1704 4312 1720 4328
rect 1672 4292 1688 4308
rect 1688 4152 1704 4168
rect 1784 4152 1800 4168
rect 1688 4132 1704 4148
rect 1768 4132 1784 4148
rect 1816 4132 1832 4148
rect 1672 4092 1688 4108
rect 1704 3832 1720 3848
rect 1704 3752 1720 3768
rect 1608 3692 1624 3708
rect 1592 3672 1608 3688
rect 1608 3632 1624 3648
rect 1448 3512 1464 3528
rect 1544 3512 1576 3528
rect 1480 3492 1496 3508
rect 1560 3492 1576 3508
rect 1448 3472 1464 3488
rect 1464 3412 1480 3428
rect 1096 3312 1112 3328
rect 1400 3312 1416 3328
rect 1432 3312 1448 3328
rect 1096 3292 1112 3308
rect 1176 3292 1192 3308
rect 1320 3272 1336 3288
rect 1368 3272 1400 3288
rect 1096 3212 1112 3228
rect 1117 3202 1153 3218
rect 1112 3172 1128 3188
rect 1160 3092 1176 3108
rect 1528 3132 1544 3148
rect 1448 3112 1464 3128
rect 1560 3312 1576 3328
rect 1240 3072 1272 3088
rect 1336 3072 1352 3088
rect 1400 3072 1416 3088
rect 1064 3052 1080 3068
rect 984 3032 1000 3048
rect 1128 2972 1144 2988
rect 1032 2952 1048 2968
rect 1496 3052 1512 3068
rect 1352 2952 1368 2968
rect 1480 2952 1496 2968
rect 824 2932 840 2948
rect 1368 2932 1384 2948
rect 728 2912 744 2928
rect 776 2912 792 2928
rect 1064 2912 1080 2928
rect 1112 2912 1128 2928
rect 712 2892 728 2908
rect 792 2892 808 2908
rect 840 2892 856 2908
rect 1384 2912 1400 2928
rect 1432 2912 1448 2928
rect 1112 2892 1128 2908
rect 1224 2892 1240 2908
rect 744 2872 760 2888
rect 760 2872 776 2888
rect 952 2872 968 2888
rect 776 2852 792 2868
rect 712 2692 728 2708
rect 696 2652 712 2668
rect 632 2612 664 2628
rect 760 2692 776 2708
rect 760 2652 776 2668
rect 728 2592 744 2608
rect 712 2572 728 2588
rect 648 2552 664 2568
rect 680 2532 696 2548
rect 616 2392 632 2408
rect 1117 2802 1153 2818
rect 792 2772 808 2788
rect 1128 2772 1144 2788
rect 952 2732 968 2748
rect 1144 2732 1160 2748
rect 888 2712 904 2728
rect 1032 2712 1048 2728
rect 840 2692 856 2708
rect 872 2692 888 2708
rect 808 2672 824 2688
rect 824 2632 840 2648
rect 696 2512 712 2528
rect 744 2512 760 2528
rect 664 2352 680 2368
rect 968 2692 984 2708
rect 1016 2692 1032 2708
rect 1080 2692 1096 2708
rect 1112 2692 1128 2708
rect 888 2652 904 2668
rect 904 2612 920 2628
rect 1032 2652 1048 2668
rect 920 2592 936 2608
rect 888 2572 904 2588
rect 920 2552 936 2568
rect 824 2532 840 2548
rect 856 2532 872 2548
rect 904 2532 920 2548
rect 696 2332 712 2348
rect 760 2332 776 2348
rect 632 2292 648 2308
rect 744 2312 760 2328
rect 536 2252 552 2268
rect 712 2252 728 2268
rect 632 2232 648 2248
rect 584 2172 600 2188
rect 616 2172 632 2188
rect 456 2132 472 2148
rect 312 2092 328 2108
rect 360 2092 376 2108
rect 264 2072 280 2088
rect 392 2072 408 2088
rect 296 1932 312 1948
rect 424 1932 440 1948
rect 328 1912 340 1928
rect 340 1912 344 1928
rect 8 1892 24 1908
rect 88 1892 104 1908
rect 168 1892 184 1908
rect 232 1892 248 1908
rect 120 1872 136 1888
rect 8 1492 24 1508
rect 120 1712 136 1728
rect 216 1852 232 1868
rect 264 1852 280 1868
rect 504 2112 520 2128
rect 552 1892 568 1908
rect 376 1852 392 1868
rect 424 1852 440 1868
rect 472 1832 488 1848
rect 552 1812 568 1828
rect 536 1792 552 1808
rect 248 1732 264 1748
rect 216 1712 232 1728
rect 232 1632 248 1648
rect 296 1752 312 1768
rect 360 1752 376 1768
rect 472 1752 488 1768
rect 312 1732 328 1748
rect 280 1712 296 1728
rect 296 1692 328 1708
rect 328 1692 344 1708
rect 264 1632 280 1648
rect 248 1572 264 1588
rect 168 1532 184 1548
rect 136 1492 152 1508
rect 232 1512 248 1528
rect 200 1492 216 1508
rect 120 1472 136 1488
rect 232 1472 248 1488
rect 184 1372 200 1388
rect 296 1572 312 1588
rect 280 1512 296 1528
rect 264 1352 280 1368
rect 56 1332 72 1348
rect 200 1332 216 1348
rect 40 712 56 728
rect 40 692 56 708
rect 72 1312 88 1328
rect 216 1312 232 1328
rect 344 1532 360 1548
rect 488 1712 504 1728
rect 728 2172 744 2188
rect 664 2112 680 2128
rect 792 2352 808 2368
rect 776 2312 792 2328
rect 776 2292 792 2308
rect 760 2232 776 2248
rect 648 2092 664 2108
rect 696 2092 712 2108
rect 744 2092 760 2108
rect 600 1932 616 1948
rect 760 1932 776 1948
rect 600 1872 616 1888
rect 664 1872 680 1888
rect 696 1852 712 1868
rect 680 1792 696 1808
rect 632 1752 648 1768
rect 600 1732 616 1748
rect 760 1832 776 1848
rect 728 1812 744 1828
rect 728 1752 744 1768
rect 856 2492 872 2508
rect 1000 2612 1016 2628
rect 1016 2572 1032 2588
rect 1112 2672 1128 2688
rect 1592 3492 1608 3508
rect 1752 3732 1768 3748
rect 1672 3672 1688 3688
rect 1736 3672 1752 3688
rect 1752 3652 1768 3668
rect 1656 3532 1672 3548
rect 1640 3492 1656 3508
rect 1672 3512 1688 3528
rect 1656 3472 1672 3488
rect 1672 3472 1688 3488
rect 1640 3392 1656 3408
rect 1912 4312 1928 4328
rect 2184 4492 2200 4508
rect 2088 4452 2104 4468
rect 2168 4452 2184 4468
rect 2232 4572 2248 4588
rect 2312 4692 2328 4708
rect 2232 4532 2248 4548
rect 2296 4532 2312 4548
rect 2120 4432 2136 4448
rect 2200 4432 2216 4448
rect 2216 4332 2232 4348
rect 2264 4332 2280 4348
rect 2216 4312 2232 4328
rect 1944 4292 1960 4308
rect 1848 4252 1864 4268
rect 1912 4252 1928 4268
rect 1880 4212 1896 4228
rect 1896 4172 1912 4188
rect 1912 4152 1944 4168
rect 1960 4152 1976 4168
rect 1896 4112 1912 4128
rect 1912 4092 1928 4108
rect 1864 3932 1880 3948
rect 1800 3892 1816 3908
rect 1912 3892 1928 3908
rect 1816 3812 1832 3828
rect 2184 4292 2200 4308
rect 2184 4272 2200 4288
rect 2088 4252 2104 4268
rect 2008 4212 2024 4228
rect 2056 4192 2072 4208
rect 2008 4172 2024 4188
rect 1960 4132 1976 4148
rect 2056 4132 2072 4148
rect 1976 4112 1992 4128
rect 2088 4112 2104 4128
rect 2040 4012 2056 4028
rect 1944 3972 1960 3988
rect 2157 4202 2193 4218
rect 2216 4192 2232 4208
rect 2152 4152 2168 4168
rect 2200 4132 2216 4148
rect 2136 4112 2152 4128
rect 2136 4072 2152 4088
rect 2120 4032 2136 4048
rect 2152 4032 2168 4048
rect 2088 3932 2104 3948
rect 1960 3892 1976 3908
rect 1960 3872 1976 3888
rect 2024 3872 2040 3888
rect 1848 3792 1864 3808
rect 1816 3592 1832 3608
rect 2024 3832 2040 3848
rect 2088 3832 2104 3848
rect 1896 3812 1912 3828
rect 2088 3812 2104 3828
rect 2216 3932 2232 3948
rect 2248 4232 2264 4248
rect 2264 4172 2280 4188
rect 2344 4672 2376 4688
rect 2376 4652 2392 4668
rect 2408 4712 2424 4728
rect 2488 4712 2504 4728
rect 2440 4692 2456 4708
rect 2440 4572 2456 4588
rect 2344 4532 2360 4548
rect 2440 4532 2456 4548
rect 2328 4492 2332 4508
rect 2332 4492 2344 4508
rect 2312 4392 2328 4408
rect 2392 4452 2408 4468
rect 2424 4372 2440 4388
rect 2520 4692 2536 4708
rect 2728 5072 2744 5088
rect 2760 5072 2776 5088
rect 2744 5012 2760 5028
rect 2840 5112 2856 5128
rect 2888 5092 2904 5108
rect 2808 5032 2824 5048
rect 2840 5032 2856 5048
rect 2776 4972 2792 4988
rect 2712 4932 2728 4948
rect 2856 4912 2872 4928
rect 2792 4892 2808 4908
rect 2728 4812 2744 4828
rect 2776 4812 2792 4828
rect 2696 4792 2712 4808
rect 2600 4752 2616 4768
rect 2680 4752 2696 4768
rect 2552 4712 2568 4728
rect 2472 4652 2504 4668
rect 2504 4612 2520 4628
rect 2536 4652 2552 4668
rect 2568 4652 2600 4668
rect 2488 4532 2504 4548
rect 2456 4512 2472 4528
rect 2472 4472 2488 4488
rect 2456 4452 2472 4468
rect 2440 4352 2456 4368
rect 2456 4312 2472 4328
rect 2328 4292 2344 4308
rect 2360 4292 2376 4308
rect 2312 4212 2328 4228
rect 2296 4152 2312 4168
rect 2280 4092 2296 4108
rect 2312 4072 2328 4088
rect 2280 4032 2296 4048
rect 2152 3892 2168 3908
rect 2184 3852 2200 3868
rect 2104 3772 2120 3788
rect 2120 3772 2136 3788
rect 2264 3832 2280 3848
rect 2157 3802 2193 3818
rect 2248 3812 2264 3828
rect 2024 3732 2040 3748
rect 2200 3732 2216 3748
rect 1896 3712 1912 3728
rect 1960 3714 1976 3728
rect 1960 3712 1976 3714
rect 1928 3512 1944 3528
rect 2248 3712 2264 3728
rect 2104 3632 2120 3648
rect 2008 3532 2024 3548
rect 2056 3532 2072 3548
rect 1832 3492 1848 3508
rect 1784 3472 1800 3488
rect 1976 3452 1992 3468
rect 1944 3372 1960 3388
rect 1752 3352 1768 3368
rect 2072 3512 2088 3528
rect 2248 3512 2264 3528
rect 2072 3492 2088 3508
rect 2120 3492 2136 3508
rect 2152 3492 2168 3508
rect 2040 3472 2056 3488
rect 2104 3452 2120 3468
rect 2056 3372 2072 3388
rect 1688 3312 1704 3328
rect 1688 3292 1704 3308
rect 1736 3292 1752 3308
rect 1640 3112 1644 3128
rect 1644 3112 1656 3128
rect 1608 3092 1624 3108
rect 1656 3092 1672 3108
rect 1592 3072 1608 3088
rect 1832 3312 1848 3328
rect 1960 3312 1976 3328
rect 1960 3292 1976 3308
rect 1768 3132 1784 3148
rect 1816 3132 1832 3148
rect 1960 3132 1976 3148
rect 1688 3112 1720 3128
rect 1736 3092 1752 3108
rect 1912 3112 1928 3128
rect 1944 3112 1960 3128
rect 1672 3072 1688 3088
rect 1736 3072 1752 3088
rect 1800 3072 1816 3088
rect 1432 2792 1448 2808
rect 1464 2792 1480 2808
rect 1336 2772 1352 2788
rect 1384 2772 1400 2788
rect 1464 2772 1480 2788
rect 1480 2712 1496 2728
rect 1144 2652 1160 2668
rect 1112 2612 1128 2628
rect 1096 2572 1112 2588
rect 1080 2552 1096 2568
rect 1240 2672 1256 2688
rect 1320 2672 1336 2688
rect 1208 2632 1224 2648
rect 1192 2612 1208 2628
rect 1160 2572 1176 2588
rect 984 2532 1000 2548
rect 1448 2592 1464 2608
rect 1272 2532 1288 2548
rect 1432 2532 1448 2548
rect 984 2512 1000 2528
rect 1064 2512 1080 2528
rect 1384 2512 1400 2528
rect 968 2492 984 2508
rect 1016 2492 1032 2508
rect 1160 2492 1176 2508
rect 1117 2402 1153 2418
rect 952 2372 968 2388
rect 1144 2372 1160 2388
rect 904 2332 920 2348
rect 952 2332 968 2348
rect 1000 2332 1016 2348
rect 1032 2312 1064 2328
rect 840 2252 856 2268
rect 984 2272 1000 2288
rect 1032 2272 1048 2288
rect 1096 2272 1112 2288
rect 856 2172 872 2188
rect 1112 2252 1128 2268
rect 968 2212 984 2228
rect 1048 2172 1064 2188
rect 1176 2472 1192 2488
rect 1256 2412 1272 2428
rect 1176 2332 1192 2348
rect 1304 2312 1320 2328
rect 1256 2292 1272 2308
rect 920 2112 936 2128
rect 1000 2112 1016 2128
rect 1128 2112 1144 2128
rect 872 2072 888 2088
rect 856 2032 872 2048
rect 808 1932 824 1948
rect 840 1932 856 1948
rect 808 1912 824 1928
rect 1032 1992 1048 2008
rect 1096 1992 1112 2008
rect 1117 2002 1153 2018
rect 1000 1952 1016 1968
rect 1096 1972 1112 1988
rect 1096 1952 1112 1968
rect 1096 1932 1112 1948
rect 920 1912 936 1928
rect 952 1912 968 1928
rect 888 1892 904 1908
rect 1000 1892 1016 1908
rect 1016 1892 1032 1908
rect 872 1872 888 1888
rect 904 1872 920 1888
rect 920 1852 936 1868
rect 1016 1832 1032 1848
rect 1080 1892 1096 1908
rect 1224 2272 1240 2288
rect 1208 2252 1240 2268
rect 1176 2152 1192 2168
rect 1176 2092 1192 2108
rect 1208 1932 1224 1948
rect 1176 1912 1192 1928
rect 1160 1872 1176 1888
rect 952 1792 968 1808
rect 1032 1792 1048 1808
rect 936 1752 952 1768
rect 776 1732 792 1748
rect 856 1732 872 1748
rect 936 1732 952 1748
rect 744 1712 760 1728
rect 824 1712 840 1728
rect 568 1692 584 1708
rect 680 1692 696 1708
rect 824 1692 840 1708
rect 856 1692 872 1708
rect 824 1672 840 1688
rect 616 1572 632 1588
rect 616 1552 632 1568
rect 568 1532 584 1548
rect 600 1532 616 1548
rect 472 1512 488 1528
rect 744 1512 760 1528
rect 552 1492 568 1508
rect 824 1492 840 1508
rect 424 1472 440 1488
rect 568 1472 584 1488
rect 600 1472 616 1488
rect 616 1452 632 1468
rect 536 1432 552 1448
rect 296 1372 312 1388
rect 408 1352 424 1368
rect 456 1352 472 1368
rect 520 1352 536 1368
rect 200 1292 216 1308
rect 264 1292 280 1308
rect 280 1292 296 1308
rect 184 1132 200 1148
rect 200 1112 216 1128
rect 264 1112 280 1128
rect 312 1172 328 1188
rect 296 1132 312 1148
rect 72 1092 88 1108
rect 216 1092 232 1108
rect 376 1312 392 1328
rect 488 1332 504 1348
rect 584 1332 600 1348
rect 392 1272 408 1288
rect 360 1172 376 1188
rect 328 1092 344 1108
rect 120 1072 136 1088
rect 376 1072 392 1088
rect 472 1272 488 1288
rect 504 1292 520 1308
rect 552 1292 568 1308
rect 600 1292 616 1308
rect 488 1252 504 1268
rect 888 1712 904 1728
rect 984 1712 1000 1728
rect 920 1692 936 1708
rect 984 1692 1000 1708
rect 1080 1832 1096 1848
rect 1528 2772 1544 2788
rect 1560 2732 1576 2748
rect 1544 2672 1560 2688
rect 1608 2912 1624 2928
rect 1656 2912 1672 2928
rect 1640 2892 1656 2908
rect 1688 2952 1704 2968
rect 1944 3092 1960 3108
rect 1928 3072 1944 3088
rect 2040 3292 2056 3308
rect 2072 3292 2088 3308
rect 2072 3272 2088 3288
rect 2152 3472 2168 3488
rect 2296 3952 2312 3968
rect 2312 3892 2328 3908
rect 2392 4192 2408 4208
rect 2408 4172 2424 4188
rect 2456 4152 2472 4168
rect 2424 4072 2440 4088
rect 2424 4012 2440 4028
rect 2488 4272 2504 4288
rect 2552 4552 2568 4568
rect 2552 4532 2568 4548
rect 2584 4532 2600 4548
rect 2520 4492 2536 4508
rect 2536 4452 2552 4468
rect 2504 4232 2520 4248
rect 2488 4092 2504 4108
rect 2536 4032 2552 4048
rect 2392 3912 2408 3928
rect 2472 3912 2488 3928
rect 2488 3912 2504 3928
rect 2344 3892 2360 3908
rect 2456 3892 2472 3908
rect 2520 3892 2536 3908
rect 2424 3872 2456 3888
rect 2680 4712 2696 4728
rect 2632 4652 2648 4668
rect 2680 4652 2696 4668
rect 2648 4632 2664 4648
rect 2616 4612 2632 4628
rect 2904 4952 2920 4968
rect 2872 4872 2904 4888
rect 2792 4732 2808 4748
rect 2808 4712 2824 4728
rect 2808 4692 2824 4708
rect 2840 4712 2856 4728
rect 2920 4912 2936 4928
rect 2984 5232 3000 5248
rect 2984 5092 3000 5108
rect 2968 5072 2984 5088
rect 3304 5272 3320 5288
rect 3165 5202 3201 5218
rect 3032 5052 3048 5068
rect 3112 5052 3128 5068
rect 3016 5012 3032 5028
rect 3112 5032 3128 5048
rect 2952 4992 2968 5008
rect 3032 4992 3048 5008
rect 3064 4932 3080 4948
rect 3096 4912 3112 4928
rect 3080 4892 3096 4908
rect 3112 4892 3128 4908
rect 2984 4872 3000 4888
rect 2936 4772 2952 4788
rect 2760 4672 2776 4688
rect 2872 4672 2888 4688
rect 2776 4572 2792 4588
rect 2872 4632 2888 4648
rect 2936 4632 2952 4648
rect 2872 4612 2888 4628
rect 2920 4592 2936 4608
rect 2616 4552 2632 4568
rect 2744 4552 2760 4568
rect 2680 4532 2696 4548
rect 2760 4532 2776 4548
rect 2824 4552 2840 4568
rect 2952 4612 2968 4628
rect 2616 4512 2632 4528
rect 2760 4512 2776 4528
rect 2568 4492 2584 4508
rect 2584 4352 2600 4368
rect 2600 4312 2616 4328
rect 2584 4292 2600 4308
rect 2568 4212 2584 4228
rect 2600 4092 2616 4108
rect 2664 4492 2680 4508
rect 2952 4492 2968 4508
rect 2840 4432 2856 4448
rect 2888 4432 2904 4448
rect 2920 4432 2936 4448
rect 2824 4392 2840 4408
rect 2712 4292 2728 4308
rect 2808 4292 2824 4308
rect 2664 4272 2680 4288
rect 2664 4232 2680 4248
rect 2744 4192 2760 4208
rect 2776 4152 2792 4168
rect 2712 4132 2728 4148
rect 2632 4112 2664 4128
rect 2696 4112 2712 4128
rect 2632 4092 2648 4108
rect 2616 4072 2632 4088
rect 2424 3852 2440 3868
rect 2536 3852 2552 3868
rect 2520 3812 2536 3828
rect 2376 3772 2392 3788
rect 2600 3952 2616 3968
rect 2584 3872 2600 3888
rect 2856 4272 2872 4288
rect 2904 4272 2920 4288
rect 2824 4132 2840 4148
rect 2872 4132 2888 4148
rect 2888 4112 2904 4128
rect 2952 4172 2968 4188
rect 2952 4132 2968 4148
rect 2792 4092 2808 4108
rect 2840 4092 2856 4108
rect 2920 4092 2936 4108
rect 3128 4732 3144 4748
rect 3432 5312 3448 5328
rect 3432 5272 3448 5288
rect 3576 5372 3592 5388
rect 3512 5352 3528 5368
rect 3640 5372 3656 5388
rect 3512 5332 3528 5348
rect 3528 5332 3544 5348
rect 3592 5332 3608 5348
rect 3624 5332 3640 5348
rect 3480 5312 3496 5328
rect 3560 5312 3576 5328
rect 3480 5272 3496 5288
rect 3592 5272 3608 5288
rect 3384 5232 3400 5248
rect 3352 5112 3368 5128
rect 3304 5032 3320 5048
rect 3368 5012 3384 5028
rect 3224 4952 3240 4968
rect 3272 4932 3288 4948
rect 3160 4912 3176 4928
rect 3224 4852 3240 4868
rect 3165 4802 3201 4818
rect 3336 4832 3352 4848
rect 3208 4752 3224 4768
rect 3384 4832 3400 4848
rect 3656 5112 3672 5128
rect 3416 4952 3432 4968
rect 3432 4932 3448 4948
rect 3432 4892 3448 4908
rect 3400 4772 3416 4788
rect 3416 4752 3432 4768
rect 3240 4732 3256 4748
rect 3368 4732 3384 4748
rect 3320 4712 3336 4728
rect 3368 4712 3384 4728
rect 3128 4692 3144 4708
rect 3208 4692 3224 4708
rect 3272 4692 3288 4708
rect 3352 4692 3368 4708
rect 3032 4632 3048 4648
rect 3064 4592 3080 4608
rect 3032 4572 3048 4588
rect 3000 4552 3016 4568
rect 3064 4552 3080 4568
rect 3000 4512 3016 4528
rect 3096 4514 3112 4528
rect 3096 4512 3112 4514
rect 3000 4492 3016 4508
rect 3192 4452 3208 4468
rect 3128 4392 3144 4408
rect 3165 4402 3201 4418
rect 3032 4312 3048 4328
rect 3000 4292 3016 4308
rect 3064 4292 3080 4308
rect 3112 4292 3128 4308
rect 3144 4312 3160 4328
rect 3064 4272 3080 4288
rect 3112 4272 3128 4288
rect 3048 4252 3064 4268
rect 3272 4652 3288 4668
rect 3272 4632 3288 4648
rect 3224 4612 3240 4628
rect 3224 4572 3240 4588
rect 3256 4532 3272 4548
rect 3288 4532 3304 4548
rect 3288 4512 3304 4528
rect 3336 4512 3352 4528
rect 3304 4492 3316 4508
rect 3316 4492 3320 4508
rect 3336 4432 3352 4448
rect 3496 4972 3512 4988
rect 3496 4952 3512 4968
rect 3688 5072 3704 5088
rect 3656 4992 3672 5008
rect 3544 4952 3560 4968
rect 3720 5232 3736 5248
rect 3800 5372 3816 5388
rect 3784 5312 3800 5328
rect 3768 5272 3784 5288
rect 3752 5232 3768 5248
rect 3832 5312 3848 5328
rect 3896 5412 3912 5428
rect 3928 5412 3944 5428
rect 3880 5292 3896 5308
rect 3928 5332 3944 5348
rect 3960 5312 3976 5328
rect 3912 5232 3928 5248
rect 4205 5402 4241 5418
rect 4360 5372 4376 5388
rect 4072 5312 4088 5328
rect 4312 5312 4328 5328
rect 4424 5312 4440 5328
rect 3992 5252 4008 5268
rect 3736 5112 3752 5128
rect 3896 5092 3912 5108
rect 3944 5092 3960 5108
rect 3736 5052 3752 5068
rect 3512 4932 3528 4948
rect 3560 4932 3576 4948
rect 3480 4892 3496 4908
rect 3496 4792 3512 4808
rect 3608 4912 3624 4928
rect 3592 4892 3608 4908
rect 3544 4792 3560 4808
rect 3640 4892 3656 4908
rect 3816 4992 3832 5008
rect 3832 4952 3848 4968
rect 3880 4952 3896 4968
rect 3816 4932 3832 4948
rect 3896 4932 3912 4948
rect 3736 4912 3752 4928
rect 3784 4912 3800 4928
rect 3864 4912 3880 4928
rect 3688 4852 3704 4868
rect 3720 4852 3736 4868
rect 3672 4812 3688 4828
rect 3640 4772 3656 4788
rect 3544 4752 3560 4768
rect 3720 4812 3736 4828
rect 3640 4732 3656 4748
rect 3688 4732 3704 4748
rect 3576 4712 3592 4728
rect 3448 4692 3464 4708
rect 3624 4692 3640 4708
rect 3704 4692 3720 4708
rect 3608 4672 3624 4688
rect 3496 4652 3512 4668
rect 3416 4632 3432 4648
rect 3448 4572 3464 4588
rect 3416 4532 3432 4548
rect 3496 4492 3512 4508
rect 3400 4412 3416 4428
rect 3432 4412 3448 4428
rect 3464 4412 3480 4428
rect 3336 4312 3352 4328
rect 3128 4232 3144 4248
rect 3048 4212 3064 4228
rect 3000 4152 3016 4168
rect 3032 4132 3048 4148
rect 3160 4172 3176 4188
rect 3256 4152 3272 4168
rect 3128 4132 3144 4148
rect 3208 4092 3224 4108
rect 3320 4172 3336 4188
rect 3400 4172 3416 4188
rect 3464 4352 3480 4368
rect 3448 4332 3464 4348
rect 3480 4312 3496 4328
rect 3480 4292 3496 4308
rect 3480 4272 3496 4288
rect 3576 4652 3592 4668
rect 3560 4572 3576 4588
rect 3544 4512 3560 4528
rect 3576 4392 3592 4408
rect 3720 4672 3736 4688
rect 3720 4652 3736 4668
rect 3672 4572 3688 4588
rect 3656 4532 3672 4548
rect 3640 4352 3656 4368
rect 3560 4332 3576 4348
rect 3528 4292 3544 4308
rect 3592 4312 3608 4328
rect 3592 4272 3608 4288
rect 3624 4272 3640 4288
rect 3512 4212 3528 4228
rect 3336 4132 3352 4148
rect 3352 4112 3368 4128
rect 3432 4112 3448 4128
rect 3448 4112 3464 4128
rect 3352 4092 3368 4108
rect 2888 4072 2904 4088
rect 2984 4072 3000 4088
rect 2760 4012 2776 4028
rect 2648 3972 2664 3988
rect 2584 3852 2600 3868
rect 2568 3812 2584 3828
rect 2552 3792 2568 3808
rect 2552 3752 2568 3768
rect 2568 3732 2584 3748
rect 2408 3712 2424 3728
rect 2520 3712 2536 3728
rect 2568 3712 2584 3728
rect 2392 3692 2408 3708
rect 2424 3692 2440 3708
rect 2360 3672 2376 3688
rect 2488 3672 2504 3688
rect 2328 3512 2344 3528
rect 2376 3512 2392 3528
rect 2296 3492 2312 3508
rect 2312 3492 2328 3508
rect 2392 3492 2408 3508
rect 2472 3492 2488 3508
rect 2296 3472 2312 3488
rect 2344 3472 2360 3488
rect 2216 3432 2232 3448
rect 2136 3392 2152 3408
rect 2157 3402 2193 3418
rect 2216 3412 2232 3428
rect 2424 3452 2440 3468
rect 2328 3412 2344 3428
rect 2472 3412 2488 3428
rect 2504 3412 2520 3428
rect 2264 3372 2280 3388
rect 2184 3352 2200 3368
rect 2456 3352 2472 3368
rect 2248 3332 2264 3348
rect 2280 3332 2296 3348
rect 2440 3332 2456 3348
rect 2760 3932 2776 3948
rect 2712 3892 2728 3908
rect 2696 3852 2712 3868
rect 2792 3752 2808 3768
rect 2616 3672 2632 3688
rect 2552 3432 2568 3448
rect 2584 3432 2600 3448
rect 2616 3492 2632 3508
rect 2616 3332 2632 3348
rect 2392 3312 2408 3328
rect 2472 3312 2488 3328
rect 2520 3312 2536 3328
rect 2968 3952 2984 3968
rect 2968 3912 2984 3928
rect 2808 3712 2824 3728
rect 2664 3692 2680 3708
rect 2808 3692 2824 3708
rect 2856 3772 2872 3788
rect 3165 4002 3201 4018
rect 3272 3972 3288 3988
rect 3320 3972 3336 3988
rect 3112 3912 3128 3928
rect 3096 3892 3112 3908
rect 3112 3892 3128 3908
rect 3160 3892 3176 3908
rect 3080 3832 3096 3848
rect 3032 3772 3048 3788
rect 3000 3752 3016 3768
rect 2920 3732 2936 3748
rect 2664 3552 2680 3568
rect 2696 3492 2712 3508
rect 2680 3472 2696 3488
rect 2760 3392 2776 3408
rect 2936 3532 2952 3548
rect 2792 3492 2808 3508
rect 3048 3732 3064 3748
rect 3080 3712 3096 3728
rect 3048 3692 3064 3708
rect 3240 3872 3256 3888
rect 3192 3832 3208 3848
rect 3144 3772 3160 3788
rect 3288 3832 3304 3848
rect 3128 3692 3144 3708
rect 3096 3632 3112 3648
rect 3165 3602 3201 3618
rect 3000 3552 3016 3568
rect 3224 3552 3240 3568
rect 3016 3532 3032 3548
rect 3160 3532 3176 3548
rect 2968 3492 2984 3508
rect 3016 3492 3032 3508
rect 2952 3472 2968 3488
rect 2808 3452 2824 3468
rect 2888 3432 2904 3448
rect 2904 3392 2920 3408
rect 2968 3352 2984 3368
rect 2952 3332 2968 3348
rect 2680 3312 2696 3328
rect 2840 3312 2856 3328
rect 2280 3292 2296 3308
rect 2344 3292 2360 3308
rect 2488 3292 2504 3308
rect 2600 3292 2616 3308
rect 2632 3292 2648 3308
rect 2696 3292 2712 3308
rect 2264 3272 2280 3288
rect 2120 3252 2136 3268
rect 2184 3252 2200 3268
rect 2008 3212 2024 3228
rect 2136 3132 2152 3148
rect 1992 3112 2008 3128
rect 2072 3112 2088 3128
rect 2008 3092 2024 3108
rect 1976 3072 1992 3088
rect 1880 2952 1896 2968
rect 1960 2952 1976 2968
rect 1752 2892 1768 2908
rect 1672 2872 1688 2888
rect 1704 2872 1720 2888
rect 1608 2772 1624 2788
rect 1576 2532 1592 2548
rect 1672 2752 1688 2768
rect 1848 2752 1864 2768
rect 1768 2732 1784 2748
rect 1848 2732 1864 2748
rect 1752 2712 1784 2728
rect 1816 2712 1832 2728
rect 1736 2672 1752 2688
rect 1768 2652 1784 2668
rect 1496 2512 1512 2528
rect 1528 2512 1544 2528
rect 1608 2512 1624 2528
rect 1672 2512 1688 2528
rect 1416 2492 1432 2508
rect 1464 2492 1480 2508
rect 1464 2452 1480 2468
rect 1432 2432 1448 2448
rect 1432 2292 1448 2308
rect 1640 2492 1656 2508
rect 1576 2452 1592 2468
rect 1512 2412 1528 2428
rect 1512 2332 1528 2348
rect 1528 2312 1544 2328
rect 1416 2272 1432 2288
rect 1464 2272 1480 2288
rect 1624 2372 1640 2388
rect 1656 2352 1672 2368
rect 1736 2592 1752 2608
rect 1576 2332 1592 2348
rect 1704 2332 1720 2348
rect 1656 2312 1672 2328
rect 1592 2272 1608 2288
rect 1320 2252 1336 2268
rect 1400 2252 1416 2268
rect 1464 2252 1480 2268
rect 1544 2252 1560 2268
rect 1320 2232 1336 2248
rect 1416 2192 1432 2208
rect 1304 2172 1320 2188
rect 1288 2132 1304 2148
rect 1432 2152 1448 2168
rect 1496 2152 1512 2168
rect 1704 2292 1720 2308
rect 1592 2232 1608 2248
rect 1624 2232 1640 2248
rect 1576 2172 1592 2188
rect 1384 2112 1400 2128
rect 1528 2112 1544 2128
rect 1592 2112 1608 2128
rect 1608 2112 1624 2128
rect 1256 2032 1272 2048
rect 1208 1892 1240 1908
rect 1208 1852 1224 1868
rect 1224 1832 1240 1848
rect 1272 1832 1288 1848
rect 1176 1812 1192 1828
rect 1080 1792 1096 1808
rect 1064 1772 1080 1788
rect 1064 1712 1080 1728
rect 1048 1692 1064 1708
rect 1176 1772 1192 1788
rect 1416 2072 1432 2088
rect 1304 1952 1320 1968
rect 1624 2092 1640 2108
rect 1592 2052 1608 2068
rect 1688 2052 1704 2068
rect 1560 2032 1576 2048
rect 1528 2012 1544 2028
rect 1512 1932 1528 1948
rect 1448 1912 1464 1928
rect 1656 1992 1672 2008
rect 1624 1932 1640 1948
rect 1400 1892 1416 1908
rect 1432 1892 1448 1908
rect 1320 1872 1336 1888
rect 1320 1852 1336 1868
rect 1304 1812 1320 1828
rect 1288 1712 1304 1728
rect 1160 1692 1176 1708
rect 1117 1602 1153 1618
rect 920 1512 936 1528
rect 1016 1512 1048 1528
rect 1080 1512 1096 1528
rect 1080 1492 1096 1508
rect 872 1452 888 1468
rect 680 1432 696 1448
rect 680 1372 696 1388
rect 744 1372 760 1388
rect 728 1332 744 1348
rect 808 1332 824 1348
rect 664 1312 680 1328
rect 568 1172 584 1188
rect 520 1132 536 1148
rect 552 1132 568 1148
rect 696 1152 712 1168
rect 632 1092 648 1108
rect 680 1092 696 1108
rect 200 1052 216 1068
rect 376 1052 408 1068
rect 184 952 200 968
rect 360 992 376 1008
rect 296 952 312 968
rect 72 912 88 928
rect 232 912 248 928
rect 216 892 232 908
rect 264 892 280 908
rect 328 892 344 908
rect 136 712 152 728
rect 216 692 248 708
rect 328 692 344 708
rect 40 632 56 648
rect 200 572 216 588
rect 56 532 72 548
rect 168 552 184 568
rect 24 512 40 528
rect 152 512 168 528
rect 8 492 24 508
rect 248 632 264 648
rect 296 592 312 608
rect 344 592 360 608
rect 232 492 264 508
rect 120 312 136 328
rect 184 312 200 328
rect 88 292 104 308
rect 120 272 136 288
rect 232 292 248 308
rect 440 952 456 968
rect 472 952 488 968
rect 600 1052 616 1068
rect 584 1012 600 1028
rect 520 992 536 1008
rect 648 1052 664 1068
rect 568 972 584 988
rect 632 972 648 988
rect 488 912 504 928
rect 504 912 520 928
rect 456 752 472 768
rect 440 712 456 728
rect 472 692 504 708
rect 456 672 472 688
rect 424 652 440 668
rect 376 532 392 548
rect 392 492 408 508
rect 360 472 376 488
rect 376 452 392 468
rect 456 592 472 608
rect 440 472 456 488
rect 312 372 328 388
rect 408 372 456 388
rect 264 272 280 288
rect 312 272 328 288
rect 280 112 296 128
rect 520 712 536 728
rect 552 912 568 928
rect 680 952 696 968
rect 616 932 632 948
rect 632 912 648 928
rect 616 892 632 908
rect 584 712 600 728
rect 488 552 504 568
rect 472 512 488 528
rect 488 512 504 528
rect 472 492 488 508
rect 504 472 520 488
rect 568 692 600 708
rect 616 692 648 708
rect 536 552 552 568
rect 568 612 584 628
rect 680 672 696 688
rect 632 632 648 648
rect 680 592 696 608
rect 584 552 600 568
rect 552 492 568 508
rect 520 452 536 468
rect 472 332 488 348
rect 568 372 584 388
rect 536 312 552 328
rect 648 512 664 528
rect 632 492 648 508
rect 632 472 648 488
rect 664 472 680 488
rect 600 372 632 388
rect 680 332 696 348
rect 728 1112 744 1128
rect 840 1312 856 1328
rect 808 1052 824 1068
rect 712 1032 728 1048
rect 712 972 728 988
rect 744 952 760 968
rect 952 1472 968 1488
rect 888 1412 904 1428
rect 936 1352 952 1368
rect 968 1332 984 1348
rect 968 1312 984 1328
rect 952 1292 968 1308
rect 984 1292 1000 1308
rect 952 1112 968 1128
rect 888 1092 904 1108
rect 952 1092 968 1108
rect 984 1092 1000 1108
rect 936 1072 952 1088
rect 888 1052 904 1068
rect 920 1052 936 1068
rect 856 992 872 1008
rect 904 972 920 988
rect 920 932 936 948
rect 792 912 808 928
rect 936 912 952 928
rect 824 892 840 908
rect 920 892 936 908
rect 808 732 824 748
rect 744 672 760 688
rect 712 532 728 548
rect 712 512 728 528
rect 792 512 808 528
rect 728 332 744 348
rect 600 312 616 328
rect 712 312 728 328
rect 584 292 600 308
rect 680 292 696 308
rect 808 312 824 328
rect 920 832 936 848
rect 904 712 920 728
rect 936 732 952 748
rect 904 672 920 688
rect 936 652 952 668
rect 984 1072 1000 1088
rect 1144 1432 1160 1448
rect 1080 1392 1096 1408
rect 1048 1352 1064 1368
rect 1016 1292 1032 1308
rect 1256 1506 1272 1508
rect 1256 1492 1272 1506
rect 1160 1392 1176 1408
rect 1192 1392 1208 1408
rect 1144 1312 1160 1328
rect 1208 1314 1224 1328
rect 1208 1312 1224 1314
rect 1224 1292 1240 1308
rect 1064 1272 1080 1288
rect 1117 1202 1153 1218
rect 1224 1172 1240 1188
rect 1160 1132 1176 1148
rect 1176 1132 1192 1148
rect 1096 1112 1112 1128
rect 1208 1112 1224 1128
rect 1192 1092 1208 1108
rect 1032 1072 1048 1088
rect 1160 1072 1176 1088
rect 1192 1072 1208 1088
rect 1000 1052 1032 1068
rect 984 992 1000 1008
rect 968 932 984 948
rect 1016 972 1032 988
rect 984 892 1000 908
rect 968 752 1000 768
rect 952 632 968 648
rect 1064 1052 1080 1068
rect 1048 912 1064 928
rect 1016 732 1032 748
rect 1016 712 1032 728
rect 1176 1032 1192 1048
rect 1192 972 1208 988
rect 1176 932 1192 948
rect 1080 912 1096 928
rect 1144 912 1160 928
rect 1288 1152 1304 1168
rect 1384 1852 1400 1868
rect 1336 1772 1352 1788
rect 1400 1772 1416 1788
rect 1320 1672 1352 1688
rect 1400 1512 1416 1528
rect 1400 1472 1416 1488
rect 1368 1432 1384 1448
rect 1384 1432 1400 1448
rect 1336 1392 1352 1408
rect 1528 1872 1544 1888
rect 1432 1792 1448 1808
rect 1512 1812 1528 1828
rect 1560 1812 1576 1828
rect 1512 1732 1528 1748
rect 1448 1712 1464 1728
rect 1480 1712 1496 1728
rect 1448 1692 1464 1708
rect 1496 1692 1512 1708
rect 1576 1714 1592 1728
rect 1576 1712 1592 1714
rect 1496 1672 1512 1688
rect 1544 1672 1560 1688
rect 1592 1652 1608 1668
rect 1448 1552 1464 1568
rect 1416 1372 1448 1388
rect 1400 1352 1416 1368
rect 1560 1512 1576 1528
rect 1528 1432 1544 1448
rect 1464 1412 1480 1428
rect 1464 1372 1480 1388
rect 1512 1372 1528 1388
rect 1416 1312 1432 1328
rect 1560 1392 1576 1408
rect 1544 1372 1560 1388
rect 1800 2532 1816 2548
rect 1752 2412 1768 2428
rect 1720 2232 1736 2248
rect 1720 2212 1736 2228
rect 1800 2492 1816 2508
rect 1880 2712 1896 2728
rect 1864 2692 1880 2708
rect 1880 2672 1896 2688
rect 1928 2632 1944 2648
rect 2056 3072 2072 3088
rect 2040 3052 2056 3068
rect 2344 3252 2360 3268
rect 2376 3252 2392 3268
rect 2376 3232 2392 3248
rect 2104 3092 2120 3108
rect 2216 3092 2232 3108
rect 2184 3072 2200 3088
rect 2072 3032 2088 3048
rect 2024 2912 2040 2928
rect 2088 2912 2104 2928
rect 2157 3002 2193 3018
rect 2232 2972 2248 2988
rect 2152 2912 2168 2928
rect 2216 2914 2232 2928
rect 2216 2912 2232 2914
rect 2264 2912 2280 2928
rect 2072 2892 2088 2908
rect 1960 2772 1976 2788
rect 2056 2772 2072 2788
rect 2168 2832 2184 2848
rect 2072 2752 2088 2768
rect 2120 2752 2136 2768
rect 2232 2752 2248 2768
rect 1976 2732 1992 2748
rect 2104 2732 2120 2748
rect 2088 2712 2104 2728
rect 2088 2692 2104 2708
rect 2008 2652 2024 2668
rect 1944 2612 1960 2628
rect 1848 2512 1864 2528
rect 1848 2492 1864 2508
rect 1992 2512 2008 2528
rect 2056 2652 2072 2668
rect 2024 2632 2040 2648
rect 2072 2592 2088 2608
rect 2072 2572 2088 2588
rect 2472 3132 2488 3148
rect 2504 3252 2520 3268
rect 2728 3232 2744 3248
rect 2760 3232 2776 3248
rect 2520 3132 2536 3148
rect 2392 3092 2408 3108
rect 2344 2972 2360 2988
rect 2408 3072 2424 3088
rect 2424 3012 2440 3028
rect 2616 3092 2632 3108
rect 2552 3072 2568 3088
rect 2712 3052 2728 3068
rect 2792 3192 2808 3208
rect 2760 3092 2776 3108
rect 2776 3072 2792 3088
rect 2600 2952 2616 2968
rect 2792 3052 2808 3068
rect 2840 3152 2856 3168
rect 2936 3152 2952 3168
rect 2824 3092 2840 3108
rect 2824 3072 2840 3088
rect 2904 3132 2920 3148
rect 2872 3092 2888 3108
rect 2888 3092 2920 3108
rect 2872 3072 2888 3088
rect 2744 2952 2760 2968
rect 2808 2952 2824 2968
rect 2840 2952 2856 2968
rect 3096 3472 3112 3488
rect 3032 3432 3048 3448
rect 3096 3392 3112 3408
rect 3080 3372 3096 3388
rect 3176 3372 3192 3388
rect 3352 3792 3368 3808
rect 3320 3752 3352 3768
rect 3288 3732 3304 3748
rect 3320 3712 3336 3728
rect 3320 3692 3336 3708
rect 3256 3632 3272 3648
rect 3272 3532 3288 3548
rect 3304 3532 3320 3548
rect 3336 3672 3352 3688
rect 3464 3852 3480 3868
rect 3384 3752 3400 3768
rect 3448 3812 3464 3828
rect 3416 3712 3432 3728
rect 3384 3652 3400 3668
rect 3304 3472 3320 3488
rect 3352 3472 3368 3488
rect 3384 3472 3400 3488
rect 3336 3432 3352 3448
rect 3272 3392 3288 3408
rect 3272 3352 3288 3368
rect 3432 3572 3448 3588
rect 3400 3432 3416 3448
rect 3368 3392 3384 3408
rect 3432 3392 3448 3408
rect 3256 3332 3272 3348
rect 3320 3332 3336 3348
rect 3256 3312 3272 3328
rect 3304 3312 3320 3328
rect 3480 3512 3496 3528
rect 3480 3492 3496 3508
rect 3640 4192 3656 4208
rect 3640 4172 3656 4188
rect 3640 4152 3656 4168
rect 3608 4132 3624 4148
rect 3816 4892 3832 4908
rect 3976 4952 3992 4968
rect 3976 4912 3992 4928
rect 4056 5132 4072 5148
rect 4120 5292 4136 5308
rect 4328 5292 4344 5308
rect 4216 5232 4232 5248
rect 4392 5132 4408 5148
rect 4360 5112 4376 5128
rect 4296 5092 4312 5108
rect 4328 5092 4344 5108
rect 4360 5092 4376 5108
rect 4232 5072 4248 5088
rect 4328 5072 4344 5088
rect 4216 5032 4232 5048
rect 4205 5002 4241 5018
rect 4168 4952 4184 4968
rect 4312 5052 4328 5068
rect 4200 4932 4216 4948
rect 4296 4932 4312 4948
rect 4104 4914 4120 4928
rect 4104 4912 4120 4914
rect 4200 4912 4216 4928
rect 4280 4912 4296 4928
rect 4312 4912 4328 4928
rect 4040 4892 4056 4908
rect 4232 4892 4248 4908
rect 3912 4872 3928 4888
rect 3928 4872 3944 4888
rect 3912 4852 3928 4868
rect 3768 4732 3784 4748
rect 3752 4692 3768 4708
rect 3816 4612 3832 4628
rect 3736 4572 3752 4588
rect 3784 4512 3800 4528
rect 3720 4492 3736 4508
rect 3704 4472 3720 4488
rect 3736 4452 3752 4468
rect 3752 4432 3768 4448
rect 3720 4352 3736 4368
rect 3704 4292 3720 4308
rect 3704 4272 3720 4288
rect 3560 4112 3576 4128
rect 3592 4112 3608 4128
rect 3656 4112 3672 4128
rect 3544 4092 3560 4108
rect 3624 4092 3640 4108
rect 3656 4092 3672 4108
rect 3512 4072 3528 4088
rect 3608 4052 3624 4068
rect 3656 4072 3672 4088
rect 3624 3972 3640 3988
rect 3560 3912 3576 3928
rect 3512 3872 3528 3888
rect 3560 3872 3576 3888
rect 3512 3832 3528 3848
rect 3528 3752 3544 3768
rect 3560 3752 3576 3768
rect 3528 3712 3544 3728
rect 3544 3632 3560 3648
rect 3784 4272 3800 4288
rect 3736 4232 3768 4248
rect 3800 4232 3816 4248
rect 3832 4512 3848 4528
rect 3880 4692 3896 4708
rect 3976 4552 3992 4568
rect 4056 4552 4072 4568
rect 4040 4532 4056 4548
rect 4120 4532 4136 4548
rect 3944 4492 3960 4508
rect 3864 4332 3880 4348
rect 3832 4292 3848 4308
rect 3960 4272 3976 4288
rect 3928 4212 3944 4228
rect 3768 4172 3784 4188
rect 3704 4152 3736 4168
rect 3688 4132 3704 4148
rect 3672 3892 3688 3908
rect 3720 4052 3736 4068
rect 3752 4032 3768 4048
rect 3784 4012 3800 4028
rect 3784 3892 3800 3908
rect 3800 3872 3816 3888
rect 3848 4112 3864 4128
rect 3864 4092 3880 4108
rect 3912 4092 3928 4108
rect 3848 4072 3864 4088
rect 3832 4032 3848 4048
rect 3864 4012 3880 4028
rect 3656 3832 3672 3848
rect 3736 3832 3752 3848
rect 3640 3752 3656 3768
rect 3672 3752 3688 3768
rect 3640 3712 3656 3728
rect 3624 3692 3640 3708
rect 3544 3612 3560 3628
rect 3576 3612 3592 3628
rect 3656 3672 3672 3688
rect 3592 3592 3608 3608
rect 3576 3552 3592 3568
rect 3752 3752 3768 3768
rect 3784 3752 3800 3768
rect 3752 3732 3768 3748
rect 3768 3632 3784 3648
rect 3704 3612 3720 3628
rect 3768 3612 3784 3628
rect 3768 3532 3784 3548
rect 3640 3492 3656 3508
rect 3672 3492 3688 3508
rect 3528 3472 3544 3488
rect 3736 3472 3752 3488
rect 3784 3492 3800 3508
rect 3752 3452 3768 3468
rect 3496 3392 3512 3408
rect 3464 3372 3480 3388
rect 3688 3372 3704 3388
rect 3944 4032 3960 4048
rect 3928 4012 3944 4028
rect 4072 4512 4088 4528
rect 4104 4512 4120 4528
rect 4168 4512 4184 4528
rect 4008 4492 4024 4508
rect 4056 4492 4072 4508
rect 4264 4732 4280 4748
rect 4312 4732 4328 4748
rect 4376 5072 4392 5088
rect 4440 5092 4456 5108
rect 4504 5412 4520 5428
rect 4536 5412 4552 5428
rect 4552 5372 4568 5388
rect 4568 5372 4584 5388
rect 4632 5372 4648 5388
rect 4728 5412 4744 5428
rect 4792 5412 4808 5428
rect 4936 5412 4952 5428
rect 5320 5412 5336 5428
rect 5368 5412 5384 5428
rect 4840 5392 4856 5408
rect 5432 5392 5448 5408
rect 5528 5352 5544 5368
rect 5576 5352 5592 5368
rect 6237 5402 6273 5418
rect 6680 5372 6696 5388
rect 6120 5352 6136 5368
rect 6392 5352 6408 5368
rect 4696 5332 4712 5348
rect 4744 5332 4760 5348
rect 4840 5332 4856 5348
rect 5064 5332 5080 5348
rect 5192 5332 5208 5348
rect 5448 5332 5464 5348
rect 5976 5332 5992 5348
rect 6008 5332 6024 5348
rect 4488 5292 4504 5308
rect 4488 5272 4504 5288
rect 4584 5312 4600 5328
rect 4664 5312 4680 5328
rect 4776 5312 4792 5328
rect 4824 5312 4840 5328
rect 4600 5292 4604 5308
rect 4604 5292 4616 5308
rect 4648 5292 4664 5308
rect 4520 5232 4536 5248
rect 4488 5132 4504 5148
rect 4472 5092 4488 5108
rect 4504 5112 4520 5128
rect 4424 5052 4440 5068
rect 4376 4992 4392 5008
rect 4360 4892 4376 4908
rect 4200 4712 4216 4728
rect 4232 4692 4248 4708
rect 4205 4602 4241 4618
rect 4248 4592 4264 4608
rect 4296 4612 4312 4628
rect 4280 4532 4296 4548
rect 4056 4472 4072 4488
rect 4120 4472 4136 4488
rect 4184 4472 4200 4488
rect 3992 4412 4008 4428
rect 4184 4432 4200 4448
rect 4104 4412 4120 4428
rect 4056 4312 4088 4328
rect 4008 4252 4024 4268
rect 4008 4232 4024 4248
rect 3976 4172 3992 4188
rect 3976 4152 3992 4168
rect 3976 4092 3992 4108
rect 3928 3972 3944 3988
rect 3848 3912 3864 3928
rect 4296 4372 4312 4388
rect 4264 4352 4280 4368
rect 4200 4312 4216 4328
rect 4168 4292 4184 4308
rect 4120 4272 4136 4288
rect 4168 4272 4184 4288
rect 4296 4272 4312 4288
rect 4264 4252 4280 4268
rect 4205 4202 4241 4218
rect 4248 4172 4264 4188
rect 4024 4132 4040 4148
rect 4024 4092 4040 4108
rect 4008 3952 4024 3968
rect 3976 3932 3992 3948
rect 3912 3912 3928 3928
rect 3896 3832 3912 3848
rect 3848 3792 3864 3808
rect 3992 3852 4008 3868
rect 4152 4132 4168 4148
rect 4136 4112 4152 4128
rect 4120 4092 4136 4108
rect 4088 4072 4104 4088
rect 4056 3952 4072 3968
rect 4088 3912 4104 3928
rect 4056 3892 4072 3908
rect 3992 3812 4008 3828
rect 3896 3772 3912 3788
rect 4104 3772 4120 3788
rect 4200 3992 4216 4008
rect 4168 3952 4184 3968
rect 4168 3892 4184 3908
rect 4280 4132 4296 4148
rect 4280 4092 4296 4108
rect 4408 4892 4424 4908
rect 4408 4812 4424 4828
rect 4456 4892 4472 4908
rect 4456 4712 4472 4728
rect 4424 4692 4440 4708
rect 4520 5072 4536 5088
rect 4648 5052 4664 5068
rect 4504 5032 4520 5048
rect 4536 5032 4552 5048
rect 4744 5292 4760 5308
rect 4808 5292 4824 5308
rect 4712 5272 4728 5288
rect 4776 5252 4792 5268
rect 4744 5112 4760 5128
rect 5176 5312 5192 5328
rect 5288 5314 5304 5328
rect 5288 5312 5304 5314
rect 5464 5312 5480 5328
rect 5640 5312 5656 5328
rect 5832 5312 5848 5328
rect 4904 5292 4920 5308
rect 4968 5252 4984 5268
rect 4968 5232 4984 5248
rect 4888 5132 4904 5148
rect 4824 5092 4840 5108
rect 4856 5092 4888 5108
rect 4696 4992 4712 5008
rect 4792 5052 4808 5068
rect 4776 5032 4792 5048
rect 4600 4952 4616 4968
rect 4792 4952 4808 4968
rect 4808 4932 4824 4948
rect 4728 4914 4744 4928
rect 4728 4912 4744 4914
rect 4568 4832 4584 4848
rect 4488 4812 4504 4828
rect 4488 4792 4504 4808
rect 4840 4992 4856 5008
rect 4968 5112 4984 5128
rect 5048 5112 5064 5128
rect 4920 5092 4936 5108
rect 4968 5092 4984 5108
rect 4872 4952 4888 4968
rect 4984 5072 5000 5088
rect 5000 4952 5016 4968
rect 4872 4932 4888 4948
rect 4984 4932 5000 4948
rect 4840 4912 4856 4928
rect 4792 4892 4808 4908
rect 4856 4892 4872 4908
rect 4728 4832 4744 4848
rect 4664 4712 4680 4728
rect 4440 4652 4456 4668
rect 4376 4592 4392 4608
rect 4344 4532 4360 4548
rect 4360 4532 4376 4548
rect 4360 4512 4376 4528
rect 4520 4672 4536 4688
rect 4536 4612 4552 4628
rect 4584 4612 4600 4628
rect 4760 4772 4776 4788
rect 4808 4712 4824 4728
rect 4744 4652 4760 4668
rect 4680 4572 4696 4588
rect 4440 4532 4456 4548
rect 4568 4532 4584 4548
rect 4408 4512 4424 4528
rect 4616 4512 4632 4528
rect 4664 4512 4680 4528
rect 4408 4492 4424 4508
rect 4488 4492 4504 4508
rect 4632 4492 4648 4508
rect 4776 4612 4792 4628
rect 4760 4572 4776 4588
rect 4776 4512 4808 4528
rect 4376 4372 4392 4388
rect 4344 4352 4360 4368
rect 4328 4172 4344 4188
rect 4616 4472 4632 4488
rect 4440 4352 4456 4368
rect 4424 4312 4440 4328
rect 4504 4312 4520 4328
rect 4408 4292 4424 4308
rect 4424 4272 4440 4288
rect 4584 4372 4600 4388
rect 4536 4352 4552 4368
rect 4552 4232 4568 4248
rect 4520 4212 4536 4228
rect 4344 4132 4360 4148
rect 4392 4132 4408 4148
rect 4456 4132 4472 4148
rect 4616 4132 4632 4148
rect 4536 4112 4552 4128
rect 4552 4112 4568 4128
rect 4584 4112 4600 4128
rect 4424 4092 4440 4108
rect 4408 4072 4424 4088
rect 4344 3952 4360 3968
rect 4296 3932 4328 3948
rect 4280 3912 4296 3928
rect 4344 3892 4360 3908
rect 4216 3852 4232 3868
rect 4264 3852 4280 3868
rect 4205 3802 4241 3818
rect 4328 3812 4344 3828
rect 4440 4032 4456 4048
rect 4472 4012 4488 4028
rect 4440 3952 4456 3968
rect 4392 3932 4408 3948
rect 4424 3932 4440 3948
rect 4424 3912 4440 3928
rect 4440 3892 4456 3908
rect 4264 3772 4280 3788
rect 4376 3772 4392 3788
rect 3912 3732 3928 3748
rect 4024 3732 4040 3748
rect 4088 3732 4104 3748
rect 4152 3732 4168 3748
rect 3896 3712 3912 3728
rect 3944 3712 3960 3728
rect 3864 3692 3880 3708
rect 3928 3672 3944 3688
rect 3864 3652 3880 3668
rect 3832 3612 3848 3628
rect 3832 3592 3848 3608
rect 3816 3572 3832 3588
rect 3832 3532 3848 3548
rect 3848 3532 3864 3548
rect 3816 3512 3832 3528
rect 3816 3432 3832 3448
rect 3384 3352 3400 3368
rect 3480 3352 3496 3368
rect 3672 3352 3688 3368
rect 3704 3332 3720 3348
rect 3448 3312 3464 3328
rect 2984 3292 3000 3308
rect 3016 3292 3032 3308
rect 3128 3292 3144 3308
rect 3240 3292 3256 3308
rect 3400 3292 3432 3308
rect 3000 3192 3016 3208
rect 3096 3252 3112 3268
rect 3165 3202 3201 3218
rect 3208 3192 3224 3208
rect 3256 3192 3272 3208
rect 3368 3132 3384 3148
rect 3080 3112 3112 3128
rect 3176 3112 3192 3128
rect 3208 3112 3224 3128
rect 3288 3112 3304 3128
rect 3352 3112 3368 3128
rect 3048 3092 3064 3108
rect 3064 3092 3080 3108
rect 2968 3052 2984 3068
rect 2920 3012 2936 3028
rect 3096 3052 3112 3068
rect 3144 3052 3160 3068
rect 3176 3052 3192 3068
rect 3064 2992 3080 3008
rect 3128 2992 3144 3008
rect 2616 2932 2632 2948
rect 2712 2932 2728 2948
rect 2760 2932 2776 2948
rect 2888 2932 2904 2948
rect 2920 2932 2936 2948
rect 3016 2932 3032 2948
rect 2472 2912 2488 2928
rect 2520 2892 2536 2908
rect 2360 2792 2376 2808
rect 2136 2692 2152 2708
rect 2232 2632 2248 2648
rect 2136 2612 2152 2628
rect 2157 2602 2193 2618
rect 2168 2572 2184 2588
rect 2120 2552 2136 2568
rect 2152 2552 2168 2568
rect 2120 2532 2136 2548
rect 2216 2532 2232 2548
rect 2520 2772 2536 2788
rect 2504 2752 2520 2768
rect 2552 2752 2568 2768
rect 2472 2732 2488 2748
rect 2376 2692 2392 2708
rect 2344 2672 2360 2688
rect 2296 2652 2312 2668
rect 2264 2592 2280 2608
rect 2328 2572 2344 2588
rect 2504 2672 2520 2688
rect 2568 2652 2584 2668
rect 2408 2612 2424 2628
rect 2312 2532 2328 2548
rect 2376 2532 2392 2548
rect 2392 2532 2408 2548
rect 2440 2532 2456 2548
rect 2488 2532 2504 2548
rect 2600 2572 2616 2588
rect 2824 2912 2840 2928
rect 3144 2932 3160 2948
rect 2664 2752 2680 2768
rect 2728 2752 2744 2768
rect 2632 2692 2648 2708
rect 2648 2632 2664 2648
rect 2648 2532 2664 2548
rect 2584 2512 2600 2528
rect 1912 2492 1928 2508
rect 2008 2492 2024 2508
rect 2280 2492 2296 2508
rect 1816 2432 1832 2448
rect 1880 2352 1896 2368
rect 1816 2306 1832 2308
rect 1816 2292 1832 2306
rect 1880 2292 1896 2308
rect 1784 2212 1800 2228
rect 1784 2152 1800 2168
rect 2360 2472 2376 2488
rect 2408 2472 2424 2488
rect 2344 2452 2360 2468
rect 2632 2492 2648 2508
rect 2584 2412 2600 2428
rect 1976 2332 1992 2348
rect 2024 2332 2040 2348
rect 2232 2332 2248 2348
rect 2376 2332 2392 2348
rect 2280 2312 2296 2328
rect 2344 2312 2360 2328
rect 2120 2292 2136 2308
rect 2296 2292 2312 2308
rect 2456 2292 2472 2308
rect 2712 2572 2728 2588
rect 2840 2852 2856 2868
rect 2776 2752 2792 2768
rect 2856 2752 2872 2768
rect 2856 2692 2872 2708
rect 2792 2612 2808 2628
rect 2776 2552 2792 2568
rect 2712 2532 2728 2548
rect 2760 2532 2776 2548
rect 2840 2652 2856 2668
rect 2904 2652 2920 2668
rect 2904 2632 2920 2648
rect 2808 2592 2824 2608
rect 2904 2592 2920 2608
rect 3224 3052 3256 3068
rect 3368 3092 3384 3108
rect 3384 3072 3400 3088
rect 3304 3052 3336 3068
rect 3432 3272 3448 3288
rect 3416 3112 3432 3128
rect 3528 3112 3544 3128
rect 3560 3272 3576 3288
rect 3736 3292 3752 3308
rect 3704 3272 3720 3288
rect 3752 3272 3768 3288
rect 3688 3152 3704 3168
rect 3784 3352 3800 3368
rect 3800 3272 3816 3288
rect 3848 3392 3864 3408
rect 3832 3292 3848 3308
rect 3784 3132 3800 3148
rect 3752 3112 3768 3128
rect 3752 3092 3768 3108
rect 3816 3192 3832 3208
rect 3896 3612 3912 3628
rect 3896 3572 3912 3588
rect 3992 3692 4008 3708
rect 4072 3672 4088 3688
rect 4072 3632 4088 3648
rect 4056 3592 4072 3608
rect 3944 3572 3960 3588
rect 3928 3552 3944 3568
rect 3896 3532 3912 3548
rect 3880 3512 3896 3528
rect 4056 3552 4072 3568
rect 3976 3532 3992 3548
rect 3992 3532 4008 3548
rect 4024 3532 4040 3548
rect 3896 3432 3912 3448
rect 4040 3512 4056 3528
rect 4088 3512 4104 3528
rect 3992 3492 4008 3508
rect 3944 3452 3960 3468
rect 3928 3432 3944 3448
rect 3912 3392 3928 3408
rect 3880 3372 3896 3388
rect 3912 3292 3928 3308
rect 3864 3252 3880 3268
rect 3800 3092 3816 3108
rect 3960 3392 3976 3408
rect 3976 3332 3992 3348
rect 3960 3292 3976 3308
rect 3928 3192 3944 3208
rect 4024 3352 4040 3368
rect 4040 3332 4056 3348
rect 3976 3272 3992 3288
rect 4072 3452 4088 3468
rect 4104 3432 4120 3448
rect 4152 3712 4168 3728
rect 4168 3712 4184 3728
rect 4248 3692 4264 3708
rect 4152 3672 4168 3688
rect 4280 3752 4296 3768
rect 4344 3752 4360 3768
rect 4408 3832 4424 3848
rect 4328 3712 4344 3728
rect 4280 3672 4296 3688
rect 4296 3632 4312 3648
rect 4344 3632 4360 3648
rect 4328 3612 4344 3628
rect 4136 3572 4152 3588
rect 4200 3572 4216 3588
rect 4296 3572 4312 3588
rect 4136 3552 4152 3568
rect 4168 3532 4184 3548
rect 4264 3532 4280 3548
rect 4312 3532 4328 3548
rect 4168 3512 4184 3528
rect 4152 3492 4168 3508
rect 4120 3352 4136 3368
rect 4072 3332 4088 3348
rect 4248 3492 4264 3508
rect 4168 3432 4184 3448
rect 4152 3412 4168 3428
rect 4376 3672 4392 3688
rect 4360 3592 4376 3608
rect 4424 3712 4440 3728
rect 4456 3692 4472 3708
rect 4488 3992 4504 4008
rect 4520 3992 4536 4008
rect 4552 4092 4568 4108
rect 4600 4092 4616 4108
rect 4536 3972 4552 3988
rect 4520 3952 4536 3968
rect 4520 3912 4536 3928
rect 4712 4452 4728 4468
rect 4744 4352 4760 4368
rect 4680 4332 4696 4348
rect 4712 4272 4728 4288
rect 4680 4172 4696 4188
rect 4664 4032 4680 4048
rect 4600 3912 4616 3928
rect 4552 3872 4568 3888
rect 4600 3872 4616 3888
rect 4632 3872 4648 3888
rect 4488 3852 4504 3868
rect 4536 3852 4552 3868
rect 4648 3852 4664 3868
rect 4568 3832 4584 3848
rect 4584 3812 4600 3828
rect 4584 3752 4600 3768
rect 4504 3692 4536 3708
rect 4360 3552 4376 3568
rect 4472 3552 4488 3568
rect 4280 3512 4296 3528
rect 4264 3432 4280 3448
rect 4205 3402 4241 3418
rect 4248 3412 4264 3428
rect 4328 3472 4344 3488
rect 4376 3472 4392 3488
rect 4392 3412 4408 3428
rect 4248 3372 4264 3388
rect 4360 3372 4376 3388
rect 4264 3352 4280 3368
rect 4360 3332 4376 3348
rect 4184 3312 4200 3328
rect 4312 3312 4328 3328
rect 4056 3292 4072 3308
rect 4056 3272 4072 3288
rect 3912 3152 3928 3168
rect 3960 3152 3976 3168
rect 3896 3112 3912 3128
rect 3928 3132 3944 3148
rect 3976 3132 3992 3148
rect 3976 3092 3992 3108
rect 3432 3072 3448 3088
rect 3464 3072 3480 3088
rect 3656 3072 3672 3088
rect 3784 3072 3800 3088
rect 3928 3072 3944 3088
rect 3400 3052 3416 3068
rect 3320 3032 3336 3048
rect 3368 3032 3384 3048
rect 3256 2972 3272 2988
rect 3256 2952 3272 2968
rect 3512 2952 3528 2968
rect 3704 3052 3720 3068
rect 3544 3032 3560 3048
rect 3656 3012 3672 3028
rect 3592 2952 3608 2968
rect 3352 2932 3368 2948
rect 3528 2932 3544 2948
rect 3608 2932 3624 2948
rect 3208 2912 3224 2928
rect 3304 2912 3320 2928
rect 3320 2912 3336 2928
rect 3608 2912 3624 2928
rect 3640 2912 3656 2928
rect 3304 2892 3320 2908
rect 3384 2892 3400 2908
rect 3576 2892 3592 2908
rect 3048 2752 3064 2768
rect 2984 2732 3000 2748
rect 3000 2692 3016 2708
rect 3080 2692 3096 2708
rect 2984 2672 3000 2688
rect 3032 2672 3048 2688
rect 2952 2652 2968 2668
rect 2936 2632 2952 2648
rect 3032 2572 3048 2588
rect 3496 2832 3512 2848
rect 3165 2802 3201 2818
rect 3592 2852 3608 2868
rect 3336 2772 3352 2788
rect 3208 2732 3224 2748
rect 3320 2672 3336 2688
rect 3112 2632 3128 2648
rect 3048 2552 3064 2568
rect 3304 2652 3320 2668
rect 3144 2592 3160 2608
rect 3144 2572 3160 2588
rect 3288 2552 3304 2568
rect 2680 2492 2696 2508
rect 2824 2492 2840 2508
rect 2776 2472 2792 2488
rect 2744 2432 2760 2448
rect 2616 2312 2632 2328
rect 2664 2312 2680 2328
rect 2616 2292 2632 2308
rect 2136 2272 2152 2288
rect 2440 2272 2456 2288
rect 1928 2252 1944 2268
rect 1896 2212 1912 2228
rect 2040 2252 2056 2268
rect 2056 2232 2072 2248
rect 1848 2192 1864 2208
rect 1944 2192 1976 2208
rect 1992 2192 2008 2208
rect 1816 2132 1832 2148
rect 1752 2092 1768 2108
rect 1752 2072 1768 2088
rect 1656 1892 1672 1908
rect 1784 1932 1800 1948
rect 1720 1872 1736 1888
rect 1704 1852 1720 1868
rect 1688 1812 1704 1828
rect 1704 1792 1720 1808
rect 1640 1732 1656 1748
rect 1624 1512 1640 1528
rect 1608 1492 1624 1508
rect 2120 2212 2136 2228
rect 2056 2172 2072 2188
rect 2008 2132 2024 2148
rect 1848 2032 1864 2048
rect 1848 1892 1864 1908
rect 1768 1872 1784 1888
rect 1832 1872 1848 1888
rect 1784 1852 1800 1868
rect 1816 1832 1832 1848
rect 1768 1792 1784 1808
rect 2280 2252 2296 2268
rect 2248 2232 2264 2248
rect 2157 2202 2193 2218
rect 2184 2152 2200 2168
rect 2136 2132 2152 2148
rect 2072 2112 2088 2128
rect 2168 2112 2184 2128
rect 2104 2092 2120 2108
rect 2200 2092 2216 2108
rect 1896 1872 1912 1888
rect 1896 1852 1912 1868
rect 2024 1852 2040 1868
rect 1880 1832 1896 1848
rect 1928 1792 1944 1808
rect 1848 1752 1864 1768
rect 1880 1752 1912 1768
rect 2008 1752 2024 1768
rect 1672 1692 1688 1708
rect 1720 1692 1752 1708
rect 1640 1432 1656 1448
rect 1592 1372 1608 1388
rect 1576 1332 1592 1348
rect 1528 1312 1544 1328
rect 1480 1292 1492 1308
rect 1492 1292 1496 1308
rect 1496 1172 1512 1188
rect 1352 1152 1368 1168
rect 1304 1132 1320 1148
rect 1336 1132 1352 1148
rect 1432 1132 1448 1148
rect 1384 1112 1400 1128
rect 1448 1112 1464 1128
rect 1416 1092 1432 1108
rect 1400 1052 1416 1068
rect 1256 992 1272 1008
rect 1240 952 1256 968
rect 1240 932 1256 948
rect 1304 932 1320 948
rect 1304 912 1320 928
rect 1352 932 1368 948
rect 1368 912 1384 928
rect 1224 892 1240 908
rect 1320 892 1332 908
rect 1332 892 1336 908
rect 1400 972 1416 988
rect 1448 1072 1464 1088
rect 1448 952 1464 968
rect 1416 932 1432 948
rect 1416 912 1432 928
rect 1176 872 1192 888
rect 1117 802 1153 818
rect 1112 772 1128 788
rect 1128 732 1144 748
rect 1032 692 1048 708
rect 1064 692 1080 708
rect 1080 672 1096 688
rect 984 652 1000 668
rect 1160 632 1176 648
rect 936 492 952 508
rect 1000 512 1016 528
rect 1096 512 1112 528
rect 1016 492 1032 508
rect 1080 492 1096 508
rect 968 472 984 488
rect 760 292 776 308
rect 824 292 840 308
rect 1032 352 1048 368
rect 1016 332 1032 348
rect 888 312 904 328
rect 1117 402 1153 418
rect 1192 832 1208 848
rect 1352 832 1368 848
rect 1192 792 1208 808
rect 1384 792 1400 808
rect 1208 672 1224 688
rect 1272 692 1288 708
rect 1256 632 1272 648
rect 1480 1012 1496 1028
rect 1496 912 1512 928
rect 1416 772 1432 788
rect 1400 752 1416 768
rect 1464 752 1480 768
rect 1496 752 1512 768
rect 1592 1192 1608 1208
rect 1592 1172 1608 1188
rect 1576 1152 1592 1168
rect 1528 1132 1544 1148
rect 1784 1672 1800 1688
rect 1848 1672 1864 1688
rect 1832 1612 1848 1628
rect 1752 1492 1768 1508
rect 1752 1452 1768 1468
rect 1832 1392 1848 1408
rect 1800 1372 1816 1388
rect 1816 1352 1832 1368
rect 1848 1352 1864 1368
rect 1976 1732 1992 1748
rect 1912 1692 1928 1708
rect 1896 1352 1912 1368
rect 1928 1492 1944 1508
rect 1992 1712 2008 1728
rect 2040 1712 2056 1728
rect 2072 1672 2088 1688
rect 2088 1652 2104 1668
rect 2152 1952 2168 1968
rect 2120 1832 2136 1848
rect 2157 1802 2193 1818
rect 2136 1752 2152 1768
rect 2104 1612 2120 1628
rect 2056 1532 2072 1548
rect 2120 1492 2136 1508
rect 1944 1452 1960 1468
rect 1992 1452 2008 1468
rect 2024 1372 2040 1388
rect 1944 1352 1960 1368
rect 1992 1352 2008 1368
rect 1784 1312 1800 1328
rect 1880 1312 1896 1328
rect 1704 1292 1720 1308
rect 1752 1292 1768 1308
rect 1832 1292 1848 1308
rect 1880 1292 1896 1308
rect 1624 1152 1640 1168
rect 1672 1152 1688 1168
rect 1880 1272 1896 1288
rect 1544 1072 1560 1088
rect 1576 1072 1592 1088
rect 1672 1072 1688 1088
rect 1784 1072 1800 1088
rect 1832 1072 1848 1088
rect 1608 1032 1624 1048
rect 1704 1032 1720 1048
rect 1544 972 1560 988
rect 1592 952 1608 968
rect 1608 912 1624 928
rect 1576 892 1592 908
rect 1608 892 1624 908
rect 1640 892 1656 908
rect 1784 932 1816 948
rect 1672 912 1704 928
rect 1672 872 1688 888
rect 1576 852 1592 868
rect 1656 852 1672 868
rect 1896 1032 1912 1048
rect 1960 1292 1976 1308
rect 1976 1272 1992 1288
rect 2008 1112 2024 1128
rect 2168 1612 2184 1628
rect 2264 1992 2280 2008
rect 2216 1912 2232 1928
rect 2232 1852 2248 1868
rect 2616 2232 2632 2248
rect 2536 2172 2552 2188
rect 2296 2132 2312 2148
rect 2456 2132 2472 2148
rect 2328 2112 2344 2128
rect 2296 2092 2312 2108
rect 2328 2012 2344 2028
rect 2504 2012 2520 2028
rect 2504 1952 2520 1968
rect 2488 1892 2504 1908
rect 2360 1852 2376 1868
rect 2312 1832 2328 1848
rect 2264 1792 2280 1808
rect 2248 1732 2264 1748
rect 2344 1732 2360 1748
rect 2232 1552 2248 1568
rect 2232 1532 2248 1548
rect 2152 1492 2168 1508
rect 2200 1492 2216 1508
rect 2232 1492 2248 1508
rect 2264 1712 2280 1728
rect 2392 1812 2408 1828
rect 2440 1872 2456 1888
rect 2456 1872 2472 1888
rect 2424 1812 2440 1828
rect 2456 1832 2472 1848
rect 2568 1912 2584 1928
rect 2536 1892 2552 1908
rect 2472 1812 2504 1828
rect 2440 1772 2456 1788
rect 2472 1752 2504 1768
rect 2456 1732 2472 1748
rect 2504 1732 2520 1748
rect 2536 1732 2552 1748
rect 2568 1872 2584 1888
rect 2600 1792 2616 1808
rect 2680 2212 2696 2228
rect 3064 2532 3080 2548
rect 3112 2532 3128 2548
rect 3224 2532 3240 2548
rect 3272 2532 3288 2548
rect 2920 2492 2936 2508
rect 2904 2472 2920 2488
rect 2824 2392 2840 2408
rect 2872 2312 2888 2328
rect 2760 2292 2776 2308
rect 2792 2232 2808 2248
rect 2792 2172 2808 2188
rect 2728 2132 2744 2148
rect 2648 2112 2664 2128
rect 2776 2152 2792 2168
rect 2744 2112 2760 2128
rect 2776 2112 2792 2128
rect 2696 2092 2712 2108
rect 2664 1972 2680 1988
rect 2744 1912 2760 1928
rect 2632 1892 2648 1908
rect 2552 1692 2568 1708
rect 2424 1652 2440 1668
rect 2600 1692 2616 1708
rect 2472 1632 2488 1648
rect 2536 1632 2552 1648
rect 2584 1632 2600 1648
rect 2264 1512 2280 1528
rect 2248 1452 2264 1468
rect 2157 1402 2193 1418
rect 2376 1612 2392 1628
rect 2520 1612 2536 1628
rect 2296 1492 2312 1508
rect 2344 1492 2360 1508
rect 2392 1492 2408 1508
rect 2440 1472 2456 1488
rect 2328 1432 2344 1448
rect 2248 1352 2264 1368
rect 2104 1312 2120 1328
rect 2296 1312 2312 1328
rect 2376 1312 2392 1328
rect 2472 1312 2488 1328
rect 2056 1152 2072 1168
rect 2072 1112 2088 1128
rect 2120 1132 2136 1148
rect 2072 1092 2088 1108
rect 2104 1092 2120 1108
rect 1928 1072 1944 1088
rect 1960 1072 1976 1088
rect 2056 1072 2072 1088
rect 1976 1052 1992 1068
rect 1960 972 1976 988
rect 1992 972 2008 988
rect 2024 972 2040 988
rect 2008 952 2024 968
rect 1896 912 1912 928
rect 1944 872 1960 888
rect 1848 852 1864 868
rect 1992 852 2008 868
rect 1704 812 1720 828
rect 1928 792 1944 808
rect 2024 792 2040 808
rect 1512 712 1528 728
rect 1288 672 1304 688
rect 1320 672 1336 688
rect 1368 672 1384 688
rect 1304 532 1320 548
rect 1240 512 1256 528
rect 1496 672 1512 688
rect 1512 552 1528 568
rect 1512 532 1528 548
rect 1336 492 1352 508
rect 1432 472 1448 488
rect 1128 352 1144 368
rect 1272 352 1288 368
rect 1384 332 1400 348
rect 1272 312 1288 328
rect 952 292 968 308
rect 1080 292 1096 308
rect 1256 292 1272 308
rect 1352 292 1368 308
rect 1016 272 1032 288
rect 1144 272 1160 288
rect 456 172 472 188
rect 648 172 664 188
rect 744 152 760 168
rect 824 152 840 168
rect 936 172 952 188
rect 1016 172 1032 188
rect 952 152 968 168
rect 1096 172 1112 188
rect 1192 172 1208 188
rect 616 132 632 148
rect 776 132 792 148
rect 824 132 840 148
rect 984 132 1000 148
rect 1080 132 1096 148
rect 1192 132 1208 148
rect 1224 132 1240 148
rect 392 112 408 128
rect 584 114 600 128
rect 584 112 600 114
rect 680 112 696 128
rect 968 112 984 128
rect 1048 112 1064 128
rect 1336 152 1352 168
rect 1288 132 1304 148
rect 1400 272 1416 288
rect 1480 332 1496 348
rect 1608 732 1624 748
rect 1800 732 1816 748
rect 1832 732 1848 748
rect 1976 732 1992 748
rect 1576 712 1592 728
rect 1576 692 1592 708
rect 1672 706 1688 708
rect 1672 692 1688 706
rect 1960 692 1976 708
rect 1624 632 1640 648
rect 1640 552 1656 568
rect 1784 592 1800 608
rect 1752 572 1768 588
rect 1768 532 1784 548
rect 1800 552 1816 568
rect 1688 512 1704 528
rect 1656 392 1672 408
rect 1560 372 1576 388
rect 1560 312 1576 328
rect 1480 292 1496 308
rect 1528 292 1544 308
rect 1464 172 1480 188
rect 1400 132 1416 148
rect 1864 592 1880 608
rect 1832 572 1848 588
rect 1992 612 2008 628
rect 1880 572 1896 588
rect 1944 552 1960 568
rect 1976 512 1992 528
rect 1832 452 1848 468
rect 1816 392 1832 408
rect 1736 292 1752 308
rect 1688 272 1704 288
rect 1848 332 1864 348
rect 1960 332 1976 348
rect 1864 312 1880 328
rect 1928 312 1944 328
rect 1880 292 1896 308
rect 1960 292 1976 308
rect 1832 172 1848 188
rect 1480 132 1496 148
rect 1800 132 1816 148
rect 2008 592 2024 608
rect 2088 1052 2104 1068
rect 2056 832 2072 848
rect 2072 812 2088 828
rect 2120 912 2136 928
rect 2104 892 2120 908
rect 2152 1292 2168 1308
rect 2312 1212 2328 1228
rect 2216 1192 2232 1208
rect 2200 1152 2216 1168
rect 2200 1132 2216 1148
rect 2248 1152 2264 1168
rect 2200 1072 2216 1088
rect 2216 1052 2232 1068
rect 2157 1002 2193 1018
rect 2152 972 2168 988
rect 2168 972 2184 988
rect 2168 932 2184 948
rect 2232 852 2248 868
rect 2232 812 2248 828
rect 2136 792 2152 808
rect 2216 752 2232 768
rect 2264 1132 2280 1148
rect 2264 1112 2280 1128
rect 2296 1112 2312 1128
rect 2296 1012 2312 1028
rect 2280 952 2296 968
rect 2280 932 2296 948
rect 2296 932 2312 948
rect 2296 912 2312 928
rect 2264 812 2280 828
rect 2072 652 2088 668
rect 2120 652 2136 668
rect 2040 632 2056 648
rect 2056 572 2072 588
rect 2072 552 2088 568
rect 2072 532 2088 548
rect 2157 602 2193 618
rect 2168 572 2184 588
rect 2136 552 2152 568
rect 2120 532 2136 548
rect 2504 1352 2520 1368
rect 2536 1552 2552 1568
rect 2536 1452 2552 1468
rect 2568 1452 2584 1468
rect 2536 1432 2552 1448
rect 2520 1312 2536 1328
rect 2488 1172 2504 1188
rect 2568 1372 2584 1388
rect 2584 1152 2600 1168
rect 2328 1092 2344 1108
rect 2440 1092 2472 1108
rect 2344 1052 2360 1068
rect 2344 992 2360 1008
rect 2328 972 2344 988
rect 2408 1052 2440 1068
rect 2392 952 2408 968
rect 2408 932 2424 948
rect 2456 1072 2472 1088
rect 2488 1052 2504 1068
rect 2456 972 2472 988
rect 2504 932 2520 948
rect 2360 912 2376 928
rect 2376 912 2392 928
rect 2424 912 2440 928
rect 2440 892 2456 908
rect 2376 832 2392 848
rect 2312 712 2328 728
rect 2360 712 2376 728
rect 2408 692 2424 708
rect 2296 552 2312 568
rect 2296 532 2312 548
rect 2232 512 2248 528
rect 2152 492 2168 508
rect 2120 392 2136 408
rect 2056 292 2072 308
rect 2248 292 2264 308
rect 2280 272 2296 288
rect 2157 202 2193 218
rect 2216 172 2232 188
rect 2296 172 2312 188
rect 1848 132 1864 148
rect 1864 132 1880 148
rect 1896 132 1912 148
rect 2120 132 2136 148
rect 1496 112 1512 128
rect 1544 112 1560 128
rect 1704 112 1720 128
rect 1880 112 1896 128
rect 1960 114 1976 128
rect 1960 112 1976 114
rect 2264 112 2280 128
rect 2360 672 2376 688
rect 2344 652 2360 668
rect 2472 752 2504 768
rect 2472 692 2488 708
rect 2424 572 2440 588
rect 2344 512 2360 528
rect 2456 512 2472 528
rect 2584 1012 2600 1028
rect 2568 972 2584 988
rect 2584 872 2600 888
rect 2536 852 2552 868
rect 2744 1872 2760 1888
rect 2712 1852 2728 1868
rect 2728 1832 2744 1848
rect 2712 1792 2728 1808
rect 2728 1752 2744 1768
rect 2840 2132 2856 2148
rect 2920 2392 2936 2408
rect 2968 2392 2984 2408
rect 2920 2292 2936 2308
rect 2968 2292 2984 2308
rect 2984 2252 3000 2268
rect 3000 2212 3016 2228
rect 3064 2492 3080 2508
rect 3256 2492 3272 2508
rect 3165 2402 3201 2418
rect 3272 2472 3288 2488
rect 3224 2332 3240 2348
rect 3064 2292 3080 2308
rect 3064 2272 3080 2288
rect 3128 2252 3144 2268
rect 3080 2212 3096 2228
rect 2920 2152 2936 2168
rect 3048 2152 3064 2168
rect 2808 2092 2824 2108
rect 2824 1992 2840 2008
rect 2840 1892 2856 1908
rect 2776 1872 2792 1888
rect 2760 1852 2776 1868
rect 2824 1852 2840 1868
rect 2680 1692 2696 1708
rect 2696 1692 2712 1708
rect 2792 1792 2824 1808
rect 2776 1732 2792 1748
rect 2744 1612 2760 1628
rect 2760 1532 2776 1548
rect 2696 1512 2712 1528
rect 2776 1512 2792 1528
rect 2776 1492 2792 1508
rect 2648 1432 2664 1448
rect 2696 1432 2712 1448
rect 2856 1872 2872 1888
rect 3032 2132 3048 2148
rect 3016 2092 3032 2108
rect 2952 2072 2968 2088
rect 3048 2052 3064 2068
rect 3048 2032 3064 2048
rect 3016 2012 3032 2028
rect 2952 1992 2968 2008
rect 2952 1952 2968 1968
rect 3144 2112 3160 2128
rect 3256 2272 3272 2288
rect 3320 2532 3336 2548
rect 3384 2732 3400 2748
rect 3352 2692 3368 2708
rect 3400 2692 3416 2708
rect 3448 2692 3464 2708
rect 3528 2692 3544 2708
rect 3432 2672 3448 2688
rect 3496 2672 3528 2688
rect 3416 2652 3432 2668
rect 3416 2632 3432 2648
rect 3464 2572 3480 2588
rect 3560 2612 3576 2628
rect 3512 2552 3528 2568
rect 3432 2532 3448 2548
rect 3320 2492 3336 2508
rect 3368 2292 3384 2308
rect 3416 2292 3432 2308
rect 3448 2512 3464 2528
rect 3464 2512 3480 2528
rect 3496 2512 3512 2528
rect 3544 2512 3560 2528
rect 3480 2312 3496 2328
rect 3544 2472 3560 2488
rect 3672 2952 3688 2968
rect 4024 3032 4040 3048
rect 4056 3032 4072 3048
rect 3864 2992 3880 3008
rect 3704 2972 3720 2988
rect 3832 2972 3848 2988
rect 3704 2952 3720 2968
rect 3720 2912 3736 2928
rect 4120 3272 4136 3288
rect 4136 3212 4152 3228
rect 4088 2972 4104 2988
rect 3880 2952 3896 2968
rect 3880 2932 3896 2948
rect 3944 2912 3960 2928
rect 3944 2892 3960 2908
rect 4040 2914 4056 2928
rect 4040 2912 4056 2914
rect 3880 2872 3896 2888
rect 3976 2872 3992 2888
rect 3752 2852 3768 2868
rect 3752 2772 3768 2788
rect 3640 2732 3656 2748
rect 3624 2692 3640 2708
rect 3672 2692 3688 2708
rect 3640 2672 3656 2688
rect 3672 2672 3688 2688
rect 3864 2672 3880 2688
rect 3624 2632 3640 2648
rect 3608 2512 3624 2528
rect 3592 2452 3608 2468
rect 3720 2632 3736 2648
rect 3752 2632 3768 2648
rect 3672 2552 3688 2568
rect 3784 2552 3800 2568
rect 3688 2532 3704 2548
rect 3704 2512 3720 2528
rect 3640 2472 3656 2488
rect 3624 2352 3640 2368
rect 3592 2312 3608 2328
rect 3464 2272 3480 2288
rect 3512 2272 3528 2288
rect 3224 2092 3240 2108
rect 3176 2052 3192 2068
rect 3165 2002 3201 2018
rect 3160 1972 3176 1988
rect 2984 1892 3000 1908
rect 2840 1792 2856 1808
rect 2872 1792 2888 1808
rect 2904 1732 2920 1748
rect 2904 1692 2920 1708
rect 2904 1612 2920 1628
rect 2824 1492 2840 1508
rect 2856 1452 2872 1468
rect 2824 1332 2840 1348
rect 2872 1332 2888 1348
rect 2696 1314 2712 1328
rect 2696 1312 2712 1314
rect 2808 1152 2824 1168
rect 2712 1092 2728 1108
rect 2696 1012 2712 1028
rect 2760 972 2776 988
rect 2536 772 2552 788
rect 2600 772 2632 788
rect 2552 692 2568 708
rect 2504 652 2520 668
rect 2488 612 2504 628
rect 2504 532 2520 548
rect 2552 612 2568 628
rect 2600 612 2616 628
rect 2472 492 2488 508
rect 2504 492 2520 508
rect 2600 552 2616 568
rect 2568 512 2584 528
rect 2696 914 2712 928
rect 2696 912 2712 914
rect 2792 912 2808 928
rect 2792 892 2808 908
rect 2744 772 2760 788
rect 2792 712 2808 728
rect 2664 672 2680 688
rect 2680 532 2696 548
rect 2648 512 2664 528
rect 2648 492 2664 508
rect 2584 472 2600 488
rect 2552 392 2568 408
rect 2344 332 2360 348
rect 2456 332 2472 348
rect 2360 312 2376 328
rect 2424 312 2440 328
rect 2376 292 2392 308
rect 2360 272 2376 288
rect 2632 312 2648 328
rect 2728 512 2744 528
rect 2792 612 2808 628
rect 2776 572 2792 588
rect 2856 1292 2872 1308
rect 2856 1252 2872 1268
rect 2840 1112 2856 1128
rect 3128 1872 3144 1888
rect 3048 1752 3064 1768
rect 3096 1732 3112 1748
rect 3080 1532 3096 1548
rect 2952 1512 2968 1528
rect 2984 1512 3000 1528
rect 3080 1512 3096 1528
rect 2952 1492 2968 1508
rect 2968 1472 2984 1488
rect 3016 1472 3032 1488
rect 3000 1452 3016 1468
rect 2952 1372 2968 1388
rect 3448 2232 3464 2248
rect 3432 2152 3448 2168
rect 3384 2132 3400 2148
rect 3272 2112 3288 2128
rect 3336 2112 3368 2128
rect 3592 2252 3608 2268
rect 3640 2172 3656 2188
rect 3512 2112 3528 2128
rect 3656 2112 3672 2128
rect 3304 2092 3320 2108
rect 3352 2092 3368 2108
rect 3496 2092 3512 2108
rect 3240 2012 3256 2028
rect 3608 2072 3624 2088
rect 3656 2072 3672 2088
rect 3304 1952 3320 1968
rect 3368 1952 3384 1968
rect 3416 1952 3432 1968
rect 3464 1952 3480 1968
rect 3288 1892 3304 1908
rect 3352 1892 3368 1908
rect 3320 1852 3336 1868
rect 3208 1812 3224 1828
rect 3240 1812 3256 1828
rect 3160 1712 3192 1728
rect 3240 1792 3256 1808
rect 3256 1752 3272 1768
rect 3240 1692 3256 1708
rect 3304 1692 3320 1708
rect 3165 1602 3201 1618
rect 3208 1612 3224 1628
rect 3336 1692 3352 1708
rect 3320 1552 3352 1568
rect 3144 1532 3160 1548
rect 3304 1532 3320 1548
rect 3464 1892 3480 1908
rect 3576 1892 3592 1908
rect 3400 1872 3416 1888
rect 3496 1872 3512 1888
rect 3528 1852 3544 1868
rect 3608 1812 3624 1828
rect 3432 1792 3448 1808
rect 3384 1752 3400 1768
rect 3416 1752 3432 1768
rect 3496 1752 3512 1768
rect 3752 2512 3768 2528
rect 4056 2852 4072 2868
rect 4104 2852 4120 2868
rect 4104 2772 4120 2788
rect 3976 2552 3992 2568
rect 3992 2532 4008 2548
rect 4088 2532 4104 2548
rect 4264 3192 4280 3208
rect 4168 3092 4184 3108
rect 4168 2872 4184 2888
rect 4205 3002 4241 3018
rect 4216 2952 4232 2968
rect 4232 2912 4248 2928
rect 4184 2852 4200 2868
rect 4184 2812 4200 2828
rect 4184 2732 4200 2748
rect 4360 3312 4376 3328
rect 4360 3272 4376 3288
rect 4344 3252 4360 3268
rect 4312 3132 4328 3148
rect 4280 3112 4296 3128
rect 4296 3092 4312 3108
rect 4280 2912 4296 2928
rect 4168 2692 4184 2708
rect 4216 2692 4232 2708
rect 4136 2632 4152 2648
rect 4120 2532 4136 2548
rect 4248 2672 4264 2688
rect 4248 2632 4264 2648
rect 4205 2602 4241 2618
rect 3880 2512 3896 2528
rect 3976 2512 3992 2528
rect 4168 2512 4184 2528
rect 3736 2492 3752 2508
rect 3848 2492 3864 2508
rect 4008 2492 4024 2508
rect 4056 2492 4072 2508
rect 3912 2472 3928 2488
rect 3896 2352 3912 2368
rect 3944 2352 3960 2368
rect 3704 2332 3720 2348
rect 3752 2332 3768 2348
rect 3816 2312 3832 2328
rect 3800 2292 3816 2308
rect 3848 2292 3864 2308
rect 3944 2292 3960 2308
rect 3720 2272 3736 2288
rect 3880 2252 3896 2268
rect 3752 2192 3768 2208
rect 3784 2192 3800 2208
rect 3752 2172 3768 2188
rect 3688 2152 3704 2168
rect 3752 2114 3768 2128
rect 3752 2112 3768 2114
rect 3880 2152 3896 2168
rect 3944 2152 3960 2168
rect 3976 2152 3992 2168
rect 3928 2112 3944 2128
rect 3992 2112 4008 2128
rect 3800 2052 3816 2068
rect 3944 2072 3960 2088
rect 3832 2012 3848 2028
rect 3928 2012 3944 2028
rect 3976 1952 3992 1968
rect 3928 1932 3944 1948
rect 3944 1912 3960 1928
rect 3944 1892 3960 1908
rect 3704 1872 3720 1888
rect 3784 1872 3800 1888
rect 3720 1852 3736 1868
rect 3752 1852 3768 1868
rect 3832 1852 3848 1868
rect 3688 1752 3704 1768
rect 3672 1732 3688 1748
rect 3528 1712 3544 1728
rect 3576 1712 3592 1728
rect 3384 1692 3400 1708
rect 3464 1692 3480 1708
rect 3528 1692 3544 1708
rect 3560 1692 3576 1708
rect 3592 1672 3608 1688
rect 3336 1512 3352 1528
rect 3368 1512 3384 1528
rect 3416 1512 3432 1528
rect 3272 1492 3288 1508
rect 3320 1492 3336 1508
rect 3208 1472 3224 1488
rect 3112 1452 3128 1468
rect 2984 1332 3000 1348
rect 3064 1332 3080 1348
rect 2952 1312 2968 1328
rect 2984 1292 3000 1308
rect 3032 1292 3048 1308
rect 2936 1272 2952 1288
rect 2920 1212 2936 1228
rect 2968 1212 2984 1228
rect 2872 1152 2888 1168
rect 2936 1152 2952 1168
rect 2952 1112 2968 1128
rect 2872 1092 2888 1108
rect 2952 1072 2968 1088
rect 2904 1052 2920 1068
rect 2872 1032 2888 1048
rect 2840 892 2856 908
rect 2824 732 2840 748
rect 2856 712 2872 728
rect 2856 692 2872 708
rect 2984 1052 3000 1068
rect 2984 1032 3000 1048
rect 3016 1012 3032 1028
rect 3000 992 3016 1008
rect 2952 932 2968 948
rect 2968 912 2984 928
rect 2936 872 2952 888
rect 2904 752 2920 768
rect 2888 672 2904 688
rect 2840 572 2856 588
rect 2968 672 2984 688
rect 3064 1112 3080 1128
rect 3032 952 3064 968
rect 3048 912 3064 928
rect 3064 892 3076 908
rect 3076 892 3080 908
rect 3048 872 3064 888
rect 2920 572 2936 588
rect 2904 532 2920 548
rect 2984 532 3000 548
rect 2808 512 2824 528
rect 2744 492 2760 508
rect 2920 492 2936 508
rect 2968 492 2984 508
rect 2760 472 2776 488
rect 2936 472 2952 488
rect 2968 472 2984 488
rect 2744 332 2760 348
rect 2584 272 2600 288
rect 2936 432 2952 448
rect 2936 352 2952 368
rect 2984 352 3000 368
rect 2872 332 2888 348
rect 2776 312 2792 328
rect 2904 312 2920 328
rect 2776 292 2792 308
rect 2824 292 2840 308
rect 3064 672 3080 688
rect 3128 1432 3144 1448
rect 3208 1412 3224 1428
rect 3256 1352 3272 1368
rect 3624 1692 3640 1708
rect 3656 1712 3672 1728
rect 3800 1832 3816 1848
rect 3912 1752 3928 1768
rect 4024 2472 4040 2488
rect 4136 2492 4152 2508
rect 4232 2492 4248 2508
rect 4104 2312 4120 2328
rect 4232 2312 4248 2328
rect 4104 2292 4120 2308
rect 4152 2272 4168 2288
rect 4056 2252 4072 2268
rect 4216 2252 4232 2268
rect 4168 2232 4184 2248
rect 4040 2132 4056 2148
rect 4136 2112 4152 2128
rect 4024 2072 4040 2088
rect 4104 2092 4120 2108
rect 4120 2092 4124 2108
rect 4124 2092 4136 2108
rect 4088 1992 4104 2008
rect 4088 1972 4120 1988
rect 4040 1952 4056 1968
rect 4008 1932 4024 1948
rect 4008 1892 4024 1908
rect 3976 1852 3992 1868
rect 4024 1852 4040 1868
rect 3912 1712 3928 1728
rect 3672 1692 3688 1708
rect 3752 1692 3768 1708
rect 3640 1552 3656 1568
rect 3768 1552 3784 1568
rect 3720 1532 3736 1548
rect 3416 1492 3432 1508
rect 3512 1506 3528 1508
rect 3512 1492 3528 1506
rect 3608 1492 3624 1508
rect 3576 1472 3592 1488
rect 3336 1432 3352 1448
rect 3448 1432 3464 1448
rect 3352 1412 3368 1428
rect 3592 1392 3608 1408
rect 3432 1372 3448 1388
rect 3480 1372 3496 1388
rect 3512 1372 3528 1388
rect 3368 1352 3384 1368
rect 3096 1312 3112 1328
rect 3144 1272 3160 1288
rect 3165 1202 3201 1218
rect 3224 1312 3240 1328
rect 3272 1312 3288 1328
rect 3256 1292 3272 1308
rect 3208 1152 3224 1168
rect 3672 1472 3688 1488
rect 3736 1452 3752 1468
rect 3640 1432 3656 1448
rect 3640 1392 3672 1408
rect 3640 1332 3656 1348
rect 3384 1312 3400 1328
rect 3304 1272 3320 1288
rect 3320 1152 3336 1168
rect 3272 1112 3288 1128
rect 3256 1092 3272 1108
rect 3304 1092 3320 1108
rect 3112 1072 3128 1088
rect 3096 912 3112 928
rect 3080 552 3096 568
rect 3032 392 3048 408
rect 3128 1012 3144 1028
rect 3192 1012 3208 1028
rect 3112 872 3128 888
rect 3160 972 3176 988
rect 3352 972 3368 988
rect 3368 952 3384 968
rect 3224 892 3240 908
rect 3165 802 3201 818
rect 3288 732 3304 748
rect 3176 692 3192 708
rect 3272 672 3288 688
rect 3512 1292 3528 1308
rect 3496 1272 3512 1288
rect 3560 1072 3576 1088
rect 3752 1312 3768 1328
rect 3864 1532 3880 1548
rect 4072 1932 4088 1948
rect 4136 1912 4152 1928
rect 4205 2202 4241 2218
rect 4184 2152 4200 2168
rect 4168 1872 4184 1888
rect 3976 1752 3992 1768
rect 4040 1772 4056 1788
rect 4008 1732 4024 1748
rect 3960 1572 3976 1588
rect 3848 1512 3864 1528
rect 3928 1512 3944 1528
rect 4008 1492 4024 1508
rect 3832 1472 3848 1488
rect 3896 1432 3912 1448
rect 3816 1352 3832 1368
rect 3944 1472 3960 1488
rect 3992 1432 4008 1448
rect 3944 1352 3960 1368
rect 3912 1332 3928 1348
rect 3880 1312 3896 1328
rect 3896 1312 3912 1328
rect 3960 1312 3976 1328
rect 3640 1272 3656 1288
rect 3704 1212 3720 1228
rect 3688 1192 3704 1208
rect 3768 1212 3784 1228
rect 3736 1152 3752 1168
rect 3640 1112 3656 1128
rect 3720 1112 3736 1128
rect 3592 1092 3608 1108
rect 3608 1072 3624 1088
rect 3640 1072 3656 1088
rect 3544 992 3560 1008
rect 3576 1032 3608 1048
rect 3544 972 3560 988
rect 3496 912 3512 928
rect 3672 1052 3688 1068
rect 3656 932 3672 948
rect 3384 892 3400 908
rect 3432 892 3448 908
rect 3464 892 3480 908
rect 3576 892 3592 908
rect 3416 732 3432 748
rect 3400 672 3416 688
rect 3368 652 3384 668
rect 3192 552 3208 568
rect 3224 532 3240 548
rect 3144 512 3160 528
rect 3256 512 3272 528
rect 3288 512 3304 528
rect 3096 352 3112 368
rect 2984 332 3000 348
rect 3016 332 3032 348
rect 2968 312 2984 328
rect 3080 312 3096 328
rect 3080 292 3096 308
rect 3096 292 3112 308
rect 2568 212 2584 228
rect 2680 212 2696 228
rect 2536 172 2552 188
rect 2696 192 2712 208
rect 2664 152 2680 168
rect 2680 152 2696 168
rect 2712 152 2728 168
rect 2904 212 2920 228
rect 3016 232 3032 248
rect 2920 192 2936 208
rect 3000 172 3016 188
rect 2760 132 2776 148
rect 2808 132 2824 148
rect 2888 132 2904 148
rect 3048 132 3064 148
rect 3144 392 3160 408
rect 3165 402 3201 418
rect 3224 392 3240 408
rect 3112 212 3128 228
rect 3128 192 3144 208
rect 3112 172 3128 188
rect 3304 372 3320 388
rect 3240 352 3256 368
rect 3288 352 3304 368
rect 3176 332 3192 348
rect 3512 872 3528 888
rect 3448 552 3464 568
rect 3432 532 3448 548
rect 3432 452 3448 468
rect 3336 412 3352 428
rect 3320 312 3336 328
rect 3240 292 3256 308
rect 3384 312 3400 328
rect 3384 292 3400 308
rect 3480 412 3496 428
rect 3416 332 3432 348
rect 3480 306 3496 308
rect 3480 292 3496 306
rect 3480 252 3496 268
rect 3400 232 3416 248
rect 3320 192 3336 208
rect 3400 192 3416 208
rect 3320 152 3336 168
rect 3256 132 3272 148
rect 3448 132 3480 148
rect 2408 112 2424 128
rect 2552 112 2568 128
rect 2744 112 2760 128
rect 3032 112 3048 128
rect 3080 112 3096 128
rect 3560 732 3576 748
rect 3528 712 3544 728
rect 3560 692 3576 708
rect 3608 692 3624 708
rect 3544 672 3560 688
rect 3544 652 3560 668
rect 3576 552 3592 568
rect 3528 512 3544 528
rect 3656 912 3672 928
rect 3640 892 3656 908
rect 3688 892 3704 908
rect 3672 872 3688 888
rect 3720 852 3736 868
rect 3704 772 3720 788
rect 3832 1292 3848 1308
rect 3800 1232 3816 1248
rect 3864 1272 3880 1288
rect 3832 1152 3848 1168
rect 3880 1152 3896 1168
rect 4024 1392 4040 1408
rect 4104 1772 4120 1788
rect 4136 1772 4152 1788
rect 4104 1732 4120 1748
rect 4232 2012 4248 2028
rect 4312 2972 4328 2988
rect 4360 3132 4376 3148
rect 4440 3492 4456 3508
rect 4424 3412 4440 3428
rect 4488 3512 4504 3528
rect 4472 3452 4488 3468
rect 4472 3292 4488 3308
rect 4456 3272 4472 3288
rect 4440 3232 4456 3248
rect 4504 3492 4520 3508
rect 4520 3472 4536 3488
rect 4504 3412 4520 3428
rect 4600 3712 4616 3728
rect 4632 3672 4648 3688
rect 4632 3612 4664 3628
rect 4680 3972 4696 3988
rect 4744 3932 4760 3948
rect 4712 3912 4728 3928
rect 4728 3892 4744 3908
rect 4680 3872 4696 3888
rect 4840 4672 4856 4688
rect 4824 4652 4840 4668
rect 4824 4532 4840 4548
rect 5032 4912 5048 4928
rect 4920 4892 4936 4908
rect 5032 4892 5048 4908
rect 5144 5272 5160 5288
rect 5192 5272 5208 5288
rect 5496 5292 5512 5308
rect 5112 5252 5128 5268
rect 5352 5252 5368 5268
rect 5213 5202 5249 5218
rect 5448 5212 5464 5228
rect 5608 5292 5624 5308
rect 5656 5292 5672 5308
rect 5576 5272 5592 5288
rect 5752 5252 5768 5268
rect 5608 5172 5624 5188
rect 5688 5172 5704 5188
rect 5576 5112 5608 5128
rect 5112 5092 5128 5108
rect 5224 5092 5240 5108
rect 5320 5092 5336 5108
rect 5192 5072 5208 5088
rect 5080 5032 5096 5048
rect 5080 5012 5096 5028
rect 5064 4872 5080 4888
rect 5080 4832 5096 4848
rect 5000 4712 5032 4728
rect 4888 4692 4904 4708
rect 4904 4672 4920 4688
rect 5000 4652 5016 4668
rect 4872 4572 4888 4588
rect 4936 4532 4952 4548
rect 4872 4512 4888 4528
rect 4920 4512 4936 4528
rect 4920 4492 4936 4508
rect 4808 4372 4824 4388
rect 4840 4352 4856 4368
rect 4840 4332 4856 4348
rect 4840 4312 4856 4328
rect 4872 4472 4888 4488
rect 4984 4452 5000 4468
rect 5048 4692 5064 4708
rect 5032 4552 5048 4568
rect 5048 4432 5064 4448
rect 5048 4352 5064 4368
rect 5032 4332 5048 4348
rect 4936 4312 4952 4328
rect 4968 4312 4984 4328
rect 4840 4292 4856 4308
rect 4856 4292 4872 4308
rect 4808 4272 4824 4288
rect 4792 4232 4808 4248
rect 4808 4114 4824 4128
rect 4808 4112 4824 4114
rect 4888 4272 4904 4288
rect 4968 4272 4984 4288
rect 5032 4272 5048 4288
rect 4872 4252 4888 4268
rect 4936 4252 4952 4268
rect 5000 4252 5016 4268
rect 4984 4212 5000 4228
rect 4872 4172 4904 4188
rect 4840 3952 4856 3968
rect 4952 4132 4968 4148
rect 4968 4132 4984 4148
rect 5016 4132 5032 4148
rect 4904 4112 4920 4128
rect 4904 4092 4920 4108
rect 5128 4752 5144 4768
rect 5480 5092 5496 5108
rect 5528 5092 5544 5108
rect 5576 5092 5592 5108
rect 5384 5072 5400 5088
rect 5480 5072 5496 5088
rect 5256 5032 5272 5048
rect 5208 4892 5224 4908
rect 5213 4802 5249 4818
rect 5448 5032 5464 5048
rect 5416 4972 5432 4988
rect 5480 4972 5496 4988
rect 5416 4952 5432 4968
rect 5352 4912 5368 4928
rect 5400 4912 5416 4928
rect 5320 4892 5336 4908
rect 5400 4892 5416 4908
rect 5480 4892 5496 4908
rect 5544 4852 5560 4868
rect 5528 4832 5544 4848
rect 5544 4772 5560 4788
rect 5592 4772 5608 4788
rect 5368 4752 5384 4768
rect 5400 4752 5416 4768
rect 5320 4732 5336 4748
rect 5208 4712 5224 4728
rect 5256 4712 5272 4728
rect 5352 4712 5368 4728
rect 5384 4712 5400 4728
rect 5304 4692 5320 4708
rect 5384 4692 5400 4708
rect 5176 4672 5192 4688
rect 5192 4652 5208 4668
rect 5288 4652 5304 4668
rect 5128 4612 5144 4628
rect 5160 4612 5176 4628
rect 5192 4552 5208 4568
rect 5208 4492 5224 4508
rect 5128 4472 5160 4488
rect 5208 4452 5224 4468
rect 5224 4452 5240 4468
rect 5213 4402 5249 4418
rect 5128 4372 5144 4388
rect 5080 4312 5096 4328
rect 5080 4292 5096 4308
rect 5160 4312 5176 4328
rect 5144 4212 5160 4228
rect 5160 4152 5176 4168
rect 5096 4132 5112 4148
rect 5064 4112 5080 4128
rect 4904 4072 4920 4088
rect 5016 4072 5032 4088
rect 5128 4052 5144 4068
rect 5000 4032 5016 4048
rect 5064 4032 5080 4048
rect 4920 3932 4936 3948
rect 4792 3912 4808 3928
rect 4824 3912 4840 3928
rect 4824 3892 4840 3908
rect 4856 3892 4872 3908
rect 4872 3872 4888 3888
rect 4840 3812 4856 3828
rect 4968 3812 4984 3828
rect 4872 3792 4888 3808
rect 4776 3772 4792 3788
rect 4776 3752 4792 3768
rect 4792 3752 4808 3768
rect 4712 3732 4728 3748
rect 4712 3712 4728 3728
rect 4696 3612 4712 3628
rect 4744 3612 4760 3628
rect 4664 3592 4680 3608
rect 4728 3532 4744 3548
rect 4584 3512 4600 3528
rect 4600 3512 4616 3528
rect 4536 3392 4552 3408
rect 4536 3312 4552 3328
rect 4520 3292 4536 3308
rect 4568 3472 4584 3488
rect 4568 3412 4584 3428
rect 4680 3512 4696 3528
rect 4968 3772 4984 3788
rect 5128 3952 5144 3968
rect 5032 3912 5048 3928
rect 4936 3672 4968 3688
rect 4824 3572 4840 3588
rect 4808 3492 4824 3508
rect 4648 3472 4664 3488
rect 4808 3472 4824 3488
rect 4744 3452 4760 3468
rect 4616 3392 4648 3408
rect 4680 3392 4696 3408
rect 4664 3372 4680 3388
rect 4600 3332 4616 3348
rect 4552 3192 4568 3208
rect 4424 3152 4440 3168
rect 4488 3152 4504 3168
rect 4440 3132 4456 3148
rect 4584 3192 4600 3208
rect 4504 3132 4520 3148
rect 4568 3132 4584 3148
rect 4552 3112 4568 3128
rect 4632 3232 4648 3248
rect 4600 3152 4616 3168
rect 4616 3132 4632 3148
rect 4424 3092 4440 3108
rect 4440 3092 4456 3108
rect 4376 3072 4392 3088
rect 4488 3072 4504 3088
rect 4600 3012 4616 3028
rect 4504 2972 4520 2988
rect 4568 2972 4584 2988
rect 4376 2914 4392 2928
rect 4376 2912 4392 2914
rect 4552 2912 4568 2928
rect 4520 2872 4536 2888
rect 4440 2852 4456 2868
rect 4568 2892 4584 2908
rect 4616 2912 4632 2928
rect 4600 2832 4616 2848
rect 4552 2812 4568 2828
rect 4488 2772 4504 2788
rect 4296 2752 4312 2768
rect 4376 2732 4392 2748
rect 4440 2732 4456 2748
rect 4328 2692 4344 2708
rect 4344 2692 4360 2708
rect 4392 2692 4408 2708
rect 4424 2692 4440 2708
rect 4296 2652 4312 2668
rect 4360 2572 4376 2588
rect 4408 2572 4424 2588
rect 4344 2532 4360 2548
rect 4344 2512 4360 2528
rect 4376 2532 4392 2548
rect 4280 2492 4296 2508
rect 4280 2472 4296 2488
rect 4328 2472 4344 2488
rect 4280 2312 4296 2328
rect 4280 2292 4296 2308
rect 4280 2212 4296 2228
rect 4344 2192 4360 2208
rect 4312 2152 4328 2168
rect 4328 2132 4344 2148
rect 4392 2132 4408 2148
rect 4584 2732 4600 2748
rect 4712 3332 4728 3348
rect 4712 3292 4728 3308
rect 4760 3252 4776 3268
rect 4856 3552 4872 3568
rect 4888 3532 4904 3548
rect 4856 3512 4872 3528
rect 4824 3372 4840 3388
rect 5016 3692 5032 3708
rect 5000 3652 5016 3668
rect 4984 3632 5000 3648
rect 4952 3532 4968 3548
rect 5000 3612 5032 3628
rect 5112 3612 5128 3628
rect 4904 3512 4920 3528
rect 4984 3512 5000 3528
rect 4936 3492 4952 3508
rect 5000 3492 5016 3508
rect 4888 3412 4904 3428
rect 5000 3372 5016 3388
rect 4840 3352 4856 3368
rect 4872 3352 4888 3368
rect 4888 3332 4904 3348
rect 4920 3332 4936 3348
rect 4792 3292 4808 3308
rect 4856 3292 4872 3308
rect 4888 3292 4904 3308
rect 4856 3272 4872 3288
rect 4872 3272 4888 3288
rect 4840 3252 4856 3268
rect 4824 3232 4840 3248
rect 4840 3152 4856 3168
rect 4696 3132 4712 3148
rect 4760 3132 4776 3148
rect 4824 3132 4840 3148
rect 4728 3112 4744 3128
rect 4648 3032 4664 3048
rect 4648 2892 4664 2908
rect 4680 3092 4696 3108
rect 4744 3092 4760 3108
rect 4744 3052 4760 3068
rect 4696 2952 4712 2968
rect 4728 2952 4744 2968
rect 4696 2932 4712 2948
rect 4696 2912 4712 2928
rect 4680 2872 4696 2888
rect 4664 2832 4680 2848
rect 4664 2752 4680 2768
rect 4536 2692 4552 2708
rect 4584 2692 4600 2708
rect 4504 2672 4520 2688
rect 4808 3012 4824 3028
rect 4808 2932 4824 2948
rect 4792 2892 4808 2908
rect 4760 2872 4776 2888
rect 4712 2812 4728 2828
rect 4680 2732 4696 2748
rect 4664 2692 4680 2708
rect 4616 2652 4632 2668
rect 4648 2652 4664 2668
rect 4520 2632 4536 2648
rect 4568 2612 4584 2628
rect 4600 2592 4616 2608
rect 4456 2532 4472 2548
rect 4520 2532 4536 2548
rect 4472 2512 4488 2528
rect 4536 2492 4552 2508
rect 4600 2492 4616 2508
rect 4440 2472 4456 2488
rect 4520 2472 4536 2488
rect 4552 2472 4568 2488
rect 4504 2452 4520 2468
rect 4808 2872 4824 2888
rect 4888 3112 4904 3128
rect 5064 3512 5080 3528
rect 5096 3492 5112 3508
rect 5080 3432 5096 3448
rect 5064 3352 5080 3368
rect 5096 3352 5112 3368
rect 5144 3712 5160 3728
rect 5320 4612 5336 4628
rect 5368 4612 5384 4628
rect 5304 4552 5320 4568
rect 5304 4472 5320 4488
rect 5448 4732 5464 4748
rect 5560 4732 5576 4748
rect 5944 5292 5960 5308
rect 5992 5292 6008 5308
rect 5912 5152 5928 5168
rect 5640 5132 5656 5148
rect 5832 5132 5848 5148
rect 5720 5092 5736 5108
rect 5800 5092 5816 5108
rect 5960 5092 5976 5108
rect 6008 5092 6024 5108
rect 5656 5032 5672 5048
rect 5480 4692 5496 4708
rect 5560 4692 5576 4708
rect 5608 4692 5624 4708
rect 5512 4672 5528 4688
rect 5448 4612 5464 4628
rect 5480 4612 5496 4628
rect 5448 4572 5464 4588
rect 5416 4552 5432 4568
rect 5384 4492 5400 4508
rect 5336 4472 5352 4488
rect 5400 4472 5416 4488
rect 5368 4452 5384 4468
rect 5384 4452 5400 4468
rect 5320 4392 5336 4408
rect 5304 4372 5320 4388
rect 5352 4192 5368 4208
rect 5432 4412 5448 4428
rect 5384 4292 5400 4308
rect 5416 4292 5432 4308
rect 5496 4552 5512 4568
rect 5464 4512 5480 4528
rect 5416 4232 5432 4248
rect 5400 4212 5416 4228
rect 5368 4152 5384 4168
rect 5208 4132 5224 4148
rect 5352 4132 5384 4148
rect 5176 4092 5208 4108
rect 5240 4052 5256 4068
rect 5213 4002 5249 4018
rect 5192 3872 5208 3888
rect 5288 4112 5304 4128
rect 5304 4112 5320 4128
rect 5176 3592 5192 3608
rect 5160 3512 5176 3528
rect 5144 3492 5160 3508
rect 4968 3292 4984 3308
rect 5000 3292 5032 3308
rect 4968 3232 4984 3248
rect 4936 3212 4952 3228
rect 4920 3112 4936 3128
rect 4968 3112 4984 3128
rect 5096 3112 5112 3128
rect 4920 3092 4936 3108
rect 5032 3092 5048 3108
rect 4856 3052 4872 3068
rect 5032 3072 5048 3088
rect 5048 3072 5064 3088
rect 5080 3072 5096 3088
rect 5032 3052 5048 3068
rect 4984 3032 5000 3048
rect 4920 2992 4936 3008
rect 4936 2952 4952 2968
rect 5000 2952 5016 2968
rect 4872 2932 4888 2948
rect 4968 2932 4984 2948
rect 4872 2912 4888 2928
rect 4920 2912 4936 2928
rect 4856 2872 4872 2888
rect 4840 2812 4856 2828
rect 4776 2792 4792 2808
rect 4776 2712 4792 2728
rect 4776 2692 4792 2708
rect 4824 2692 4840 2708
rect 4728 2672 4744 2688
rect 4744 2652 4760 2668
rect 4744 2632 4760 2648
rect 4712 2572 4728 2588
rect 4632 2552 4648 2568
rect 4712 2532 4728 2548
rect 4664 2512 4680 2528
rect 4648 2492 4664 2508
rect 4616 2452 4632 2468
rect 4744 2452 4760 2468
rect 4664 2432 4680 2448
rect 4920 2872 4936 2888
rect 4888 2832 4904 2848
rect 4936 2772 4952 2788
rect 4904 2732 4920 2748
rect 4888 2712 4904 2728
rect 4856 2632 4872 2648
rect 4792 2612 4808 2628
rect 4808 2532 4824 2548
rect 4792 2512 4808 2528
rect 4792 2492 4808 2508
rect 4568 2372 4584 2388
rect 4440 2292 4456 2308
rect 4712 2292 4728 2308
rect 4936 2692 4952 2708
rect 4968 2872 4984 2888
rect 4968 2852 4984 2868
rect 5016 2832 5032 2848
rect 5080 2992 5096 3008
rect 5064 2972 5080 2988
rect 5160 3472 5176 3488
rect 5256 3692 5272 3708
rect 5224 3632 5240 3648
rect 5213 3602 5249 3618
rect 5208 3572 5224 3588
rect 5192 3412 5208 3428
rect 5176 3352 5192 3368
rect 5256 3352 5272 3368
rect 5240 3232 5256 3248
rect 5192 3192 5208 3208
rect 5213 3202 5249 3218
rect 5160 3172 5176 3188
rect 5144 3032 5160 3048
rect 5128 2932 5144 2948
rect 5128 2752 5144 2768
rect 5064 2692 5080 2708
rect 5112 2692 5128 2708
rect 4952 2592 4968 2608
rect 4952 2572 4968 2588
rect 4920 2552 4936 2568
rect 4968 2532 4984 2548
rect 4952 2512 4968 2528
rect 4952 2432 4968 2448
rect 5000 2432 5016 2448
rect 4872 2392 4888 2408
rect 4872 2372 4888 2388
rect 4424 2272 4440 2288
rect 4696 2272 4712 2288
rect 4584 2252 4600 2268
rect 4632 2252 4648 2268
rect 4536 2192 4552 2208
rect 4568 2192 4584 2208
rect 4472 2172 4488 2188
rect 4456 2112 4472 2128
rect 4632 2232 4648 2248
rect 4520 2112 4536 2128
rect 4600 2112 4616 2128
rect 4456 2092 4472 2108
rect 4504 2092 4520 2108
rect 4536 2092 4552 2108
rect 4312 2052 4328 2068
rect 4248 1972 4264 1988
rect 4328 1972 4344 1988
rect 4232 1932 4248 1948
rect 4248 1932 4280 1948
rect 4328 1892 4344 1908
rect 4280 1872 4296 1888
rect 4248 1832 4264 1848
rect 4205 1802 4241 1818
rect 4216 1772 4232 1788
rect 4104 1712 4120 1728
rect 4120 1712 4136 1728
rect 4184 1712 4200 1728
rect 4120 1552 4152 1568
rect 4296 1792 4312 1808
rect 4376 2072 4392 2088
rect 4440 2072 4456 2088
rect 4456 2072 4472 2088
rect 4376 2012 4392 2028
rect 4424 2012 4440 2028
rect 4568 2072 4584 2088
rect 4520 1972 4536 1988
rect 4536 1952 4552 1968
rect 4472 1932 4488 1948
rect 4488 1912 4504 1928
rect 4520 1912 4536 1928
rect 4456 1892 4472 1908
rect 4376 1872 4392 1888
rect 4360 1832 4376 1848
rect 4424 1812 4440 1828
rect 4344 1772 4360 1788
rect 4312 1732 4328 1748
rect 4376 1732 4392 1748
rect 4248 1712 4264 1728
rect 4424 1712 4440 1728
rect 4216 1692 4232 1708
rect 4328 1692 4344 1708
rect 4232 1672 4248 1688
rect 4248 1672 4264 1688
rect 4312 1672 4328 1688
rect 4264 1572 4280 1588
rect 4408 1672 4424 1688
rect 4328 1632 4344 1648
rect 4376 1632 4392 1648
rect 4408 1632 4424 1648
rect 4440 1632 4456 1648
rect 4392 1572 4408 1588
rect 4264 1532 4296 1548
rect 4104 1512 4120 1528
rect 4168 1512 4184 1528
rect 4088 1492 4104 1508
rect 4344 1472 4360 1488
rect 4072 1452 4088 1468
rect 4264 1452 4280 1468
rect 4312 1452 4328 1468
rect 4312 1432 4328 1448
rect 4056 1412 4072 1428
rect 4088 1412 4104 1428
rect 4008 1372 4056 1388
rect 4008 1352 4024 1368
rect 4024 1312 4056 1328
rect 4072 1312 4088 1328
rect 4205 1402 4241 1418
rect 4248 1412 4264 1428
rect 4248 1352 4280 1368
rect 4152 1332 4168 1348
rect 4280 1332 4296 1348
rect 4168 1312 4184 1328
rect 4312 1312 4328 1328
rect 4392 1312 4408 1328
rect 4424 1552 4440 1568
rect 4440 1532 4456 1548
rect 4488 1832 4504 1848
rect 4504 1772 4520 1788
rect 4584 2052 4600 2068
rect 4632 2132 4648 2148
rect 4776 2192 4792 2208
rect 4760 2152 4776 2168
rect 4696 2132 4712 2148
rect 4664 2112 4680 2128
rect 4824 2072 4840 2088
rect 4632 2052 4648 2068
rect 4808 2052 4824 2068
rect 4728 2012 4744 2028
rect 4840 1972 4856 1988
rect 4792 1932 4808 1948
rect 4824 1932 4840 1948
rect 4600 1912 4616 1928
rect 4664 1912 4680 1928
rect 4760 1912 4776 1928
rect 4600 1892 4616 1908
rect 4632 1892 4648 1908
rect 4872 1912 4888 1928
rect 4776 1872 4792 1888
rect 4680 1852 4696 1868
rect 4712 1852 4728 1868
rect 4584 1812 4600 1828
rect 4648 1792 4680 1808
rect 4552 1732 4568 1748
rect 4616 1732 4632 1748
rect 4696 1732 4712 1748
rect 4568 1712 4584 1728
rect 4632 1712 4648 1728
rect 4648 1712 4664 1728
rect 4696 1712 4712 1728
rect 4536 1692 4552 1708
rect 4568 1692 4584 1708
rect 4664 1692 4680 1708
rect 4808 1792 4824 1808
rect 4760 1732 4776 1748
rect 4744 1692 4760 1708
rect 4664 1672 4680 1688
rect 4776 1672 4792 1688
rect 4616 1652 4632 1668
rect 4744 1652 4760 1668
rect 4584 1612 4600 1628
rect 4680 1552 4696 1568
rect 4728 1552 4744 1568
rect 4504 1532 4520 1548
rect 4664 1532 4680 1548
rect 4472 1512 4488 1528
rect 4616 1512 4632 1528
rect 4456 1472 4472 1488
rect 4552 1472 4568 1488
rect 4440 1412 4456 1428
rect 4584 1452 4600 1468
rect 4648 1412 4664 1428
rect 4584 1392 4600 1408
rect 4456 1312 4472 1328
rect 4552 1312 4568 1328
rect 4600 1312 4616 1328
rect 4280 1292 4296 1308
rect 4504 1292 4520 1308
rect 4552 1292 4568 1308
rect 3912 1272 3928 1288
rect 3992 1272 4008 1288
rect 4056 1272 4072 1288
rect 4072 1272 4088 1288
rect 3928 1252 3944 1268
rect 3992 1252 4008 1268
rect 4008 1252 4024 1268
rect 3816 1112 3832 1128
rect 3848 1112 3880 1128
rect 3928 1112 3944 1128
rect 3976 1152 3992 1168
rect 3784 1092 3800 1108
rect 3816 1092 3832 1108
rect 3864 1092 3880 1108
rect 3784 1072 3800 1088
rect 3784 1052 3800 1068
rect 3816 1052 3832 1068
rect 3848 972 3864 988
rect 3848 952 3864 968
rect 3832 932 3848 948
rect 3848 912 3864 928
rect 3768 872 3784 888
rect 3800 892 3816 908
rect 3864 892 3880 908
rect 3736 752 3752 768
rect 3640 712 3656 728
rect 3736 712 3752 728
rect 3832 872 3848 888
rect 3896 1072 3912 1088
rect 4200 1272 4216 1288
rect 4344 1272 4360 1288
rect 4104 1252 4120 1268
rect 4232 1232 4248 1248
rect 4104 1152 4120 1168
rect 4312 1132 4328 1148
rect 4056 1112 4072 1128
rect 4088 1112 4104 1128
rect 4280 1112 4296 1128
rect 3992 1072 4008 1088
rect 3960 1052 3976 1068
rect 4088 1092 4104 1108
rect 4136 1092 4152 1108
rect 4184 1092 4200 1108
rect 4264 1092 4280 1108
rect 4056 1072 4072 1088
rect 4088 1072 4104 1088
rect 4120 1052 4136 1068
rect 4248 1052 4264 1068
rect 4312 1052 4328 1068
rect 3976 1012 3992 1028
rect 4008 1012 4024 1028
rect 3944 932 3960 948
rect 3912 912 3928 928
rect 3928 912 3944 928
rect 3960 892 3976 908
rect 3896 872 3912 888
rect 3960 852 3976 868
rect 3912 832 3928 848
rect 4024 992 4040 1008
rect 4072 952 4088 968
rect 4104 952 4120 968
rect 4056 912 4088 928
rect 4120 912 4136 928
rect 3992 892 4008 908
rect 3992 872 4008 888
rect 4024 872 4040 888
rect 3848 772 3864 788
rect 3848 752 3864 768
rect 3896 752 3912 768
rect 3832 732 3848 748
rect 4024 772 4040 788
rect 3816 712 3832 728
rect 3848 712 3864 728
rect 4205 1002 4241 1018
rect 4248 952 4264 968
rect 4200 912 4216 928
rect 4264 912 4280 928
rect 4184 892 4200 908
rect 4232 892 4248 908
rect 4056 792 4072 808
rect 4120 872 4136 888
rect 4312 912 4328 928
rect 4328 892 4344 908
rect 4360 1212 4376 1228
rect 4376 1152 4392 1168
rect 4440 1232 4456 1248
rect 4408 1172 4424 1188
rect 4360 1132 4376 1148
rect 4392 1132 4408 1148
rect 4392 1112 4408 1128
rect 4504 1272 4520 1288
rect 4472 1212 4488 1228
rect 4632 1312 4648 1328
rect 4520 1252 4536 1268
rect 4616 1252 4632 1268
rect 4552 1232 4568 1248
rect 4520 1212 4536 1228
rect 4504 1192 4520 1208
rect 4440 1152 4472 1168
rect 4536 1192 4552 1208
rect 4664 1372 4680 1388
rect 4680 1332 4696 1348
rect 4680 1312 4696 1328
rect 4680 1272 4696 1288
rect 4552 1152 4568 1168
rect 4664 1152 4680 1168
rect 4504 1112 4520 1128
rect 4520 1112 4536 1128
rect 4792 1512 4808 1528
rect 4712 1472 4728 1488
rect 4728 1472 4744 1488
rect 4728 1452 4744 1468
rect 4408 1072 4424 1088
rect 4456 1072 4472 1088
rect 4376 1032 4392 1048
rect 4408 992 4424 1008
rect 4248 872 4280 888
rect 4344 852 4360 868
rect 4312 812 4328 828
rect 4136 752 4152 768
rect 4280 752 4296 768
rect 4088 732 4104 748
rect 4120 732 4136 748
rect 4248 732 4264 748
rect 4328 732 4344 748
rect 4104 712 4120 728
rect 4328 712 4344 728
rect 3816 692 3848 708
rect 3896 692 3912 708
rect 3992 692 4008 708
rect 4040 692 4056 708
rect 4120 692 4136 708
rect 3720 672 3736 688
rect 3800 672 3816 688
rect 3688 652 3704 668
rect 3704 652 3720 668
rect 3784 652 3800 668
rect 3784 632 3800 648
rect 3768 552 3784 568
rect 3720 532 3736 548
rect 3768 532 3784 548
rect 3704 512 3720 528
rect 3624 492 3640 508
rect 3704 412 3736 428
rect 3704 392 3720 408
rect 3688 352 3704 368
rect 3608 332 3624 348
rect 3656 272 3672 288
rect 3640 212 3656 228
rect 3544 192 3576 208
rect 3624 192 3640 208
rect 3528 152 3544 168
rect 3544 132 3560 148
rect 3752 332 3768 348
rect 3848 652 3864 668
rect 3816 512 3832 528
rect 3816 492 3832 508
rect 3800 392 3816 408
rect 4040 672 4056 688
rect 4104 672 4120 688
rect 3976 632 3992 648
rect 3896 572 3912 588
rect 3928 572 3944 588
rect 3896 552 3912 568
rect 3864 532 3880 548
rect 3864 512 3880 528
rect 3848 432 3864 448
rect 3944 532 3960 548
rect 3912 352 3928 368
rect 3816 292 3832 308
rect 3880 292 3896 308
rect 3992 412 4008 428
rect 4056 572 4072 588
rect 4264 672 4280 688
rect 4152 652 4168 668
rect 4296 632 4312 648
rect 4205 602 4241 618
rect 4264 612 4280 628
rect 4200 572 4216 588
rect 4296 572 4312 588
rect 4104 552 4120 568
rect 4312 552 4328 568
rect 4104 532 4120 548
rect 4152 532 4168 548
rect 4328 532 4344 548
rect 4520 1092 4536 1108
rect 4504 1052 4520 1068
rect 4488 1012 4504 1028
rect 4488 972 4504 988
rect 4536 1032 4552 1048
rect 4504 952 4520 968
rect 4456 932 4472 948
rect 4520 932 4536 948
rect 4552 932 4568 948
rect 4632 1072 4648 1088
rect 4616 1012 4632 1028
rect 4600 952 4616 968
rect 4488 912 4504 928
rect 4520 912 4536 928
rect 4584 912 4600 928
rect 4648 992 4664 1008
rect 4632 932 4648 948
rect 4408 872 4440 888
rect 4472 872 4488 888
rect 4376 832 4392 848
rect 4392 712 4408 728
rect 4376 692 4392 708
rect 4392 672 4408 688
rect 4472 652 4488 668
rect 4408 632 4424 648
rect 4392 612 4408 628
rect 4408 592 4424 608
rect 4520 892 4536 908
rect 4584 872 4600 888
rect 4584 732 4600 748
rect 4520 692 4536 708
rect 4616 692 4632 708
rect 4600 672 4616 688
rect 4440 532 4456 548
rect 4472 532 4488 548
rect 4520 532 4536 548
rect 4104 492 4120 508
rect 4072 392 4088 408
rect 4104 392 4120 408
rect 4024 352 4040 368
rect 4072 332 4088 348
rect 3784 272 3800 288
rect 3832 272 3848 288
rect 3816 252 3832 268
rect 3864 252 3880 268
rect 3672 172 3688 188
rect 3656 152 3672 168
rect 3848 152 3864 168
rect 3976 232 3992 248
rect 3992 172 4008 188
rect 3944 152 3960 168
rect 4088 272 4104 288
rect 4392 492 4408 508
rect 4296 472 4312 488
rect 4152 292 4184 308
rect 4312 352 4328 368
rect 4376 352 4392 368
rect 4408 352 4424 368
rect 4296 292 4312 308
rect 4328 332 4344 348
rect 4376 332 4392 348
rect 4168 272 4184 288
rect 4264 272 4280 288
rect 4376 272 4392 288
rect 4200 252 4216 268
rect 4360 252 4376 268
rect 4120 232 4136 248
rect 4232 232 4248 248
rect 4205 202 4241 218
rect 4104 172 4120 188
rect 4232 152 4248 168
rect 3224 112 3240 128
rect 3320 114 3336 128
rect 3320 112 3336 114
rect 3592 112 3608 128
rect 3656 114 3672 128
rect 3656 112 3672 114
rect 4056 112 4072 128
rect 4216 112 4232 128
rect 4312 112 4328 128
rect 312 92 328 108
rect 392 92 408 108
rect 424 92 440 108
rect 680 92 696 108
rect 728 92 744 108
rect 1256 92 1272 108
rect 1288 92 1304 108
rect 1496 92 1512 108
rect 1560 92 1576 108
rect 1864 92 1880 108
rect 2184 92 2200 108
rect 2280 92 2296 108
rect 2312 92 2328 108
rect 2744 92 2760 108
rect 2792 92 2808 108
rect 3144 92 3160 108
rect 3224 92 3240 108
rect 3560 92 3592 108
rect 4024 92 4040 108
rect 4072 92 4088 108
rect 4392 92 4408 108
rect 1117 2 1153 18
rect 3165 2 3201 18
rect 4024 12 4040 28
rect 4424 292 4440 308
rect 4568 632 4584 648
rect 4696 1112 4712 1128
rect 4808 1472 4824 1488
rect 4952 2412 4968 2428
rect 5000 2332 5016 2348
rect 4968 2312 4984 2328
rect 4920 2172 4936 2188
rect 4952 2152 4968 2168
rect 4920 2132 4936 2148
rect 5048 2372 5064 2388
rect 5112 2512 5128 2528
rect 5144 2712 5160 2728
rect 5160 2632 5176 2648
rect 5256 3052 5272 3068
rect 5240 2872 5256 2888
rect 5213 2802 5249 2818
rect 5256 2792 5272 2808
rect 5208 2712 5224 2728
rect 5304 3872 5320 3888
rect 5320 3872 5336 3888
rect 5320 3812 5336 3828
rect 5288 3732 5304 3748
rect 5416 4152 5432 4168
rect 5400 4052 5416 4068
rect 5448 4112 5464 4128
rect 5480 4452 5496 4468
rect 5608 4652 5624 4668
rect 5656 5012 5672 5028
rect 5640 4952 5656 4968
rect 5640 4932 5656 4948
rect 5720 5012 5736 5028
rect 5672 4972 5688 4988
rect 5688 4972 5704 4988
rect 5848 5012 5864 5028
rect 5816 4992 5832 5008
rect 5672 4772 5688 4788
rect 5656 4732 5672 4748
rect 6136 5332 6152 5348
rect 6312 5332 6328 5348
rect 6360 5332 6376 5348
rect 6584 5332 6600 5348
rect 6648 5332 6664 5348
rect 6744 5332 6760 5348
rect 6104 5312 6120 5328
rect 6536 5312 6552 5328
rect 6056 5292 6072 5308
rect 6120 5292 6136 5308
rect 6056 5212 6072 5228
rect 5928 4992 5944 5008
rect 5912 4972 5944 4988
rect 5832 4952 5848 4968
rect 5752 4832 5768 4848
rect 5800 4832 5816 4848
rect 5944 4952 5960 4968
rect 6040 5052 6056 5068
rect 5864 4912 5880 4928
rect 5912 4912 5928 4928
rect 5896 4892 5912 4908
rect 6024 4892 6040 4908
rect 5896 4872 5912 4888
rect 5848 4772 5864 4788
rect 5832 4752 5848 4768
rect 5752 4732 5768 4748
rect 5768 4732 5784 4748
rect 5816 4732 5832 4748
rect 5688 4712 5704 4728
rect 5544 4612 5560 4628
rect 5624 4612 5640 4628
rect 5528 4532 5544 4548
rect 5576 4572 5592 4588
rect 5592 4572 5608 4588
rect 5640 4572 5656 4588
rect 5560 4552 5576 4568
rect 5576 4552 5592 4568
rect 5656 4552 5672 4568
rect 5512 4412 5528 4428
rect 5528 4312 5544 4328
rect 5528 4292 5544 4308
rect 5496 4212 5512 4228
rect 5496 4192 5512 4208
rect 5512 4152 5528 4168
rect 5480 4112 5496 4128
rect 5560 4332 5576 4348
rect 5752 4692 5768 4708
rect 5688 4312 5704 4328
rect 5576 4152 5592 4168
rect 5544 4092 5560 4108
rect 5464 4052 5480 4068
rect 5528 4052 5544 4068
rect 5432 3952 5448 3968
rect 5528 3952 5544 3968
rect 5352 3892 5368 3908
rect 5384 3892 5400 3908
rect 5448 3912 5464 3928
rect 5432 3892 5448 3908
rect 5496 3872 5512 3888
rect 5512 3872 5528 3888
rect 5512 3852 5528 3868
rect 5416 3832 5432 3848
rect 5400 3812 5416 3828
rect 5352 3712 5368 3728
rect 5464 3752 5480 3768
rect 5496 3752 5512 3768
rect 5624 4212 5640 4228
rect 5672 4212 5688 4228
rect 5800 4612 5816 4628
rect 5752 4552 5768 4568
rect 5944 4832 5960 4848
rect 5832 4692 5848 4708
rect 5816 4572 5832 4588
rect 5800 4512 5816 4528
rect 5816 4512 5832 4528
rect 5880 4672 5896 4688
rect 5928 4652 5944 4668
rect 5880 4572 5896 4588
rect 5864 4532 5880 4548
rect 5848 4512 5864 4528
rect 5832 4492 5848 4508
rect 5736 4472 5752 4488
rect 5768 4472 5784 4488
rect 5816 4472 5832 4488
rect 5848 4452 5864 4468
rect 5848 4352 5864 4368
rect 5912 4492 5928 4508
rect 5928 4472 5944 4488
rect 5896 4372 5912 4388
rect 5880 4332 5896 4348
rect 5816 4272 5832 4288
rect 5832 4272 5848 4288
rect 5624 4132 5640 4148
rect 5704 4132 5720 4148
rect 5704 4112 5720 4128
rect 5752 4112 5768 4128
rect 5592 3972 5608 3988
rect 5560 3932 5576 3948
rect 5752 4072 5784 4088
rect 5640 4052 5656 4068
rect 5624 3912 5640 3928
rect 5720 3912 5736 3928
rect 5688 3872 5704 3888
rect 5592 3852 5608 3868
rect 5576 3752 5592 3768
rect 5512 3732 5528 3748
rect 5560 3732 5576 3748
rect 5592 3732 5608 3748
rect 5624 3732 5640 3748
rect 5432 3712 5448 3728
rect 5336 3692 5352 3708
rect 5368 3692 5384 3708
rect 5416 3692 5432 3708
rect 5448 3652 5464 3668
rect 5448 3632 5464 3648
rect 5336 3612 5352 3628
rect 5384 3612 5400 3628
rect 5304 3572 5320 3588
rect 5288 3452 5304 3468
rect 5320 3492 5336 3508
rect 5320 3472 5336 3488
rect 5416 3452 5432 3468
rect 5304 3392 5320 3408
rect 5288 3292 5304 3308
rect 5288 3212 5304 3228
rect 5352 3332 5368 3348
rect 5528 3452 5544 3468
rect 5656 3692 5672 3708
rect 5656 3652 5672 3668
rect 5592 3592 5608 3608
rect 5704 3792 5720 3808
rect 5704 3732 5720 3748
rect 5896 4272 5912 4288
rect 5928 4272 5944 4288
rect 5880 4252 5896 4268
rect 5800 4232 5816 4248
rect 5864 4212 5880 4228
rect 5848 4192 5864 4208
rect 5848 4112 5864 4128
rect 5784 3952 5800 3968
rect 5832 3912 5848 3928
rect 5800 3892 5816 3908
rect 5800 3812 5816 3828
rect 5784 3772 5800 3788
rect 5848 3892 5864 3908
rect 5976 4752 5992 4768
rect 6072 5112 6088 5128
rect 6120 5112 6136 5128
rect 6504 5112 6520 5128
rect 6280 5092 6296 5108
rect 6536 5092 6552 5108
rect 6104 5072 6120 5088
rect 6328 5072 6344 5088
rect 6440 5072 6456 5088
rect 6488 5072 6504 5088
rect 6504 5072 6520 5088
rect 6136 4952 6152 4968
rect 6136 4812 6152 4828
rect 6237 5002 6273 5018
rect 6280 4952 6296 4968
rect 6408 5012 6424 5028
rect 6168 4912 6184 4928
rect 6216 4912 6232 4928
rect 6200 4892 6216 4908
rect 6392 4892 6408 4908
rect 6360 4872 6376 4888
rect 6232 4852 6248 4868
rect 6232 4812 6248 4828
rect 6168 4792 6184 4808
rect 6152 4732 6168 4748
rect 6104 4712 6120 4728
rect 6472 5052 6488 5068
rect 6568 5052 6584 5068
rect 6936 5372 6952 5388
rect 7224 5352 7240 5368
rect 6808 5332 6824 5348
rect 6904 5332 6920 5348
rect 7208 5332 7224 5348
rect 6872 5312 6888 5328
rect 7064 5312 7080 5328
rect 7224 5312 7240 5328
rect 7304 5312 7320 5328
rect 7048 5292 7064 5308
rect 6888 5272 6904 5288
rect 6968 5272 6984 5288
rect 7128 5272 7144 5288
rect 7160 5232 7176 5248
rect 7272 5192 7288 5208
rect 7320 5132 7336 5148
rect 7320 5112 7336 5128
rect 6872 5092 6888 5108
rect 6968 5092 6984 5108
rect 7144 5092 7160 5108
rect 7192 5092 7208 5108
rect 7304 5092 7320 5108
rect 6824 5072 6840 5088
rect 6792 5052 6808 5068
rect 6904 5052 6920 5068
rect 7016 5052 7032 5068
rect 6616 5032 6632 5048
rect 6696 5012 6712 5028
rect 6568 4972 6584 4988
rect 6712 4972 6728 4988
rect 6824 4972 6840 4988
rect 6488 4932 6504 4948
rect 6536 4932 6552 4948
rect 6472 4912 6488 4928
rect 6440 4832 6456 4848
rect 6552 4792 6568 4808
rect 6408 4772 6424 4788
rect 6440 4772 6456 4788
rect 6696 4932 6712 4948
rect 6760 4932 6776 4948
rect 6744 4912 6760 4928
rect 6648 4892 6664 4908
rect 6680 4892 6696 4908
rect 6808 4892 6824 4908
rect 6872 4892 6888 4908
rect 6952 4972 6968 4988
rect 6936 4912 6952 4928
rect 6632 4832 6648 4848
rect 6488 4732 6504 4748
rect 6472 4712 6488 4728
rect 6056 4692 6072 4708
rect 6136 4692 6152 4708
rect 6296 4692 6312 4708
rect 6424 4692 6440 4708
rect 5960 4672 5976 4688
rect 6216 4672 6232 4688
rect 5960 4652 5976 4668
rect 5960 4632 5976 4648
rect 5960 4592 5976 4608
rect 6088 4652 6104 4668
rect 6152 4652 6168 4668
rect 6120 4612 6136 4628
rect 6120 4572 6136 4588
rect 6040 4532 6056 4548
rect 6072 4532 6088 4548
rect 5960 4512 5976 4528
rect 6216 4632 6232 4648
rect 6237 4602 6273 4618
rect 6184 4552 6200 4568
rect 6088 4512 6104 4528
rect 6216 4512 6232 4528
rect 6056 4472 6072 4488
rect 6088 4472 6104 4488
rect 6120 4472 6136 4488
rect 5976 4392 5992 4408
rect 6040 4372 6056 4388
rect 5960 4352 5976 4368
rect 6056 4352 6072 4368
rect 6024 4312 6040 4328
rect 5976 4252 5992 4268
rect 5896 4212 5912 4228
rect 5944 4212 5960 4228
rect 5992 4132 6008 4148
rect 5912 4112 5928 4128
rect 6120 4452 6136 4468
rect 6136 4392 6152 4408
rect 6104 4312 6120 4328
rect 6120 4312 6136 4328
rect 6088 4252 6104 4268
rect 6072 4172 6088 4188
rect 6072 4152 6088 4168
rect 5896 4092 5912 4108
rect 5960 3892 5976 3908
rect 5912 3872 5928 3888
rect 5864 3852 5880 3868
rect 5880 3792 5896 3808
rect 5816 3752 5832 3768
rect 5976 3752 5992 3768
rect 5816 3732 5832 3748
rect 5896 3732 5912 3748
rect 5896 3692 5912 3708
rect 5688 3632 5704 3648
rect 5720 3632 5736 3648
rect 5800 3632 5816 3648
rect 5704 3572 5720 3588
rect 5752 3572 5768 3588
rect 5704 3532 5720 3548
rect 5640 3452 5656 3468
rect 5560 3412 5576 3428
rect 5416 3372 5432 3388
rect 5544 3372 5560 3388
rect 5416 3352 5432 3368
rect 5400 3312 5416 3328
rect 5432 3332 5448 3348
rect 5448 3312 5464 3328
rect 5496 3312 5512 3328
rect 5368 3292 5384 3308
rect 5368 3132 5384 3148
rect 5288 3112 5320 3128
rect 5384 3112 5400 3128
rect 5400 3072 5416 3088
rect 5416 3052 5432 3068
rect 5528 3292 5544 3308
rect 5624 3312 5640 3328
rect 5608 3292 5624 3308
rect 5576 3272 5592 3288
rect 5528 3252 5544 3268
rect 5512 3232 5528 3248
rect 5768 3532 5784 3548
rect 5784 3532 5800 3548
rect 5720 3512 5736 3528
rect 5752 3512 5768 3528
rect 5736 3492 5752 3508
rect 5768 3452 5784 3468
rect 5816 3592 5832 3608
rect 6056 4092 6072 4108
rect 6104 4052 6120 4068
rect 6088 4032 6104 4048
rect 6072 3992 6088 4008
rect 6088 3972 6104 3988
rect 6072 3932 6088 3948
rect 6200 4492 6216 4508
rect 6184 4472 6200 4488
rect 6168 4452 6184 4468
rect 6376 4672 6392 4688
rect 6312 4552 6328 4568
rect 6280 4452 6296 4468
rect 6232 4412 6248 4428
rect 6264 4352 6280 4368
rect 6168 4332 6184 4348
rect 6200 4332 6216 4348
rect 6216 4332 6232 4348
rect 6184 4312 6200 4328
rect 6328 4472 6344 4488
rect 6456 4532 6472 4548
rect 6376 4512 6392 4528
rect 6472 4512 6488 4528
rect 6440 4492 6456 4508
rect 6584 4752 6600 4768
rect 6664 4872 6680 4888
rect 6856 4872 6872 4888
rect 6664 4832 6680 4848
rect 6728 4832 6744 4848
rect 6696 4812 6712 4828
rect 6680 4792 6696 4808
rect 6552 4692 6568 4708
rect 6504 4652 6520 4668
rect 6520 4512 6536 4528
rect 6504 4492 6520 4508
rect 6392 4472 6408 4488
rect 6504 4472 6520 4488
rect 6344 4432 6360 4448
rect 6328 4412 6344 4428
rect 6296 4392 6312 4408
rect 6280 4312 6296 4328
rect 6152 4292 6168 4308
rect 6168 4192 6184 4208
rect 6424 4332 6440 4348
rect 6408 4312 6424 4328
rect 6456 4312 6472 4328
rect 6344 4292 6360 4308
rect 6392 4292 6408 4308
rect 6312 4272 6328 4288
rect 6328 4272 6344 4288
rect 6216 4252 6232 4268
rect 6440 4252 6456 4268
rect 6360 4232 6376 4248
rect 6568 4672 6584 4688
rect 6616 4732 6632 4748
rect 6728 4772 6744 4788
rect 6984 4872 7000 4888
rect 6936 4852 6952 4868
rect 6792 4792 6808 4808
rect 6776 4772 6792 4788
rect 6648 4712 6664 4728
rect 6632 4672 6648 4688
rect 6584 4612 6600 4628
rect 6584 4572 6600 4588
rect 6616 4552 6632 4568
rect 6632 4512 6648 4528
rect 6936 4752 6952 4768
rect 7128 5072 7144 5088
rect 7096 5052 7112 5068
rect 7032 5032 7048 5048
rect 7032 4972 7048 4988
rect 7176 5072 7192 5088
rect 7160 5032 7176 5048
rect 7304 5072 7320 5088
rect 7240 5052 7256 5068
rect 7288 5052 7304 5068
rect 7192 4992 7208 5008
rect 7208 4972 7224 4988
rect 7160 4914 7176 4928
rect 7160 4912 7176 4914
rect 7096 4872 7112 4888
rect 7000 4852 7016 4868
rect 6984 4832 7000 4848
rect 6968 4772 6984 4788
rect 6984 4752 7016 4768
rect 6792 4712 6808 4728
rect 6808 4712 6824 4728
rect 6696 4672 6712 4688
rect 6808 4692 6824 4708
rect 6760 4652 6776 4668
rect 6808 4652 6824 4668
rect 6712 4632 6728 4648
rect 6856 4712 6872 4728
rect 6872 4712 6888 4728
rect 6936 4692 6952 4708
rect 7064 4732 7080 4748
rect 7048 4712 7064 4728
rect 6920 4632 6936 4648
rect 6760 4612 6776 4628
rect 6824 4612 6840 4628
rect 6696 4552 6712 4568
rect 6744 4552 6760 4568
rect 6744 4532 6760 4548
rect 6632 4492 6648 4508
rect 6648 4492 6664 4508
rect 6680 4492 6696 4508
rect 6712 4492 6728 4508
rect 6872 4592 6888 4608
rect 6792 4572 6808 4588
rect 6792 4552 6808 4568
rect 6952 4552 6968 4568
rect 6808 4512 6824 4528
rect 6856 4512 6872 4528
rect 6568 4472 6584 4488
rect 6632 4452 6648 4468
rect 6680 4452 6696 4468
rect 6760 4452 6776 4468
rect 6712 4432 6728 4448
rect 6552 4392 6568 4408
rect 6648 4392 6664 4408
rect 6760 4372 6776 4388
rect 6952 4512 6968 4528
rect 6904 4492 6920 4508
rect 6840 4472 6856 4488
rect 6872 4472 6888 4488
rect 6920 4472 6936 4488
rect 6808 4432 6824 4448
rect 6680 4352 6696 4368
rect 6792 4352 6808 4368
rect 6568 4292 6584 4308
rect 6648 4272 6664 4288
rect 6216 4212 6232 4228
rect 6237 4202 6273 4218
rect 6280 4212 6296 4228
rect 6408 4212 6424 4228
rect 6520 4212 6536 4228
rect 6280 4152 6296 4168
rect 6264 4132 6280 4148
rect 6520 4192 6536 4208
rect 6424 4172 6440 4188
rect 6456 4172 6472 4188
rect 6296 4132 6312 4148
rect 6424 4132 6440 4148
rect 6200 4112 6216 4128
rect 6344 4112 6360 4128
rect 6200 4072 6216 4088
rect 6296 4012 6312 4028
rect 6216 3972 6232 3988
rect 6120 3932 6136 3948
rect 6152 3932 6168 3948
rect 6120 3892 6136 3908
rect 6104 3872 6120 3888
rect 6088 3792 6104 3808
rect 6328 3972 6344 3988
rect 6280 3892 6296 3908
rect 6120 3852 6136 3868
rect 6216 3872 6232 3888
rect 6200 3772 6216 3788
rect 6104 3732 6120 3748
rect 6168 3732 6184 3748
rect 6056 3692 6072 3708
rect 6008 3652 6024 3668
rect 5832 3552 5848 3568
rect 5912 3532 5928 3548
rect 5848 3412 5864 3428
rect 5880 3372 5896 3388
rect 5768 3352 5784 3368
rect 5848 3352 5864 3368
rect 5896 3352 5912 3368
rect 5832 3332 5848 3348
rect 5704 3312 5720 3328
rect 5672 3272 5688 3288
rect 5640 3232 5656 3248
rect 5672 3232 5688 3248
rect 5688 3212 5704 3228
rect 5768 3292 5784 3308
rect 5752 3252 5768 3268
rect 5864 3292 5880 3308
rect 5848 3272 5864 3288
rect 5800 3232 5816 3248
rect 5576 3152 5608 3168
rect 5624 3152 5640 3168
rect 5480 3132 5496 3148
rect 5480 3092 5496 3108
rect 5448 3072 5464 3088
rect 5432 2992 5448 3008
rect 5400 2952 5416 2968
rect 5448 2932 5464 2948
rect 5496 2932 5512 2948
rect 5384 2912 5400 2928
rect 5288 2852 5304 2868
rect 5368 2732 5384 2748
rect 5304 2712 5320 2728
rect 5336 2712 5352 2728
rect 5256 2672 5272 2688
rect 5240 2652 5256 2668
rect 5240 2612 5256 2628
rect 5272 2592 5288 2608
rect 5272 2552 5288 2568
rect 5320 2652 5336 2668
rect 5320 2612 5336 2628
rect 5448 2892 5464 2908
rect 5416 2872 5432 2888
rect 5400 2732 5416 2748
rect 5384 2572 5400 2588
rect 5352 2552 5368 2568
rect 5288 2512 5304 2528
rect 5304 2512 5320 2528
rect 5176 2412 5192 2428
rect 5213 2402 5249 2418
rect 5128 2332 5144 2348
rect 5208 2312 5224 2328
rect 5528 3112 5544 3128
rect 5544 3092 5560 3108
rect 5720 3132 5736 3148
rect 5832 3132 5848 3148
rect 5592 3112 5608 3128
rect 5576 3072 5592 3088
rect 5624 3092 5640 3108
rect 5640 3092 5656 3108
rect 5608 3052 5624 3068
rect 5576 2952 5592 2968
rect 5544 2932 5560 2948
rect 5576 2932 5592 2948
rect 5704 3092 5720 3108
rect 5688 3052 5704 3068
rect 5704 2952 5720 2968
rect 5656 2912 5672 2928
rect 5512 2892 5528 2908
rect 5576 2872 5592 2888
rect 5528 2852 5544 2868
rect 5496 2832 5512 2848
rect 5480 2812 5496 2828
rect 5432 2712 5464 2728
rect 5416 2612 5432 2628
rect 5416 2592 5432 2608
rect 5368 2432 5384 2448
rect 5320 2312 5336 2328
rect 5176 2292 5192 2308
rect 5016 2212 5032 2228
rect 5064 2212 5080 2228
rect 5016 2192 5032 2208
rect 5128 2272 5144 2288
rect 5112 2232 5128 2248
rect 5144 2252 5160 2268
rect 5096 2152 5112 2168
rect 5096 2112 5112 2128
rect 5000 2092 5016 2108
rect 5032 2032 5048 2048
rect 5144 2032 5160 2048
rect 4968 1932 4984 1948
rect 4888 1852 4904 1868
rect 4888 1772 4904 1788
rect 4984 1912 5000 1928
rect 4952 1832 4968 1848
rect 4984 1852 5000 1868
rect 5000 1812 5016 1828
rect 4904 1752 4936 1768
rect 4968 1752 4984 1768
rect 4984 1732 5000 1748
rect 4920 1712 4936 1728
rect 4984 1712 5000 1728
rect 4840 1692 4856 1708
rect 5256 2272 5272 2288
rect 5272 2272 5288 2288
rect 5208 2152 5224 2168
rect 5213 2002 5249 2018
rect 5176 1892 5192 1908
rect 5112 1852 5128 1868
rect 5192 1852 5208 1868
rect 5096 1792 5112 1808
rect 5016 1772 5032 1788
rect 5176 1832 5192 1848
rect 5176 1792 5192 1808
rect 5192 1772 5208 1788
rect 5224 1752 5240 1768
rect 5112 1732 5128 1748
rect 5080 1712 5096 1728
rect 5096 1712 5112 1728
rect 5144 1712 5160 1728
rect 4872 1632 4888 1648
rect 5032 1692 5048 1708
rect 4904 1552 4920 1568
rect 4952 1512 4968 1528
rect 4856 1492 4872 1508
rect 5016 1672 5032 1688
rect 5064 1672 5080 1688
rect 5192 1672 5208 1688
rect 5176 1632 5192 1648
rect 5224 1632 5240 1648
rect 5048 1572 5064 1588
rect 5064 1512 5080 1528
rect 5064 1492 5080 1508
rect 5112 1612 5128 1628
rect 5160 1532 5176 1548
rect 5048 1472 5064 1488
rect 5096 1472 5112 1488
rect 4760 1452 4776 1468
rect 4824 1452 4840 1468
rect 4824 1412 4840 1428
rect 4920 1412 4936 1428
rect 4872 1392 4888 1408
rect 4920 1392 4936 1408
rect 4968 1392 4984 1408
rect 4840 1332 4856 1348
rect 4888 1332 4904 1348
rect 4760 1292 4776 1308
rect 4824 1172 4840 1188
rect 4984 1172 5000 1188
rect 4792 1152 4808 1168
rect 4792 1132 4808 1148
rect 5096 1452 5112 1468
rect 5213 1602 5249 1618
rect 5192 1492 5208 1508
rect 5384 2352 5400 2368
rect 5672 2892 5704 2908
rect 5688 2872 5704 2888
rect 5704 2872 5720 2888
rect 5672 2852 5688 2868
rect 5640 2772 5656 2788
rect 5480 2672 5496 2688
rect 5624 2712 5640 2728
rect 5640 2712 5656 2728
rect 5736 3092 5752 3108
rect 5784 3112 5800 3128
rect 5768 3072 5784 3088
rect 5880 3212 5896 3228
rect 5880 3192 5896 3208
rect 5848 3092 5864 3108
rect 5816 3072 5832 3088
rect 5800 3012 5816 3028
rect 5752 2912 5768 2928
rect 5800 2892 5816 2908
rect 6088 3392 6104 3408
rect 5944 3372 5960 3388
rect 5992 3372 6008 3388
rect 6152 3712 6168 3728
rect 6168 3692 6184 3708
rect 6152 3612 6168 3628
rect 6152 3532 6168 3548
rect 6120 3412 6136 3428
rect 6184 3672 6200 3688
rect 6237 3802 6273 3818
rect 6232 3752 6248 3768
rect 6360 4012 6376 4028
rect 6440 4012 6456 4028
rect 6616 4172 6632 4188
rect 6536 4152 6552 4168
rect 6552 4132 6568 4148
rect 6648 4132 6664 4148
rect 6712 4332 6728 4348
rect 6728 4332 6744 4348
rect 6776 4332 6792 4348
rect 6792 4332 6808 4348
rect 6792 4292 6808 4308
rect 6984 4692 7000 4708
rect 7000 4672 7016 4688
rect 6984 4532 7000 4548
rect 6824 4272 6840 4288
rect 6744 4232 6760 4248
rect 6872 4312 6888 4328
rect 6888 4292 6904 4308
rect 6936 4292 6952 4308
rect 6856 4252 6872 4268
rect 6728 4212 6744 4228
rect 6712 4152 6728 4168
rect 6600 4112 6616 4128
rect 6664 4112 6696 4128
rect 6488 4052 6504 4068
rect 6536 4052 6552 4068
rect 6456 3952 6472 3968
rect 6344 3932 6360 3948
rect 6392 3906 6408 3908
rect 6392 3892 6408 3906
rect 6520 3972 6536 3988
rect 6616 4072 6632 4088
rect 6584 3972 6600 3988
rect 6584 3892 6600 3908
rect 6840 4092 6856 4108
rect 6776 3992 6792 4008
rect 6808 3952 6824 3968
rect 6632 3932 6648 3948
rect 6744 3932 6760 3948
rect 6792 3932 6808 3948
rect 6664 3912 6680 3928
rect 6616 3872 6632 3888
rect 6568 3832 6584 3848
rect 6488 3792 6504 3808
rect 6456 3752 6472 3768
rect 6264 3692 6280 3708
rect 6248 3672 6264 3688
rect 6200 3652 6232 3668
rect 6184 3612 6200 3628
rect 6264 3592 6280 3608
rect 6232 3552 6248 3568
rect 6200 3532 6216 3548
rect 6312 3532 6328 3548
rect 6344 3532 6360 3548
rect 6408 3692 6424 3708
rect 6376 3672 6392 3688
rect 6408 3672 6424 3688
rect 6280 3512 6296 3528
rect 6360 3512 6376 3528
rect 6200 3472 6216 3488
rect 5928 3292 5944 3308
rect 5944 3272 5960 3288
rect 5944 3252 5960 3268
rect 6024 3252 6040 3268
rect 6056 3252 6072 3268
rect 5928 3212 5944 3228
rect 5896 3112 5912 3128
rect 5896 3092 5912 3108
rect 5896 3072 5912 3088
rect 5864 3012 5880 3028
rect 5880 2912 5896 2928
rect 5720 2832 5736 2848
rect 5784 2832 5800 2848
rect 5736 2792 5752 2808
rect 5688 2712 5704 2728
rect 5752 2712 5784 2728
rect 5848 2792 5864 2808
rect 5864 2752 5880 2768
rect 5912 2952 5928 2968
rect 5944 3092 5960 3108
rect 5960 3092 5976 3108
rect 5976 3052 5992 3068
rect 6152 3232 6168 3248
rect 6232 3452 6248 3468
rect 6237 3402 6273 3418
rect 6392 3492 6408 3508
rect 6408 3472 6424 3488
rect 6328 3412 6344 3428
rect 6392 3392 6408 3408
rect 6280 3352 6296 3368
rect 6328 3352 6344 3368
rect 6360 3352 6376 3368
rect 6440 3652 6456 3668
rect 6424 3352 6440 3368
rect 6344 3312 6360 3328
rect 6408 3312 6424 3328
rect 6392 3292 6408 3308
rect 6200 3212 6216 3228
rect 6168 3192 6184 3208
rect 6088 3112 6104 3128
rect 6376 3112 6392 3128
rect 6424 3252 6440 3268
rect 6472 3512 6488 3528
rect 6536 3752 6552 3768
rect 6632 3832 6648 3848
rect 6680 3832 6696 3848
rect 6600 3812 6616 3828
rect 6616 3792 6632 3808
rect 6744 3892 6760 3908
rect 6920 4212 6936 4228
rect 6904 4172 6920 4188
rect 6968 4332 6984 4348
rect 7080 4652 7096 4668
rect 7064 4512 7080 4528
rect 7080 4492 7096 4508
rect 7032 4412 7048 4428
rect 7048 4352 7064 4368
rect 7080 4352 7096 4368
rect 7288 4992 7304 5008
rect 7272 4912 7288 4928
rect 7176 4832 7192 4848
rect 7240 4832 7256 4848
rect 7128 4752 7144 4768
rect 7128 4712 7144 4728
rect 7128 4692 7144 4708
rect 7144 4612 7160 4628
rect 7128 4552 7144 4568
rect 7208 4632 7224 4648
rect 7192 4572 7208 4588
rect 7272 4552 7288 4568
rect 7160 4472 7176 4488
rect 7160 4392 7176 4408
rect 7240 4514 7256 4528
rect 7240 4512 7256 4514
rect 7032 4332 7048 4348
rect 7112 4332 7128 4348
rect 7176 4332 7192 4348
rect 7000 4312 7016 4328
rect 6968 4212 6984 4228
rect 6984 4132 7000 4148
rect 6872 3992 6888 4008
rect 6840 3932 6856 3948
rect 6952 4012 6968 4028
rect 6968 3992 7000 4008
rect 6936 3952 6952 3968
rect 6968 3952 6984 3968
rect 6904 3932 6920 3948
rect 6872 3892 6888 3908
rect 6808 3872 6824 3888
rect 6760 3852 6776 3868
rect 6728 3832 6744 3848
rect 6760 3832 6776 3848
rect 6696 3732 6712 3748
rect 6584 3672 6600 3688
rect 6664 3592 6680 3608
rect 6584 3532 6600 3548
rect 6504 3492 6520 3508
rect 6552 3492 6568 3508
rect 6536 3472 6552 3488
rect 6536 3452 6552 3468
rect 6488 3412 6504 3428
rect 6472 3292 6488 3308
rect 6504 3292 6520 3308
rect 6632 3472 6648 3488
rect 6584 3452 6600 3468
rect 6632 3452 6648 3468
rect 6648 3432 6664 3448
rect 6728 3712 6744 3728
rect 6856 3712 6872 3728
rect 6712 3432 6728 3448
rect 6696 3392 6712 3408
rect 6840 3612 6856 3628
rect 6760 3532 6776 3548
rect 6824 3512 6840 3528
rect 6824 3492 6840 3508
rect 6776 3472 6792 3488
rect 6760 3372 6776 3388
rect 6632 3332 6648 3348
rect 6696 3332 6712 3348
rect 6744 3332 6760 3348
rect 6616 3312 6632 3328
rect 6680 3312 6696 3328
rect 6712 3312 6728 3328
rect 6568 3292 6584 3308
rect 6472 3252 6488 3268
rect 6728 3252 6744 3268
rect 6456 3192 6472 3208
rect 6744 3232 6760 3248
rect 6648 3172 6664 3188
rect 6680 3172 6696 3188
rect 6728 3152 6744 3168
rect 6936 3892 6952 3908
rect 6888 3832 6904 3848
rect 6952 3832 6968 3848
rect 6952 3792 6968 3808
rect 6888 3752 6904 3768
rect 7080 4252 7096 4268
rect 7032 4212 7048 4228
rect 7016 4112 7032 4128
rect 7016 4092 7032 4108
rect 7032 4072 7048 4088
rect 7016 3992 7032 4008
rect 7016 3972 7032 3988
rect 7000 3952 7016 3968
rect 7000 3932 7016 3948
rect 7048 3932 7064 3948
rect 7112 4292 7128 4308
rect 7128 4292 7144 4308
rect 7112 4272 7128 4288
rect 7128 4232 7144 4248
rect 7192 4312 7208 4328
rect 7208 4292 7224 4308
rect 7176 4272 7192 4288
rect 7224 4272 7240 4288
rect 7272 4272 7288 4288
rect 7160 4212 7176 4228
rect 7208 4212 7224 4228
rect 7256 4212 7272 4228
rect 7160 4172 7176 4188
rect 7128 4152 7144 4168
rect 7192 4152 7208 4168
rect 7304 4692 7320 4708
rect 7112 4052 7128 4068
rect 7064 3912 7080 3928
rect 7096 3912 7112 3928
rect 7048 3892 7064 3908
rect 7032 3872 7048 3888
rect 7096 3872 7112 3888
rect 7032 3852 7048 3868
rect 7128 3912 7144 3928
rect 7176 3912 7192 3928
rect 7160 3872 7176 3888
rect 6968 3752 6984 3768
rect 6936 3712 6952 3728
rect 6920 3692 6936 3708
rect 7048 3692 7064 3708
rect 6936 3592 6968 3608
rect 6984 3592 7000 3608
rect 6936 3552 6952 3568
rect 6872 3492 6888 3508
rect 7048 3552 7064 3568
rect 7144 3792 7160 3808
rect 7128 3732 7144 3748
rect 7144 3552 7160 3568
rect 7000 3532 7016 3548
rect 7064 3512 7080 3528
rect 7112 3512 7128 3528
rect 7016 3492 7032 3508
rect 6936 3452 6952 3468
rect 6904 3412 6920 3428
rect 6808 3292 6824 3308
rect 6792 3212 6808 3228
rect 6520 3132 6536 3148
rect 6776 3132 6792 3148
rect 6104 3092 6120 3108
rect 6152 3092 6168 3108
rect 6456 3092 6472 3108
rect 6184 3072 6200 3088
rect 6248 3072 6264 3088
rect 6248 3052 6264 3068
rect 6328 3072 6344 3088
rect 6264 3032 6280 3048
rect 6216 3012 6232 3028
rect 6237 3002 6273 3018
rect 6104 2952 6120 2968
rect 6152 2952 6168 2968
rect 5928 2912 5944 2928
rect 6056 2932 6072 2948
rect 6136 2932 6152 2948
rect 6344 2932 6360 2948
rect 6104 2912 6120 2928
rect 6264 2912 6280 2928
rect 6312 2912 6328 2928
rect 5992 2892 6008 2908
rect 5896 2872 5912 2888
rect 6024 2872 6040 2888
rect 5880 2732 5896 2748
rect 6328 2872 6344 2888
rect 6040 2812 6056 2828
rect 6328 2812 6344 2828
rect 6200 2792 6216 2808
rect 6024 2732 6040 2748
rect 5928 2712 5944 2728
rect 5800 2692 5816 2708
rect 5864 2692 5880 2708
rect 5608 2672 5624 2688
rect 5624 2672 5640 2688
rect 5880 2672 5896 2688
rect 5912 2672 5928 2688
rect 5528 2652 5544 2668
rect 5560 2652 5576 2668
rect 5528 2632 5544 2648
rect 5880 2632 5896 2648
rect 5560 2612 5576 2628
rect 5512 2592 5544 2608
rect 5656 2592 5672 2608
rect 5496 2552 5512 2568
rect 5496 2532 5512 2548
rect 5640 2552 5656 2568
rect 5480 2512 5496 2528
rect 5544 2512 5560 2528
rect 5528 2452 5544 2468
rect 5704 2572 5720 2588
rect 5704 2532 5720 2548
rect 5592 2452 5608 2468
rect 5560 2352 5592 2368
rect 5496 2332 5512 2348
rect 5416 2312 5432 2328
rect 5368 2292 5384 2308
rect 5400 2292 5416 2308
rect 5352 2272 5368 2288
rect 5384 2272 5400 2288
rect 5432 2272 5448 2288
rect 5304 2252 5320 2268
rect 5288 2232 5304 2248
rect 5272 2152 5288 2168
rect 5272 2072 5288 2088
rect 5320 1892 5336 1908
rect 5368 2172 5384 2188
rect 5448 2212 5464 2228
rect 5400 2152 5416 2168
rect 5608 2392 5624 2408
rect 5592 2332 5608 2348
rect 5496 2292 5512 2308
rect 5480 2232 5496 2248
rect 5480 2192 5496 2208
rect 5464 2172 5480 2188
rect 5496 2152 5512 2168
rect 5480 2132 5496 2148
rect 5384 2112 5400 2128
rect 5400 2112 5416 2128
rect 5384 2092 5400 2108
rect 5368 1872 5384 1888
rect 5288 1832 5304 1848
rect 5352 1772 5368 1788
rect 5304 1732 5320 1748
rect 5352 1732 5368 1748
rect 5368 1732 5384 1748
rect 5272 1692 5288 1708
rect 5288 1692 5320 1708
rect 5288 1532 5304 1548
rect 5272 1492 5288 1508
rect 5256 1472 5272 1488
rect 5256 1392 5272 1408
rect 5112 1352 5128 1368
rect 5176 1352 5192 1368
rect 5080 1332 5096 1348
rect 5208 1332 5224 1348
rect 5000 1152 5016 1168
rect 4712 1092 4728 1108
rect 4696 1072 4712 1088
rect 4680 1032 4696 1048
rect 4936 1112 4952 1128
rect 4856 1092 4872 1108
rect 4936 1092 4952 1108
rect 5144 1106 5160 1108
rect 5144 1092 5160 1106
rect 4760 1072 4776 1088
rect 4760 1052 4776 1068
rect 4744 1012 4760 1028
rect 4808 1032 4824 1048
rect 4856 1032 4872 1048
rect 4808 972 4824 988
rect 4840 932 4856 948
rect 4680 912 4696 928
rect 4760 912 4776 928
rect 4808 912 4824 928
rect 4696 892 4712 908
rect 4744 892 4760 908
rect 4776 892 4792 908
rect 4808 892 4824 908
rect 4904 1072 4920 1088
rect 4936 1072 4952 1088
rect 4968 1072 4984 1088
rect 4888 1052 4904 1068
rect 5016 1052 5048 1068
rect 4872 1012 4888 1028
rect 4920 992 4936 1008
rect 4904 912 4920 928
rect 4888 892 4904 908
rect 4968 972 4984 988
rect 4744 872 4760 888
rect 4664 712 4680 728
rect 4664 692 4680 708
rect 4664 672 4680 688
rect 4632 612 4648 628
rect 4568 572 4584 588
rect 4664 572 4680 588
rect 4552 552 4568 568
rect 4696 552 4712 568
rect 4632 532 4648 548
rect 4584 512 4600 528
rect 4632 512 4648 528
rect 4728 514 4744 528
rect 4728 512 4744 514
rect 4536 492 4552 508
rect 4824 672 4840 688
rect 4776 652 4792 668
rect 4648 312 4664 328
rect 4632 292 4648 308
rect 4520 272 4536 288
rect 4504 252 4520 268
rect 4536 192 4552 208
rect 4616 192 4632 208
rect 4424 152 4456 168
rect 4488 152 4504 168
rect 4440 112 4456 128
rect 4600 112 4616 128
rect 4472 92 4488 108
rect 4680 272 4696 288
rect 4856 572 4872 588
rect 4920 792 4936 808
rect 4904 732 4920 748
rect 4936 752 4952 768
rect 5016 932 5032 948
rect 5064 1012 5080 1028
rect 5213 1202 5249 1218
rect 5384 1452 5400 1468
rect 5368 1372 5384 1388
rect 5352 1332 5368 1348
rect 5384 1312 5400 1328
rect 5464 2092 5480 2108
rect 5416 1932 5432 1948
rect 5768 2532 5784 2548
rect 5672 2492 5688 2508
rect 5720 2492 5736 2508
rect 5736 2452 5752 2468
rect 5784 2432 5816 2448
rect 5656 2352 5672 2368
rect 5640 2312 5656 2328
rect 5720 2292 5736 2308
rect 5704 2272 5720 2288
rect 5672 2252 5688 2268
rect 5608 2232 5624 2248
rect 5592 2172 5608 2188
rect 5560 2132 5576 2148
rect 5528 2112 5544 2128
rect 5592 2112 5608 2128
rect 5624 2152 5640 2168
rect 5736 2172 5752 2188
rect 6008 2712 6024 2728
rect 6104 2692 6120 2708
rect 6152 2692 6168 2708
rect 5976 2652 5992 2668
rect 6088 2672 6104 2688
rect 6120 2672 6136 2688
rect 6232 2672 6248 2688
rect 6168 2652 6184 2668
rect 6008 2592 6024 2608
rect 6008 2572 6024 2588
rect 5960 2512 5976 2528
rect 5864 2452 5880 2468
rect 5848 2432 5864 2448
rect 5848 2412 5864 2428
rect 5832 2332 5848 2348
rect 5912 2332 5928 2348
rect 5912 2312 5928 2328
rect 5880 2292 5896 2308
rect 5864 2272 5880 2288
rect 5944 2272 5960 2288
rect 5848 2212 5864 2228
rect 5912 2212 5928 2228
rect 5656 2132 5672 2148
rect 5704 2132 5720 2148
rect 5816 2132 5832 2148
rect 5688 2112 5704 2128
rect 5800 2114 5816 2128
rect 5800 2112 5816 2114
rect 5608 2072 5624 2088
rect 5560 1952 5576 1968
rect 5432 1892 5448 1908
rect 5592 1892 5608 1908
rect 5448 1872 5464 1888
rect 5528 1872 5544 1888
rect 5464 1852 5480 1868
rect 5464 1832 5480 1848
rect 5496 1792 5512 1808
rect 5592 1852 5608 1868
rect 5544 1832 5560 1848
rect 5560 1792 5576 1808
rect 5592 1792 5608 1808
rect 5576 1772 5592 1788
rect 5480 1752 5496 1768
rect 5432 1732 5448 1748
rect 5576 1732 5592 1748
rect 5608 1772 5624 1788
rect 5432 1712 5448 1728
rect 5496 1712 5512 1728
rect 5464 1692 5480 1708
rect 5592 1692 5608 1708
rect 5528 1672 5544 1688
rect 5448 1612 5464 1628
rect 5480 1532 5496 1548
rect 5416 1512 5432 1528
rect 5544 1512 5548 1528
rect 5548 1512 5560 1528
rect 5512 1492 5528 1508
rect 5560 1492 5576 1508
rect 5576 1472 5592 1488
rect 5528 1452 5560 1468
rect 5448 1392 5464 1408
rect 5416 1372 5432 1388
rect 5416 1352 5432 1368
rect 5496 1332 5512 1348
rect 5464 1312 5480 1328
rect 5512 1292 5528 1308
rect 5480 1192 5496 1208
rect 5464 1132 5480 1148
rect 5432 1112 5448 1128
rect 5464 1112 5480 1128
rect 5240 1092 5256 1108
rect 5272 1092 5288 1108
rect 5320 1092 5336 1108
rect 5448 1092 5464 1108
rect 5336 1072 5352 1088
rect 5208 1052 5224 1068
rect 5080 972 5096 988
rect 5096 952 5112 968
rect 5176 952 5192 968
rect 5080 932 5096 948
rect 5016 872 5032 888
rect 5000 732 5016 748
rect 5000 712 5016 728
rect 4968 672 4984 688
rect 4920 652 4936 668
rect 4872 552 4888 568
rect 4920 552 4936 568
rect 4872 532 4888 548
rect 4792 492 4808 508
rect 4840 492 4856 508
rect 4904 512 4920 528
rect 4824 412 4840 428
rect 4744 292 4760 308
rect 4872 432 4888 448
rect 4920 292 4936 308
rect 4760 272 4776 288
rect 4856 272 4872 288
rect 4712 152 4728 168
rect 4728 132 4744 148
rect 4792 112 4808 128
rect 4728 92 4744 108
rect 4792 92 4808 108
rect 4872 172 4888 188
rect 4984 632 5000 648
rect 4952 572 4968 588
rect 4984 492 5000 508
rect 5064 832 5080 848
rect 5176 932 5192 948
rect 5112 912 5128 928
rect 5112 852 5128 868
rect 5096 732 5112 748
rect 5048 712 5064 728
rect 5080 712 5096 728
rect 5112 712 5128 728
rect 5048 692 5064 708
rect 5096 672 5112 688
rect 5112 672 5128 688
rect 5032 552 5048 568
rect 5160 732 5176 748
rect 5128 632 5144 648
rect 5112 532 5128 548
rect 5032 312 5048 328
rect 5128 312 5144 328
rect 5016 292 5032 308
rect 5080 292 5096 308
rect 5240 972 5256 988
rect 5352 972 5368 988
rect 5368 952 5384 968
rect 5304 914 5320 928
rect 5304 912 5320 914
rect 5213 802 5249 818
rect 5240 732 5256 748
rect 5400 912 5416 928
rect 5400 892 5416 908
rect 5624 1692 5640 1708
rect 5656 1972 5672 1988
rect 5752 1906 5768 1908
rect 5752 1892 5768 1906
rect 5928 2172 5944 2188
rect 6008 2512 6024 2528
rect 5976 2492 5992 2508
rect 5992 2492 6008 2508
rect 6136 2612 6152 2628
rect 6237 2602 6273 2618
rect 6184 2532 6200 2548
rect 6376 3052 6392 3068
rect 6424 3052 6440 3068
rect 6456 3032 6472 3048
rect 6728 3112 6744 3128
rect 6760 3112 6776 3128
rect 6488 2932 6504 2948
rect 6440 2912 6456 2928
rect 6440 2752 6456 2768
rect 6392 2712 6408 2728
rect 6472 2572 6488 2588
rect 6360 2552 6376 2568
rect 6408 2552 6424 2568
rect 6136 2512 6152 2528
rect 6200 2512 6216 2528
rect 6296 2512 6312 2528
rect 6072 2492 6088 2508
rect 6200 2492 6216 2508
rect 6328 2492 6344 2508
rect 6056 2472 6072 2488
rect 6088 2472 6104 2488
rect 6040 2432 6072 2448
rect 6024 2352 6040 2368
rect 6024 2292 6040 2308
rect 6040 2232 6056 2248
rect 6008 2172 6024 2188
rect 5960 2112 5976 2128
rect 6024 2112 6040 2128
rect 6136 2472 6152 2488
rect 6120 2392 6136 2408
rect 6072 2372 6088 2388
rect 6120 2372 6136 2388
rect 6088 2352 6104 2368
rect 6072 2332 6088 2348
rect 6216 2472 6232 2488
rect 6216 2432 6232 2448
rect 6248 2392 6264 2408
rect 6136 2312 6152 2328
rect 6136 2292 6152 2308
rect 6168 2292 6184 2308
rect 6104 2252 6120 2268
rect 6168 2252 6184 2268
rect 6136 2172 6152 2188
rect 6104 2112 6120 2128
rect 6056 2072 6072 2088
rect 5992 2052 6008 2068
rect 5976 2032 5992 2048
rect 6040 2032 6056 2048
rect 5928 1972 5944 1988
rect 5928 1932 5944 1948
rect 6072 2052 6088 2068
rect 6152 2112 6168 2128
rect 6200 2312 6216 2328
rect 6232 2312 6248 2328
rect 6472 2512 6488 2528
rect 6440 2492 6456 2508
rect 6360 2452 6376 2468
rect 6344 2412 6360 2428
rect 6296 2352 6312 2368
rect 6392 2372 6424 2388
rect 6488 2412 6504 2428
rect 6424 2312 6440 2328
rect 6472 2312 6504 2328
rect 6632 3032 6648 3048
rect 6648 2972 6664 2988
rect 6680 2952 6696 2968
rect 6568 2932 6584 2948
rect 6792 3092 6808 3108
rect 6568 2912 6584 2928
rect 6584 2912 6600 2928
rect 6664 2912 6680 2928
rect 6712 2912 6744 2928
rect 6776 2992 6792 3008
rect 6824 3112 6840 3128
rect 6904 3312 6920 3328
rect 6824 3092 6840 3108
rect 6808 2972 6824 2988
rect 6568 2892 6584 2908
rect 6760 2892 6776 2908
rect 6648 2772 6664 2788
rect 6616 2732 6632 2748
rect 6520 2692 6536 2708
rect 6584 2592 6600 2608
rect 6568 2552 6584 2568
rect 6568 2532 6584 2548
rect 6600 2512 6616 2528
rect 6520 2492 6536 2508
rect 6536 2472 6552 2488
rect 6520 2392 6536 2408
rect 6536 2352 6552 2368
rect 6680 2752 6696 2768
rect 6696 2612 6712 2628
rect 6808 2572 6824 2588
rect 6728 2532 6744 2548
rect 6776 2532 6792 2548
rect 6648 2512 6664 2528
rect 6616 2492 6632 2508
rect 6840 3052 6856 3068
rect 6840 2952 6856 2968
rect 6968 3412 6984 3428
rect 6952 3312 6968 3328
rect 7080 3492 7096 3508
rect 7032 3392 7048 3408
rect 7112 3472 7128 3488
rect 7144 3432 7160 3448
rect 7096 3352 7112 3368
rect 7160 3352 7176 3368
rect 6984 3332 7000 3348
rect 7128 3332 7144 3348
rect 6904 3272 6920 3288
rect 6952 3272 6968 3288
rect 6904 3232 6920 3248
rect 6872 3132 6888 3148
rect 6888 2952 6904 2968
rect 6936 3172 6952 3188
rect 6968 3132 6984 3148
rect 6936 3112 6952 3128
rect 6936 2932 6952 2948
rect 6872 2912 6888 2928
rect 6968 2914 6984 2928
rect 6968 2912 6984 2914
rect 6904 2892 6920 2908
rect 6920 2812 6936 2828
rect 6984 2812 7000 2828
rect 6856 2772 6872 2788
rect 6984 2772 7000 2788
rect 6904 2692 6920 2708
rect 6872 2632 6888 2648
rect 6840 2572 6856 2588
rect 6952 2572 6968 2588
rect 6856 2552 6872 2568
rect 6920 2552 6936 2568
rect 6728 2512 6744 2528
rect 6696 2412 6712 2428
rect 6744 2412 6760 2428
rect 6600 2372 6616 2388
rect 6632 2352 6648 2368
rect 6568 2312 6584 2328
rect 6600 2312 6616 2328
rect 6552 2292 6568 2308
rect 6360 2272 6376 2288
rect 6584 2272 6600 2288
rect 6328 2252 6344 2268
rect 6184 2232 6200 2248
rect 6216 2192 6232 2208
rect 6237 2202 6273 2218
rect 6200 2172 6216 2188
rect 6312 2132 6328 2148
rect 6360 2132 6376 2148
rect 6216 2112 6232 2128
rect 6120 2072 6136 2088
rect 6200 2072 6216 2088
rect 6232 2072 6248 2088
rect 6072 1952 6088 1968
rect 6104 1952 6120 1968
rect 5864 1892 5880 1908
rect 5944 1892 5960 1908
rect 5848 1872 5864 1888
rect 5944 1872 5960 1888
rect 5992 1872 6008 1888
rect 5752 1772 5768 1788
rect 5704 1732 5720 1748
rect 5640 1632 5656 1648
rect 5624 1452 5640 1468
rect 5640 1452 5656 1468
rect 5592 1372 5608 1388
rect 5576 1252 5592 1268
rect 5544 1212 5560 1228
rect 5528 1112 5544 1128
rect 5512 1092 5528 1108
rect 5464 932 5480 948
rect 5480 932 5496 948
rect 5512 932 5528 948
rect 5560 1072 5576 1088
rect 5832 1832 5848 1848
rect 5672 1712 5688 1728
rect 5656 1332 5672 1348
rect 5640 1312 5656 1328
rect 5656 1272 5672 1288
rect 5816 1712 5832 1728
rect 5736 1692 5752 1708
rect 5800 1692 5816 1708
rect 5880 1732 5896 1748
rect 5752 1672 5768 1688
rect 5720 1652 5736 1668
rect 5816 1652 5832 1668
rect 5768 1632 5800 1648
rect 5720 1612 5736 1628
rect 5736 1512 5752 1528
rect 5688 1472 5704 1488
rect 5752 1452 5768 1468
rect 5736 1392 5752 1408
rect 5752 1352 5768 1368
rect 5768 1312 5784 1328
rect 5736 1292 5752 1308
rect 5752 1292 5768 1308
rect 5672 1212 5688 1228
rect 5704 1212 5720 1228
rect 5624 1172 5640 1188
rect 5640 1132 5656 1148
rect 5608 1012 5624 1028
rect 5688 1092 5704 1108
rect 5640 952 5656 968
rect 5688 952 5704 968
rect 5560 932 5576 948
rect 5800 1532 5816 1548
rect 6040 1692 6056 1708
rect 5976 1652 5992 1668
rect 5880 1612 5896 1628
rect 5960 1612 5976 1628
rect 5960 1572 5976 1588
rect 5896 1552 5912 1568
rect 5800 1492 5816 1508
rect 5832 1492 5848 1508
rect 5816 1372 5832 1388
rect 5816 1292 5832 1308
rect 5864 1532 5880 1548
rect 6040 1552 6056 1568
rect 5992 1532 6008 1548
rect 6104 1912 6120 1928
rect 6200 1992 6216 2008
rect 6184 1932 6200 1948
rect 6504 2152 6520 2168
rect 6552 2152 6568 2168
rect 6520 2132 6536 2148
rect 6552 2132 6568 2148
rect 6456 2092 6488 2108
rect 6376 2012 6392 2028
rect 6280 1952 6296 1968
rect 6344 1952 6360 1968
rect 6440 1952 6456 1968
rect 6296 1932 6312 1948
rect 6328 1912 6344 1928
rect 6344 1912 6360 1928
rect 6168 1832 6184 1848
rect 6104 1812 6120 1828
rect 6120 1792 6136 1808
rect 6088 1772 6104 1788
rect 6344 1852 6360 1868
rect 6200 1832 6216 1848
rect 6237 1802 6273 1818
rect 6168 1772 6184 1788
rect 6264 1772 6280 1788
rect 6232 1752 6248 1768
rect 6168 1712 6184 1728
rect 6104 1692 6120 1708
rect 6296 1752 6312 1768
rect 6296 1712 6312 1728
rect 6280 1692 6296 1708
rect 6088 1672 6104 1688
rect 6184 1672 6200 1688
rect 6216 1672 6232 1688
rect 6168 1652 6184 1668
rect 6072 1632 6088 1648
rect 6104 1552 6120 1568
rect 6072 1532 6088 1548
rect 5992 1512 6008 1528
rect 6056 1512 6072 1528
rect 5976 1492 5992 1508
rect 5880 1472 5896 1488
rect 5912 1452 5928 1468
rect 5880 1432 5896 1448
rect 5896 1352 5912 1368
rect 5944 1352 5960 1368
rect 5864 1332 5880 1348
rect 5784 1272 5800 1288
rect 5848 1252 5864 1268
rect 5880 1212 5896 1228
rect 5992 1472 6008 1488
rect 5864 1132 5880 1148
rect 5816 1112 5832 1128
rect 5736 1092 5752 1108
rect 5784 1072 5800 1088
rect 5768 1012 5784 1028
rect 5752 952 5768 968
rect 5704 932 5720 948
rect 5528 912 5544 928
rect 5448 892 5464 908
rect 5448 772 5464 788
rect 5432 752 5448 768
rect 5352 692 5368 708
rect 5208 672 5224 688
rect 5352 632 5368 648
rect 5448 632 5464 648
rect 5384 592 5400 608
rect 5432 592 5448 608
rect 5320 572 5336 588
rect 5224 552 5256 568
rect 5384 552 5400 568
rect 5336 532 5352 548
rect 5240 512 5256 528
rect 5320 512 5336 528
rect 5208 492 5224 508
rect 5288 492 5304 508
rect 5213 402 5249 418
rect 5192 272 5208 288
rect 4952 252 4968 268
rect 5000 252 5016 268
rect 4952 132 4968 148
rect 4952 112 4968 128
rect 4856 12 4872 28
rect 4920 12 4952 28
rect 4968 12 4984 28
rect 5048 132 5064 148
rect 5032 92 5048 108
rect 5208 172 5224 188
rect 5080 132 5096 148
rect 5128 112 5144 128
rect 5064 52 5080 68
rect 5096 52 5112 68
rect 5176 52 5192 68
rect 5064 12 5080 28
rect 5112 32 5128 48
rect 5160 32 5176 48
rect 5416 492 5432 508
rect 5368 432 5384 448
rect 5560 812 5576 828
rect 5544 712 5560 728
rect 5576 712 5592 728
rect 5592 692 5608 708
rect 5592 672 5608 688
rect 5512 632 5528 648
rect 5528 612 5544 628
rect 5512 532 5528 548
rect 5464 452 5480 468
rect 5432 312 5448 328
rect 5464 312 5480 328
rect 5336 306 5352 308
rect 5336 292 5352 306
rect 5400 292 5416 308
rect 5416 292 5432 308
rect 5368 252 5384 268
rect 5448 292 5464 308
rect 5448 272 5464 288
rect 5448 132 5464 148
rect 5336 114 5352 128
rect 5336 112 5352 114
rect 5400 112 5416 128
rect 5720 872 5736 888
rect 5960 1172 5976 1188
rect 5912 1112 5928 1128
rect 5896 1072 5912 1088
rect 5960 1092 5976 1108
rect 5880 1052 5896 1068
rect 5928 1032 5944 1048
rect 5992 1012 6008 1028
rect 5976 952 5992 968
rect 5784 932 5800 948
rect 5800 932 5816 948
rect 5848 932 5864 948
rect 5864 932 5880 948
rect 5976 932 5992 948
rect 5800 912 5816 928
rect 5832 912 5848 928
rect 5992 912 6008 928
rect 5656 732 5672 748
rect 5624 712 5640 728
rect 5608 592 5624 608
rect 5704 692 5720 708
rect 5544 532 5560 548
rect 5560 492 5576 508
rect 5576 432 5592 448
rect 5592 352 5608 368
rect 5528 272 5544 288
rect 5496 172 5528 188
rect 5704 592 5720 608
rect 5656 492 5668 508
rect 5668 492 5672 508
rect 5656 372 5672 388
rect 5624 292 5640 308
rect 5576 232 5592 248
rect 5544 172 5560 188
rect 5576 132 5592 148
rect 5592 132 5608 148
rect 5400 92 5416 108
rect 5464 92 5480 108
rect 5192 32 5208 48
rect 5272 32 5288 48
rect 5320 32 5336 48
rect 5400 32 5416 48
rect 5192 12 5208 28
rect 5213 2 5249 18
rect 5304 12 5320 28
rect 5352 12 5368 28
rect 5720 352 5736 368
rect 5784 592 5800 608
rect 5768 572 5784 588
rect 5960 852 5976 868
rect 6040 1492 6056 1508
rect 6088 1492 6104 1508
rect 6120 1352 6136 1368
rect 6088 1312 6104 1328
rect 6104 1292 6120 1308
rect 6152 1292 6168 1308
rect 6024 1212 6040 1228
rect 6024 1172 6040 1188
rect 6072 1152 6088 1168
rect 6040 1112 6056 1128
rect 6024 1072 6040 1088
rect 6040 952 6056 968
rect 6120 1212 6136 1228
rect 6120 1092 6136 1108
rect 6184 1472 6200 1488
rect 6216 1452 6232 1468
rect 6264 1452 6280 1468
rect 6216 1432 6232 1448
rect 6200 1352 6216 1368
rect 6237 1402 6273 1418
rect 6440 1912 6456 1928
rect 6424 1852 6440 1868
rect 6424 1772 6440 1788
rect 6648 2292 6664 2308
rect 6632 2272 6648 2288
rect 6584 2092 6600 2108
rect 6488 1972 6504 1988
rect 6552 1892 6568 1908
rect 6632 2232 6648 2248
rect 6632 2212 6648 2228
rect 6680 2112 6696 2128
rect 6712 2372 6728 2388
rect 6728 2312 6744 2328
rect 6664 2092 6680 2108
rect 6696 2092 6712 2108
rect 6696 2072 6712 2088
rect 6840 2352 6856 2368
rect 6824 2332 6840 2348
rect 6760 2312 6776 2328
rect 6792 2292 6808 2308
rect 7144 3312 7160 3328
rect 7208 3832 7224 3848
rect 7192 3772 7208 3788
rect 7256 3812 7272 3828
rect 7224 3732 7240 3748
rect 7176 3332 7192 3348
rect 7240 3332 7256 3348
rect 7064 3292 7080 3308
rect 7112 3292 7128 3308
rect 7048 3272 7064 3288
rect 7064 3252 7080 3268
rect 7176 3232 7192 3248
rect 7160 3192 7176 3208
rect 7128 3152 7144 3168
rect 7064 3132 7080 3148
rect 7080 3112 7096 3128
rect 7096 3072 7112 3088
rect 7112 2992 7128 3008
rect 7096 2972 7112 2988
rect 7208 3092 7224 3108
rect 7208 3072 7224 3088
rect 7192 2992 7208 3008
rect 7096 2932 7112 2948
rect 7128 2932 7144 2948
rect 7080 2892 7096 2908
rect 7112 2892 7128 2908
rect 7208 2912 7224 2928
rect 7240 2912 7256 2928
rect 7224 2892 7240 2908
rect 7144 2872 7160 2888
rect 7176 2872 7192 2888
rect 7160 2792 7176 2808
rect 7096 2752 7112 2768
rect 7112 2712 7128 2728
rect 7080 2692 7096 2708
rect 7112 2692 7128 2708
rect 7128 2692 7144 2708
rect 7064 2612 7080 2628
rect 7096 2612 7112 2628
rect 7080 2572 7096 2588
rect 7032 2552 7048 2568
rect 7016 2532 7032 2548
rect 6872 2512 6888 2528
rect 6904 2512 6920 2528
rect 6968 2512 6984 2528
rect 6920 2492 6936 2508
rect 6952 2492 6968 2508
rect 6984 2472 7000 2488
rect 6904 2452 6920 2468
rect 6968 2412 6984 2428
rect 6904 2392 6920 2408
rect 6888 2372 6904 2388
rect 7032 2492 7048 2508
rect 7032 2432 7048 2448
rect 7064 2432 7080 2448
rect 6920 2372 6936 2388
rect 6936 2352 6952 2368
rect 6856 2292 6872 2308
rect 6872 2292 6888 2308
rect 6776 2212 6792 2228
rect 6824 2152 6840 2168
rect 6808 2112 6824 2128
rect 6760 2072 6776 2088
rect 6840 2132 6856 2148
rect 6808 2072 6824 2088
rect 6792 2032 6808 2048
rect 6712 1992 6744 2008
rect 6632 1972 6648 1988
rect 6664 1892 6680 1908
rect 6600 1872 6616 1888
rect 6632 1872 6648 1888
rect 6712 1872 6728 1888
rect 6552 1852 6568 1868
rect 6584 1852 6600 1868
rect 6504 1832 6520 1848
rect 6408 1732 6424 1748
rect 6456 1732 6472 1748
rect 6520 1732 6536 1748
rect 6392 1712 6408 1728
rect 6424 1712 6440 1728
rect 6376 1692 6392 1708
rect 6456 1692 6472 1708
rect 6488 1712 6504 1728
rect 6472 1612 6488 1628
rect 6424 1592 6440 1608
rect 6360 1572 6376 1588
rect 6408 1572 6424 1588
rect 6312 1492 6328 1508
rect 6392 1492 6408 1508
rect 6344 1452 6360 1468
rect 6296 1312 6312 1328
rect 6264 1292 6280 1308
rect 6328 1292 6344 1308
rect 6360 1332 6376 1348
rect 6536 1532 6552 1548
rect 6568 1672 6584 1688
rect 6600 1712 6616 1728
rect 6600 1692 6616 1708
rect 6584 1632 6600 1648
rect 6440 1472 6456 1488
rect 6440 1412 6456 1428
rect 6424 1332 6440 1348
rect 6408 1312 6424 1328
rect 6216 1192 6232 1208
rect 6184 1152 6200 1168
rect 6264 1132 6280 1148
rect 6312 1132 6328 1148
rect 6200 1092 6216 1108
rect 6552 1392 6568 1408
rect 6488 1312 6504 1328
rect 6552 1312 6568 1328
rect 6472 1272 6488 1288
rect 6376 1212 6392 1228
rect 6376 1152 6392 1168
rect 6424 1152 6440 1168
rect 6536 1272 6552 1288
rect 6680 1752 6696 1768
rect 6648 1672 6664 1688
rect 6616 1592 6632 1608
rect 6712 1592 6728 1608
rect 6616 1572 6632 1588
rect 6696 1552 6712 1568
rect 6648 1512 6664 1528
rect 6600 1492 6616 1508
rect 6680 1492 6696 1508
rect 6680 1332 6696 1348
rect 6712 1472 6728 1488
rect 6712 1452 6728 1468
rect 6616 1312 6632 1328
rect 6632 1312 6648 1328
rect 6696 1312 6712 1328
rect 6664 1292 6680 1308
rect 6584 1272 6600 1288
rect 6680 1272 6696 1288
rect 6568 1252 6584 1268
rect 6632 1232 6648 1248
rect 6504 1212 6520 1228
rect 6552 1172 6568 1188
rect 6520 1152 6536 1168
rect 6392 1132 6408 1148
rect 6488 1132 6504 1148
rect 6584 1132 6600 1148
rect 6616 1132 6632 1148
rect 6280 1112 6296 1128
rect 6360 1112 6376 1128
rect 6456 1112 6472 1128
rect 6504 1112 6520 1128
rect 6616 1112 6632 1128
rect 6408 1092 6424 1108
rect 6440 1092 6456 1108
rect 6168 1032 6184 1048
rect 6200 1032 6216 1048
rect 6264 1032 6280 1048
rect 6237 1002 6273 1018
rect 6200 932 6216 948
rect 6392 1032 6408 1048
rect 6440 972 6456 988
rect 6424 952 6440 968
rect 6088 912 6104 928
rect 6152 912 6168 928
rect 6184 914 6200 928
rect 6184 912 6200 914
rect 6296 912 6312 928
rect 6680 1112 6696 1128
rect 6568 1092 6584 1108
rect 6632 1092 6648 1108
rect 6504 1052 6520 1068
rect 6568 1052 6584 1068
rect 6584 1032 6600 1048
rect 6552 1012 6568 1028
rect 6568 952 6584 968
rect 6008 812 6024 828
rect 5880 732 5896 748
rect 5976 732 5992 748
rect 6024 712 6036 728
rect 6036 712 6040 728
rect 6008 692 6024 708
rect 5928 672 5944 688
rect 5960 672 5976 688
rect 5848 592 5864 608
rect 6088 692 6104 708
rect 5976 552 5992 568
rect 6072 532 6088 548
rect 5832 492 5848 508
rect 5976 492 5992 508
rect 6040 492 6056 508
rect 5800 432 5816 448
rect 5704 332 5720 348
rect 5736 332 5752 348
rect 5688 312 5704 328
rect 5672 292 5688 308
rect 5816 332 5832 348
rect 5672 272 5688 288
rect 5800 272 5816 288
rect 6344 752 6360 768
rect 6120 732 6136 748
rect 6232 712 6248 728
rect 6312 712 6328 728
rect 6120 692 6136 708
rect 6088 512 6120 528
rect 6280 672 6296 688
rect 6237 602 6273 618
rect 6392 732 6408 748
rect 6392 712 6408 728
rect 6424 712 6440 728
rect 6504 932 6520 948
rect 6488 912 6504 928
rect 6456 892 6472 908
rect 6568 732 6584 748
rect 6376 692 6392 708
rect 6424 692 6440 708
rect 6440 692 6456 708
rect 6136 572 6152 588
rect 6168 552 6184 568
rect 6120 492 6136 508
rect 6136 492 6152 508
rect 6200 492 6216 508
rect 6104 472 6120 488
rect 6072 352 6088 368
rect 6008 312 6024 328
rect 5832 292 5848 308
rect 5928 292 5944 308
rect 5976 292 6008 308
rect 5912 272 5928 288
rect 6232 452 6248 468
rect 6296 472 6328 488
rect 6280 432 6296 448
rect 6296 332 6312 348
rect 6280 312 6296 328
rect 6168 292 6184 308
rect 6024 272 6040 288
rect 6136 272 6152 288
rect 6168 272 6184 288
rect 6312 272 6328 288
rect 5880 252 5896 268
rect 5832 132 5848 148
rect 5768 112 5784 128
rect 5816 112 5832 128
rect 5816 92 5832 108
rect 5992 92 6008 108
rect 5736 32 5752 48
rect 6088 252 6104 268
rect 6152 252 6168 268
rect 6120 172 6136 188
rect 6136 132 6152 148
rect 6237 202 6273 218
rect 6184 152 6200 168
rect 6248 152 6264 168
rect 6200 132 6216 148
rect 6168 112 6184 128
rect 6168 92 6184 108
rect 6264 12 6280 28
rect 6376 552 6392 568
rect 6360 512 6376 528
rect 6360 492 6376 508
rect 6456 552 6472 568
rect 6440 532 6456 548
rect 6584 512 6600 528
rect 6392 472 6408 488
rect 6424 472 6440 488
rect 6424 352 6440 368
rect 6376 312 6392 328
rect 6344 292 6360 308
rect 6392 292 6408 308
rect 6456 332 6472 348
rect 6520 312 6536 328
rect 6440 272 6456 288
rect 6376 252 6392 268
rect 6408 92 6424 108
rect 6488 252 6504 268
rect 6568 212 6584 228
rect 6504 172 6520 188
rect 6536 152 6552 168
rect 6504 132 6520 148
rect 6824 1992 6840 2008
rect 6904 2112 6920 2128
rect 6872 2092 6888 2108
rect 6904 2052 6920 2068
rect 6888 1992 6904 2008
rect 6840 1952 6856 1968
rect 6744 1912 6760 1928
rect 6776 1912 6792 1928
rect 6792 1892 6808 1908
rect 6872 1912 6888 1928
rect 6808 1872 6824 1888
rect 6744 1852 6760 1868
rect 6872 1832 6888 1848
rect 6904 1772 6920 1788
rect 6840 1732 6856 1748
rect 6760 1712 6776 1728
rect 6808 1632 6824 1648
rect 6856 1632 6872 1648
rect 6872 1572 6888 1588
rect 6776 1512 6792 1528
rect 6904 1512 6920 1528
rect 6824 1492 6840 1508
rect 6792 1472 6808 1488
rect 7032 2332 7048 2348
rect 7176 2672 7192 2688
rect 7176 2652 7192 2668
rect 7160 2572 7176 2588
rect 7144 2552 7160 2568
rect 7112 2512 7128 2528
rect 7096 2492 7112 2508
rect 7096 2472 7112 2488
rect 7128 2452 7144 2468
rect 7096 2372 7112 2388
rect 6952 2292 6968 2308
rect 6968 2292 6984 2308
rect 6952 2112 6968 2128
rect 7048 2312 7064 2328
rect 7080 2312 7096 2328
rect 7096 2272 7112 2288
rect 7000 2212 7016 2228
rect 7064 2212 7080 2228
rect 6984 2092 7000 2108
rect 6952 2072 6968 2088
rect 7016 2112 7032 2128
rect 7112 2112 7128 2128
rect 7064 2092 7080 2108
rect 7112 2092 7128 2108
rect 7160 2392 7176 2408
rect 7144 2352 7160 2368
rect 7208 2772 7224 2788
rect 7272 3792 7288 3808
rect 7352 5052 7368 5068
rect 7352 4992 7368 5008
rect 7336 4492 7352 4508
rect 7384 5072 7400 5088
rect 7400 5052 7416 5068
rect 7416 4932 7432 4948
rect 7432 4692 7448 4708
rect 7400 4632 7416 4648
rect 7400 4532 7416 4548
rect 7400 4472 7416 4488
rect 7336 4452 7352 4468
rect 7368 4452 7384 4468
rect 7368 4432 7384 4448
rect 7384 4332 7400 4348
rect 7368 4052 7384 4068
rect 7352 4032 7368 4048
rect 7336 3912 7352 3928
rect 7304 3812 7320 3828
rect 7336 3812 7352 3828
rect 7384 3812 7400 3828
rect 7352 3772 7368 3788
rect 7368 3712 7384 3728
rect 7352 3692 7368 3708
rect 7288 3612 7304 3628
rect 7272 3392 7288 3408
rect 7336 3392 7352 3408
rect 7272 3312 7304 3328
rect 7336 3312 7352 3328
rect 7352 3212 7368 3228
rect 7336 3092 7352 3108
rect 7400 3732 7416 3748
rect 7384 3452 7400 3468
rect 7384 3332 7400 3348
rect 7336 3072 7352 3088
rect 7304 2892 7320 2908
rect 7288 2772 7304 2788
rect 7240 2692 7256 2708
rect 7288 2672 7304 2688
rect 7208 2632 7224 2648
rect 7240 2572 7256 2588
rect 7336 2912 7352 2928
rect 7336 2892 7352 2908
rect 7320 2612 7336 2628
rect 7304 2572 7320 2588
rect 7272 2512 7288 2528
rect 7256 2472 7272 2488
rect 7240 2452 7256 2468
rect 7224 2432 7240 2448
rect 7288 2372 7304 2388
rect 7192 2332 7208 2348
rect 7272 2312 7288 2328
rect 7224 2292 7240 2308
rect 7208 2252 7224 2268
rect 7240 2132 7256 2148
rect 7144 2112 7160 2128
rect 7144 2092 7160 2108
rect 7048 2072 7064 2088
rect 6968 2052 6984 2068
rect 7032 2052 7048 2068
rect 7064 2052 7080 2068
rect 7032 1952 7048 1968
rect 7080 1992 7112 2008
rect 7064 1912 7080 1928
rect 7128 1952 7144 1968
rect 7176 2032 7192 2048
rect 7160 1992 7192 2008
rect 7048 1892 7064 1908
rect 7160 1892 7176 1908
rect 6936 1872 6952 1888
rect 7000 1852 7016 1868
rect 7272 1912 7288 1928
rect 7224 1892 7240 1908
rect 7160 1832 7192 1848
rect 7064 1772 7080 1788
rect 7016 1752 7032 1768
rect 6936 1732 6952 1748
rect 6984 1732 7000 1748
rect 6968 1712 6984 1728
rect 7000 1692 7016 1708
rect 7016 1532 7032 1548
rect 7016 1492 7032 1508
rect 6920 1452 6936 1468
rect 6744 1432 6760 1448
rect 6776 1432 6792 1448
rect 6824 1432 6840 1448
rect 6744 1412 6760 1428
rect 6744 1352 6760 1368
rect 6744 1332 6760 1348
rect 6792 1392 6808 1408
rect 6936 1372 6952 1388
rect 6856 1332 6872 1348
rect 6904 1332 6920 1348
rect 6728 1292 6744 1308
rect 6840 1292 6856 1308
rect 6808 1272 6824 1288
rect 6760 1252 6776 1268
rect 6664 1032 6680 1048
rect 6744 1012 6760 1028
rect 6680 992 6696 1008
rect 6840 1132 6856 1148
rect 6888 1232 6904 1248
rect 6904 1172 6920 1188
rect 6936 1332 6952 1348
rect 6952 1312 6968 1328
rect 6920 1152 6936 1168
rect 6936 1132 6952 1148
rect 6792 1112 6796 1128
rect 6796 1112 6808 1128
rect 6872 1112 6888 1128
rect 6888 1092 6904 1108
rect 6952 1092 6968 1108
rect 6824 1072 6840 1088
rect 6840 1032 6856 1048
rect 6808 992 6824 1008
rect 6744 972 6760 988
rect 6904 972 6920 988
rect 6936 972 6952 988
rect 6968 972 6984 988
rect 6632 952 6648 968
rect 6776 952 6792 968
rect 7048 1572 7064 1588
rect 7128 1632 7144 1648
rect 7144 1572 7160 1588
rect 7048 1552 7064 1568
rect 7096 1552 7112 1568
rect 7112 1532 7128 1548
rect 7096 1512 7112 1528
rect 7080 1492 7096 1508
rect 7128 1492 7144 1508
rect 7032 1452 7048 1468
rect 7080 1452 7096 1468
rect 7064 1392 7080 1408
rect 7080 1372 7096 1388
rect 7064 1272 7080 1288
rect 7000 1192 7016 1208
rect 7016 1112 7032 1128
rect 7032 1092 7048 1108
rect 7064 1092 7080 1108
rect 7032 1012 7048 1028
rect 7096 1012 7112 1028
rect 6984 952 7000 968
rect 6984 932 7000 948
rect 7000 932 7016 948
rect 6888 912 6904 928
rect 6968 912 6984 928
rect 7000 912 7016 928
rect 6744 872 6760 888
rect 6728 812 6744 828
rect 6696 732 6712 748
rect 6680 692 6696 708
rect 6648 672 6664 688
rect 6680 532 6696 548
rect 6600 492 6632 508
rect 6680 492 6696 508
rect 6648 332 6664 348
rect 6664 292 6680 308
rect 6760 712 6776 728
rect 6776 672 6792 688
rect 6744 532 6760 548
rect 7064 992 7080 1008
rect 6888 732 6920 748
rect 7032 712 7048 728
rect 7016 672 7032 688
rect 6904 652 6920 668
rect 7032 632 7048 648
rect 7144 1372 7160 1388
rect 7128 1352 7144 1368
rect 7208 1812 7224 1828
rect 7256 1812 7272 1828
rect 7240 1772 7256 1788
rect 7304 2292 7320 2308
rect 7384 2912 7400 2928
rect 7400 2872 7416 2888
rect 7368 2772 7384 2788
rect 7368 2452 7384 2468
rect 7384 2412 7400 2428
rect 7384 2392 7400 2408
rect 7304 2192 7320 2208
rect 7304 2172 7320 2188
rect 7416 2352 7432 2368
rect 7352 2312 7368 2328
rect 7384 2192 7400 2208
rect 7400 2172 7416 2188
rect 7368 1972 7384 1988
rect 7352 1952 7368 1968
rect 7320 1932 7336 1948
rect 7336 1912 7352 1928
rect 7304 1892 7320 1908
rect 7304 1732 7320 1748
rect 7416 1992 7432 2008
rect 7384 1892 7400 1908
rect 7368 1752 7384 1768
rect 7416 1752 7432 1768
rect 7176 1712 7192 1728
rect 7272 1712 7288 1728
rect 7256 1692 7272 1708
rect 7176 1672 7192 1688
rect 7208 1632 7224 1648
rect 7384 1732 7400 1748
rect 7416 1732 7432 1748
rect 7384 1712 7400 1728
rect 7352 1672 7368 1688
rect 7272 1592 7288 1608
rect 7224 1512 7240 1528
rect 7352 1512 7368 1528
rect 7336 1492 7352 1508
rect 7352 1492 7368 1508
rect 7384 1492 7400 1508
rect 7208 1472 7224 1488
rect 7368 1472 7384 1488
rect 7176 1392 7192 1408
rect 7192 1352 7208 1368
rect 7224 1392 7240 1408
rect 7336 1452 7352 1468
rect 7368 1452 7384 1468
rect 7400 1272 7416 1288
rect 7192 1172 7208 1188
rect 7224 1172 7240 1188
rect 7192 1152 7208 1168
rect 7128 1112 7144 1128
rect 7160 1112 7176 1128
rect 7368 1112 7384 1128
rect 7128 1092 7144 1108
rect 7192 1092 7208 1108
rect 7256 1092 7272 1108
rect 7336 1092 7352 1108
rect 7384 1092 7400 1108
rect 7144 1072 7160 1088
rect 7112 972 7128 988
rect 7112 912 7128 928
rect 7080 852 7096 868
rect 7096 732 7112 748
rect 7144 712 7160 728
rect 7128 692 7144 708
rect 7320 1072 7336 1088
rect 7208 1052 7224 1068
rect 7272 1052 7288 1068
rect 7224 1012 7240 1028
rect 7288 992 7304 1008
rect 7240 972 7256 988
rect 7304 972 7320 988
rect 7400 972 7416 988
rect 7304 952 7320 968
rect 7224 932 7240 948
rect 7224 912 7240 928
rect 7208 892 7224 908
rect 7352 892 7368 908
rect 7384 792 7400 808
rect 7176 692 7192 708
rect 7176 652 7192 668
rect 7160 552 7176 568
rect 7128 532 7144 548
rect 6712 312 6728 328
rect 6696 292 6712 308
rect 6808 472 6824 488
rect 6808 452 6824 468
rect 6824 412 6840 428
rect 7000 512 7016 528
rect 7048 512 7064 528
rect 7112 512 7128 528
rect 6968 492 6984 508
rect 7016 492 7032 508
rect 7032 492 7048 508
rect 7080 492 7096 508
rect 7112 492 7128 508
rect 7144 472 7160 488
rect 7064 452 7080 468
rect 6984 312 7000 328
rect 7032 312 7048 328
rect 6872 292 6888 308
rect 6920 292 6936 308
rect 6952 292 6968 308
rect 6872 272 6888 288
rect 6808 152 6824 168
rect 6744 132 6760 148
rect 6936 232 6952 248
rect 7032 292 7048 308
rect 7000 232 7016 248
rect 6952 212 6968 228
rect 7016 212 7032 228
rect 6968 152 6984 168
rect 6600 112 6616 128
rect 6648 112 6664 128
rect 6648 92 6664 108
rect 6824 92 6840 108
rect 6568 32 6584 48
rect 7128 192 7144 208
rect 7288 672 7304 688
rect 7192 612 7208 628
rect 7192 572 7208 588
rect 7256 632 7272 648
rect 7224 572 7240 588
rect 7208 532 7224 548
rect 7432 552 7448 568
rect 7320 512 7336 528
rect 7432 512 7448 528
rect 7208 312 7224 328
rect 7176 292 7192 308
rect 7304 492 7320 508
rect 7288 472 7304 488
rect 7288 312 7304 328
rect 7320 292 7336 308
rect 7368 292 7384 308
rect 7192 272 7208 288
rect 7384 272 7400 288
rect 7336 212 7352 228
rect 7144 172 7160 188
rect 7384 172 7400 188
rect 7224 152 7240 168
rect 7176 132 7192 148
rect 7192 132 7208 148
rect 6936 112 6952 128
rect 7032 112 7048 128
rect 7256 114 7272 128
rect 7256 112 7272 114
rect 6904 12 6920 28
<< metal3 >>
rect 3064 5417 3080 5423
rect 3128 5417 3160 5423
rect 3912 5417 3928 5423
rect 3080 5397 3128 5403
rect 4808 5397 4840 5403
rect 5368 5397 5432 5403
rect 120 5377 296 5383
rect 392 5377 664 5383
rect 680 5377 856 5383
rect 1960 5377 2056 5383
rect 2072 5377 2424 5383
rect 3208 5377 3384 5383
rect 3592 5377 3640 5383
rect 3656 5377 3800 5383
rect 4376 5377 4552 5383
rect 4584 5377 4632 5383
rect 4648 5377 5064 5383
rect 6696 5377 6936 5383
rect 1288 5357 1400 5363
rect 1416 5357 1512 5363
rect 3528 5357 5528 5363
rect 5544 5357 5576 5363
rect 6136 5357 6200 5363
rect 6216 5357 6392 5363
rect 7213 5357 7224 5363
rect 40 5337 56 5343
rect 840 5337 1032 5343
rect 1064 5337 1320 5343
rect 1400 5337 1496 5343
rect 1688 5337 1736 5343
rect 1848 5337 1992 5343
rect 2376 5337 2616 5343
rect 3016 5337 3512 5343
rect 3544 5337 3592 5343
rect 3640 5337 3928 5343
rect 3944 5337 4696 5343
rect 4712 5337 4744 5343
rect 4856 5337 5064 5343
rect 5208 5337 5448 5343
rect 6024 5337 6136 5343
rect 6376 5337 6584 5343
rect 6600 5337 6648 5343
rect 6664 5337 6744 5343
rect 6824 5337 6904 5343
rect 7128 5337 7208 5343
rect 7069 5328 7075 5332
rect 56 5317 184 5323
rect 248 5317 520 5323
rect 536 5317 600 5323
rect 808 5317 872 5323
rect 904 5317 936 5323
rect 1160 5317 1208 5323
rect 1224 5317 1288 5323
rect 1448 5317 1480 5323
rect 1976 5317 2296 5323
rect 2424 5317 2472 5323
rect 2488 5317 2504 5323
rect 3448 5317 3480 5323
rect 3576 5317 3784 5323
rect 3848 5317 3960 5323
rect 3976 5317 4072 5323
rect 4328 5317 4424 5323
rect 4600 5317 4664 5323
rect 4792 5317 4824 5323
rect 5192 5317 5288 5323
rect 5656 5317 5832 5323
rect 6120 5317 6536 5323
rect 6856 5317 6872 5323
rect 7112 5317 7224 5323
rect 24 5297 88 5303
rect 664 5297 760 5303
rect 776 5297 1064 5303
rect 1336 5297 1368 5303
rect 1384 5297 1448 5303
rect 1496 5297 1624 5303
rect 1720 5297 1832 5303
rect 1928 5297 2120 5303
rect 2136 5297 2568 5303
rect 2824 5297 2872 5303
rect 2888 5297 3880 5303
rect 4136 5297 4328 5303
rect 4504 5297 4600 5303
rect 4664 5297 4744 5303
rect 4824 5297 4904 5303
rect 5512 5297 5608 5303
rect 5624 5297 5656 5303
rect 5672 5297 5944 5303
rect 5960 5297 5992 5303
rect 6008 5297 6056 5303
rect 6072 5297 6120 5303
rect 7064 5297 7144 5303
rect 1448 5277 1976 5283
rect 1992 5277 2024 5283
rect 2184 5277 2392 5283
rect 3320 5277 3432 5283
rect 3496 5277 3592 5283
rect 3608 5277 3768 5283
rect 4728 5277 5144 5283
rect 5208 5277 5576 5283
rect 6904 5277 6968 5283
rect 6984 5277 7128 5283
rect 968 5257 1960 5263
rect 4008 5257 4776 5263
rect 4984 5257 5112 5263
rect 5368 5257 5752 5263
rect 2760 5237 2984 5243
rect 3000 5237 3384 5243
rect 3736 5237 3752 5243
rect 3928 5237 4216 5243
rect 4536 5237 4968 5243
rect 7176 5237 7304 5243
rect 1464 5217 2312 5223
rect 2328 5217 2360 5223
rect 2376 5217 2584 5223
rect 1416 5197 1464 5203
rect 1480 5197 1496 5203
rect 1512 5197 2712 5203
rect 5464 5217 6056 5223
rect 5261 5197 7272 5203
rect 2296 5177 2488 5183
rect 5261 5183 5267 5197
rect 3544 5177 5267 5183
rect 5624 5177 5688 5183
rect 504 5157 680 5163
rect 4584 5157 5912 5163
rect 5928 5157 6120 5163
rect 296 5137 408 5143
rect 536 5137 568 5143
rect 584 5137 728 5143
rect 744 5137 776 5143
rect 1080 5137 1704 5143
rect 2472 5137 2536 5143
rect 4072 5137 4392 5143
rect 4504 5137 4888 5143
rect 5656 5137 5832 5143
rect 7336 5137 7352 5143
rect 392 5117 488 5123
rect 632 5117 648 5123
rect 664 5117 840 5123
rect 1192 5117 1368 5123
rect 1624 5117 1720 5123
rect 1816 5117 1848 5123
rect 2312 5117 2440 5123
rect 2456 5117 2840 5123
rect 3368 5117 3656 5123
rect 3672 5117 3736 5123
rect 4376 5117 4504 5123
rect 4760 5117 4824 5123
rect 4984 5117 5048 5123
rect 5608 5117 6008 5123
rect 6024 5117 6072 5123
rect 6088 5117 6120 5123
rect 6520 5117 7192 5123
rect 7208 5117 7320 5123
rect 408 5097 616 5103
rect 792 5097 904 5103
rect 1352 5097 1384 5103
rect 1400 5097 1704 5103
rect 1720 5097 1752 5103
rect 1864 5097 1960 5103
rect 2184 5097 2248 5103
rect 2472 5097 2504 5103
rect 2600 5097 2632 5103
rect 2904 5097 2984 5103
rect 3960 5097 3976 5103
rect 4344 5097 4360 5103
rect 4376 5097 4440 5103
rect 4456 5097 4472 5103
rect 4840 5097 4856 5103
rect 4888 5097 4920 5103
rect 4936 5097 4968 5103
rect 5128 5097 5224 5103
rect 5240 5097 5320 5103
rect 5496 5097 5528 5103
rect 5592 5097 5720 5103
rect 5816 5097 5960 5103
rect 6024 5097 6280 5103
rect 6296 5097 6536 5103
rect 6888 5097 6968 5103
rect 6984 5097 7144 5103
rect 7208 5097 7304 5103
rect 3693 5088 3699 5092
rect 408 5077 504 5083
rect 616 5077 632 5083
rect 744 5077 904 5083
rect 1048 5077 1128 5083
rect 1144 5077 1544 5083
rect 1560 5077 1704 5083
rect 1992 5077 2392 5083
rect 2520 5077 2728 5083
rect 2776 5077 2968 5083
rect 4248 5077 4328 5083
rect 4344 5077 4376 5083
rect 4536 5077 4568 5083
rect 5000 5077 5192 5083
rect 5400 5077 5480 5083
rect 6040 5077 6051 5083
rect 3117 5068 3123 5072
rect 4797 5068 4803 5072
rect 6045 5068 6051 5077
rect 6120 5077 6328 5083
rect 6456 5077 6488 5083
rect 6520 5077 6824 5083
rect 7144 5077 7176 5083
rect 7192 5077 7304 5083
rect 7320 5077 7384 5083
rect 632 5057 808 5063
rect 1656 5057 1784 5063
rect 1800 5057 1880 5063
rect 1896 5057 2088 5063
rect 2104 5057 2376 5063
rect 2664 5057 3032 5063
rect 3224 5057 3736 5063
rect 3752 5057 4312 5063
rect 4440 5057 4648 5063
rect 6488 5057 6568 5063
rect 6920 5057 7016 5063
rect 7032 5057 7096 5063
rect 7256 5057 7288 5063
rect 7368 5057 7400 5063
rect 424 5037 456 5043
rect 472 5037 632 5043
rect 728 5037 776 5043
rect 824 5037 968 5043
rect 984 5037 1000 5043
rect 1496 5037 1544 5043
rect 1560 5037 1672 5043
rect 1896 5037 2072 5043
rect 2152 5037 2328 5043
rect 2552 5037 2808 5043
rect 2824 5037 2840 5043
rect 3128 5037 3304 5043
rect 4200 5037 4216 5043
rect 4520 5037 4536 5043
rect 4792 5037 5080 5043
rect 5272 5037 5448 5043
rect 5672 5037 6616 5043
rect 6632 5037 6968 5043
rect 7048 5037 7160 5043
rect 376 5017 2008 5023
rect 2232 5017 2456 5023
rect 2616 5017 2680 5023
rect 2712 5017 2744 5023
rect 3032 5017 3368 5023
rect 2392 4997 2952 5003
rect 3048 4997 3656 5003
rect 5096 5017 5656 5023
rect 5736 5017 5848 5023
rect 4392 4997 4696 5003
rect 4712 4997 4840 5003
rect 5325 4997 5816 5003
rect 88 4977 232 4983
rect 776 4977 840 4983
rect 1272 4977 1352 4983
rect 1688 4977 1864 4983
rect 1880 4977 2008 4983
rect 2088 4977 2376 4983
rect 2440 4977 2456 4983
rect 2568 4977 2600 4983
rect 5325 4983 5331 4997
rect 5832 4997 5928 5003
rect 6424 5017 6696 5023
rect 6493 4997 7192 5003
rect 3512 4977 5331 4983
rect 5432 4977 5480 4983
rect 5496 4977 5672 4983
rect 5704 4977 5912 4983
rect 6493 4983 6499 4997
rect 7304 4997 7352 5003
rect 5944 4977 6499 4983
rect 6584 4977 6712 4983
rect 6840 4977 6952 4983
rect 6968 4977 7032 4983
rect 7048 4977 7208 4983
rect 24 4957 72 4963
rect 296 4957 456 4963
rect 2328 4957 2664 4963
rect 2680 4957 2904 4963
rect 2920 4957 3224 4963
rect 3432 4957 3496 4963
rect 3560 4957 3832 4963
rect 3848 4957 3880 4963
rect 3992 4957 4168 4963
rect 4616 4957 4792 4963
rect 4888 4957 5000 4963
rect 5432 4957 5640 4963
rect 5848 4957 5944 4963
rect 6152 4957 6280 4963
rect 216 4937 296 4943
rect 312 4937 504 4943
rect 520 4937 536 4943
rect 696 4937 808 4943
rect 1160 4937 1400 4943
rect 1960 4937 2232 4943
rect 2360 4937 2424 4943
rect 2728 4937 3064 4943
rect 3288 4937 3432 4943
rect 3528 4937 3560 4943
rect 3832 4937 3896 4943
rect 3912 4937 4088 4943
rect 4109 4937 4200 4943
rect 4109 4928 4115 4937
rect 4312 4937 4696 4943
rect 4824 4937 4872 4943
rect 5000 4937 5448 4943
rect 5656 4937 6040 4943
rect 6232 4937 6488 4943
rect 6504 4937 6536 4943
rect 6712 4937 6760 4943
rect 6776 4937 7416 4943
rect 6221 4928 6227 4932
rect 88 4917 104 4923
rect 200 4917 792 4923
rect 824 4917 952 4923
rect 968 4917 1192 4923
rect 1208 4917 1272 4923
rect 1288 4917 1560 4923
rect 1592 4917 1656 4923
rect 2008 4917 2056 4923
rect 2072 4917 2120 4923
rect 2408 4917 2456 4923
rect 2872 4917 2920 4923
rect 2936 4917 3096 4923
rect 3176 4917 3608 4923
rect 3752 4917 3784 4923
rect 3880 4917 3976 4923
rect 4216 4917 4280 4923
rect 4328 4917 4472 4923
rect 4744 4917 4840 4923
rect 5048 4917 5352 4923
rect 5368 4917 5400 4923
rect 5880 4917 5912 4923
rect 5928 4917 6168 4923
rect 6184 4917 6216 4923
rect 6280 4917 6472 4923
rect 6488 4917 6504 4923
rect 6760 4917 6936 4923
rect 7176 4917 7272 4923
rect 40 4897 136 4903
rect 152 4897 184 4903
rect 456 4897 504 4903
rect 952 4897 1432 4903
rect 1624 4897 1752 4903
rect 2088 4897 2360 4903
rect 2376 4897 2392 4903
rect 2408 4897 2472 4903
rect 2488 4897 2584 4903
rect 2600 4897 2792 4903
rect 3096 4897 3112 4903
rect 3448 4897 3480 4903
rect 3496 4897 3592 4903
rect 3608 4897 3640 4903
rect 4056 4897 4232 4903
rect 4376 4897 4408 4903
rect 4424 4897 4456 4903
rect 4840 4897 4856 4903
rect 4872 4897 4920 4903
rect 5048 4897 5208 4903
rect 5416 4897 5480 4903
rect 5912 4897 6024 4903
rect 6216 4897 6392 4903
rect 6664 4897 6680 4903
rect 6696 4897 6808 4903
rect 6824 4897 6872 4903
rect 6888 4897 7032 4903
rect 904 4877 1880 4883
rect 1896 4877 1944 4883
rect 2120 4877 2296 4883
rect 2312 4877 2872 4883
rect 3000 4877 3912 4883
rect 3944 4877 4344 4883
rect 5080 4877 5896 4883
rect 5912 4877 6360 4883
rect 6680 4877 6856 4883
rect 7000 4877 7096 4883
rect 1416 4857 1480 4863
rect 3112 4857 3224 4863
rect 3704 4857 3720 4863
rect 3928 4857 5496 4863
rect 5560 4857 6232 4863
rect 6248 4857 6840 4863
rect 6952 4857 7000 4863
rect 792 4837 872 4843
rect 888 4837 1592 4843
rect 1608 4837 1768 4843
rect 1784 4837 1816 4843
rect 3352 4837 3384 4843
rect 3416 4837 4568 4843
rect 4584 4837 4728 4843
rect 5544 4837 5752 4843
rect 5768 4837 5800 4843
rect 5816 4837 5944 4843
rect 5960 4837 6440 4843
rect 6648 4837 6664 4843
rect 6744 4837 6984 4843
rect 7192 4837 7240 4843
rect 72 4797 1016 4803
rect 1032 4797 1096 4803
rect 1256 4817 1272 4823
rect 1288 4817 1416 4823
rect 2552 4817 2728 4823
rect 2744 4817 2776 4823
rect 1165 4797 2696 4803
rect 1165 4783 1171 4797
rect 3688 4817 3720 4823
rect 4424 4817 4488 4823
rect 3512 4797 3544 4803
rect 4504 4797 4536 4803
rect 5272 4817 6136 4823
rect 6248 4817 6696 4823
rect 6184 4797 6552 4803
rect 6696 4797 6792 4803
rect 584 4777 1171 4783
rect 2952 4777 3400 4783
rect 3656 4777 3848 4783
rect 4776 4777 5544 4783
rect 5608 4777 5672 4783
rect 5864 4777 6408 4783
rect 6456 4777 6616 4783
rect 6632 4777 6728 4783
rect 6792 4777 6968 4783
rect 680 4757 1288 4763
rect 1512 4757 1608 4763
rect 2024 4757 2600 4763
rect 2696 4757 3208 4763
rect 3432 4757 3544 4763
rect 5144 4757 5368 4763
rect 5416 4757 5832 4763
rect 5992 4757 6584 4763
rect 6952 4757 6984 4763
rect 7016 4757 7128 4763
rect 872 4737 968 4743
rect 984 4737 1032 4743
rect 1480 4737 2536 4743
rect 2808 4737 3112 4743
rect 3629 4737 3640 4743
rect 3704 4737 3768 4743
rect 5336 4737 5400 4743
rect 5464 4737 5560 4743
rect 5672 4737 5752 4743
rect 5784 4737 5816 4743
rect 5880 4737 6152 4743
rect 6504 4737 6616 4743
rect 6632 4737 7064 4743
rect 4461 4728 4467 4732
rect 152 4717 264 4723
rect 648 4717 888 4723
rect 904 4717 936 4723
rect 952 4717 1576 4723
rect 1832 4717 1928 4723
rect 1976 4717 2024 4723
rect 2136 4717 2264 4723
rect 2424 4717 2488 4723
rect 2568 4717 2680 4723
rect 2824 4717 2840 4723
rect 3112 4717 3320 4723
rect 3384 4717 3395 4723
rect 4216 4717 4227 4723
rect 4680 4717 4808 4723
rect 4824 4717 5000 4723
rect 5032 4717 5208 4723
rect 5272 4717 5352 4723
rect 5400 4717 5688 4723
rect 6120 4717 6472 4723
rect 6664 4717 6792 4723
rect 6824 4717 6856 4723
rect 6888 4717 7048 4723
rect 7144 4717 7491 4723
rect 3709 4708 3715 4712
rect 4429 4708 4435 4712
rect 248 4697 280 4703
rect 296 4697 504 4703
rect 584 4697 648 4703
rect 760 4697 904 4703
rect 952 4697 984 4703
rect 1096 4697 1208 4703
rect 1320 4697 1336 4703
rect 1496 4697 1528 4703
rect 1544 4697 1576 4703
rect 1704 4697 1864 4703
rect 1912 4697 1960 4703
rect 2024 4697 2056 4703
rect 2120 4697 2248 4703
rect 2328 4697 2440 4703
rect 2536 4697 2808 4703
rect 3144 4697 3208 4703
rect 3224 4697 3272 4703
rect 3464 4697 3624 4703
rect 3768 4697 3880 4703
rect 4904 4697 5048 4703
rect 5320 4697 5384 4703
rect 5469 4697 5480 4703
rect 5576 4697 5608 4703
rect 5768 4697 5832 4703
rect 6072 4697 6136 4703
rect 6312 4697 6424 4703
rect 6440 4697 6552 4703
rect 6824 4697 6936 4703
rect 6952 4697 6984 4703
rect 7016 4697 7128 4703
rect 7320 4697 7432 4703
rect 1357 4688 1363 4692
rect 3725 4688 3731 4692
rect 4525 4688 4531 4692
rect 392 4677 568 4683
rect 1240 4677 1304 4683
rect 1432 4677 1448 4683
rect 1576 4677 1720 4683
rect 1896 4677 2344 4683
rect 2376 4677 2552 4683
rect 2584 4677 2760 4683
rect 2888 4677 3576 4683
rect 4856 4677 4904 4683
rect 5192 4677 5512 4683
rect 5896 4677 5960 4683
rect 6232 4677 6376 4683
rect 6584 4677 6632 4683
rect 6648 4677 6696 4683
rect 6728 4677 7000 4683
rect 2573 4668 2579 4672
rect 24 4657 200 4663
rect 440 4657 696 4663
rect 904 4657 952 4663
rect 1000 4657 1208 4663
rect 1240 4657 1304 4663
rect 1336 4657 1368 4663
rect 1480 4657 1491 4663
rect 2392 4657 2472 4663
rect 2504 4657 2536 4663
rect 2648 4657 2675 4663
rect 104 4637 312 4643
rect 504 4637 664 4643
rect 680 4637 776 4643
rect 1016 4637 1384 4643
rect 1944 4637 2648 4643
rect 2669 4643 2675 4657
rect 2696 4657 3240 4663
rect 3288 4657 3496 4663
rect 3512 4657 3576 4663
rect 3704 4657 3720 4663
rect 4456 4657 4744 4663
rect 4840 4657 5000 4663
rect 5208 4657 5288 4663
rect 5304 4657 5608 4663
rect 5624 4657 5928 4663
rect 5976 4657 6088 4663
rect 6168 4657 6504 4663
rect 6776 4657 6808 4663
rect 7048 4657 7080 4663
rect 2669 4637 2872 4643
rect 2952 4637 3032 4643
rect 3048 4637 3096 4643
rect 3112 4637 3272 4643
rect 3432 4637 4408 4643
rect 4472 4637 5960 4643
rect 5992 4637 6216 4643
rect 6728 4637 6920 4643
rect 6936 4637 7208 4643
rect 7224 4637 7400 4643
rect 1000 4617 1048 4623
rect 1368 4617 1384 4623
rect 1768 4617 1800 4623
rect 1816 4617 2136 4623
rect 24 4597 520 4603
rect 536 4597 792 4603
rect 1032 4597 1240 4603
rect 1256 4597 1368 4603
rect 1416 4597 1560 4603
rect 2520 4617 2616 4623
rect 2888 4617 2952 4623
rect 3240 4617 3816 4623
rect 2936 4597 3064 4603
rect 4312 4617 4536 4623
rect 4552 4617 4584 4623
rect 4792 4617 5128 4623
rect 5176 4617 5320 4623
rect 5336 4617 5368 4623
rect 5400 4617 5448 4623
rect 5496 4617 5544 4623
rect 5560 4617 5624 4623
rect 5816 4617 6120 4623
rect 4264 4597 4376 4603
rect 4424 4597 5960 4603
rect 6600 4617 6760 4623
rect 6776 4617 6824 4623
rect 6840 4617 7144 4623
rect 6296 4597 6872 4603
rect 120 4577 296 4583
rect 312 4577 328 4583
rect 600 4577 696 4583
rect 1208 4577 1256 4583
rect 1384 4577 1496 4583
rect 1672 4577 2056 4583
rect 2077 4583 2083 4592
rect 2077 4577 2088 4583
rect 2152 4577 2232 4583
rect 2456 4577 2776 4583
rect 3048 4577 3224 4583
rect 3240 4577 3448 4583
rect 3576 4577 3672 4583
rect 3752 4577 4083 4583
rect 1032 4557 1144 4563
rect 1176 4557 1912 4563
rect 1928 4557 1944 4563
rect 1960 4557 2552 4563
rect 2568 4557 2616 4563
rect 2760 4557 2824 4563
rect 3016 4557 3064 4563
rect 3992 4557 4056 4563
rect 4077 4563 4083 4577
rect 4696 4577 4760 4583
rect 4888 4577 5448 4583
rect 5480 4577 5576 4583
rect 5832 4577 5880 4583
rect 6136 4577 6408 4583
rect 6600 4577 6792 4583
rect 4077 4557 5032 4563
rect 5208 4557 5256 4563
rect 5320 4557 5416 4563
rect 5512 4557 5560 4563
rect 5592 4557 5656 4563
rect 5768 4557 6184 4563
rect 6328 4557 6616 4563
rect 6712 4557 6744 4563
rect 6808 4557 6952 4563
rect 7144 4557 7272 4563
rect 488 4537 632 4543
rect 680 4537 728 4543
rect 872 4537 1128 4543
rect 1144 4537 1224 4543
rect 1336 4537 1384 4543
rect 1496 4537 1720 4543
rect 2184 4537 2232 4543
rect 2312 4537 2344 4543
rect 2456 4537 2488 4543
rect 2568 4537 2584 4543
rect 2696 4537 2760 4543
rect 3272 4537 3288 4543
rect 3432 4537 3656 4543
rect 4056 4537 4120 4543
rect 4296 4537 4344 4543
rect 4456 4537 4568 4543
rect 4584 4537 4792 4543
rect 4808 4537 4824 4543
rect 4952 4537 5528 4543
rect 5544 4537 5864 4543
rect 5880 4537 6040 4543
rect 6088 4537 6200 4543
rect 6472 4537 6664 4543
rect 6760 4537 6984 4543
rect 7144 4537 7400 4543
rect 88 4517 168 4523
rect 248 4517 424 4523
rect 632 4517 664 4523
rect 712 4517 728 4523
rect 856 4517 872 4523
rect 1016 4517 1032 4523
rect 1064 4517 1192 4523
rect 1288 4517 1320 4523
rect 1352 4517 1416 4523
rect 1432 4517 1704 4523
rect 1720 4517 2456 4523
rect 2472 4517 2616 4523
rect 2632 4517 2760 4523
rect 3016 4517 3096 4523
rect 3304 4517 3336 4523
rect 3560 4517 3784 4523
rect 3848 4517 4072 4523
rect 4184 4517 4360 4523
rect 4392 4517 4408 4523
rect 4632 4517 4664 4523
rect 4765 4517 4776 4523
rect 4808 4517 4872 4523
rect 4936 4517 5464 4523
rect 5480 4517 5800 4523
rect 5832 4517 5848 4523
rect 5976 4517 6088 4523
rect 6392 4517 6472 4523
rect 6536 4517 6616 4523
rect 6648 4517 6808 4523
rect 6968 4517 7064 4523
rect 893 4508 899 4512
rect 40 4497 72 4503
rect 728 4497 888 4503
rect 952 4497 968 4503
rect 984 4497 1032 4503
rect 1144 4497 1464 4503
rect 1848 4497 1976 4503
rect 2008 4497 2088 4503
rect 2104 4497 2184 4503
rect 2216 4497 2328 4503
rect 2392 4497 2520 4503
rect 2584 4497 2664 4503
rect 2968 4497 3000 4503
rect 3320 4497 3496 4503
rect 3704 4497 3715 4503
rect 3709 4488 3715 4497
rect 3736 4497 3944 4503
rect 4072 4497 4408 4503
rect 4504 4497 4632 4503
rect 5224 4497 5384 4503
rect 5400 4497 5832 4503
rect 5928 4497 6200 4503
rect 6456 4497 6504 4503
rect 6536 4497 6632 4503
rect 6728 4497 6739 4503
rect 6920 4497 7080 4503
rect 7288 4497 7336 4503
rect 7448 4497 7491 4503
rect 568 4477 776 4483
rect 952 4477 984 4483
rect 1000 4477 1080 4483
rect 1096 4477 1672 4483
rect 1688 4477 2472 4483
rect 3896 4477 4056 4483
rect 4136 4477 4184 4483
rect 4200 4477 4616 4483
rect 4888 4477 5128 4483
rect 5160 4477 5304 4483
rect 5352 4477 5400 4483
rect 5784 4477 5816 4483
rect 5944 4477 6056 4483
rect 6072 4477 6088 4483
rect 6200 4477 6328 4483
rect 6408 4477 6504 4483
rect 6685 4483 6691 4492
rect 6584 4477 6840 4483
rect 6888 4477 6920 4483
rect 6936 4477 7160 4483
rect 7176 4477 7400 4483
rect 392 4457 904 4463
rect 920 4457 952 4463
rect 1048 4457 1800 4463
rect 1864 4457 2088 4463
rect 2184 4457 2392 4463
rect 2472 4457 2536 4463
rect 3208 4457 3448 4463
rect 3752 4457 4712 4463
rect 5000 4457 5208 4463
rect 5240 4457 5368 4463
rect 5400 4457 5480 4463
rect 5864 4457 6120 4463
rect 6184 4457 6280 4463
rect 6648 4457 6680 4463
rect 7352 4457 7368 4463
rect 776 4437 2072 4443
rect 2136 4437 2200 4443
rect 2856 4437 2888 4443
rect 2904 4437 2920 4443
rect 3352 4437 3752 4443
rect 3912 4437 4184 4443
rect 4200 4437 4824 4443
rect 5064 4437 6344 4443
rect 6728 4437 6808 4443
rect 7224 4437 7368 4443
rect 1272 4417 1352 4423
rect 1560 4417 1704 4423
rect 1720 4417 1784 4423
rect 1368 4397 1528 4403
rect 1544 4397 1656 4403
rect 1672 4397 2312 4403
rect 2344 4397 2824 4403
rect 2840 4397 3128 4403
rect 3416 4417 3432 4423
rect 3480 4417 3992 4423
rect 4008 4417 4104 4423
rect 3453 4397 3576 4403
rect 1304 4377 1368 4383
rect 1848 4377 2248 4383
rect 2264 4377 2424 4383
rect 3453 4383 3459 4397
rect 3592 4397 3656 4403
rect 5448 4417 5512 4423
rect 5528 4417 6232 4423
rect 6248 4417 6328 4423
rect 6360 4417 7032 4423
rect 5336 4397 5512 4403
rect 5992 4397 6115 4403
rect 2440 4377 3459 4383
rect 4392 4377 4584 4383
rect 4824 4377 5128 4383
rect 5320 4377 5784 4383
rect 5912 4377 6035 4383
rect 376 4357 856 4363
rect 1064 4357 1256 4363
rect 1880 4357 2440 4363
rect 2600 4357 3464 4363
rect 3656 4357 3720 4363
rect 3736 4357 4264 4363
rect 4280 4357 4344 4363
rect 4360 4357 4440 4363
rect 4456 4357 4536 4363
rect 4552 4357 4744 4363
rect 4856 4357 5048 4363
rect 5864 4357 5960 4363
rect 5976 4357 6008 4363
rect 6029 4363 6035 4377
rect 6109 4383 6115 4397
rect 6152 4397 6296 4403
rect 6568 4397 6648 4403
rect 7016 4397 7160 4403
rect 6056 4377 6099 4383
rect 6109 4377 6760 4383
rect 6029 4357 6056 4363
rect 6093 4363 6099 4377
rect 6093 4357 6264 4363
rect 6696 4357 6792 4363
rect 7064 4357 7080 4363
rect 600 4337 696 4343
rect 712 4337 808 4343
rect 840 4337 1816 4343
rect 2232 4337 2264 4343
rect 3464 4337 3560 4343
rect 3880 4337 4584 4343
rect 4696 4337 4840 4343
rect 5021 4337 5032 4343
rect 5512 4337 5560 4343
rect 5896 4337 6136 4343
rect 6184 4337 6200 4343
rect 6232 4337 6360 4343
rect 6440 4337 6648 4343
rect 6664 4337 6712 4343
rect 6744 4337 6776 4343
rect 6808 4337 6920 4343
rect 6936 4337 6968 4343
rect 7048 4337 7112 4343
rect 7336 4337 7384 4343
rect 24 4317 72 4323
rect 88 4317 216 4323
rect 536 4317 728 4323
rect 904 4317 952 4323
rect 1000 4317 1080 4323
rect 1112 4317 1176 4323
rect 1192 4317 1336 4323
rect 1352 4317 1448 4323
rect 1544 4317 1560 4323
rect 1592 4317 1672 4323
rect 1720 4317 1912 4323
rect 2088 4317 2216 4323
rect 2472 4317 2600 4323
rect 3048 4317 3144 4323
rect 3352 4317 3480 4323
rect 3608 4317 3619 4323
rect 4216 4317 4424 4323
rect 4440 4317 4504 4323
rect 4856 4317 4936 4323
rect 5096 4317 5160 4323
rect 5544 4317 5688 4323
rect 5704 4317 6024 4323
rect 6056 4317 6104 4323
rect 6136 4317 6184 4323
rect 6296 4317 6408 4323
rect 6424 4317 6456 4323
rect 6888 4317 7000 4323
rect 7069 4317 7192 4323
rect 765 4308 771 4312
rect 88 4297 168 4303
rect 328 4297 360 4303
rect 488 4297 632 4303
rect 728 4297 760 4303
rect 872 4297 984 4303
rect 1048 4297 1160 4303
rect 1192 4297 1544 4303
rect 1560 4297 1608 4303
rect 1688 4297 1944 4303
rect 2200 4297 2328 4303
rect 2376 4297 2584 4303
rect 2728 4297 2808 4303
rect 3016 4297 3064 4303
rect 3080 4297 3112 4303
rect 3496 4297 3512 4303
rect 3720 4297 3832 4303
rect 3864 4297 4120 4303
rect 4136 4297 4168 4303
rect 4424 4297 4840 4303
rect 4872 4297 5080 4303
rect 5096 4297 5384 4303
rect 5800 4297 6152 4303
rect 6216 4297 6344 4303
rect 6408 4297 6568 4303
rect 6808 4297 6888 4303
rect 7069 4303 7075 4317
rect 7208 4317 7491 4323
rect 6952 4297 7075 4303
rect 7096 4297 7112 4303
rect 7144 4297 7208 4303
rect 4125 4288 4131 4292
rect 632 4277 664 4283
rect 680 4277 808 4283
rect 856 4277 904 4283
rect 920 4277 1016 4283
rect 1080 4277 1160 4283
rect 1176 4277 1208 4283
rect 1256 4277 1288 4283
rect 1320 4277 1432 4283
rect 1448 4277 1608 4283
rect 1624 4277 2184 4283
rect 2200 4277 2360 4283
rect 2504 4277 2664 4283
rect 2680 4277 2856 4283
rect 2920 4277 3064 4283
rect 3128 4277 3480 4283
rect 3640 4277 3704 4283
rect 3800 4277 3960 4283
rect 4184 4277 4296 4283
rect 4440 4277 4451 4283
rect 4728 4277 4808 4283
rect 4984 4277 5032 4283
rect 5048 4277 5320 4283
rect 5336 4277 5816 4283
rect 5848 4277 5896 4283
rect 6056 4277 6312 4283
rect 6344 4277 6424 4283
rect 6440 4277 6648 4283
rect 6840 4277 7112 4283
rect 7128 4277 7176 4283
rect 7240 4277 7272 4283
rect 13 4268 19 4272
rect 616 4257 1352 4263
rect 1368 4257 1736 4263
rect 1864 4257 1912 4263
rect 2104 4257 3048 4263
rect 4024 4257 4264 4263
rect 4888 4257 4936 4263
rect 5896 4257 5976 4263
rect 6104 4257 6200 4263
rect 6232 4257 6440 4263
rect 6872 4257 7032 4263
rect 7048 4257 7080 4263
rect 120 4237 296 4243
rect 312 4237 840 4243
rect 904 4237 1016 4243
rect 1240 4237 1512 4243
rect 1736 4237 2248 4243
rect 2264 4237 2504 4243
rect 2520 4237 2664 4243
rect 3144 4237 3736 4243
rect 3768 4237 3800 4243
rect 3816 4237 4008 4243
rect 4568 4237 4792 4243
rect 4824 4237 5416 4243
rect 5816 4237 6360 4243
rect 6760 4237 7128 4243
rect 408 4217 1864 4223
rect 1896 4217 2008 4223
rect 888 4197 1016 4203
rect 1272 4197 1720 4203
rect 1752 4197 2056 4203
rect 2328 4217 2568 4223
rect 3064 4217 3400 4223
rect 3528 4217 3928 4223
rect 2232 4197 2392 4203
rect 2760 4197 3608 4203
rect 3656 4197 4104 4203
rect 4280 4217 4520 4223
rect 4536 4217 4984 4223
rect 5096 4217 5144 4223
rect 5416 4217 5496 4223
rect 5512 4217 5624 4223
rect 5640 4217 5672 4223
rect 5880 4217 5896 4223
rect 5960 4217 6216 4223
rect 5368 4197 5496 4203
rect 5864 4197 6168 4203
rect 6296 4217 6408 4223
rect 6536 4217 6728 4223
rect 6744 4217 6920 4223
rect 6936 4217 6968 4223
rect 7048 4217 7160 4223
rect 7224 4217 7256 4223
rect 6424 4197 6520 4203
rect 200 4177 296 4183
rect 376 4177 440 4183
rect 456 4177 888 4183
rect 904 4177 1144 4183
rect 1160 4177 1896 4183
rect 2024 4177 2264 4183
rect 2280 4177 2408 4183
rect 2968 4177 3160 4183
rect 3336 4177 3400 4183
rect 3656 4177 3768 4183
rect 3992 4177 4248 4183
rect 4344 4177 4680 4183
rect 4696 4177 4872 4183
rect 4904 4177 6072 4183
rect 6104 4177 6424 4183
rect 6472 4177 6616 4183
rect 6632 4177 6904 4183
rect 6920 4177 7160 4183
rect 1016 4157 1048 4163
rect 1208 4157 1688 4163
rect 1800 4157 1912 4163
rect 1944 4157 1960 4163
rect 1976 4157 2152 4163
rect 2312 4157 2456 4163
rect 2792 4157 3000 4163
rect 3272 4157 3640 4163
rect 3736 4157 3976 4163
rect 4488 4157 5160 4163
rect 5384 4157 5416 4163
rect 5528 4157 5576 4163
rect 6088 4157 6264 4163
rect 6296 4157 6536 4163
rect 6552 4157 6712 4163
rect 6984 4157 7128 4163
rect 7144 4157 7192 4163
rect 104 4137 232 4143
rect 1048 4137 1192 4143
rect 1208 4137 1368 4143
rect 1704 4137 1768 4143
rect 1976 4137 2056 4143
rect 2072 4137 2200 4143
rect 2376 4137 2568 4143
rect 2584 4137 2712 4143
rect 2840 4137 2872 4143
rect 2888 4137 2952 4143
rect 3144 4137 3336 4143
rect 3624 4137 3688 4143
rect 3704 4137 4024 4143
rect 4040 4137 4152 4143
rect 4296 4137 4344 4143
rect 4408 4137 4456 4143
rect 4632 4137 4952 4143
rect 4984 4137 5016 4143
rect 5112 4137 5208 4143
rect 5224 4137 5352 4143
rect 5384 4137 5400 4143
rect 5528 4137 5624 4143
rect 5640 4137 5704 4143
rect 5720 4137 5992 4143
rect 6072 4137 6264 4143
rect 6440 4137 6552 4143
rect 6600 4137 6648 4143
rect 1821 4128 1827 4132
rect 232 4117 264 4123
rect 504 4117 568 4123
rect 776 4117 984 4123
rect 1144 4117 1155 4123
rect 1149 4108 1155 4117
rect 1176 4117 1288 4123
rect 1480 4117 1624 4123
rect 1912 4117 1976 4123
rect 2104 4117 2136 4123
rect 2488 4117 2499 4123
rect 2493 4108 2499 4117
rect 2664 4117 2696 4123
rect 2952 4117 3128 4123
rect 3144 4117 3352 4123
rect 3368 4117 3432 4123
rect 3464 4117 3560 4123
rect 3608 4117 3656 4123
rect 3864 4117 4136 4123
rect 4152 4117 4536 4123
rect 4568 4117 4584 4123
rect 4824 4117 4904 4123
rect 5080 4117 5288 4123
rect 5320 4117 5448 4123
rect 5720 4117 5752 4123
rect 5864 4117 5912 4123
rect 5928 4117 6184 4123
rect 6216 4117 6344 4123
rect 6616 4117 6664 4123
rect 7032 4117 7080 4123
rect 1608 4097 1624 4103
rect 1640 4097 1672 4103
rect 1928 4097 2280 4103
rect 2616 4097 2632 4103
rect 2648 4097 2792 4103
rect 2808 4097 2840 4103
rect 2856 4097 2920 4103
rect 3224 4097 3352 4103
rect 3560 4097 3624 4103
rect 3672 4097 3864 4103
rect 3928 4097 3976 4103
rect 4040 4097 4120 4103
rect 4136 4097 4280 4103
rect 4440 4097 4552 4103
rect 4616 4097 4696 4103
rect 4856 4097 4904 4103
rect 5208 4097 5544 4103
rect 6072 4097 6584 4103
rect 6605 4097 6840 4103
rect 397 4088 403 4092
rect 925 4088 931 4092
rect 4413 4088 4419 4092
rect 1080 4077 1640 4083
rect 2152 4077 2312 4083
rect 2440 4077 2616 4083
rect 2904 4077 2984 4083
rect 3528 4077 3656 4083
rect 3864 4077 4088 4083
rect 5032 4077 5432 4083
rect 5448 4077 5752 4083
rect 6605 4083 6611 4097
rect 7032 4097 7491 4103
rect 6216 4077 6611 4083
rect 6632 4077 6760 4083
rect 6776 4077 7032 4083
rect 40 4057 200 4063
rect 216 4057 2792 4063
rect 3352 4057 3608 4063
rect 3640 4057 3720 4063
rect 4120 4057 5128 4063
rect 5256 4057 5400 4063
rect 5480 4057 5528 4063
rect 5544 4057 5608 4063
rect 5656 4057 5784 4063
rect 6120 4057 6488 4063
rect 6552 4057 7112 4063
rect 616 4037 856 4043
rect 872 4037 2120 4043
rect 2168 4037 2280 4043
rect 2552 4037 3736 4043
rect 3768 4037 3832 4043
rect 3848 4037 3944 4043
rect 3960 4037 4440 4043
rect 4472 4037 4664 4043
rect 5016 4037 5064 4043
rect 6104 4037 6632 4043
rect 6648 4037 7352 4043
rect 344 3997 408 4003
rect 424 3997 456 4003
rect 2056 4017 2360 4023
rect 2440 4017 2760 4023
rect 3800 4017 3864 4023
rect 3880 4017 3928 4023
rect 3944 4017 4472 4023
rect 4216 3997 4456 4003
rect 4504 3997 4520 4003
rect 6232 4017 6296 4023
rect 6456 4017 6600 4023
rect 6088 3997 6776 4003
rect 6888 3997 6968 4003
rect 7000 3997 7016 4003
rect 40 3977 536 3983
rect 552 3977 584 3983
rect 600 3977 728 3983
rect 1960 3977 2648 3983
rect 3288 3977 3320 3983
rect 3640 3977 3928 3983
rect 3944 3977 4408 3983
rect 4696 3977 4840 3983
rect 5608 3977 6088 3983
rect 6184 3977 6216 3983
rect 6344 3977 6520 3983
rect 6536 3977 6584 3983
rect 6616 3977 7016 3983
rect 4525 3968 4531 3972
rect 1032 3957 1464 3963
rect 1480 3957 1512 3963
rect 2312 3957 2600 3963
rect 2616 3957 2632 3963
rect 4024 3957 4056 3963
rect 4072 3957 4168 3963
rect 4360 3957 4440 3963
rect 4856 3957 5128 3963
rect 5448 3957 5528 3963
rect 5800 3957 6456 3963
rect 6824 3957 6936 3963
rect 6984 3957 7000 3963
rect 824 3937 1016 3943
rect 1032 3937 1064 3943
rect 1144 3937 1320 3943
rect 1464 3937 1864 3943
rect 1949 3937 2088 3943
rect 936 3917 968 3923
rect 984 3917 1064 3923
rect 1080 3917 1208 3923
rect 1949 3923 1955 3937
rect 2232 3937 2744 3943
rect 2776 3937 3960 3943
rect 3992 3937 4296 3943
rect 4328 3937 4392 3943
rect 4440 3937 4520 3943
rect 4760 3937 4920 3943
rect 5080 3937 5560 3943
rect 6088 3937 6120 3943
rect 6136 3937 6152 3943
rect 6360 3937 6632 3943
rect 6760 3937 6792 3943
rect 7016 3937 7048 3943
rect 1464 3917 1955 3923
rect 2984 3917 3112 3923
rect 3576 3917 3848 3923
rect 3864 3917 3912 3923
rect 4104 3917 4280 3923
rect 4296 3917 4424 3923
rect 4616 3917 4627 3923
rect 4728 3917 4792 3923
rect 4840 3917 5032 3923
rect 5464 3917 5624 3923
rect 5736 3917 5832 3923
rect 6680 3917 7064 3923
rect 7080 3917 7096 3923
rect 7144 3917 7176 3923
rect 7192 3917 7336 3923
rect 1965 3908 1971 3912
rect 2349 3908 2355 3912
rect 216 3897 280 3903
rect 392 3897 424 3903
rect 456 3897 488 3903
rect 600 3897 744 3903
rect 984 3897 1048 3903
rect 1080 3897 1192 3903
rect 1416 3897 1432 3903
rect 1448 3897 1544 3903
rect 1816 3897 1912 3903
rect 2168 3897 2312 3903
rect 2360 3897 2456 3903
rect 2536 3897 2712 3903
rect 3128 3897 3160 3903
rect 3688 3897 3784 3903
rect 4072 3897 4168 3903
rect 4328 3897 4344 3903
rect 4456 3897 4728 3903
rect 5368 3897 5384 3903
rect 5416 3897 5432 3903
rect 5816 3897 5848 3903
rect 5976 3897 6120 3903
rect 6296 3897 6392 3903
rect 6600 3897 6744 3903
rect 6760 3897 6872 3903
rect 6952 3897 7048 3903
rect 7064 3897 7080 3903
rect 509 3888 515 3892
rect 3101 3888 3107 3892
rect 4877 3888 4883 3892
rect 5517 3888 5523 3892
rect 104 3877 200 3883
rect 360 3877 392 3883
rect 536 3877 632 3883
rect 920 3877 984 3883
rect 1000 3877 1160 3883
rect 1512 3877 1640 3883
rect 1976 3877 2024 3883
rect 2173 3877 2424 3883
rect 696 3857 888 3863
rect 968 3857 1368 3863
rect 2173 3863 2179 3877
rect 3256 3877 3512 3883
rect 3528 3877 3560 3883
rect 3816 3877 3832 3883
rect 4264 3877 4552 3883
rect 4616 3877 4632 3883
rect 4696 3877 4728 3883
rect 5208 3877 5304 3883
rect 5336 3877 5496 3883
rect 5704 3877 5912 3883
rect 6120 3877 6216 3883
rect 6632 3877 6808 3883
rect 7048 3877 7096 3883
rect 7112 3877 7160 3883
rect 1400 3857 2179 3863
rect 2200 3857 2211 3863
rect 2440 3857 2536 3863
rect 2600 3857 2696 3863
rect 3480 3857 3992 3863
rect 4232 3857 4264 3863
rect 4280 3857 4488 3863
rect 4552 3857 4595 3863
rect 200 3837 296 3843
rect 632 3837 872 3843
rect 888 3837 984 3843
rect 1720 3837 2024 3843
rect 2104 3837 2264 3843
rect 3096 3837 3192 3843
rect 3208 3837 3288 3843
rect 3528 3837 3656 3843
rect 3672 3837 3736 3843
rect 3752 3837 3896 3843
rect 4424 3837 4568 3843
rect 4589 3843 4595 3857
rect 4664 3857 5512 3863
rect 5608 3857 5864 3863
rect 6776 3857 7032 3863
rect 4589 3837 4888 3843
rect 5432 3837 5816 3843
rect 6584 3837 6632 3843
rect 6648 3837 6680 3843
rect 6744 3837 6760 3843
rect 6904 3837 6952 3843
rect 6968 3837 7208 3843
rect 7224 3837 7416 3843
rect 1016 3817 1528 3823
rect 1544 3817 1816 3823
rect 1912 3817 2088 3823
rect 264 3797 1000 3803
rect 1272 3797 1544 3803
rect 1864 3797 2088 3803
rect 2264 3817 2520 3823
rect 2584 3817 3448 3823
rect 3704 3817 3992 3823
rect 2568 3797 3352 3803
rect 3736 3797 3848 3803
rect 4344 3817 4536 3823
rect 4552 3817 4584 3823
rect 4856 3817 4968 3823
rect 5336 3817 5400 3823
rect 5416 3817 5800 3823
rect 4584 3797 4872 3803
rect 4904 3797 5704 3803
rect 5896 3797 6088 3803
rect 6616 3817 6856 3823
rect 7272 3817 7304 3823
rect 7352 3817 7384 3823
rect 6504 3797 6616 3803
rect 6648 3797 6952 3803
rect 7160 3797 7272 3803
rect 312 3777 504 3783
rect 920 3777 1064 3783
rect 1976 3777 2104 3783
rect 2136 3777 2376 3783
rect 2872 3777 2888 3783
rect 3048 3777 3144 3783
rect 3912 3777 4104 3783
rect 4120 3777 4264 3783
rect 4280 3777 4376 3783
rect 4984 3777 5784 3783
rect 5800 3777 6200 3783
rect 6216 3777 7192 3783
rect 7208 3777 7352 3783
rect 184 3757 456 3763
rect 1208 3757 1496 3763
rect 1544 3757 1624 3763
rect 2568 3757 2776 3763
rect 3016 3757 3320 3763
rect 3352 3757 3384 3763
rect 3544 3757 3560 3763
rect 3656 3757 3672 3763
rect 3768 3757 3784 3763
rect 3960 3757 4280 3763
rect 4296 3757 4344 3763
rect 4600 3757 4776 3763
rect 5512 3757 5576 3763
rect 5832 3757 5976 3763
rect 6136 3757 6232 3763
rect 6472 3757 6536 3763
rect 6904 3757 6968 3763
rect 2797 3748 2803 3752
rect 7405 3748 7411 3752
rect 264 3737 312 3743
rect 376 3737 408 3743
rect 808 3737 904 3743
rect 1656 3737 1752 3743
rect 2040 3737 2200 3743
rect 2936 3737 3048 3743
rect 3304 3737 3752 3743
rect 3768 3737 3912 3743
rect 4040 3737 4088 3743
rect 4168 3737 4696 3743
rect 5304 3737 5512 3743
rect 5576 3737 5592 3743
rect 5656 3737 5704 3743
rect 5832 3737 5896 3743
rect 5912 3737 6104 3743
rect 6184 3737 6696 3743
rect 7144 3737 7224 3743
rect 152 3717 200 3723
rect 296 3717 536 3723
rect 728 3717 808 3723
rect 920 3717 1032 3723
rect 1064 3717 1112 3723
rect 1128 3717 1336 3723
rect 1448 3717 1480 3723
rect 1544 3717 1560 3723
rect 1912 3717 1960 3723
rect 2264 3717 2408 3723
rect 2536 3717 2568 3723
rect 2792 3717 2808 3723
rect 2824 3717 3080 3723
rect 3336 3717 3416 3723
rect 3464 3717 3528 3723
rect 3544 3717 3640 3723
rect 3912 3717 3944 3723
rect 3965 3717 4152 3723
rect 40 3697 200 3703
rect 696 3697 920 3703
rect 952 3697 1016 3703
rect 1032 3697 1096 3703
rect 1112 3697 1288 3703
rect 2408 3697 2424 3703
rect 2680 3697 2808 3703
rect 3064 3697 3128 3703
rect 3336 3697 3624 3703
rect 3965 3703 3971 3717
rect 4184 3717 4312 3723
rect 4344 3717 4424 3723
rect 4616 3717 4712 3723
rect 5160 3717 5352 3723
rect 5448 3717 5896 3723
rect 6168 3717 6696 3723
rect 6712 3717 6728 3723
rect 6872 3717 6936 3723
rect 6952 3717 7368 3723
rect 3880 3697 3971 3703
rect 4008 3697 4248 3703
rect 4472 3697 4504 3703
rect 4536 3697 5016 3703
rect 5272 3697 5336 3703
rect 5352 3697 5368 3703
rect 5384 3697 5416 3703
rect 5672 3697 5896 3703
rect 6072 3697 6168 3703
rect 6280 3697 6408 3703
rect 6936 3697 7048 3703
rect 381 3688 387 3692
rect 184 3677 264 3683
rect 904 3677 968 3683
rect 1096 3677 1592 3683
rect 1608 3677 1672 3683
rect 2376 3677 2488 3683
rect 2632 3677 3336 3683
rect 3672 3677 3928 3683
rect 4088 3677 4152 3683
rect 4296 3677 4376 3683
rect 4648 3677 4936 3683
rect 4984 3677 6184 3683
rect 6264 3677 6376 3683
rect 6424 3677 6584 3683
rect 568 3657 1240 3663
rect 1352 3657 1752 3663
rect 3400 3657 3704 3663
rect 3880 3657 5000 3663
rect 5464 3657 5656 3663
rect 5672 3657 6008 3663
rect 6024 3657 6200 3663
rect 6232 3657 6440 3663
rect 24 3637 56 3643
rect 72 3637 328 3643
rect 984 3637 1544 3643
rect 1624 3637 2104 3643
rect 3112 3637 3256 3643
rect 3560 3637 3768 3643
rect 3784 3637 4072 3643
rect 4088 3637 4296 3643
rect 4360 3637 4408 3643
rect 4424 3637 4984 3643
rect 5240 3637 5448 3643
rect 5464 3637 5688 3643
rect 5736 3637 5800 3643
rect 200 3617 424 3623
rect 1544 3617 3128 3623
rect 1832 3597 3144 3603
rect 3560 3617 3576 3623
rect 3720 3617 3768 3623
rect 3848 3617 3896 3623
rect 3912 3617 4328 3623
rect 4360 3617 4632 3623
rect 4664 3617 4696 3623
rect 4760 3617 5000 3623
rect 5032 3617 5112 3623
rect 3608 3597 3832 3603
rect 4072 3597 4360 3603
rect 4840 3597 5176 3603
rect 5352 3617 5368 3623
rect 5400 3617 6152 3623
rect 6200 3617 6760 3623
rect 6776 3617 6840 3623
rect 7304 3617 7384 3623
rect 5608 3597 5816 3603
rect 6184 3597 6264 3603
rect 6680 3597 6936 3603
rect 6968 3597 6984 3603
rect 1448 3577 3432 3583
rect 3448 3577 3800 3583
rect 3832 3577 3896 3583
rect 3960 3577 4136 3583
rect 4216 3577 4296 3583
rect 4376 3577 4824 3583
rect 5224 3577 5304 3583
rect 5512 3577 5704 3583
rect 7485 3583 7491 3603
rect 5768 3577 7491 3583
rect 824 3557 1000 3563
rect 1208 3557 1384 3563
rect 2680 3557 3000 3563
rect 3240 3557 3576 3563
rect 3944 3557 4056 3563
rect 4152 3557 4296 3563
rect 4376 3557 4472 3563
rect 4488 3557 4856 3563
rect 5848 3557 6232 3563
rect 6952 3557 7048 3563
rect 7160 3557 7491 3563
rect 136 3537 264 3543
rect 1112 3537 1160 3543
rect 1176 3537 1352 3543
rect 1448 3537 1656 3543
rect 2024 3537 2056 3543
rect 2072 3537 2328 3543
rect 2952 3537 3016 3543
rect 3176 3537 3272 3543
rect 3320 3537 3384 3543
rect 3469 3537 3768 3543
rect 152 3517 200 3523
rect 312 3517 584 3523
rect 856 3517 936 3523
rect 1400 3517 1448 3523
rect 1576 3517 1672 3523
rect 1944 3517 2072 3523
rect 2264 3517 2328 3523
rect 3469 3523 3475 3537
rect 3784 3537 3832 3543
rect 3864 3537 3896 3543
rect 4008 3537 4024 3543
rect 4040 3537 4168 3543
rect 4280 3537 4312 3543
rect 4717 3537 4728 3543
rect 4904 3537 4952 3543
rect 5720 3537 5768 3543
rect 5800 3537 5912 3543
rect 5928 3537 6152 3543
rect 6216 3537 6312 3543
rect 6360 3537 6552 3543
rect 6600 3537 6760 3543
rect 6776 3537 7000 3543
rect 2392 3517 3475 3523
rect 3496 3517 3512 3523
rect 3832 3517 3880 3523
rect 4056 3517 4088 3523
rect 4184 3517 4280 3523
rect 4312 3517 4488 3523
rect 4504 3517 4584 3523
rect 4872 3517 4904 3523
rect 5000 3517 5064 3523
rect 5176 3517 5592 3523
rect 5736 3517 5752 3523
rect 5784 3517 6280 3523
rect 6376 3517 6472 3523
rect 6840 3517 6952 3523
rect 6968 3517 7064 3523
rect 7128 3517 7491 3523
rect 6557 3508 6563 3512
rect 40 3497 88 3503
rect 104 3497 152 3503
rect 440 3497 456 3503
rect 616 3497 792 3503
rect 808 3497 856 3503
rect 1304 3497 1384 3503
rect 1496 3497 1560 3503
rect 1608 3497 1640 3503
rect 1656 3497 1832 3503
rect 2088 3497 2120 3503
rect 2168 3497 2296 3503
rect 2328 3497 2392 3503
rect 2488 3497 2616 3503
rect 2712 3497 2792 3503
rect 3032 3497 3464 3503
rect 3496 3497 3640 3503
rect 3688 3497 3784 3503
rect 3800 3497 3992 3503
rect 4168 3497 4248 3503
rect 4456 3497 4504 3503
rect 4536 3497 4728 3503
rect 4744 3497 4808 3503
rect 4952 3497 5000 3503
rect 5016 3497 5032 3503
rect 5112 3497 5144 3503
rect 5160 3497 5320 3503
rect 5528 3497 5736 3503
rect 6168 3497 6392 3503
rect 6408 3497 6504 3503
rect 6840 3497 6856 3503
rect 7032 3497 7080 3503
rect 24 3477 72 3483
rect 88 3477 136 3483
rect 312 3477 360 3483
rect 376 3477 552 3483
rect 1464 3477 1656 3483
rect 1688 3477 1784 3483
rect 2056 3477 2152 3483
rect 2312 3477 2344 3483
rect 2456 3477 2680 3483
rect 2696 3477 2936 3483
rect 2968 3477 3096 3483
rect 3320 3477 3352 3483
rect 3544 3477 3736 3483
rect 3928 3477 4328 3483
rect 4344 3477 4376 3483
rect 4536 3477 4568 3483
rect 4664 3477 4771 3483
rect 253 3468 259 3472
rect 472 3457 488 3463
rect 776 3457 920 3463
rect 936 3457 1320 3463
rect 1336 3457 1352 3463
rect 1992 3457 2104 3463
rect 2120 3457 2424 3463
rect 2824 3457 3608 3463
rect 3784 3457 3944 3463
rect 4488 3457 4744 3463
rect 4765 3463 4771 3477
rect 5336 3477 6200 3483
rect 6552 3477 6632 3483
rect 6792 3477 7112 3483
rect 4765 3457 5107 3463
rect 1768 3437 2216 3443
rect 2568 3437 2584 3443
rect 2904 3437 3032 3443
rect 3048 3437 3336 3443
rect 3416 3437 3816 3443
rect 3912 3437 3928 3443
rect 3944 3437 4104 3443
rect 4120 3437 4168 3443
rect 4184 3437 4264 3443
rect 4296 3437 5080 3443
rect 5101 3443 5107 3457
rect 5304 3457 5352 3463
rect 5368 3457 5416 3463
rect 5496 3457 5528 3463
rect 5656 3457 5768 3463
rect 6248 3457 6360 3463
rect 6376 3457 6536 3463
rect 6600 3457 6632 3463
rect 7000 3457 7384 3463
rect 5101 3437 6648 3443
rect 6728 3437 7144 3443
rect 216 3417 296 3423
rect 392 3417 440 3423
rect 568 3417 776 3423
rect 792 3417 856 3423
rect 872 3417 936 3423
rect 984 3417 1128 3423
rect 1144 3417 1224 3423
rect 1240 3417 1416 3423
rect 1432 3417 1464 3423
rect 216 3397 264 3403
rect 920 3397 952 3403
rect 1656 3397 2136 3403
rect 2232 3417 2328 3423
rect 2344 3417 2472 3423
rect 2520 3417 4152 3423
rect 2776 3397 2904 3403
rect 3112 3397 3256 3403
rect 3288 3397 3368 3403
rect 3384 3397 3432 3403
rect 3512 3397 3848 3403
rect 3928 3397 3944 3403
rect 4264 3417 4392 3423
rect 4408 3417 4424 3423
rect 4440 3417 4504 3423
rect 4584 3417 4888 3423
rect 5208 3417 5560 3423
rect 5864 3417 5944 3423
rect 5960 3417 6120 3423
rect 4552 3397 4616 3403
rect 4648 3397 4680 3403
rect 5320 3397 6088 3403
rect 6344 3417 6488 3423
rect 6920 3417 6968 3423
rect 7064 3397 7272 3403
rect 7288 3397 7336 3403
rect 1240 3377 1368 3383
rect 1960 3377 2056 3383
rect 2072 3377 2264 3383
rect 3096 3377 3176 3383
rect 3352 3377 3464 3383
rect 3480 3377 3688 3383
rect 3896 3377 4248 3383
rect 4376 3377 4664 3383
rect 4840 3377 5000 3383
rect 5432 3377 5544 3383
rect 5560 3377 5864 3383
rect 5896 3377 5944 3383
rect 5960 3377 5992 3383
rect 6264 3377 6760 3383
rect 744 3357 1752 3363
rect 2200 3357 2456 3363
rect 2984 3357 3272 3363
rect 3688 3357 3784 3363
rect 3800 3357 4024 3363
rect 4136 3357 4232 3363
rect 4536 3357 4840 3363
rect 4856 3357 4872 3363
rect 5112 3357 5176 3363
rect 5192 3357 5256 3363
rect 5784 3357 5848 3363
rect 5912 3357 6280 3363
rect 6296 3357 6328 3363
rect 6376 3357 6424 3363
rect 7112 3357 7160 3363
rect 7176 3357 7443 3363
rect 3389 3348 3395 3352
rect 248 3337 392 3343
rect 408 3337 520 3343
rect 536 3337 1192 3343
rect 1272 3337 1288 3343
rect 1304 3337 2248 3343
rect 2296 3337 2440 3343
rect 2456 3337 2616 3343
rect 2632 3337 2952 3343
rect 3272 3337 3320 3343
rect 3485 3343 3491 3352
rect 3485 3337 3496 3343
rect 3736 3337 3912 3343
rect 3928 3337 3976 3343
rect 4056 3337 4072 3343
rect 4376 3337 4600 3343
rect 4616 3337 4648 3343
rect 4728 3337 4888 3343
rect 4936 3337 5352 3343
rect 5880 3337 6632 3343
rect 6712 3337 6744 3343
rect 7000 3337 7128 3343
rect 7192 3337 7240 3343
rect 7256 3337 7384 3343
rect 7437 3343 7443 3357
rect 7437 3337 7491 3343
rect 2253 3328 2259 3332
rect 5437 3328 5443 3332
rect 5837 3328 5843 3332
rect 40 3317 56 3323
rect 168 3317 216 3323
rect 280 3317 408 3323
rect 424 3317 456 3323
rect 600 3317 696 3323
rect 952 3317 1096 3323
rect 1416 3317 1432 3323
rect 1576 3317 1688 3323
rect 1848 3317 1960 3323
rect 2376 3317 2392 3323
rect 2488 3317 2520 3323
rect 2536 3317 2680 3323
rect 2696 3317 2840 3323
rect 3272 3317 3304 3323
rect 3384 3317 3448 3323
rect 3464 3317 4184 3323
rect 4328 3317 4360 3323
rect 4552 3317 4712 3323
rect 4728 3317 5400 3323
rect 5464 3317 5496 3323
rect 5640 3317 5704 3323
rect 6333 3317 6344 3323
rect 6424 3317 6616 3323
rect 6696 3317 6712 3323
rect 6920 3317 6952 3323
rect 7096 3317 7144 3323
rect 7160 3317 7272 3323
rect 7304 3317 7336 3323
rect 232 3297 760 3303
rect 1112 3297 1176 3303
rect 1704 3297 1736 3303
rect 1976 3297 2040 3303
rect 2088 3297 2280 3303
rect 2360 3297 2488 3303
rect 2504 3297 2600 3303
rect 2616 3297 2632 3303
rect 2712 3297 2968 3303
rect 3000 3297 3016 3303
rect 3032 3297 3128 3303
rect 3144 3297 3240 3303
rect 3256 3297 3400 3303
rect 3432 3297 3720 3303
rect 3752 3297 3763 3303
rect 3976 3297 4056 3303
rect 4488 3297 4520 3303
rect 4760 3297 4792 3303
rect 4872 3297 4888 3303
rect 4904 3297 4968 3303
rect 4984 3297 5000 3303
rect 5304 3297 5368 3303
rect 5544 3297 5608 3303
rect 5784 3297 5864 3303
rect 5944 3297 6200 3303
rect 6408 3297 6472 3303
rect 6520 3297 6568 3303
rect 6584 3297 6808 3303
rect 7080 3297 7112 3303
rect 7448 3297 7491 3303
rect 1336 3277 1368 3283
rect 1400 3277 2072 3283
rect 2104 3277 2264 3283
rect 2280 3277 3123 3283
rect 2136 3257 2184 3263
rect 2200 3257 2344 3263
rect 2392 3257 2504 3263
rect 2717 3257 3096 3263
rect 136 3237 184 3243
rect 200 3237 376 3243
rect 648 3237 696 3243
rect 2717 3243 2723 3257
rect 3117 3263 3123 3277
rect 3576 3277 3704 3283
rect 3768 3277 3800 3283
rect 3837 3283 3843 3292
rect 3837 3277 3976 3283
rect 4072 3277 4120 3283
rect 4376 3277 4456 3283
rect 4472 3277 4856 3283
rect 5592 3277 5672 3283
rect 5864 3277 5944 3283
rect 5960 3277 6904 3283
rect 6968 3277 7048 3283
rect 3117 3257 3864 3263
rect 3992 3257 4344 3263
rect 4776 3257 4840 3263
rect 5544 3257 5752 3263
rect 5848 3257 5944 3263
rect 6040 3257 6056 3263
rect 6072 3257 6424 3263
rect 6488 3257 6728 3263
rect 6760 3257 7064 3263
rect 2392 3237 2723 3243
rect 2744 3237 2760 3243
rect 3149 3237 4440 3243
rect 3149 3223 3155 3237
rect 4648 3237 4824 3243
rect 4840 3237 4968 3243
rect 5229 3237 5240 3243
rect 5528 3237 5640 3243
rect 5688 3237 5800 3243
rect 5928 3237 6152 3243
rect 6168 3237 6568 3243
rect 6584 3237 6744 3243
rect 6920 3237 7176 3243
rect 2024 3217 3155 3223
rect 2808 3197 3000 3203
rect 4152 3217 4936 3223
rect 4952 3217 5192 3223
rect 3224 3197 3256 3203
rect 3832 3197 3928 3203
rect 4200 3197 4264 3203
rect 4600 3197 4808 3203
rect 4824 3197 5192 3203
rect 5304 3217 5688 3223
rect 5704 3217 5880 3223
rect 5896 3217 5928 3223
rect 6216 3217 6792 3223
rect 7032 3217 7352 3223
rect 5448 3197 5880 3203
rect 6184 3197 6200 3203
rect 6472 3197 7160 3203
rect 568 3177 824 3183
rect 1032 3177 1112 3183
rect 2376 3177 5128 3183
rect 5144 3177 5160 3183
rect 5208 3177 6648 3183
rect 6696 3177 6936 3183
rect 472 3157 1000 3163
rect 2856 3157 2936 3163
rect 3704 3157 3912 3163
rect 3976 3157 4424 3163
rect 4504 3157 4600 3163
rect 4856 3157 5576 3163
rect 5608 3157 5624 3163
rect 6744 3157 7128 3163
rect 488 3137 552 3143
rect 1544 3137 1768 3143
rect 1784 3137 1816 3143
rect 1976 3137 2136 3143
rect 2488 3137 2520 3143
rect 2536 3137 2904 3143
rect 3384 3137 3784 3143
rect 3944 3137 3976 3143
rect 3992 3137 4184 3143
rect 4328 3137 4360 3143
rect 4456 3137 4504 3143
rect 4520 3137 4568 3143
rect 4584 3137 4616 3143
rect 4632 3137 4696 3143
rect 4776 3137 4824 3143
rect 5384 3137 5480 3143
rect 5736 3137 5832 3143
rect 5864 3137 6520 3143
rect 6536 3137 6776 3143
rect 6888 3137 6968 3143
rect 6984 3137 7064 3143
rect 72 3117 104 3123
rect 376 3117 504 3123
rect 712 3117 744 3123
rect 776 3117 840 3123
rect 1016 3117 1048 3123
rect 1464 3117 1640 3123
rect 1720 3117 1912 3123
rect 1928 3117 1944 3123
rect 1960 3117 1992 3123
rect 2088 3117 2888 3123
rect 2904 3117 3080 3123
rect 3112 3117 3176 3123
rect 3192 3117 3208 3123
rect 3304 3117 3352 3123
rect 3432 3117 3528 3123
rect 3912 3117 4072 3123
rect 4088 3117 4280 3123
rect 4296 3117 4552 3123
rect 4568 3117 4728 3123
rect 4904 3117 4920 3123
rect 4984 3117 5096 3123
rect 5112 3117 5288 3123
rect 5320 3117 5384 3123
rect 5544 3117 5592 3123
rect 5608 3117 5784 3123
rect 5800 3117 5896 3123
rect 6104 3117 6376 3123
rect 6840 3117 6936 3123
rect 7064 3117 7080 3123
rect 200 3097 232 3103
rect 424 3097 616 3103
rect 632 3097 904 3103
rect 920 3097 968 3103
rect 984 3097 1160 3103
rect 1624 3097 1656 3103
rect 1752 3097 1944 3103
rect 2024 3097 2104 3103
rect 2120 3097 2216 3103
rect 2232 3097 2392 3103
rect 2605 3097 2616 3103
rect 2776 3097 2824 3103
rect 2840 3097 2872 3103
rect 2920 3097 3048 3103
rect 3080 3097 3352 3103
rect 3384 3097 3752 3103
rect 3768 3097 3800 3103
rect 3992 3097 4168 3103
rect 4312 3097 4424 3103
rect 4456 3097 4515 3103
rect 24 3077 248 3083
rect 264 3077 456 3083
rect 472 3077 488 3083
rect 792 3077 952 3083
rect 1064 3077 1240 3083
rect 1272 3077 1336 3083
rect 1352 3077 1400 3083
rect 1608 3077 1672 3083
rect 1752 3077 1800 3083
rect 1944 3077 1976 3083
rect 1992 3077 2056 3083
rect 2200 3077 2392 3083
rect 2424 3077 2552 3083
rect 2888 3077 3384 3083
rect 3400 3077 3432 3083
rect 3480 3077 3656 3083
rect 3800 3077 3928 3083
rect 4152 3077 4376 3083
rect 4392 3077 4488 3083
rect 4509 3083 4515 3097
rect 4696 3097 4744 3103
rect 4808 3097 4920 3103
rect 5048 3097 5464 3103
rect 5496 3097 5544 3103
rect 5560 3097 5624 3103
rect 5656 3097 5704 3103
rect 5720 3097 5736 3103
rect 5752 3097 5848 3103
rect 5912 3097 5944 3103
rect 5976 3097 6104 3103
rect 6168 3097 6456 3103
rect 6808 3097 6824 3103
rect 7224 3097 7336 3103
rect 4509 3077 5032 3083
rect 5064 3077 5080 3083
rect 5096 3077 5256 3083
rect 5416 3077 5448 3083
rect 5592 3077 5768 3083
rect 5784 3077 5816 3083
rect 5912 3077 6184 3083
rect 6264 3077 6328 3083
rect 7112 3077 7208 3083
rect 7341 3068 7347 3072
rect 600 3057 1064 3063
rect 1512 3057 2040 3063
rect 2728 3057 2792 3063
rect 2984 3057 3096 3063
rect 3160 3057 3176 3063
rect 3192 3057 3224 3063
rect 3256 3057 3304 3063
rect 3336 3057 3400 3063
rect 3416 3057 3704 3063
rect 4760 3057 4856 3063
rect 5016 3057 5032 3063
rect 5272 3057 5416 3063
rect 5624 3057 5688 3063
rect 5704 3057 5976 3063
rect 6264 3057 6376 3063
rect 6440 3057 6840 3063
rect 205 3048 211 3052
rect 520 3037 984 3043
rect 1000 3037 2072 3043
rect 3336 3037 3368 3043
rect 3528 3037 3544 3043
rect 4040 3037 4056 3043
rect 4664 3037 4984 3043
rect 5000 3037 5144 3043
rect 5864 3037 6264 3043
rect 6472 3037 6552 3043
rect 6568 3037 6632 3043
rect 40 3017 88 3023
rect 312 2997 760 3003
rect 776 2997 1352 3003
rect 2936 3017 3656 3023
rect 3080 2997 3128 3003
rect 3672 2997 3864 3003
rect 4616 3017 4808 3023
rect 5816 3017 5864 3023
rect 5880 3017 6216 3023
rect 4936 2997 5080 3003
rect 5448 2997 5944 3003
rect 6792 2997 7112 3003
rect 7128 2997 7192 3003
rect 216 2977 376 2983
rect 392 2977 680 2983
rect 696 2977 1128 2983
rect 1144 2977 1752 2983
rect 2248 2977 2344 2983
rect 2360 2977 3256 2983
rect 3720 2977 3832 2983
rect 3848 2977 4088 2983
rect 4328 2977 4504 2983
rect 4520 2977 4568 2983
rect 4760 2977 5064 2983
rect 5272 2977 6632 2983
rect 6824 2977 7096 2983
rect 312 2957 488 2963
rect 1048 2957 1352 2963
rect 1368 2957 1480 2963
rect 1704 2957 1880 2963
rect 1896 2957 1960 2963
rect 2616 2957 2744 2963
rect 2824 2957 2840 2963
rect 3272 2957 3512 2963
rect 3528 2957 3592 2963
rect 3720 2957 3864 2963
rect 3896 2957 4216 2963
rect 4712 2957 4728 2963
rect 4952 2957 5000 2963
rect 5416 2957 5576 2963
rect 5592 2957 5704 2963
rect 5928 2957 6104 2963
rect 6120 2957 6152 2963
rect 6200 2957 6648 2963
rect 6664 2957 6680 2963
rect 6856 2957 6888 2963
rect 280 2937 371 2943
rect 365 2928 371 2937
rect 568 2937 824 2943
rect 1384 2937 2616 2943
rect 2728 2937 2760 2943
rect 2776 2937 2888 2943
rect 2936 2937 3016 2943
rect 3160 2937 3352 2943
rect 3368 2937 3528 2943
rect 3624 2937 3880 2943
rect 4472 2937 4696 2943
rect 4888 2937 4968 2943
rect 5464 2937 5496 2943
rect 5512 2937 5544 2943
rect 5560 2937 5576 2943
rect 5656 2937 6056 2943
rect 6072 2937 6136 2943
rect 6360 2937 6488 2943
rect 6584 2937 6936 2943
rect 7112 2937 7128 2943
rect 168 2917 216 2923
rect 248 2917 264 2923
rect 472 2917 728 2923
rect 744 2917 776 2923
rect 1080 2917 1112 2923
rect 1128 2917 1384 2923
rect 1400 2917 1432 2923
rect 1448 2917 1608 2923
rect 1624 2917 1656 2923
rect 1672 2917 2024 2923
rect 2040 2917 2088 2923
rect 2168 2917 2216 2923
rect 2280 2917 2472 2923
rect 2488 2917 2824 2923
rect 3224 2917 3304 2923
rect 3336 2917 3608 2923
rect 3656 2917 3720 2923
rect 3960 2917 4040 2923
rect 4200 2917 4232 2923
rect 4296 2917 4376 2923
rect 4568 2917 4616 2923
rect 4712 2917 4872 2923
rect 4936 2917 4947 2923
rect 5400 2917 5656 2923
rect 5672 2917 5752 2923
rect 6120 2917 6264 2923
rect 6328 2917 6440 2923
rect 6536 2917 6568 2923
rect 6600 2917 6664 2923
rect 6680 2917 6712 2923
rect 6888 2917 6968 2923
rect 7224 2917 7240 2923
rect 7352 2917 7384 2923
rect 200 2897 392 2903
rect 520 2897 568 2903
rect 584 2897 680 2903
rect 728 2897 792 2903
rect 808 2897 840 2903
rect 1128 2897 1224 2903
rect 1656 2897 1752 2903
rect 2088 2897 2520 2903
rect 3320 2897 3384 2903
rect 3592 2897 3944 2903
rect 3960 2897 4120 2903
rect 4584 2897 4648 2903
rect 4808 2897 5448 2903
rect 5464 2897 5512 2903
rect 5528 2897 5672 2903
rect 5704 2897 5800 2903
rect 5816 2897 5992 2903
rect 6584 2897 6760 2903
rect 6776 2897 6904 2903
rect 7096 2897 7112 2903
rect 7240 2897 7304 2903
rect 136 2877 616 2883
rect 776 2877 952 2883
rect 1688 2877 1704 2883
rect 3720 2877 3880 2883
rect 3992 2877 4168 2883
rect 4184 2877 4520 2883
rect 4696 2877 4760 2883
rect 4776 2877 4808 2883
rect 4872 2877 4920 2883
rect 4984 2877 5240 2883
rect 5592 2877 5688 2883
rect 5720 2877 5896 2883
rect 6040 2877 6328 2883
rect 7160 2877 7176 2883
rect 7272 2877 7400 2883
rect 792 2857 824 2863
rect 2856 2857 3336 2863
rect 3608 2857 3752 2863
rect 4072 2857 4104 2863
rect 4120 2857 4184 2863
rect 4200 2857 4440 2863
rect 4456 2857 4968 2863
rect 5304 2857 5528 2863
rect 2184 2837 3208 2843
rect 3512 2837 4600 2843
rect 4680 2837 4888 2843
rect 4904 2837 5016 2843
rect 5032 2837 5496 2843
rect 5512 2837 5720 2843
rect 1448 2797 1464 2803
rect 1480 2797 2360 2803
rect 4200 2817 4552 2823
rect 4728 2817 4840 2823
rect 5496 2817 6040 2823
rect 6344 2817 6920 2823
rect 6936 2817 6984 2823
rect 5272 2797 5736 2803
rect 5768 2797 5848 2803
rect 7000 2797 7160 2803
rect 605 2783 611 2792
rect 6205 2788 6211 2792
rect 605 2777 616 2783
rect 1144 2777 1176 2783
rect 1352 2777 1384 2783
rect 1496 2777 1528 2783
rect 1544 2777 1608 2783
rect 1976 2777 2040 2783
rect 2536 2777 2824 2783
rect 2840 2777 3336 2783
rect 3768 2777 4104 2783
rect 4504 2777 4936 2783
rect 5176 2777 5640 2783
rect 5656 2777 6008 2783
rect 6664 2777 6856 2783
rect 6872 2777 6984 2783
rect 7000 2777 7208 2783
rect 7224 2777 7288 2783
rect 1688 2757 1848 2763
rect 2061 2763 2067 2772
rect 2056 2757 2067 2763
rect 2088 2757 2120 2763
rect 2248 2757 2504 2763
rect 2520 2757 2552 2763
rect 2568 2757 2664 2763
rect 2680 2757 2728 2763
rect 2792 2757 2856 2763
rect 3064 2757 4296 2763
rect 4680 2757 5128 2763
rect 5144 2757 5864 2763
rect 6456 2757 6680 2763
rect 152 2737 264 2743
rect 968 2737 1144 2743
rect 1576 2737 1768 2743
rect 1864 2737 1976 2743
rect 2093 2737 2104 2743
rect 2488 2737 2984 2743
rect 3224 2737 3384 2743
rect 3656 2737 4184 2743
rect 4456 2737 4584 2743
rect 4600 2737 4680 2743
rect 4920 2737 5368 2743
rect 5416 2737 5880 2743
rect 6040 2737 6616 2743
rect 6696 2737 7491 2743
rect 24 2717 200 2723
rect 440 2717 520 2723
rect 1048 2717 1480 2723
rect 1496 2717 1720 2723
rect 1784 2717 1816 2723
rect 1896 2717 1907 2723
rect 2392 2717 4691 2723
rect 248 2697 280 2703
rect 376 2697 504 2703
rect 552 2697 632 2703
rect 728 2697 760 2703
rect 776 2697 840 2703
rect 888 2697 968 2703
rect 984 2697 1016 2703
rect 1128 2697 1864 2703
rect 1880 2697 2088 2703
rect 2104 2697 2136 2703
rect 2152 2697 2376 2703
rect 2648 2697 2776 2703
rect 2792 2697 2856 2703
rect 3016 2697 3080 2703
rect 3368 2697 3400 2703
rect 3464 2697 3528 2703
rect 3640 2697 3672 2703
rect 4184 2697 4216 2703
rect 4360 2697 4392 2703
rect 4440 2697 4536 2703
rect 4600 2697 4664 2703
rect 4685 2703 4691 2717
rect 4792 2717 4888 2723
rect 4920 2717 5144 2723
rect 5224 2717 5304 2723
rect 5352 2717 5432 2723
rect 5464 2717 5624 2723
rect 5656 2717 5672 2723
rect 5704 2717 5752 2723
rect 5784 2717 5928 2723
rect 6024 2717 6248 2723
rect 6408 2717 6488 2723
rect 7128 2717 7176 2723
rect 4685 2697 4776 2703
rect 4952 2697 5064 2703
rect 5080 2697 5112 2703
rect 5128 2697 5800 2703
rect 5816 2697 5848 2703
rect 6120 2697 6152 2703
rect 6536 2697 6904 2703
rect 6920 2697 7016 2703
rect 7096 2697 7112 2703
rect 7144 2697 7240 2703
rect 7448 2697 7491 2703
rect 301 2688 307 2692
rect 7293 2688 7299 2692
rect 504 2677 808 2683
rect 824 2677 1112 2683
rect 1336 2677 1544 2683
rect 1752 2677 1880 2683
rect 1896 2677 1992 2683
rect 2360 2677 2504 2683
rect 3000 2677 3032 2683
rect 3336 2677 3432 2683
rect 3528 2677 3640 2683
rect 3688 2677 3864 2683
rect 4264 2677 4440 2683
rect 4520 2677 4696 2683
rect 5272 2677 5480 2683
rect 5528 2677 5608 2683
rect 5640 2677 5880 2683
rect 5901 2677 5912 2683
rect 6104 2677 6120 2683
rect 6136 2677 6232 2683
rect 6248 2677 7176 2683
rect -51 2657 8 2663
rect 104 2657 568 2663
rect 712 2657 760 2663
rect 904 2657 1032 2663
rect 1160 2657 1768 2663
rect 1784 2657 2008 2663
rect 2072 2657 2296 2663
rect 2584 2657 2840 2663
rect 2920 2657 2952 2663
rect 3320 2657 3416 2663
rect 3432 2657 4296 2663
rect 4632 2657 4648 2663
rect 5336 2657 5528 2663
rect 5576 2657 5976 2663
rect 6184 2657 6995 2663
rect 264 2637 376 2643
rect 584 2637 824 2643
rect 840 2637 1208 2643
rect 1224 2637 1928 2643
rect 1944 2637 2024 2643
rect 2040 2637 2232 2643
rect 2664 2637 2904 2643
rect 2952 2637 3112 2643
rect 3128 2637 3416 2643
rect 3432 2637 3624 2643
rect 3736 2637 3752 2643
rect 4152 2637 4248 2643
rect 4536 2637 4728 2643
rect 4760 2637 4856 2643
rect 4872 2637 5160 2643
rect 5544 2637 5784 2643
rect 5896 2637 6312 2643
rect 6808 2637 6872 2643
rect 6989 2643 6995 2657
rect 7192 2657 7491 2663
rect 6989 2637 7208 2643
rect 7224 2637 7432 2643
rect 568 2617 632 2623
rect 664 2617 904 2623
rect 920 2617 1000 2623
rect 1016 2617 1112 2623
rect 1128 2617 1192 2623
rect 1960 2617 2136 2623
rect -51 2597 104 2603
rect 120 2597 184 2603
rect 392 2597 728 2603
rect 744 2597 920 2603
rect 936 2597 1448 2603
rect 1464 2597 1736 2603
rect 1752 2597 2072 2603
rect 2424 2617 2792 2623
rect 2808 2617 3064 2623
rect 3080 2617 3560 2623
rect 2824 2597 2904 2603
rect 2920 2597 3144 2603
rect 4584 2617 4792 2623
rect 5256 2617 5320 2623
rect 5432 2617 5560 2623
rect 5592 2617 6136 2623
rect 4616 2597 4952 2603
rect 5288 2597 5384 2603
rect 5544 2597 5656 2603
rect 5672 2597 6008 2603
rect 6712 2617 7064 2623
rect 7112 2617 7320 2623
rect 7389 2617 7491 2623
rect 7389 2603 7395 2617
rect 6600 2597 7395 2603
rect 24 2577 712 2583
rect 728 2577 888 2583
rect 1032 2577 1096 2583
rect 1112 2577 1160 2583
rect 2088 2577 2168 2583
rect 2184 2577 2328 2583
rect 2616 2577 2712 2583
rect 3048 2577 3144 2583
rect 4376 2577 4408 2583
rect 4424 2577 4712 2583
rect 4968 2577 5384 2583
rect 5405 2577 5704 2583
rect -51 2557 8 2563
rect 40 2557 451 2563
rect 296 2537 360 2543
rect 445 2543 451 2557
rect 472 2557 648 2563
rect 664 2557 920 2563
rect 1096 2557 2120 2563
rect 2168 2557 2776 2563
rect 3064 2557 3288 2563
rect 3304 2557 3512 2563
rect 3800 2557 3976 2563
rect 4440 2557 4632 2563
rect 4936 2557 5256 2563
rect 5288 2557 5352 2563
rect 5405 2563 5411 2577
rect 6024 2577 6120 2583
rect 6136 2577 6472 2583
rect 6520 2577 6808 2583
rect 6824 2577 6840 2583
rect 6968 2577 7080 2583
rect 7096 2577 7160 2583
rect 7176 2577 7240 2583
rect 7256 2577 7304 2583
rect 7469 2577 7491 2583
rect 5368 2557 5411 2563
rect 5512 2557 5640 2563
rect 6376 2557 6408 2563
rect 6424 2557 6568 2563
rect 6872 2557 6920 2563
rect 6936 2557 7032 2563
rect 7469 2563 7475 2577
rect 7160 2557 7475 2563
rect 445 2537 680 2543
rect 696 2537 824 2543
rect 840 2537 856 2543
rect 920 2537 984 2543
rect 1288 2537 1432 2543
rect 1592 2537 1640 2543
rect 1656 2537 1800 2543
rect 2136 2537 2216 2543
rect 2328 2537 2376 2543
rect 2408 2537 2440 2543
rect 2504 2537 2648 2543
rect 2728 2537 2760 2543
rect 3080 2537 3112 2543
rect 3240 2537 3272 2543
rect 3336 2537 3416 2543
rect 3448 2537 3688 2543
rect 3704 2537 3992 2543
rect 4104 2537 4120 2543
rect 4360 2537 4376 2543
rect 4472 2537 4520 2543
rect 4824 2537 4968 2543
rect 5720 2537 5768 2543
rect 5789 2537 6184 2543
rect 381 2528 387 2532
rect 4461 2528 4467 2532
rect -51 2517 24 2523
rect 344 2517 371 2523
rect 152 2497 216 2503
rect 312 2497 344 2503
rect 365 2503 371 2517
rect 408 2517 456 2523
rect 664 2517 696 2523
rect 712 2517 744 2523
rect 1000 2517 1064 2523
rect 1400 2517 1496 2523
rect 1512 2517 1528 2523
rect 1624 2517 1672 2523
rect 1864 2517 1992 2523
rect 2600 2517 2904 2523
rect 2920 2517 3432 2523
rect 3480 2517 3496 2523
rect 3560 2517 3592 2523
rect 3624 2517 3704 2523
rect 3720 2517 3752 2523
rect 3768 2517 3880 2523
rect 3992 2517 4168 2523
rect 4264 2517 4344 2523
rect 4360 2517 4424 2523
rect 4488 2517 4664 2523
rect 4680 2517 4776 2523
rect 4808 2517 4952 2523
rect 5128 2517 5288 2523
rect 5320 2517 5464 2523
rect 5789 2523 5795 2537
rect 6200 2537 6552 2543
rect 6584 2537 6728 2543
rect 6744 2537 6776 2543
rect 6904 2537 7016 2543
rect 7064 2537 7491 2543
rect 5560 2517 5795 2523
rect 5976 2517 6008 2523
rect 6024 2517 6136 2523
rect 6152 2517 6200 2523
rect 6216 2517 6296 2523
rect 6488 2517 6600 2523
rect 6888 2517 6904 2523
rect 6984 2517 7048 2523
rect 7064 2517 7112 2523
rect 7160 2517 7272 2523
rect 365 2497 584 2503
rect 872 2497 968 2503
rect 984 2497 1016 2503
rect 1432 2497 1464 2503
rect 1480 2497 1640 2503
rect 1656 2497 1784 2503
rect 1816 2497 1848 2503
rect 1864 2497 1912 2503
rect 2024 2497 2280 2503
rect 2648 2497 2680 2503
rect 2696 2497 2824 2503
rect 2936 2497 3064 2503
rect 3272 2497 3320 2503
rect 3752 2497 3848 2503
rect 4024 2497 4056 2503
rect 4072 2497 4136 2503
rect 4152 2497 4232 2503
rect 4248 2497 4280 2503
rect 4552 2497 4600 2503
rect 4808 2497 5576 2503
rect 5688 2497 5720 2503
rect 5736 2497 5976 2503
rect 6088 2497 6200 2503
rect 6344 2497 6440 2503
rect 6456 2497 6520 2503
rect 6632 2497 6920 2503
rect 6968 2497 6979 2503
rect 7048 2497 7096 2503
rect 7448 2497 7491 2503
rect -51 2477 56 2483
rect 72 2477 136 2483
rect 168 2477 264 2483
rect 1192 2477 2360 2483
rect 2376 2477 2408 2483
rect 2792 2477 2904 2483
rect 3288 2477 3544 2483
rect 3656 2477 3912 2483
rect 3928 2477 4024 2483
rect 4296 2477 4328 2483
rect 4344 2477 4440 2483
rect 4536 2477 4552 2483
rect 4664 2477 6056 2483
rect 6104 2477 6136 2483
rect 6232 2477 6536 2483
rect 7000 2477 7080 2483
rect 7240 2477 7256 2483
rect 1480 2457 1576 2463
rect 2360 2457 3592 2463
rect 4520 2457 4616 2463
rect 4632 2457 4744 2463
rect 5544 2457 5592 2463
rect 5752 2457 5864 2463
rect 6376 2457 6744 2463
rect 6920 2457 7128 2463
rect 7256 2457 7368 2463
rect 88 2437 136 2443
rect 152 2437 312 2443
rect 1832 2437 2744 2443
rect 4680 2437 4840 2443
rect 4856 2437 4952 2443
rect 4968 2437 5000 2443
rect 5384 2437 5784 2443
rect 5816 2437 5848 2443
rect 6072 2437 6216 2443
rect 6536 2437 7032 2443
rect 7080 2437 7224 2443
rect 344 2397 616 2403
rect 1272 2417 1512 2423
rect 1784 2417 2584 2423
rect 2840 2397 2920 2403
rect 2936 2397 2968 2403
rect 4968 2417 5176 2423
rect 4557 2397 4872 2403
rect 968 2377 1144 2383
rect 4557 2383 4563 2397
rect 5864 2417 6344 2423
rect 6504 2417 6696 2423
rect 6760 2417 6968 2423
rect 7096 2417 7384 2423
rect 5624 2397 6120 2403
rect 6264 2397 6520 2403
rect 6920 2397 7160 2403
rect 1640 2377 4563 2383
rect 4584 2377 4872 2383
rect 4888 2377 5048 2383
rect 5912 2377 6072 2383
rect 6136 2377 6392 2383
rect 6424 2377 6600 2383
rect 6728 2377 6888 2383
rect 6936 2377 7096 2383
rect 7133 2377 7288 2383
rect 680 2357 792 2363
rect 1672 2357 1880 2363
rect 3640 2357 3896 2363
rect 3912 2357 3944 2363
rect 5400 2357 5560 2363
rect 5592 2357 5656 2363
rect 6040 2357 6088 2363
rect 6104 2357 6296 2363
rect 6312 2357 6536 2363
rect 6552 2357 6632 2363
rect 6648 2357 6840 2363
rect 6856 2357 6936 2363
rect 7133 2363 7139 2377
rect 6952 2357 7139 2363
rect 7160 2357 7416 2363
rect 712 2337 760 2343
rect 776 2337 904 2343
rect 920 2337 952 2343
rect 1016 2337 1176 2343
rect 1528 2337 1576 2343
rect 1592 2337 1704 2343
rect 1720 2337 1976 2343
rect 1992 2337 2024 2343
rect 2248 2337 2376 2343
rect 2392 2337 3224 2343
rect 3720 2337 3752 2343
rect 5016 2337 5128 2343
rect 5144 2337 5496 2343
rect 5512 2337 5528 2343
rect 5848 2337 5912 2343
rect 6088 2337 6824 2343
rect 7048 2337 7192 2343
rect 264 2317 280 2323
rect 424 2317 456 2323
rect 760 2317 776 2323
rect 1320 2317 1528 2323
rect 2296 2317 2344 2323
rect 2360 2317 2616 2323
rect 2632 2317 2664 2323
rect 2888 2317 3480 2323
rect 3608 2317 3816 2323
rect 4008 2317 4104 2323
rect 4248 2317 4280 2323
rect 5224 2317 5320 2323
rect 5336 2317 5416 2323
rect 5928 2317 6136 2323
rect 6216 2317 6232 2323
rect 6440 2317 6472 2323
rect 6504 2317 6568 2323
rect 6616 2317 6696 2323
rect 6744 2317 6760 2323
rect 7096 2317 7208 2323
rect 7224 2317 7272 2323
rect 4973 2308 4979 2312
rect 5645 2308 5651 2312
rect 7053 2308 7059 2312
rect 7357 2308 7363 2312
rect 152 2297 232 2303
rect 280 2297 424 2303
rect 440 2297 632 2303
rect 648 2297 776 2303
rect 792 2297 1256 2303
rect 1448 2297 1704 2303
rect 1832 2297 1880 2303
rect 2136 2297 2296 2303
rect 2472 2297 2616 2303
rect 2776 2297 2920 2303
rect 2984 2297 3064 2303
rect 3384 2297 3416 2303
rect 3432 2297 3800 2303
rect 3816 2297 3848 2303
rect 3960 2297 4104 2303
rect 4296 2297 4440 2303
rect 4632 2297 4648 2303
rect 4664 2297 4712 2303
rect 4984 2297 5176 2303
rect 5352 2297 5368 2303
rect 5416 2297 5496 2303
rect 5736 2297 5880 2303
rect 6013 2297 6024 2303
rect 6184 2297 6552 2303
rect 6568 2297 6648 2303
rect 6664 2297 6792 2303
rect 6808 2297 6856 2303
rect 6888 2297 6952 2303
rect 6984 2297 7048 2303
rect 7240 2297 7304 2303
rect 472 2277 984 2283
rect 1000 2277 1032 2283
rect 1112 2277 1208 2283
rect 1432 2277 1464 2283
rect 2152 2277 2440 2283
rect 3080 2277 3256 2283
rect 3528 2277 3720 2283
rect 4168 2277 4424 2283
rect 4712 2277 4872 2283
rect 5144 2277 5256 2283
rect 5288 2277 5352 2283
rect 5400 2277 5432 2283
rect 5448 2277 5704 2283
rect 5720 2277 5864 2283
rect 5880 2277 5944 2283
rect 5976 2277 6360 2283
rect 6600 2277 6632 2283
rect 1229 2268 1235 2272
rect 24 2257 200 2263
rect 216 2257 376 2263
rect 552 2257 712 2263
rect 856 2257 1112 2263
rect 1128 2257 1208 2263
rect 1336 2257 1400 2263
rect 1480 2257 1544 2263
rect 1597 2263 1603 2272
rect 1592 2257 1603 2263
rect 1944 2257 2040 2263
rect 2056 2257 2280 2263
rect 2296 2257 2984 2263
rect 3000 2257 3128 2263
rect 3608 2257 3880 2263
rect 3896 2257 4056 2263
rect 4072 2257 4216 2263
rect 4232 2257 4584 2263
rect 4648 2257 5144 2263
rect 5320 2257 5672 2263
rect 6120 2257 6168 2263
rect 6184 2257 6328 2263
rect 6824 2257 7208 2263
rect 232 2237 296 2243
rect 312 2237 632 2243
rect 648 2237 760 2243
rect 776 2237 1320 2243
rect 1608 2237 1624 2243
rect 2072 2237 2248 2243
rect 2264 2237 2616 2243
rect 2808 2237 3448 2243
rect 4184 2237 4552 2243
rect 4568 2237 4632 2243
rect 5128 2237 5288 2243
rect 5496 2237 5608 2243
rect 6056 2237 6184 2243
rect 6200 2237 6632 2243
rect 984 2217 1720 2223
rect 1736 2217 1784 2223
rect 1912 2217 2120 2223
rect 1432 2197 1832 2203
rect 1864 2197 1944 2203
rect 1976 2197 1992 2203
rect 2696 2217 3000 2223
rect 3016 2217 3080 2223
rect 3768 2197 3784 2203
rect 4296 2217 4808 2223
rect 5032 2217 5064 2223
rect 5080 2217 5448 2223
rect 5464 2217 5848 2223
rect 5864 2217 5912 2223
rect 4360 2197 4536 2203
rect 4584 2197 4776 2203
rect 5032 2197 5480 2203
rect 5560 2197 6216 2203
rect 6648 2217 6776 2223
rect 6792 2217 7000 2223
rect 7016 2217 7064 2223
rect 7320 2197 7384 2203
rect 312 2177 344 2183
rect 360 2177 584 2183
rect 632 2177 728 2183
rect 744 2177 856 2183
rect 1064 2177 1304 2183
rect 1592 2177 2056 2183
rect 2552 2177 2792 2183
rect 3656 2177 3752 2183
rect 4488 2177 4920 2183
rect 5384 2177 5464 2183
rect 5480 2177 5592 2183
rect 5752 2177 5928 2183
rect 5944 2177 6008 2183
rect 6024 2177 6136 2183
rect 6216 2177 6504 2183
rect 7320 2177 7400 2183
rect 216 2157 408 2163
rect 424 2157 744 2163
rect 1192 2157 1432 2163
rect 1512 2157 1704 2163
rect 1800 2157 2184 2163
rect 2792 2157 2920 2163
rect 2936 2157 3048 2163
rect 3064 2157 3432 2163
rect 3704 2157 3880 2163
rect 3960 2157 3976 2163
rect 4200 2157 4312 2163
rect 4776 2157 4952 2163
rect 4968 2157 5096 2163
rect 5112 2157 5208 2163
rect 5288 2157 5400 2163
rect 5512 2157 5624 2163
rect 6520 2157 6552 2163
rect 6840 2157 7032 2163
rect 184 2137 456 2143
rect 1832 2137 2008 2143
rect 2024 2137 2136 2143
rect 2312 2137 2456 2143
rect 2744 2137 2771 2143
rect 1293 2128 1299 2132
rect 152 2117 232 2123
rect 520 2117 664 2123
rect 936 2117 1000 2123
rect 1144 2117 1176 2123
rect 1400 2117 1512 2123
rect 1544 2117 1592 2123
rect 1624 2117 1848 2123
rect 2088 2117 2099 2123
rect 2184 2117 2328 2123
rect 2664 2117 2744 2123
rect 2765 2123 2771 2137
rect 3048 2137 3384 2143
rect 4056 2137 4328 2143
rect 4344 2137 4392 2143
rect 4648 2137 4696 2143
rect 4936 2137 5480 2143
rect 5672 2137 5704 2143
rect 5832 2137 6312 2143
rect 6376 2137 6520 2143
rect 6568 2137 6792 2143
rect 6856 2137 7208 2143
rect 7224 2137 7240 2143
rect 7256 2137 7288 2143
rect 2845 2128 2851 2132
rect 2765 2117 2776 2123
rect 3160 2117 3272 2123
rect 3288 2117 3336 2123
rect 3368 2117 3512 2123
rect 3672 2117 3752 2123
rect 3944 2117 3992 2123
rect 4008 2117 4136 2123
rect 4472 2117 4520 2123
rect 4616 2117 4664 2123
rect 5000 2117 5096 2123
rect 5112 2117 5160 2123
rect 5192 2117 5384 2123
rect 5544 2117 5592 2123
rect 5608 2117 5624 2123
rect 5704 2117 5800 2123
rect 5976 2117 6024 2123
rect 6040 2117 6104 2123
rect 6168 2117 6216 2123
rect 6232 2117 6344 2123
rect 6360 2117 6680 2123
rect 6696 2117 6808 2123
rect 6824 2117 6888 2123
rect 6968 2117 7016 2123
rect 7032 2117 7112 2123
rect 7128 2117 7144 2123
rect 7160 2117 7336 2123
rect 328 2097 360 2103
rect 376 2097 616 2103
rect 664 2097 696 2103
rect 712 2097 744 2103
rect 1192 2097 1496 2103
rect 1512 2097 1624 2103
rect 1768 2097 2104 2103
rect 2216 2097 2296 2103
rect 2712 2097 2808 2103
rect 2824 2097 3016 2103
rect 3032 2097 3224 2103
rect 3320 2097 3352 2103
rect 3512 2097 4104 2103
rect 4136 2097 4456 2103
rect 4552 2097 5000 2103
rect 5400 2097 5416 2103
rect 5480 2097 6456 2103
rect 6488 2097 6584 2103
rect 6600 2097 6664 2103
rect 6712 2097 6872 2103
rect 6888 2097 6984 2103
rect 7080 2097 7112 2103
rect 7160 2097 7491 2103
rect 4509 2088 4515 2092
rect 24 2077 264 2083
rect 280 2077 392 2083
rect 888 2077 1416 2083
rect 1432 2077 1752 2083
rect 2104 2077 2952 2083
rect 2968 2077 3416 2083
rect 3624 2077 3656 2083
rect 3960 2077 4024 2083
rect 4392 2077 4440 2083
rect 4584 2077 4712 2083
rect 4840 2077 5272 2083
rect 5624 2077 6056 2083
rect 6136 2077 6200 2083
rect 6248 2077 6696 2083
rect 6776 2077 6808 2083
rect 6968 2077 7048 2083
rect 1608 2057 1688 2063
rect 1704 2057 3048 2063
rect 3192 2057 3800 2063
rect 4328 2057 4584 2063
rect 4648 2057 4808 2063
rect 6008 2057 6072 2063
rect 6920 2057 6968 2063
rect 7048 2057 7064 2063
rect 872 2037 1064 2043
rect 1080 2037 1256 2043
rect 1576 2037 1848 2043
rect 3064 2037 5032 2043
rect 5160 2037 5960 2043
rect 5992 2037 6040 2043
rect 6808 2037 7176 2043
rect 1048 1997 1080 2003
rect 1544 2017 2328 2023
rect 2520 2017 3016 2023
rect 1672 1997 2264 2003
rect 2840 1997 2952 2003
rect 3256 2017 3832 2023
rect 3848 2017 3928 2023
rect 4248 2017 4376 2023
rect 4440 2017 4728 2023
rect 4104 1997 5176 2003
rect 5656 2017 6376 2023
rect 6216 1997 6712 2003
rect 6744 1997 6824 2003
rect 6904 1997 7080 2003
rect 7112 1997 7160 2003
rect 7192 1997 7416 2003
rect 1112 1977 2664 1983
rect 3176 1977 4088 1983
rect 4120 1977 4248 1983
rect 4344 1977 4504 1983
rect 4536 1977 4840 1983
rect 5496 1977 5656 1983
rect 5944 1977 6488 1983
rect 6504 1977 6632 1983
rect 6648 1977 7368 1983
rect 1016 1957 1080 1963
rect 1112 1957 1304 1963
rect 2168 1957 2504 1963
rect 2968 1957 3304 1963
rect 3320 1957 3368 1963
rect 3384 1957 3416 1963
rect 3432 1957 3464 1963
rect 3992 1957 4040 1963
rect 4056 1957 4536 1963
rect 5576 1957 5864 1963
rect 6088 1957 6104 1963
rect 6296 1957 6344 1963
rect 6456 1957 6840 1963
rect 7064 1957 7128 1963
rect 7144 1957 7352 1963
rect 7448 1957 7491 1963
rect 7037 1948 7043 1952
rect 168 1937 296 1943
rect 312 1937 424 1943
rect 616 1937 760 1943
rect 856 1937 1096 1943
rect 1224 1937 1512 1943
rect 1528 1937 1624 1943
rect 1720 1937 1784 1943
rect 3944 1937 4008 1943
rect 4088 1937 4232 1943
rect 4280 1937 4472 1943
rect 4488 1937 4536 1943
rect 4808 1937 4824 1943
rect 4840 1937 4968 1943
rect 5432 1937 5928 1943
rect 6200 1937 6296 1943
rect 7192 1937 7320 1943
rect 7336 1937 7491 1943
rect 344 1917 808 1923
rect 824 1917 920 1923
rect 968 1917 1016 1923
rect 1032 1917 1176 1923
rect 1480 1917 2216 1923
rect 2584 1917 2744 1923
rect 3960 1917 4024 1923
rect 4040 1917 4136 1923
rect 4152 1917 4280 1923
rect 4504 1917 4520 1923
rect 4616 1917 4664 1923
rect 4776 1917 4872 1923
rect 4888 1917 4984 1923
rect 6120 1917 6328 1923
rect 6456 1917 6744 1923
rect 6792 1917 6872 1923
rect 7080 1917 7272 1923
rect 7485 1917 7491 1937
rect 6349 1908 6355 1912
rect 24 1897 88 1903
rect 104 1897 168 1903
rect 248 1897 552 1903
rect 589 1897 888 1903
rect 589 1883 595 1897
rect 904 1897 1000 1903
rect 1032 1897 1080 1903
rect 1096 1897 1208 1903
rect 1416 1897 1432 1903
rect 1672 1897 1683 1903
rect 1864 1897 2488 1903
rect 2552 1897 2632 1903
rect 2856 1897 2984 1903
rect 3304 1897 3352 1903
rect 3480 1897 3576 1903
rect 3960 1897 3992 1903
rect 4264 1897 4328 1903
rect 4472 1897 4600 1903
rect 4920 1897 5176 1903
rect 5309 1897 5320 1903
rect 5448 1897 5544 1903
rect 5768 1897 5864 1903
rect 6904 1897 7048 1903
rect 7064 1897 7160 1903
rect 7240 1897 7304 1903
rect 7320 1897 7384 1903
rect 136 1877 595 1883
rect 616 1877 664 1883
rect 920 1877 1160 1883
rect 1176 1877 1320 1883
rect 1544 1877 1720 1883
rect 1784 1877 1832 1883
rect 1864 1877 1896 1883
rect 1912 1877 2440 1883
rect 2472 1877 2568 1883
rect 2760 1877 2776 1883
rect 2792 1877 2856 1883
rect 3144 1877 3400 1883
rect 3512 1877 3704 1883
rect 3800 1877 4152 1883
rect 4184 1877 4280 1883
rect 4392 1877 4696 1883
rect 4712 1877 4776 1883
rect 4797 1877 5368 1883
rect 232 1857 264 1863
rect 280 1857 376 1863
rect 440 1857 696 1863
rect 936 1857 1208 1863
rect 1400 1857 1688 1863
rect 1720 1857 1784 1863
rect 2040 1857 2232 1863
rect 2376 1857 2712 1863
rect 2776 1857 2824 1863
rect 3336 1857 3528 1863
rect 3544 1857 3720 1863
rect 3768 1857 3832 1863
rect 3848 1857 3976 1863
rect 4040 1857 4520 1863
rect 4584 1857 4680 1863
rect 4797 1863 4803 1877
rect 5464 1877 5528 1883
rect 5864 1877 5944 1883
rect 5960 1877 5992 1883
rect 6008 1877 6584 1883
rect 6616 1877 6632 1883
rect 6728 1877 6792 1883
rect 6824 1877 6936 1883
rect 4728 1857 4803 1863
rect 4904 1857 4984 1863
rect 5128 1857 5192 1863
rect 5480 1857 5592 1863
rect 6360 1857 6424 1863
rect 6568 1857 6584 1863
rect 6760 1857 6952 1863
rect 6968 1857 7000 1863
rect 488 1837 760 1843
rect 1032 1837 1080 1843
rect 1096 1837 1224 1843
rect 1288 1837 1800 1843
rect 1832 1837 1880 1843
rect 1896 1837 2120 1843
rect 2328 1837 2456 1843
rect 2744 1837 3784 1843
rect 3816 1837 4248 1843
rect 4376 1837 4488 1843
rect 4504 1837 4952 1843
rect 5192 1837 5288 1843
rect 5480 1837 5512 1843
rect 5528 1837 5544 1843
rect 5848 1837 6168 1843
rect 6216 1837 6504 1843
rect 6888 1837 7160 1843
rect 312 1817 552 1823
rect 568 1817 728 1823
rect 1192 1817 1304 1823
rect 1528 1817 1560 1823
rect 1704 1817 2136 1823
rect 552 1797 680 1803
rect 968 1797 1032 1803
rect 1048 1797 1080 1803
rect 1448 1797 1704 1803
rect 1944 1797 2120 1803
rect 2440 1817 2472 1823
rect 2504 1817 3208 1823
rect 3256 1817 3608 1823
rect 2280 1797 2600 1803
rect 2728 1797 2792 1803
rect 2824 1797 2840 1803
rect 2888 1797 3240 1803
rect 4440 1817 4568 1823
rect 4600 1817 5000 1823
rect 5021 1817 6104 1823
rect 4312 1797 4648 1803
rect 4680 1797 4808 1803
rect 5021 1803 5027 1817
rect 4840 1797 5027 1803
rect 5112 1797 5176 1803
rect 5192 1797 5288 1803
rect 5512 1797 5560 1803
rect 5608 1797 5640 1803
rect 6136 1797 6200 1803
rect 7224 1817 7256 1823
rect 1080 1777 1176 1783
rect 1192 1777 1336 1783
rect 1416 1777 2435 1783
rect 312 1757 360 1763
rect 488 1757 632 1763
rect 744 1757 936 1763
rect 1864 1757 1880 1763
rect 1912 1757 2008 1763
rect 2152 1757 2360 1763
rect 2429 1763 2435 1777
rect 2456 1777 4040 1783
rect 4120 1777 4136 1783
rect 4232 1777 4344 1783
rect 4520 1777 4744 1783
rect 4760 1777 4888 1783
rect 5032 1777 5192 1783
rect 5416 1777 5576 1783
rect 5640 1777 5752 1783
rect 5768 1777 6056 1783
rect 6072 1777 6088 1783
rect 6184 1777 6264 1783
rect 6296 1777 6424 1783
rect 6920 1777 7064 1783
rect 2429 1757 2472 1763
rect 2504 1757 2728 1763
rect 3064 1757 3256 1763
rect 3400 1757 3416 1763
rect 3432 1757 3496 1763
rect 3704 1757 3912 1763
rect 3992 1757 4792 1763
rect 4808 1757 4904 1763
rect 4936 1757 4968 1763
rect 4984 1757 5224 1763
rect 5400 1757 5480 1763
rect 5496 1757 5736 1763
rect 5752 1757 6232 1763
rect 6696 1757 7016 1763
rect 7320 1757 7368 1763
rect 7384 1757 7416 1763
rect 264 1737 312 1743
rect 792 1737 856 1743
rect 952 1737 1512 1743
rect 1656 1737 1976 1743
rect 1992 1737 2248 1743
rect 2472 1737 2504 1743
rect 2792 1737 2888 1743
rect 2920 1737 3096 1743
rect 3112 1737 3672 1743
rect 3688 1737 4008 1743
rect 4120 1737 4312 1743
rect 4392 1737 4552 1743
rect 4600 1737 4616 1743
rect 4712 1737 4760 1743
rect 4973 1737 4984 1743
rect 5128 1737 5304 1743
rect 5336 1737 5352 1743
rect 5384 1737 5432 1743
rect 5592 1737 5704 1743
rect 5896 1737 6408 1743
rect 6424 1737 6440 1743
rect 6472 1737 6520 1743
rect 6776 1737 6840 1743
rect 6952 1737 6984 1743
rect 7320 1737 7384 1743
rect 749 1728 755 1732
rect 136 1717 216 1723
rect 296 1717 488 1723
rect 632 1717 744 1723
rect 840 1717 888 1723
rect 1000 1717 1064 1723
rect 1304 1717 1448 1723
rect 1496 1717 1576 1723
rect 1608 1717 1784 1723
rect 1800 1717 1992 1723
rect 2008 1717 2040 1723
rect 2280 1717 3160 1723
rect 3192 1717 3523 1723
rect 344 1697 568 1703
rect 696 1697 824 1703
rect 872 1697 920 1703
rect 1000 1697 1048 1703
rect 1176 1697 1448 1703
rect 1464 1697 1496 1703
rect 1512 1697 1672 1703
rect 1688 1697 1720 1703
rect 1752 1697 1912 1703
rect 1928 1697 2552 1703
rect 2616 1697 2680 1703
rect 2712 1697 2904 1703
rect 3256 1697 3304 1703
rect 3352 1697 3384 1703
rect 3400 1697 3464 1703
rect 3517 1703 3523 1717
rect 3544 1717 3576 1723
rect 3672 1717 3912 1723
rect 3944 1717 4104 1723
rect 4136 1717 4184 1723
rect 4264 1717 4424 1723
rect 4584 1717 4632 1723
rect 4664 1717 4696 1723
rect 5000 1717 5080 1723
rect 5128 1717 5144 1723
rect 5512 1717 5672 1723
rect 5832 1717 6168 1723
rect 6184 1717 6296 1723
rect 6440 1717 6488 1723
rect 6616 1717 6760 1723
rect 6984 1717 7176 1723
rect 7288 1717 7368 1723
rect 6381 1708 6387 1712
rect 3517 1697 3528 1703
rect 3576 1697 3624 1703
rect 3688 1697 3752 1703
rect 3944 1697 4216 1703
rect 4232 1697 4328 1703
rect 4552 1697 4568 1703
rect 4680 1697 4691 1703
rect 4728 1697 4744 1703
rect 4856 1697 5032 1703
rect 5480 1697 5592 1703
rect 5640 1697 5736 1703
rect 5752 1697 5800 1703
rect 6056 1697 6104 1703
rect 6120 1697 6280 1703
rect 6472 1697 6600 1703
rect 7016 1697 7256 1703
rect 5197 1688 5203 1692
rect 1352 1677 1496 1683
rect 1512 1677 1544 1683
rect 1800 1677 1848 1683
rect 1864 1677 2072 1683
rect 3608 1677 4232 1683
rect 4264 1677 4312 1683
rect 4328 1677 4408 1683
rect 4792 1677 4824 1683
rect 5053 1677 5064 1683
rect 5544 1677 5752 1683
rect 6104 1677 6184 1683
rect 6232 1677 6376 1683
rect 6584 1677 6648 1683
rect 7192 1677 7352 1683
rect 1608 1657 2088 1663
rect 2440 1657 4616 1663
rect 4712 1657 4744 1663
rect 5736 1657 5816 1663
rect 5992 1657 6168 1663
rect 248 1637 264 1643
rect 2488 1637 2536 1643
rect 2552 1637 2584 1643
rect 2600 1637 2744 1643
rect 4344 1637 4376 1643
rect 4424 1637 4440 1643
rect 4456 1637 4872 1643
rect 5192 1637 5224 1643
rect 5800 1637 6072 1643
rect 6088 1637 6584 1643
rect 6824 1637 6856 1643
rect 6872 1637 7064 1643
rect 7080 1637 7128 1643
rect 7144 1637 7208 1643
rect 1848 1617 2104 1623
rect 2120 1617 2168 1623
rect 2184 1617 2376 1623
rect 2392 1617 2520 1623
rect 2536 1617 2744 1623
rect 2760 1617 2904 1623
rect 3224 1617 4584 1623
rect 4744 1617 5112 1623
rect 5464 1617 5720 1623
rect 5736 1617 5880 1623
rect 5976 1617 6472 1623
rect 6632 1597 6712 1603
rect 6728 1597 7272 1603
rect 264 1577 296 1583
rect 312 1577 616 1583
rect 2264 1577 3960 1583
rect 4152 1577 4264 1583
rect 4408 1577 4616 1583
rect 4632 1577 5048 1583
rect 5880 1577 5960 1583
rect 6376 1577 6408 1583
rect 6424 1577 6616 1583
rect 6632 1577 6872 1583
rect 7064 1577 7144 1583
rect 632 1557 1448 1563
rect 1464 1557 2232 1563
rect 2552 1557 3320 1563
rect 3352 1557 3640 1563
rect 3784 1557 4120 1563
rect 4152 1557 4424 1563
rect 4552 1557 4680 1563
rect 4744 1557 4904 1563
rect 6056 1557 6104 1563
rect 6712 1557 7048 1563
rect 184 1537 344 1543
rect 584 1537 600 1543
rect 2072 1537 2232 1543
rect 2776 1537 3080 1543
rect 3160 1537 3304 1543
rect 3736 1537 3864 1543
rect 4456 1537 4504 1543
rect 4680 1537 5016 1543
rect 5176 1537 5288 1543
rect 5304 1537 5480 1543
rect 5544 1537 5800 1543
rect 5880 1537 5992 1543
rect 6088 1537 6536 1543
rect 7032 1537 7112 1543
rect 248 1517 280 1523
rect 488 1517 744 1523
rect 760 1517 920 1523
rect 936 1517 1016 1523
rect 1048 1517 1080 1523
rect 1192 1517 1400 1523
rect 1576 1517 1624 1523
rect 2024 1517 2264 1523
rect 2712 1517 2776 1523
rect 2968 1517 2984 1523
rect 3096 1517 3336 1523
rect 3384 1517 3416 1523
rect 3864 1517 3928 1523
rect 4136 1517 4168 1523
rect 4184 1517 4472 1523
rect 4808 1517 4952 1523
rect 5432 1517 5544 1523
rect 5752 1517 5992 1523
rect 6216 1517 6648 1523
rect 6792 1517 6904 1523
rect 7112 1517 7224 1523
rect 4109 1508 4115 1512
rect 6061 1508 6067 1512
rect 24 1497 136 1503
rect 152 1497 200 1503
rect 568 1497 824 1503
rect 1096 1497 1256 1503
rect 1624 1497 1752 1503
rect 1944 1497 2120 1503
rect 2168 1497 2200 1503
rect 2216 1497 2232 1503
rect 2248 1497 2296 1503
rect 2360 1497 2392 1503
rect 2408 1497 2776 1503
rect 2792 1497 2824 1503
rect 2968 1497 3256 1503
rect 3288 1497 3320 1503
rect 3432 1497 3512 1503
rect 3624 1497 4008 1503
rect 4120 1497 4856 1503
rect 4888 1497 5064 1503
rect 5080 1497 5192 1503
rect 5288 1497 5512 1503
rect 5528 1497 5560 1503
rect 5848 1497 5976 1503
rect 5992 1497 6040 1503
rect 6072 1497 6088 1503
rect 6328 1497 6392 1503
rect 6616 1497 6680 1503
rect 6920 1497 7016 1503
rect 7096 1497 7128 1503
rect 7144 1497 7256 1503
rect 7272 1497 7336 1503
rect 7368 1497 7384 1503
rect 136 1477 232 1483
rect 440 1477 568 1483
rect 664 1477 952 1483
rect 1416 1477 2440 1483
rect 2984 1477 3016 1483
rect 3032 1477 3208 1483
rect 3592 1477 3672 1483
rect 3848 1477 3944 1483
rect 3976 1477 4344 1483
rect 4472 1477 4483 1483
rect 4568 1477 4712 1483
rect 5064 1477 5096 1483
rect 5272 1477 5576 1483
rect 5704 1477 5880 1483
rect 5944 1477 5992 1483
rect 6200 1477 6440 1483
rect 6728 1477 6792 1483
rect 7224 1477 7368 1483
rect 632 1457 872 1463
rect 1768 1457 1944 1463
rect 1960 1457 1992 1463
rect 2264 1457 2536 1463
rect 2584 1457 2856 1463
rect 3016 1457 3112 1463
rect 3752 1457 4072 1463
rect 4280 1457 4296 1463
rect 4328 1457 4584 1463
rect 4744 1457 4760 1463
rect 4840 1457 5096 1463
rect 5112 1457 5176 1463
rect 5400 1457 5528 1463
rect 5560 1457 5624 1463
rect 5656 1457 5752 1463
rect 5928 1457 6216 1463
rect 6280 1457 6344 1463
rect 6728 1457 6920 1463
rect 7048 1457 7080 1463
rect 7304 1457 7336 1463
rect 7384 1457 7395 1463
rect 552 1437 680 1443
rect 1160 1437 1368 1443
rect 1544 1437 1640 1443
rect 2072 1437 2328 1443
rect 2552 1437 2648 1443
rect 2712 1437 3128 1443
rect 3144 1437 3336 1443
rect 3464 1437 3640 1443
rect 4008 1437 4312 1443
rect 4376 1437 5880 1443
rect 6232 1437 6712 1443
rect 6760 1437 6776 1443
rect 6792 1437 6824 1443
rect 840 1417 888 1423
rect 904 1417 1464 1423
rect 1480 1417 1976 1423
rect 1096 1397 1160 1403
rect 1208 1397 1336 1403
rect 1352 1397 1560 1403
rect 3224 1417 3352 1423
rect 3368 1417 3896 1423
rect 4072 1417 4088 1423
rect 3608 1397 3640 1403
rect 3672 1397 4024 1403
rect 4264 1417 4440 1423
rect 4664 1417 4824 1423
rect 4600 1397 4792 1403
rect 4936 1397 4968 1403
rect 5272 1397 5448 1403
rect 6456 1417 6744 1423
rect 6568 1397 6792 1403
rect 6808 1397 7064 1403
rect 7080 1397 7176 1403
rect 7229 1388 7235 1392
rect 200 1377 296 1383
rect 312 1377 680 1383
rect 760 1377 1416 1383
rect 1448 1377 1464 1383
rect 1480 1377 1512 1383
rect 1560 1377 1592 1383
rect 1816 1377 2024 1383
rect 2584 1377 2952 1383
rect 3448 1377 3480 1383
rect 3528 1377 4008 1383
rect 4056 1377 4664 1383
rect 5384 1377 5416 1383
rect 5608 1377 5816 1383
rect 5848 1377 6936 1383
rect 7096 1377 7144 1383
rect 7160 1377 7224 1383
rect 280 1357 408 1363
rect 424 1357 456 1363
rect 472 1357 520 1363
rect 952 1357 1032 1363
rect 1416 1357 1816 1363
rect 1832 1357 1848 1363
rect 1912 1357 1944 1363
rect 2008 1357 2248 1363
rect 2520 1357 2840 1363
rect 3272 1357 3368 1363
rect 3592 1357 3816 1363
rect 3832 1357 3944 1363
rect 4024 1357 4248 1363
rect 4280 1357 4728 1363
rect 5128 1357 5176 1363
rect 5432 1357 5752 1363
rect 5912 1357 5944 1363
rect 5960 1357 6120 1363
rect 6136 1357 6200 1363
rect 6216 1357 6456 1363
rect 6760 1357 7128 1363
rect 7144 1357 7192 1363
rect 72 1337 200 1343
rect 216 1337 488 1343
rect 600 1337 728 1343
rect 744 1337 808 1343
rect 1592 1337 2808 1343
rect 2893 1343 2899 1352
rect 2888 1337 2899 1343
rect 2909 1337 2984 1343
rect 88 1317 216 1323
rect 344 1317 376 1323
rect 856 1317 968 1323
rect 1160 1317 1208 1323
rect 1432 1317 1528 1323
rect 1720 1317 1784 1323
rect 1896 1317 2104 1323
rect 2312 1317 2376 1323
rect 2488 1317 2520 1323
rect 2909 1323 2915 1337
rect 3080 1337 3640 1343
rect 4296 1337 4504 1343
rect 4696 1337 4840 1343
rect 4904 1337 5080 1343
rect 5096 1337 5208 1343
rect 5224 1337 5352 1343
rect 5512 1337 5656 1343
rect 5672 1337 5864 1343
rect 6376 1337 6424 1343
rect 6440 1337 6680 1343
rect 6696 1337 6744 1343
rect 6872 1337 6904 1343
rect 6952 1337 6968 1343
rect 3069 1328 3075 1332
rect 4605 1328 4611 1332
rect 2712 1317 2915 1323
rect 2968 1317 3048 1323
rect 3112 1317 3224 1323
rect 3240 1317 3272 1323
rect 3288 1317 3384 1323
rect 3512 1317 3752 1323
rect 3768 1317 3880 1323
rect 3912 1317 3928 1323
rect 3976 1317 3992 1323
rect 4008 1317 4024 1323
rect 4056 1317 4072 1323
rect 4184 1317 4312 1323
rect 4408 1317 4456 1323
rect 4472 1317 4552 1323
rect 4648 1317 4680 1323
rect 5368 1317 5384 1323
rect 5400 1317 5464 1323
rect 5656 1317 5768 1323
rect 5784 1317 6088 1323
rect 6312 1317 6408 1323
rect 6504 1317 6552 1323
rect 6568 1317 6616 1323
rect 6648 1317 6696 1323
rect 6968 1317 6984 1323
rect 216 1297 264 1303
rect 296 1297 504 1303
rect 520 1297 552 1303
rect 568 1297 600 1303
rect 968 1297 984 1303
rect 1000 1297 1016 1303
rect 1496 1297 1704 1303
rect 1768 1297 1832 1303
rect 1896 1297 1960 1303
rect 2168 1297 2840 1303
rect 2872 1297 2984 1303
rect 3000 1297 3032 1303
rect 3048 1297 3256 1303
rect 3293 1297 3512 1303
rect 408 1277 472 1283
rect 488 1277 1064 1283
rect 1080 1277 1880 1283
rect 1992 1277 2920 1283
rect 3293 1283 3299 1297
rect 3848 1297 4120 1303
rect 4488 1297 4504 1303
rect 4568 1297 4760 1303
rect 5528 1297 5736 1303
rect 5768 1297 5816 1303
rect 6120 1297 6152 1303
rect 6168 1297 6264 1303
rect 6280 1297 6328 1303
rect 6680 1297 6728 1303
rect 6797 1297 6840 1303
rect 3160 1277 3299 1283
rect 3320 1277 3496 1283
rect 3512 1277 3640 1283
rect 3880 1277 3912 1283
rect 3928 1277 3960 1283
rect 4008 1277 4056 1283
rect 4088 1277 4200 1283
rect 4333 1277 4344 1283
rect 4520 1277 4680 1283
rect 5672 1277 5784 1283
rect 6488 1277 6536 1283
rect 6552 1277 6584 1283
rect 6797 1283 6803 1297
rect 6696 1277 6803 1283
rect 6824 1277 7048 1283
rect 504 1257 2856 1263
rect 3944 1257 3992 1263
rect 4024 1257 4104 1263
rect 5592 1257 5848 1263
rect 6584 1257 6760 1263
rect 3816 1237 4232 1243
rect 4264 1237 4440 1243
rect 4456 1237 4552 1243
rect 5752 1237 6632 1243
rect 1736 1217 2312 1223
rect 2936 1217 2968 1223
rect 1608 1197 2216 1203
rect 3720 1217 3768 1223
rect 4376 1217 4440 1223
rect 4488 1217 4520 1223
rect 3704 1197 4504 1203
rect 4552 1197 4888 1203
rect 5560 1217 5672 1223
rect 5720 1217 5880 1223
rect 6040 1217 6120 1223
rect 6136 1217 6168 1223
rect 6392 1217 6504 1223
rect 6520 1217 6968 1223
rect 5496 1197 5656 1203
rect 5672 1197 6216 1203
rect 6248 1197 7000 1203
rect 328 1177 360 1183
rect 376 1177 568 1183
rect 1240 1177 1496 1183
rect 1512 1177 1592 1183
rect 2040 1177 2488 1183
rect 2504 1177 3752 1183
rect 4424 1177 4824 1183
rect 5000 1177 5624 1183
rect 5976 1177 6024 1183
rect 6568 1177 6904 1183
rect 7208 1177 7224 1183
rect 712 1157 1288 1163
rect 1304 1157 1352 1163
rect 1592 1157 1608 1163
rect 1640 1157 1672 1163
rect 2072 1157 2147 1163
rect 200 1137 296 1143
rect 312 1137 520 1143
rect 568 1137 1160 1143
rect 1192 1137 1288 1143
rect 1320 1137 1336 1143
rect 1352 1137 1432 1143
rect 1448 1137 1528 1143
rect 1544 1137 2120 1143
rect 2141 1143 2147 1157
rect 2216 1157 2248 1163
rect 2264 1157 2584 1163
rect 2600 1157 2808 1163
rect 2888 1157 2936 1163
rect 3224 1157 3320 1163
rect 3752 1157 3832 1163
rect 3896 1157 3976 1163
rect 4120 1157 4360 1163
rect 4392 1157 4440 1163
rect 4472 1157 4536 1163
rect 4568 1157 4664 1163
rect 4808 1157 5000 1163
rect 5432 1157 6072 1163
rect 6200 1157 6376 1163
rect 6392 1157 6408 1163
rect 6440 1157 6520 1163
rect 6936 1157 7192 1163
rect 2141 1137 2200 1143
rect 2280 1137 4296 1143
rect 4328 1137 4360 1143
rect 4376 1137 4392 1143
rect 4408 1137 4792 1143
rect 5480 1137 5640 1143
rect 5880 1137 6264 1143
rect 6328 1137 6392 1143
rect 6504 1137 6584 1143
rect 6632 1137 6840 1143
rect 6952 1137 6984 1143
rect 216 1117 264 1123
rect 744 1117 952 1123
rect 1080 1117 1096 1123
rect 1112 1117 1208 1123
rect 1224 1117 1384 1123
rect 1400 1117 1448 1123
rect 1464 1117 2008 1123
rect 2088 1117 2248 1123
rect 2280 1117 2296 1123
rect 2856 1117 2952 1123
rect 3080 1117 3272 1123
rect 3656 1117 3720 1123
rect 3832 1117 3848 1123
rect 3880 1117 3928 1123
rect 4072 1117 4083 1123
rect 4104 1117 4280 1123
rect 4296 1117 4392 1123
rect 4536 1117 4696 1123
rect 4952 1117 4963 1123
rect 5304 1117 5432 1123
rect 5480 1117 5528 1123
rect 5752 1117 5816 1123
rect 5928 1117 6040 1123
rect 6376 1117 6456 1123
rect 6520 1117 6616 1123
rect 6696 1117 6792 1123
rect 7032 1117 7080 1123
rect 7144 1117 7160 1123
rect 7352 1117 7368 1123
rect 88 1097 216 1103
rect 344 1097 632 1103
rect 696 1097 888 1103
rect 968 1097 984 1103
rect 1208 1097 1320 1103
rect 1336 1097 1416 1103
rect 1432 1097 2072 1103
rect 2120 1097 2328 1103
rect 2344 1097 2440 1103
rect 2472 1097 2483 1103
rect 2728 1097 2872 1103
rect 3272 1097 3304 1103
rect 3608 1097 3784 1103
rect 3832 1097 3864 1103
rect 4104 1097 4136 1103
rect 4173 1097 4184 1103
rect 4280 1097 4520 1103
rect 4568 1097 4712 1103
rect 4872 1097 4936 1103
rect 5160 1097 5240 1103
rect 5288 1097 5320 1103
rect 5336 1097 5448 1103
rect 5528 1097 5688 1103
rect 5752 1097 5816 1103
rect 6136 1097 6200 1103
rect 6216 1097 6408 1103
rect 6456 1097 6568 1103
rect 6648 1097 6888 1103
rect 6904 1097 6952 1103
rect 7048 1097 7064 1103
rect 7144 1097 7192 1103
rect 7272 1097 7320 1103
rect 7368 1097 7384 1103
rect 136 1077 376 1083
rect 632 1077 936 1083
rect 1000 1077 1032 1083
rect 1176 1077 1192 1083
rect 1464 1077 1544 1083
rect 1688 1077 1784 1083
rect 1848 1077 1928 1083
rect 2072 1077 2200 1083
rect 2472 1077 2920 1083
rect 3128 1077 3560 1083
rect 3576 1077 3608 1083
rect 3800 1077 3896 1083
rect 4008 1077 4040 1083
rect 4072 1077 4088 1083
rect 4109 1077 4408 1083
rect 1069 1068 1075 1072
rect 216 1057 376 1063
rect 824 1057 888 1063
rect 936 1057 1000 1063
rect 1032 1057 1048 1063
rect 1080 1057 1400 1063
rect 1992 1057 2088 1063
rect 2360 1057 2392 1063
rect 2440 1057 2488 1063
rect 2920 1057 2984 1063
rect 3688 1057 3768 1063
rect 3800 1057 3816 1063
rect 4109 1063 4115 1077
rect 4472 1077 4632 1083
rect 4648 1077 4696 1083
rect 4712 1077 4760 1083
rect 4952 1077 4968 1083
rect 5352 1077 5560 1083
rect 5800 1077 5896 1083
rect 6040 1077 6824 1083
rect 6840 1077 7144 1083
rect 7160 1077 7320 1083
rect 4909 1068 4915 1072
rect 3976 1057 4115 1063
rect 4136 1057 4147 1063
rect 4264 1057 4312 1063
rect 4520 1057 4760 1063
rect 4776 1057 4888 1063
rect 5048 1057 5208 1063
rect 5896 1057 6392 1063
rect 6408 1057 6504 1063
rect 6584 1057 7208 1063
rect 7224 1057 7272 1063
rect 728 1037 1176 1043
rect 1448 1037 1608 1043
rect 1720 1037 1896 1043
rect 1912 1037 2872 1043
rect 3000 1037 3576 1043
rect 3608 1037 4376 1043
rect 4392 1037 4536 1043
rect 4696 1037 4808 1043
rect 4872 1037 5928 1043
rect 6184 1037 6200 1043
rect 6280 1037 6392 1043
rect 6600 1037 6664 1043
rect 6856 1037 7000 1043
rect 600 1017 1480 1023
rect 376 997 392 1003
rect 536 997 840 1003
rect 872 997 984 1003
rect 1272 997 2147 1003
rect 2312 1017 2584 1023
rect 2712 1017 3016 1023
rect 3032 1017 3128 1023
rect 3144 1017 3192 1023
rect 3992 1017 4008 1023
rect 584 977 632 983
rect 728 977 824 983
rect 920 977 1016 983
rect 1208 977 1384 983
rect 1416 977 1544 983
rect 1581 977 1960 983
rect 200 957 296 963
rect 312 957 440 963
rect 488 957 680 963
rect 696 957 744 963
rect 909 957 1240 963
rect 909 943 915 957
rect 1581 963 1587 977
rect 2008 977 2024 983
rect 2141 983 2147 997
rect 2968 997 3000 1003
rect 3560 997 3592 1003
rect 4504 1017 4616 1023
rect 4760 1017 4872 1023
rect 4888 1017 5064 1023
rect 5624 1017 5768 1023
rect 6008 1017 6184 1023
rect 4424 997 4531 1003
rect 2141 977 2152 983
rect 2184 977 2312 983
rect 2344 977 2456 983
rect 2584 977 2760 983
rect 3176 977 3352 983
rect 3368 977 3544 983
rect 3864 977 4488 983
rect 4525 983 4531 997
rect 4552 997 4648 1003
rect 4936 997 6200 1003
rect 6568 1017 6707 1023
rect 6296 997 6680 1003
rect 6701 1003 6707 1017
rect 6760 1017 7032 1023
rect 7112 1017 7224 1023
rect 6701 997 6808 1003
rect 6824 997 7064 1003
rect 7080 997 7288 1003
rect 4525 977 4808 983
rect 4984 977 5080 983
rect 5096 977 5240 983
rect 5384 977 6440 983
rect 6733 977 6744 983
rect 6765 977 6904 983
rect 1464 957 1587 963
rect 1608 957 1848 963
rect 1864 957 2008 963
rect 2024 957 2280 963
rect 2296 957 2392 963
rect 3064 957 3368 963
rect 3629 957 3848 963
rect 632 937 915 943
rect 936 937 968 943
rect 1192 937 1240 943
rect 1368 937 1416 943
rect 1576 937 1784 943
rect 1816 937 2120 943
rect 2184 937 2280 943
rect 2312 937 2408 943
rect 2424 937 2504 943
rect 3629 943 3635 957
rect 3933 957 4072 963
rect 2968 937 3635 943
rect 3645 937 3656 943
rect 88 917 232 923
rect 520 917 552 923
rect 568 917 632 923
rect 808 917 936 923
rect 1160 917 1304 923
rect 1320 917 1368 923
rect 1432 917 1496 923
rect 1624 917 1672 923
rect 1912 917 2120 923
rect 2136 917 2296 923
rect 2312 917 2360 923
rect 2392 917 2424 923
rect 2712 917 2792 923
rect 2872 917 2968 923
rect 3064 917 3096 923
rect 3645 923 3651 937
rect 3933 943 3939 957
rect 4120 957 4232 963
rect 4264 957 4504 963
rect 5112 957 5176 963
rect 5192 957 5368 963
rect 5656 957 5688 963
rect 5768 957 5976 963
rect 6056 957 6424 963
rect 6493 957 6568 963
rect 3848 937 3939 943
rect 3960 937 4456 943
rect 4536 937 4552 943
rect 4648 937 4840 943
rect 5032 937 5080 943
rect 5496 937 5512 943
rect 5576 937 5704 943
rect 5816 937 5848 943
rect 5992 937 6200 943
rect 6493 943 6499 957
rect 6765 963 6771 977
rect 6984 977 7112 983
rect 7320 977 7400 983
rect 6648 957 6771 963
rect 6792 957 6984 963
rect 7000 957 7304 963
rect 6216 937 6499 943
rect 6520 937 6888 943
rect 6904 937 6984 943
rect 7016 937 7224 943
rect 3512 917 3651 923
rect 3672 917 3736 923
rect 3864 917 3912 923
rect 3944 917 4056 923
rect 4088 917 4120 923
rect 4216 917 4264 923
rect 4328 917 4488 923
rect 4536 917 4584 923
rect 4696 917 4760 923
rect 4824 917 4904 923
rect 4952 917 5112 923
rect 5320 917 5400 923
rect 5544 917 5800 923
rect 5848 917 5992 923
rect 6168 917 6184 923
rect 6216 917 6296 923
rect 6504 917 6520 923
rect 6904 917 6968 923
rect 232 897 264 903
rect 296 897 328 903
rect 840 897 920 903
rect 936 897 984 903
rect 1240 897 1288 903
rect 1336 897 1560 903
rect 1592 897 1608 903
rect 1656 897 2104 903
rect 2408 897 2440 903
rect 2760 897 2792 903
rect 2808 897 2840 903
rect 3080 897 3224 903
rect 3400 897 3432 903
rect 3656 897 3688 903
rect 3816 897 3864 903
rect 4008 897 4184 903
rect 4248 897 4328 903
rect 4536 897 4552 903
rect 4760 897 4776 903
rect 5416 897 5448 903
rect 5592 897 6456 903
rect 7224 897 7352 903
rect 4429 888 4435 892
rect 1192 877 1672 883
rect 1960 877 2328 883
rect 2600 877 2936 883
rect 3064 877 3112 883
rect 3640 877 3672 883
rect 3784 877 3832 883
rect 3912 877 3992 883
rect 4008 877 4024 883
rect 4040 877 4120 883
rect 4280 877 4408 883
rect 5032 877 5720 883
rect 5736 877 6744 883
rect 1592 857 1640 863
rect 1672 857 1848 863
rect 2008 857 2216 863
rect 2248 857 2536 863
rect 3752 857 3960 863
rect 3992 857 4248 863
rect 4360 857 4440 863
rect 5048 857 5112 863
rect 5480 857 5960 863
rect 5992 857 7080 863
rect 936 837 1192 843
rect 1368 837 2056 843
rect 2392 837 3907 843
rect 1720 817 2072 823
rect 2088 817 2232 823
rect 2280 817 3144 823
rect 3901 823 3907 837
rect 3928 837 4376 843
rect 5080 837 5267 843
rect 1208 797 1384 803
rect 1400 797 1928 803
rect 2040 797 2136 803
rect 3901 817 4312 823
rect 5261 823 5267 837
rect 3768 797 4056 803
rect 4072 797 4920 803
rect 5261 817 5560 823
rect 6024 817 6728 823
rect 5272 797 7384 803
rect 1128 777 1416 783
rect 2552 777 2600 783
rect 2632 777 2744 783
rect 3720 777 3848 783
rect 3912 777 4024 783
rect 5176 777 5448 783
rect 472 757 968 763
rect 1000 757 1400 763
rect 1416 757 1464 763
rect 1512 757 2216 763
rect 2504 757 2904 763
rect 3752 757 3848 763
rect 4008 757 4136 763
rect 4152 757 4280 763
rect 4952 757 5112 763
rect 5448 757 6344 763
rect 824 737 936 743
rect 1032 737 1128 743
rect 1624 737 1800 743
rect 1816 737 1832 743
rect 1992 737 2008 743
rect 2840 737 3288 743
rect 3432 737 3560 743
rect 3848 737 4088 743
rect 4136 737 4248 743
rect 4600 737 4904 743
rect 5016 737 5032 743
rect 5112 737 5160 743
rect 5176 737 5240 743
rect 5672 737 5880 743
rect 5992 737 6120 743
rect 6408 737 6568 743
rect 6712 737 6888 743
rect 6920 737 6968 743
rect 6984 737 7096 743
rect 56 717 136 723
rect 456 717 520 723
rect 536 717 584 723
rect 920 717 1016 723
rect 1528 717 1576 723
rect 2328 717 2360 723
rect 2808 717 2856 723
rect 3544 717 3640 723
rect 3752 717 3816 723
rect 3864 717 4104 723
rect 4248 717 4328 723
rect 4344 717 4392 723
rect 4680 717 5000 723
rect 5016 717 5048 723
rect 5096 717 5112 723
rect 5560 717 5576 723
rect 5592 717 5624 723
rect 6040 717 6232 723
rect 6328 717 6392 723
rect 6440 717 6760 723
rect 7048 717 7144 723
rect 56 697 216 703
rect 344 697 472 703
rect 504 697 568 703
rect 600 697 616 703
rect 648 697 1032 703
rect 1048 697 1064 703
rect 1080 697 1272 703
rect 1592 697 1672 703
rect 1976 697 2024 703
rect 2424 697 2472 703
rect 2488 697 2552 703
rect 2872 697 3176 703
rect 3480 697 3560 703
rect 3576 697 3608 703
rect 3624 697 3736 703
rect 3848 697 3896 703
rect 4056 697 4120 703
rect 4392 697 4520 703
rect 4632 697 4664 703
rect 5064 697 5352 703
rect 5608 697 5704 703
rect 6024 697 6088 703
rect 6104 697 6120 703
rect 6392 697 6424 703
rect 6456 697 6680 703
rect 7144 697 7176 703
rect 472 677 616 683
rect 696 677 744 683
rect 920 677 1080 683
rect 1224 677 1288 683
rect 1304 677 1320 683
rect 1384 677 1496 683
rect 2376 677 2664 683
rect 2904 677 2968 683
rect 2984 677 3064 683
rect 3288 677 3400 683
rect 3560 677 3720 683
rect 3816 677 4040 683
rect 4120 677 4264 683
rect 4408 677 4600 683
rect 4680 677 4824 683
rect 4984 677 5096 683
rect 5128 677 5208 683
rect 5608 677 5928 683
rect 5944 677 5960 683
rect 5976 677 6280 683
rect 6296 677 6648 683
rect 6664 677 6776 683
rect 7032 677 7288 683
rect 440 657 936 663
rect 952 657 984 663
rect 2088 657 2120 663
rect 2360 657 2504 663
rect 3384 657 3544 663
rect 3720 657 3784 663
rect 3864 657 4152 663
rect 4488 657 4776 663
rect 4936 657 6904 663
rect 7192 657 7208 663
rect 56 637 248 643
rect 264 637 632 643
rect 968 637 1160 643
rect 1176 637 1256 643
rect 1640 637 2040 643
rect 3736 637 3784 643
rect 3800 637 3976 643
rect 4312 637 4408 643
rect 4584 637 4984 643
rect 5144 637 5352 643
rect 5464 637 5512 643
rect 7048 637 7256 643
rect 584 617 600 623
rect 312 597 344 603
rect 360 597 456 603
rect 472 597 680 603
rect 1800 597 1864 603
rect 1880 597 2008 603
rect 2504 617 2552 623
rect 2616 617 2792 623
rect 4280 617 4392 623
rect 4648 617 5528 623
rect 4424 597 4680 603
rect 5400 597 5432 603
rect 5464 597 5608 603
rect 5624 597 5704 603
rect 5800 597 5848 603
rect 6824 617 6920 623
rect 6936 617 7192 623
rect 216 577 584 583
rect 1768 577 1832 583
rect 1848 577 1880 583
rect 2072 577 2168 583
rect 2184 577 2424 583
rect 2792 577 2840 583
rect 2856 577 2920 583
rect 3880 577 3896 583
rect 3944 577 4056 583
rect 4072 577 4195 583
rect 184 557 488 563
rect 552 557 584 563
rect 760 557 952 563
rect 968 557 1512 563
rect 1656 557 1800 563
rect 1960 557 2072 563
rect 2093 557 2136 563
rect 72 537 376 543
rect 392 537 616 543
rect 632 537 712 543
rect 1528 537 1768 543
rect 1784 537 2056 543
rect 2093 543 2099 557
rect 2312 557 2600 563
rect 3096 557 3192 563
rect 3208 557 3416 563
rect 3592 557 3768 563
rect 3912 557 4104 563
rect 4189 563 4195 577
rect 4216 577 4296 583
rect 4328 577 4568 583
rect 4680 577 4856 583
rect 4872 577 4952 583
rect 5357 577 5768 583
rect 4189 557 4312 563
rect 4568 557 4696 563
rect 4888 557 4920 563
rect 5048 557 5224 563
rect 5357 563 5363 577
rect 5784 577 6136 583
rect 7208 577 7224 583
rect 5256 557 5363 563
rect 5400 557 5795 563
rect 2088 537 2099 543
rect 2136 537 2296 543
rect 2520 537 2680 543
rect 2920 537 2984 543
rect 3000 537 3224 543
rect 3448 537 3720 543
rect 3736 537 3768 543
rect 3880 537 3944 543
rect 4120 537 4152 543
rect 4344 537 4440 543
rect 4488 537 4520 543
rect 4648 537 4739 543
rect 1309 528 1315 532
rect 4733 528 4739 537
rect 4888 537 5112 543
rect 5128 537 5336 543
rect 5352 537 5512 543
rect 5528 537 5544 543
rect 5789 543 5795 557
rect 5992 557 6168 563
rect 6392 557 6456 563
rect 7176 557 7432 563
rect 5789 537 6072 543
rect 6200 537 6440 543
rect 6456 537 6680 543
rect 7144 537 7208 543
rect 6749 528 6755 532
rect 40 517 152 523
rect 168 517 472 523
rect 504 517 648 523
rect 728 517 744 523
rect 808 517 1000 523
rect 1112 517 1240 523
rect 1704 517 1976 523
rect 1992 517 2232 523
rect 2472 517 2568 523
rect 2664 517 2728 523
rect 2824 517 3144 523
rect 3160 517 3256 523
rect 3304 517 3528 523
rect 3720 517 3816 523
rect 4536 517 4584 523
rect 4600 517 4632 523
rect 4920 517 5240 523
rect 5336 517 6088 523
rect 6120 517 6360 523
rect 6376 517 6584 523
rect 7016 517 7048 523
rect 7064 517 7112 523
rect 7128 517 7320 523
rect 7448 517 7491 523
rect 3869 508 3875 512
rect 24 497 232 503
rect 264 497 392 503
rect 488 497 552 503
rect 568 497 632 503
rect 952 497 1016 503
rect 1096 497 1336 503
rect 2488 497 2504 503
rect 2664 497 2744 503
rect 2936 497 2968 503
rect 3640 497 3816 503
rect 4120 497 4392 503
rect 4552 497 4792 503
rect 4808 497 4840 503
rect 4856 497 4984 503
rect 5224 497 5288 503
rect 5304 497 5416 503
rect 5576 497 5656 503
rect 5848 497 5976 503
rect 5992 497 6040 503
rect 6056 497 6120 503
rect 6152 497 6200 503
rect 6376 497 6600 503
rect 6632 497 6680 503
rect 6984 497 7016 503
rect 7048 497 7080 503
rect 7128 497 7304 503
rect 376 477 440 483
rect 456 477 504 483
rect 648 477 664 483
rect 984 477 1432 483
rect 2600 477 2760 483
rect 2776 477 2936 483
rect 2984 477 4296 483
rect 4312 477 5768 483
rect 6120 477 6296 483
rect 6328 477 6392 483
rect 6408 477 6424 483
rect 6824 477 7144 483
rect 7160 477 7288 483
rect 392 457 520 463
rect 1848 457 3432 463
rect 3448 457 5464 463
rect 6248 457 6808 463
rect 6888 457 7064 463
rect 2952 437 3848 443
rect 4264 437 4872 443
rect 5384 437 5576 443
rect 5816 437 6280 443
rect 1672 397 1816 403
rect 1832 397 2120 403
rect 2136 397 2552 403
rect 3048 397 3144 403
rect 3352 417 3480 423
rect 3496 417 3704 423
rect 3736 417 3992 423
rect 4616 417 4824 423
rect 3240 397 3704 403
rect 3816 397 4072 403
rect 4088 397 4104 403
rect 5784 417 6824 423
rect 328 377 408 383
rect 584 377 600 383
rect 1416 377 1560 383
rect 1576 377 3304 383
rect 3320 377 5656 383
rect 840 357 1032 363
rect 1144 357 1272 363
rect 2952 357 2984 363
rect 3112 357 3240 363
rect 3256 357 3288 363
rect 3304 357 3672 363
rect 3704 357 3912 363
rect 4040 357 4312 363
rect 4392 357 4408 363
rect 5608 357 5720 363
rect 6088 357 6424 363
rect 488 337 680 343
rect 744 337 1016 343
rect 1032 337 1096 343
rect 1400 337 1480 343
rect 1864 337 1960 343
rect 2360 337 2456 343
rect 2760 337 2872 343
rect 3000 337 3016 343
rect 3032 337 3176 343
rect 3432 337 3608 343
rect 3624 337 3752 343
rect 4088 337 4328 343
rect 4344 337 4376 343
rect 4392 337 5176 343
rect 5720 337 5736 343
rect 5752 337 5816 343
rect 6312 337 6440 343
rect 6472 337 6648 343
rect 136 317 184 323
rect 200 317 536 323
rect 616 317 712 323
rect 824 317 888 323
rect 1288 317 1560 323
rect 1880 317 1928 323
rect 1944 317 2360 323
rect 2376 317 2424 323
rect 2648 317 2776 323
rect 2920 317 2968 323
rect 3096 317 3320 323
rect 3336 317 3384 323
rect 3432 317 4648 323
rect 5192 317 5432 323
rect 5448 317 5464 323
rect 5704 317 6008 323
rect 6024 317 6280 323
rect 6392 317 6520 323
rect 6728 317 6984 323
rect 7048 317 7208 323
rect 7304 317 7491 323
rect 5133 308 5139 312
rect 104 297 232 303
rect 600 297 680 303
rect 776 297 824 303
rect 968 297 1080 303
rect 1272 297 1352 303
rect 1368 297 1480 303
rect 1496 297 1528 303
rect 1752 297 1880 303
rect 1976 297 2056 303
rect 2264 297 2376 303
rect 2792 297 2824 303
rect 2840 297 3080 303
rect 3112 297 3240 303
rect 3400 297 3480 303
rect 3832 297 3880 303
rect 3896 297 4152 303
rect 4184 297 4296 303
rect 4440 297 4632 303
rect 4648 297 4744 303
rect 4904 297 4920 303
rect 5032 297 5080 303
rect 5352 297 5400 303
rect 5432 297 5448 303
rect 5464 297 5624 303
rect 5688 297 5832 303
rect 5944 297 5976 303
rect 6008 297 6168 303
rect 6360 297 6392 303
rect 6456 297 6664 303
rect 6712 297 6872 303
rect 6936 297 6952 303
rect 7048 297 7176 303
rect 7336 297 7368 303
rect 136 277 264 283
rect 1032 277 1144 283
rect 1416 277 1688 283
rect 2296 277 2360 283
rect 2376 277 2584 283
rect 3672 277 3784 283
rect 3800 277 3832 283
rect 4104 277 4168 283
rect 4184 277 4264 283
rect 4280 277 4376 283
rect 4536 277 4680 283
rect 4696 277 4760 283
rect 4776 277 4856 283
rect 5208 277 5448 283
rect 5544 277 5672 283
rect 5688 277 5800 283
rect 5832 277 5912 283
rect 5928 277 6024 283
rect 6152 277 6168 283
rect 6328 277 6440 283
rect 6888 277 7192 283
rect 7336 277 7384 283
rect 3496 257 3816 263
rect 3880 257 4200 263
rect 4376 257 4504 263
rect 4968 257 5000 263
rect 5384 257 5880 263
rect 5896 257 6088 263
rect 6104 257 6152 263
rect 6168 257 6376 263
rect 6392 257 6488 263
rect 2952 237 3016 243
rect 3032 237 3400 243
rect 3992 237 4120 243
rect 4136 237 4232 243
rect 5592 237 6920 243
rect 6952 237 7000 243
rect 2584 217 2680 223
rect 2696 217 2904 223
rect 2920 217 3112 223
rect 3608 217 3640 223
rect 2712 197 2920 203
rect 3144 197 3320 203
rect 3416 197 3544 203
rect 3576 197 3624 203
rect 4264 197 4536 203
rect 4552 197 4616 203
rect 6584 217 6952 223
rect 7032 217 7336 223
rect 7133 188 7139 192
rect 472 177 648 183
rect 952 177 1016 183
rect 1112 177 1192 183
rect 1480 177 1832 183
rect 2232 177 2296 183
rect 2312 177 2536 183
rect 3016 177 3112 183
rect 3128 177 3672 183
rect 4008 177 4104 183
rect 4120 177 4872 183
rect 5224 177 5496 183
rect 5528 177 5544 183
rect 6136 177 6504 183
rect 7288 177 7384 183
rect 760 157 824 163
rect 840 157 952 163
rect 968 157 1336 163
rect 2696 157 2712 163
rect 3336 157 3528 163
rect 3544 157 3656 163
rect 3672 157 3848 163
rect 3864 157 3944 163
rect 4456 157 4488 163
rect 4728 157 6184 163
rect 6200 157 6248 163
rect 6552 157 6808 163
rect 6824 157 6968 163
rect 7149 157 7155 172
rect 7229 148 7235 152
rect 632 137 776 143
rect 840 137 984 143
rect 1096 137 1192 143
rect 1240 137 1288 143
rect 1496 137 1800 143
rect 1816 137 1848 143
rect 1912 137 2120 143
rect 2776 137 2808 143
rect 2904 137 3048 143
rect 3272 137 3448 143
rect 3560 137 4616 143
rect 4632 137 4728 143
rect 4968 137 5048 143
rect 5464 137 5576 143
rect 5608 137 5832 143
rect 6152 137 6200 143
rect 6520 137 6744 143
rect 5085 128 5091 132
rect 7197 128 7203 132
rect 296 117 392 123
rect 600 117 680 123
rect 984 117 1048 123
rect 1064 117 1496 123
rect 1560 117 1704 123
rect 1896 117 1960 123
rect 2280 117 2408 123
rect 2568 117 2744 123
rect 3048 117 3080 123
rect 3240 117 3320 123
rect 3608 117 3656 123
rect 4072 117 4216 123
rect 4456 117 4600 123
rect 4808 117 4952 123
rect 5352 117 5400 123
rect 5784 117 5816 123
rect 5832 117 6168 123
rect 6616 117 6648 123
rect 6664 117 6936 123
rect 6952 117 7032 123
rect 5037 108 5043 112
rect 328 97 392 103
rect 440 97 680 103
rect 696 97 728 103
rect 1272 97 1288 103
rect 1512 97 1544 103
rect 1880 97 2184 103
rect 2200 97 2280 103
rect 2296 97 2312 103
rect 2760 97 2792 103
rect 2808 97 3144 103
rect 3160 97 3224 103
rect 3240 97 3560 103
rect 4040 97 4072 103
rect 4408 97 4472 103
rect 4488 97 4520 103
rect 4536 97 4728 103
rect 4744 97 4792 103
rect 5416 97 5464 103
rect 5832 97 5992 103
rect 6184 97 6408 103
rect 6664 97 6824 103
rect 5080 57 5096 63
rect 5128 57 5176 63
rect 5128 37 5160 43
rect 5208 37 5272 43
rect 5336 37 5400 43
rect 5752 37 6568 43
rect 4952 17 4968 23
rect 5080 17 5112 23
rect 5144 17 5192 23
rect 5336 17 5352 23
rect 6280 17 6904 23
<< m4contact >>
rect 2158 5402 2186 5418
rect 4206 5402 4234 5418
rect 4504 5412 4520 5428
rect 4536 5412 4552 5428
rect 4728 5412 4744 5428
rect 4808 5412 4824 5428
rect 4936 5412 4952 5428
rect 5320 5412 5336 5428
rect 5368 5412 5384 5428
rect 4792 5392 4808 5408
rect 5352 5392 5368 5408
rect 6238 5402 6266 5418
rect 5064 5372 5080 5388
rect 6664 5372 6680 5388
rect 6200 5352 6216 5368
rect 7224 5352 7240 5368
rect 24 5332 40 5348
rect 5992 5332 6008 5348
rect 6152 5332 6168 5348
rect 6296 5332 6312 5348
rect 7064 5332 7080 5348
rect 7112 5332 7128 5348
rect 3096 5312 3112 5328
rect 5448 5312 5464 5328
rect 6840 5312 6856 5328
rect 7096 5312 7112 5328
rect 7288 5312 7304 5328
rect 760 5292 776 5308
rect 7144 5292 7160 5308
rect 4504 5272 4520 5288
rect 7304 5232 7320 5248
rect 1118 5202 1146 5218
rect 3166 5202 3194 5218
rect 5214 5202 5242 5218
rect 1240 5172 1256 5188
rect 3528 5172 3544 5188
rect 4568 5152 4584 5168
rect 6120 5152 6136 5168
rect 2536 5132 2552 5148
rect 7352 5132 7368 5148
rect 4824 5112 4840 5128
rect 6008 5112 6024 5128
rect 6504 5112 6520 5128
rect 7192 5112 7208 5128
rect 3688 5092 3704 5108
rect 3880 5092 3896 5108
rect 3976 5092 3992 5108
rect 4296 5092 4312 5108
rect 3112 5072 3128 5088
rect 4568 5072 4584 5088
rect 4792 5072 4808 5088
rect 6024 5072 6040 5088
rect 808 5052 824 5068
rect 1432 5052 1448 5068
rect 1880 5052 1896 5068
rect 3208 5052 3224 5068
rect 6792 5052 6808 5068
rect 4184 5032 4200 5048
rect 6968 5032 6984 5048
rect 2008 5012 2024 5028
rect 1960 4992 1976 5008
rect 2158 5002 2186 5018
rect 3832 4992 3848 5008
rect 4206 5002 4234 5018
rect 2792 4972 2808 4988
rect 6238 5002 6266 5018
rect 1880 4952 1896 4968
rect 504 4932 520 4948
rect 4088 4932 4104 4948
rect 4696 4932 4712 4948
rect 5448 4932 5464 4948
rect 6040 4932 6056 4948
rect 6216 4932 6232 4948
rect 808 4912 824 4928
rect 4472 4912 4488 4928
rect 5416 4912 5432 4928
rect 6264 4912 6280 4928
rect 6504 4912 6520 4928
rect 872 4892 888 4908
rect 1432 4892 1448 4908
rect 3128 4892 3144 4908
rect 3832 4892 3848 4908
rect 4808 4892 4840 4908
rect 5320 4892 5336 4908
rect 7032 4892 7048 4908
rect 4344 4872 4360 4888
rect 6648 4872 6664 4888
rect 3096 4852 3112 4868
rect 5496 4852 5512 4868
rect 6840 4852 6856 4868
rect 7000 4852 7016 4868
rect 3400 4832 3416 4848
rect 5080 4832 5096 4848
rect 1118 4802 1146 4818
rect 1240 4812 1256 4828
rect 2536 4812 2552 4828
rect 3166 4802 3194 4818
rect 4536 4792 4552 4808
rect 5214 4802 5242 4818
rect 5256 4812 5272 4828
rect 3848 4772 3864 4788
rect 6616 4772 6632 4788
rect 1288 4752 1304 4768
rect 2008 4752 2024 4768
rect 2536 4732 2552 4748
rect 3112 4732 3128 4748
rect 3256 4732 3272 4748
rect 3352 4732 3368 4748
rect 3640 4732 3656 4748
rect 4248 4732 4264 4748
rect 4296 4732 4312 4748
rect 4456 4732 4472 4748
rect 5400 4732 5416 4748
rect 5768 4732 5784 4748
rect 5864 4732 5880 4748
rect 1576 4712 1592 4728
rect 3096 4712 3112 4728
rect 3368 4712 3384 4728
rect 3592 4712 3608 4728
rect 3704 4712 3720 4728
rect 4200 4712 4216 4728
rect 4424 4712 4440 4728
rect 6792 4712 6808 4728
rect 1336 4692 1368 4708
rect 1384 4692 1400 4708
rect 3336 4692 3352 4708
rect 3720 4692 3736 4708
rect 4248 4692 4264 4708
rect 4520 4692 4536 4708
rect 5480 4692 5496 4708
rect 7000 4692 7016 4708
rect 1016 4672 1032 4688
rect 2552 4672 2584 4688
rect 3576 4672 3592 4688
rect 3624 4672 3640 4688
rect 6712 4672 6728 4688
rect 888 4652 904 4668
rect 1208 4652 1224 4668
rect 1304 4652 1320 4668
rect 1464 4652 1480 4668
rect 1976 4652 1992 4668
rect 2584 4652 2600 4668
rect 3240 4652 3256 4668
rect 3688 4652 3704 4668
rect 7032 4652 7048 4668
rect 3096 4632 3112 4648
rect 4408 4632 4424 4648
rect 4456 4632 4472 4648
rect 5976 4632 5992 4648
rect 1384 4612 1400 4628
rect 8 4592 24 4608
rect 1016 4592 1032 4608
rect 1368 4592 1384 4608
rect 2158 4602 2186 4618
rect 4206 4602 4234 4618
rect 5384 4612 5400 4628
rect 4408 4592 4424 4608
rect 6238 4602 6266 4618
rect 6280 4592 6296 4608
rect 2056 4572 2072 4588
rect 2088 4572 2104 4588
rect 5464 4572 5480 4588
rect 5608 4572 5640 4588
rect 6408 4572 6424 4588
rect 7176 4572 7192 4588
rect 5256 4552 5272 4568
rect 6616 4552 6632 4568
rect 1976 4532 1992 4548
rect 2168 4532 2184 4548
rect 4792 4532 4808 4548
rect 6056 4532 6072 4548
rect 6200 4532 6216 4548
rect 6664 4532 6680 4548
rect 7128 4532 7144 4548
rect 600 4512 616 4528
rect 888 4512 904 4528
rect 1320 4512 1352 4528
rect 1704 4512 1720 4528
rect 4120 4512 4136 4528
rect 4376 4512 4392 4528
rect 4776 4512 4792 4528
rect 5864 4512 5880 4528
rect 6200 4512 6216 4528
rect 6616 4512 6632 4528
rect 6840 4512 6856 4528
rect 7224 4512 7240 4528
rect 1464 4492 1480 4508
rect 1480 4492 1496 4508
rect 1592 4492 1608 4508
rect 1816 4492 1832 4508
rect 2200 4492 2216 4508
rect 2376 4492 2392 4508
rect 3688 4492 3704 4508
rect 4008 4492 4024 4508
rect 4936 4492 4952 4508
rect 6520 4492 6536 4508
rect 6664 4492 6680 4508
rect 6712 4492 6728 4508
rect 7272 4492 7288 4508
rect 7432 4492 7448 4508
rect 3880 4472 3896 4488
rect 5752 4472 5768 4488
rect 6136 4472 6152 4488
rect 7160 4472 7176 4488
rect 3448 4452 3464 4468
rect 6760 4452 6776 4468
rect 2072 4432 2088 4448
rect 3896 4432 3912 4448
rect 4824 4432 4840 4448
rect 7208 4432 7224 4448
rect 1118 4402 1146 4418
rect 1256 4412 1272 4428
rect 1544 4412 1560 4428
rect 1352 4392 1368 4408
rect 2328 4392 2344 4408
rect 3166 4402 3194 4418
rect 1288 4372 1304 4388
rect 2248 4372 2264 4388
rect 3656 4392 3672 4408
rect 5214 4402 5242 4418
rect 6344 4412 6360 4428
rect 5512 4392 5528 4408
rect 4312 4372 4328 4388
rect 5784 4372 5800 4388
rect 1864 4352 1880 4368
rect 6008 4352 6024 4368
rect 7000 4392 7016 4408
rect 1816 4332 1832 4348
rect 4584 4332 4600 4348
rect 5032 4332 5048 4348
rect 5496 4332 5512 4348
rect 6136 4332 6152 4348
rect 6360 4332 6376 4348
rect 6648 4332 6664 4348
rect 6920 4332 6936 4348
rect 7176 4332 7192 4348
rect 7320 4332 7336 4348
rect 1080 4312 1096 4328
rect 1464 4312 1480 4328
rect 1560 4312 1576 4328
rect 1576 4312 1592 4328
rect 2072 4312 2088 4328
rect 3592 4312 3608 4328
rect 4040 4312 4056 4328
rect 4088 4312 4104 4328
rect 4984 4312 5000 4328
rect 6040 4312 6056 4328
rect 760 4292 776 4308
rect 1000 4292 1016 4308
rect 1160 4292 1192 4308
rect 1960 4292 1976 4308
rect 2344 4292 2360 4308
rect 3512 4292 3528 4308
rect 3848 4292 3864 4308
rect 4120 4292 4136 4308
rect 5432 4292 5448 4308
rect 5512 4292 5528 4308
rect 5784 4292 5800 4308
rect 6200 4292 6216 4308
rect 7080 4292 7096 4308
rect 8 4272 24 4288
rect 904 4272 920 4288
rect 1016 4272 1032 4288
rect 2360 4272 2376 4288
rect 3608 4272 3624 4288
rect 4424 4272 4440 4288
rect 4888 4272 4904 4288
rect 5320 4272 5336 4288
rect 5928 4272 5944 4288
rect 6040 4272 6056 4288
rect 6424 4272 6440 4288
rect 1352 4252 1368 4268
rect 1736 4252 1752 4268
rect 5000 4252 5016 4268
rect 6200 4252 6216 4268
rect 7032 4252 7048 4268
rect 1720 4232 1736 4248
rect 4008 4232 4024 4248
rect 4808 4232 4824 4248
rect 1864 4212 1880 4228
rect 872 4192 888 4208
rect 1256 4192 1272 4208
rect 1720 4192 1752 4208
rect 2158 4202 2186 4218
rect 3400 4212 3416 4228
rect 3608 4192 3624 4208
rect 4104 4192 4120 4208
rect 4206 4202 4234 4218
rect 4264 4212 4280 4228
rect 5080 4212 5096 4228
rect 6238 4202 6266 4218
rect 6408 4192 6424 4208
rect 888 4172 904 4188
rect 6088 4172 6104 4188
rect 1000 4152 1016 4168
rect 3688 4152 3704 4168
rect 4472 4152 4488 4168
rect 6264 4152 6280 4168
rect 6968 4152 6984 4168
rect 1192 4132 1208 4148
rect 2360 4132 2376 4148
rect 2568 4132 2584 4148
rect 3048 4132 3064 4148
rect 5400 4132 5416 4148
rect 5512 4132 5528 4148
rect 6056 4132 6072 4148
rect 6280 4132 6296 4148
rect 6584 4132 6600 4148
rect 6984 4132 7000 4148
rect 744 4112 760 4128
rect 1128 4112 1144 4128
rect 1816 4112 1832 4128
rect 2472 4112 2488 4128
rect 2632 4112 2648 4128
rect 2904 4112 2920 4128
rect 2936 4112 2952 4128
rect 3128 4112 3144 4128
rect 3832 4112 3848 4128
rect 5496 4112 5512 4128
rect 6184 4112 6200 4128
rect 7080 4112 7096 4128
rect 392 4092 408 4108
rect 920 4092 936 4108
rect 4408 4092 4424 4108
rect 4696 4092 4712 4108
rect 4840 4092 4856 4108
rect 5176 4092 5192 4108
rect 5912 4092 5928 4108
rect 6584 4092 6600 4108
rect 4888 4072 4904 4088
rect 5432 4072 5448 4088
rect 6760 4072 6776 4088
rect 24 4052 40 4068
rect 2792 4052 2808 4068
rect 3336 4052 3352 4068
rect 3624 4052 3640 4068
rect 4104 4052 4120 4068
rect 5608 4052 5624 4068
rect 5784 4052 5800 4068
rect 7368 4052 7384 4068
rect 600 4032 616 4048
rect 3736 4032 3752 4048
rect 4456 4032 4472 4048
rect 6632 4032 6648 4048
rect 1000 4012 1016 4028
rect 1118 4002 1146 4018
rect 2360 4012 2376 4028
rect 3166 4002 3194 4018
rect 4456 3992 4472 4008
rect 5214 4002 5242 4018
rect 6216 4012 6232 4028
rect 6360 4012 6376 4028
rect 6600 4012 6616 4028
rect 6952 4012 6968 4028
rect 4408 3972 4424 3988
rect 4520 3972 4536 3988
rect 4536 3972 4552 3988
rect 4840 3972 4856 3988
rect 6168 3972 6184 3988
rect 6600 3972 6616 3988
rect 2632 3952 2648 3968
rect 2968 3952 2984 3968
rect 1064 3912 1080 3928
rect 2744 3932 2760 3948
rect 3960 3932 3976 3948
rect 4520 3932 4536 3948
rect 5064 3932 5080 3948
rect 6856 3932 6872 3948
rect 6920 3932 6936 3948
rect 1960 3912 1976 3928
rect 2344 3912 2360 3928
rect 2376 3912 2392 3928
rect 2504 3912 2520 3928
rect 4504 3912 4520 3928
rect 4600 3912 4616 3928
rect 424 3892 440 3908
rect 920 3892 936 3908
rect 4312 3892 4328 3908
rect 4840 3892 4856 3908
rect 4856 3892 4872 3908
rect 4872 3892 4888 3908
rect 5400 3892 5416 3908
rect 5512 3892 5528 3908
rect 7080 3892 7096 3908
rect 504 3872 520 3888
rect 904 3872 920 3888
rect 1160 3872 1176 3888
rect 392 3852 408 3868
rect 1368 3852 1384 3868
rect 2440 3872 2456 3888
rect 2584 3872 2600 3888
rect 3096 3872 3112 3888
rect 3832 3872 3848 3888
rect 4248 3872 4264 3888
rect 4728 3872 4744 3888
rect 2184 3852 2200 3868
rect 6136 3852 6152 3868
rect 4888 3832 4904 3848
rect 5816 3832 5832 3848
rect 7416 3832 7432 3848
rect 1256 3792 1272 3808
rect 2088 3792 2104 3808
rect 2158 3802 2186 3818
rect 3688 3812 3704 3828
rect 3720 3792 3736 3808
rect 4206 3802 4234 3818
rect 4536 3812 4552 3828
rect 4568 3792 4584 3808
rect 4888 3792 4904 3808
rect 6238 3802 6266 3818
rect 6856 3812 6872 3828
rect 6632 3792 6648 3808
rect 1960 3772 1976 3788
rect 2888 3772 2904 3788
rect 4792 3772 4808 3788
rect 1704 3752 1720 3768
rect 2776 3752 2792 3768
rect 3944 3752 3960 3768
rect 4808 3752 4824 3768
rect 5480 3752 5496 3768
rect 6120 3752 6136 3768
rect 7400 3752 7416 3768
rect 1160 3732 1176 3748
rect 2584 3732 2600 3748
rect 2792 3732 2808 3748
rect 4696 3732 4712 3748
rect 5608 3732 5624 3748
rect 5640 3732 5656 3748
rect 1432 3712 1448 3728
rect 1496 3712 1512 3728
rect 2776 3712 2792 3728
rect 3448 3712 3464 3728
rect 376 3692 392 3708
rect 1016 3692 1032 3708
rect 1608 3692 1624 3708
rect 2440 3692 2456 3708
rect 4312 3712 4328 3728
rect 4584 3712 4600 3728
rect 5896 3712 5912 3728
rect 6696 3712 6712 3728
rect 7368 3692 7384 3708
rect 1736 3672 1752 3688
rect 4968 3672 4984 3688
rect 3704 3652 3720 3668
rect 1544 3632 1560 3648
rect 4408 3632 4424 3648
rect 1118 3602 1146 3618
rect 3128 3612 3144 3628
rect 3144 3592 3160 3608
rect 3166 3602 3194 3618
rect 4344 3612 4360 3628
rect 4680 3592 4696 3608
rect 4824 3592 4840 3608
rect 5214 3602 5242 3618
rect 5368 3612 5384 3628
rect 6760 3612 6776 3628
rect 7384 3612 7400 3628
rect 6168 3592 6184 3608
rect 3800 3572 3816 3588
rect 4360 3572 4376 3588
rect 5496 3572 5512 3588
rect 776 3552 792 3568
rect 1000 3552 1016 3568
rect 4296 3552 4312 3568
rect 5816 3552 5832 3568
rect 1432 3532 1448 3548
rect 2328 3532 2344 3548
rect 3384 3532 3400 3548
rect 824 3512 840 3528
rect 1464 3512 1480 3528
rect 1544 3512 1560 3528
rect 4728 3532 4744 3548
rect 5784 3532 5800 3548
rect 6552 3532 6568 3548
rect 3512 3512 3528 3528
rect 4024 3512 4040 3528
rect 4296 3512 4312 3528
rect 4616 3512 4632 3528
rect 4664 3512 4680 3528
rect 5592 3512 5608 3528
rect 5768 3512 5784 3528
rect 6552 3512 6568 3528
rect 6952 3512 6968 3528
rect 2968 3492 2984 3508
rect 3464 3492 3480 3508
rect 4520 3492 4536 3508
rect 4728 3492 4744 3508
rect 5032 3492 5048 3508
rect 5512 3492 5528 3508
rect 6152 3492 6168 3508
rect 6856 3492 6872 3508
rect 248 3472 264 3488
rect 2440 3472 2456 3488
rect 2936 3472 2952 3488
rect 3368 3472 3384 3488
rect 3912 3472 3928 3488
rect 3608 3452 3624 3468
rect 3768 3452 3784 3468
rect 4072 3452 4088 3468
rect 4808 3472 4824 3488
rect 5176 3472 5192 3488
rect 6424 3472 6440 3488
rect 1752 3432 1768 3448
rect 4280 3432 4296 3448
rect 5352 3452 5368 3468
rect 5480 3452 5496 3468
rect 6360 3452 6376 3468
rect 6920 3452 6936 3468
rect 6984 3452 7000 3468
rect 2158 3402 2186 3418
rect 3256 3392 3272 3408
rect 3944 3392 3960 3408
rect 4206 3402 4234 3418
rect 5944 3412 5960 3428
rect 6238 3402 6266 3418
rect 6408 3392 6424 3408
rect 6712 3392 6728 3408
rect 7048 3392 7064 3408
rect 1224 3372 1240 3388
rect 3336 3372 3352 3388
rect 5864 3372 5880 3388
rect 6248 3372 6264 3388
rect 4232 3352 4264 3368
rect 4520 3352 4536 3368
rect 5080 3352 5096 3368
rect 5400 3352 5416 3368
rect 5896 3352 5912 3368
rect 1288 3332 1304 3348
rect 3384 3332 3400 3348
rect 3496 3332 3512 3348
rect 3704 3332 3720 3348
rect 3720 3332 3736 3348
rect 3912 3332 3928 3348
rect 4648 3332 4664 3348
rect 4696 3332 4712 3348
rect 4904 3332 4920 3348
rect 5864 3332 5880 3348
rect 2248 3312 2264 3328
rect 2360 3312 2376 3328
rect 3368 3312 3384 3328
rect 4712 3312 4728 3328
rect 5432 3312 5448 3328
rect 5832 3312 5848 3328
rect 6344 3312 6360 3328
rect 7080 3312 7096 3328
rect 2968 3292 2984 3308
rect 3720 3292 3736 3308
rect 3736 3292 3752 3308
rect 3912 3292 3928 3308
rect 4728 3292 4760 3308
rect 6200 3292 6216 3308
rect 7432 3292 7448 3308
rect 2088 3272 2104 3288
rect 376 3232 392 3248
rect 3416 3272 3432 3288
rect 4872 3272 4888 3288
rect 3976 3252 3992 3268
rect 5832 3252 5848 3268
rect 6744 3252 6760 3268
rect 1080 3212 1096 3228
rect 1118 3202 1146 3218
rect 5240 3232 5256 3248
rect 5912 3232 5928 3248
rect 6568 3232 6584 3248
rect 3166 3202 3194 3218
rect 5192 3212 5208 3228
rect 4184 3192 4200 3208
rect 4552 3192 4568 3208
rect 4808 3192 4824 3208
rect 5214 3202 5242 3218
rect 7016 3212 7032 3228
rect 5432 3192 5448 3208
rect 6200 3192 6216 3208
rect 2360 3172 2376 3188
rect 5128 3172 5144 3188
rect 5192 3172 5208 3188
rect 4184 3132 4200 3148
rect 5848 3132 5864 3148
rect 2888 3112 2904 3128
rect 3768 3112 3784 3128
rect 4072 3112 4088 3128
rect 6712 3112 6728 3128
rect 6760 3112 6776 3128
rect 7048 3112 7064 3128
rect 24 3092 40 3108
rect 2616 3092 2632 3108
rect 2888 3092 2904 3108
rect 3352 3092 3368 3108
rect 248 3072 264 3088
rect 2392 3072 2408 3088
rect 2792 3072 2824 3088
rect 4136 3072 4152 3088
rect 4664 3092 4680 3108
rect 4792 3092 4808 3108
rect 5464 3092 5480 3108
rect 5256 3072 5272 3088
rect 200 3052 216 3068
rect 5000 3052 5016 3068
rect 7336 3052 7352 3068
rect 3512 3032 3528 3048
rect 5848 3032 5864 3048
rect 6552 3032 6568 3048
rect 296 2992 312 3008
rect 1352 2992 1368 3008
rect 2158 3002 2186 3018
rect 2440 3012 2456 3028
rect 3656 2992 3672 3008
rect 4206 3002 4234 3018
rect 5944 2992 5960 3008
rect 6238 3002 6266 3018
rect 376 2972 392 2988
rect 1752 2972 1768 2988
rect 4744 2972 4760 2988
rect 5256 2972 5272 2988
rect 6632 2972 6648 2988
rect 3688 2952 3704 2968
rect 3864 2952 3880 2968
rect 6184 2952 6200 2968
rect 6648 2952 6664 2968
rect 1352 2932 1368 2948
rect 4456 2932 4472 2948
rect 4792 2932 4808 2948
rect 5112 2932 5128 2948
rect 5640 2932 5656 2948
rect 2840 2912 2856 2928
rect 4184 2912 4200 2928
rect 4920 2912 4936 2928
rect 5896 2912 5912 2928
rect 5944 2912 5960 2928
rect 6520 2912 6536 2928
rect 6584 2912 6600 2928
rect 6744 2912 6760 2928
rect 4120 2892 4136 2908
rect 7336 2892 7352 2908
rect 744 2872 760 2888
rect 3704 2872 3720 2888
rect 5400 2872 5416 2888
rect 7256 2872 7272 2888
rect 824 2852 840 2868
rect 3336 2852 3352 2868
rect 5688 2852 5704 2868
rect 3208 2832 3224 2848
rect 4664 2832 4680 2848
rect 5784 2832 5800 2848
rect 1118 2802 1146 2818
rect 3166 2802 3194 2818
rect 4776 2792 4792 2808
rect 5214 2802 5242 2818
rect 5752 2792 5768 2808
rect 6984 2792 7000 2808
rect 616 2772 632 2788
rect 776 2772 792 2788
rect 1176 2772 1192 2788
rect 1480 2772 1496 2788
rect 2040 2772 2056 2788
rect 2824 2772 2840 2788
rect 5160 2772 5176 2788
rect 6008 2772 6024 2788
rect 6200 2772 6216 2788
rect 7352 2772 7368 2788
rect 2040 2752 2056 2768
rect 7080 2752 7096 2768
rect 2104 2732 2120 2748
rect 4360 2732 4376 2748
rect 6680 2732 6696 2748
rect 200 2712 216 2728
rect 872 2712 888 2728
rect 1720 2712 1736 2728
rect 1752 2712 1768 2728
rect 1880 2712 1896 2728
rect 2104 2712 2120 2728
rect 2376 2712 2392 2728
rect 1096 2692 1112 2708
rect 2776 2692 2792 2708
rect 4328 2692 4344 2708
rect 4584 2692 4600 2708
rect 4904 2712 4920 2728
rect 5672 2712 5688 2728
rect 6248 2712 6264 2728
rect 6488 2712 6504 2728
rect 7176 2712 7192 2728
rect 4808 2692 4824 2708
rect 5848 2692 5864 2708
rect 5864 2692 5880 2708
rect 6520 2692 6536 2708
rect 7016 2692 7032 2708
rect 7288 2692 7304 2708
rect 7432 2692 7448 2708
rect 296 2672 312 2688
rect 1240 2672 1256 2688
rect 1736 2672 1752 2688
rect 1992 2672 2008 2688
rect 4440 2672 4456 2688
rect 4696 2672 4712 2688
rect 4728 2672 4744 2688
rect 5512 2672 5528 2688
rect 5608 2672 5624 2688
rect 5912 2672 5928 2688
rect 8 2652 24 2668
rect 4312 2652 4328 2668
rect 4744 2652 4760 2668
rect 5224 2652 5240 2668
rect 392 2632 408 2648
rect 4728 2632 4744 2648
rect 5784 2632 5800 2648
rect 6312 2632 6328 2648
rect 6792 2632 6808 2648
rect 7432 2632 7448 2648
rect 2158 2602 2186 2618
rect 3064 2612 3080 2628
rect 2264 2592 2280 2608
rect 4206 2602 4234 2618
rect 5576 2612 5592 2628
rect 5384 2592 5416 2608
rect 6238 2602 6266 2618
rect 8 2572 24 2588
rect 3464 2572 3480 2588
rect 8 2552 24 2568
rect 408 2532 424 2548
rect 456 2552 472 2568
rect 3656 2552 3672 2568
rect 4424 2552 4440 2568
rect 5256 2552 5272 2568
rect 6120 2572 6136 2588
rect 6504 2572 6520 2588
rect 1640 2532 1656 2548
rect 3416 2532 3432 2548
rect 4712 2532 4728 2548
rect 5480 2532 5496 2548
rect 376 2512 392 2528
rect 648 2512 664 2528
rect 2904 2512 2920 2528
rect 3432 2512 3448 2528
rect 3592 2512 3608 2528
rect 4248 2512 4264 2528
rect 4424 2512 4440 2528
rect 4456 2512 4472 2528
rect 4776 2512 4792 2528
rect 5464 2512 5480 2528
rect 6552 2532 6568 2548
rect 6888 2532 6904 2548
rect 7048 2532 7064 2548
rect 6632 2512 6648 2528
rect 6712 2512 6728 2528
rect 7048 2512 7064 2528
rect 7144 2512 7160 2528
rect 1160 2492 1176 2508
rect 1784 2492 1800 2508
rect 4664 2492 4680 2508
rect 5576 2492 5592 2508
rect 6952 2492 6968 2508
rect 7432 2492 7448 2508
rect 4648 2472 4664 2488
rect 7080 2472 7096 2488
rect 7224 2472 7240 2488
rect 4504 2452 4520 2468
rect 6744 2452 6760 2468
rect 1432 2432 1448 2448
rect 4840 2432 4856 2448
rect 6520 2432 6536 2448
rect 328 2392 344 2408
rect 1118 2402 1146 2418
rect 1768 2412 1784 2428
rect 3166 2402 3194 2418
rect 5214 2402 5242 2418
rect 7080 2412 7096 2428
rect 7384 2392 7400 2408
rect 5896 2372 5912 2388
rect 7144 2352 7160 2368
rect 5528 2332 5544 2348
rect 5608 2332 5624 2348
rect 7032 2332 7048 2348
rect 1016 2312 1032 2328
rect 1064 2312 1080 2328
rect 1640 2312 1656 2328
rect 3992 2312 4008 2328
rect 6488 2312 6504 2328
rect 6696 2312 6712 2328
rect 7208 2312 7224 2328
rect 4616 2292 4632 2308
rect 4648 2292 4664 2308
rect 4968 2292 4984 2308
rect 5336 2292 5352 2308
rect 5640 2292 5656 2308
rect 6024 2292 6040 2308
rect 6120 2292 6136 2308
rect 6952 2292 6968 2308
rect 7048 2292 7064 2308
rect 7352 2292 7368 2308
rect 1208 2272 1224 2288
rect 1224 2272 1240 2288
rect 3464 2272 3480 2288
rect 4680 2272 4696 2288
rect 4872 2272 4888 2288
rect 5960 2272 5976 2288
rect 7096 2272 7112 2288
rect 1576 2252 1592 2268
rect 6808 2252 6824 2268
rect 1720 2232 1736 2248
rect 4552 2232 4568 2248
rect 1832 2192 1848 2208
rect 2158 2202 2186 2218
rect 4206 2202 4234 2218
rect 4808 2212 4824 2228
rect 5544 2192 5560 2208
rect 6238 2202 6266 2218
rect 6504 2172 6520 2188
rect 408 2152 424 2168
rect 744 2152 760 2168
rect 1704 2152 1720 2168
rect 7032 2152 7048 2168
rect 328 2112 344 2128
rect 1176 2112 1192 2128
rect 1288 2112 1320 2128
rect 1512 2112 1528 2128
rect 1608 2112 1624 2128
rect 1848 2112 1864 2128
rect 2072 2112 2088 2128
rect 5576 2132 5592 2148
rect 6792 2132 6808 2148
rect 7208 2132 7224 2148
rect 7288 2132 7304 2148
rect 2840 2112 2872 2128
rect 4984 2112 5000 2128
rect 5160 2112 5192 2128
rect 5624 2112 5640 2128
rect 6344 2112 6360 2128
rect 6888 2112 6904 2128
rect 7336 2112 7352 2128
rect 616 2092 632 2108
rect 1496 2092 1512 2108
rect 5416 2092 5432 2108
rect 2088 2072 2104 2088
rect 3416 2072 3432 2088
rect 4504 2072 4520 2088
rect 4712 2072 4728 2088
rect 1064 2032 1080 2048
rect 1544 2032 1560 2048
rect 5960 2032 5976 2048
rect 1080 1992 1096 2008
rect 1118 2002 1146 2018
rect 3166 2002 3194 2018
rect 5176 1992 5192 2008
rect 5214 2002 5242 2018
rect 5640 2012 5656 2028
rect 4104 1972 4120 1988
rect 4504 1972 4520 1988
rect 5480 1972 5496 1988
rect 1080 1952 1096 1968
rect 5864 1952 5880 1968
rect 7048 1952 7064 1968
rect 7432 1952 7448 1968
rect 808 1932 824 1948
rect 1704 1932 1720 1948
rect 4248 1932 4264 1948
rect 4536 1932 4552 1948
rect 7032 1932 7048 1948
rect 7176 1932 7192 1948
rect 1016 1912 1032 1928
rect 1464 1912 1480 1928
rect 4024 1912 4040 1928
rect 4280 1912 4296 1928
rect 6328 1912 6344 1928
rect 7272 1912 7288 1928
rect 7336 1912 7352 1928
rect 1656 1892 1672 1908
rect 3992 1892 4008 1908
rect 4248 1892 4264 1908
rect 4456 1892 4472 1908
rect 4648 1892 4664 1908
rect 4904 1892 4920 1908
rect 5320 1892 5336 1908
rect 5544 1892 5560 1908
rect 5576 1892 5592 1908
rect 5944 1892 5960 1908
rect 6344 1892 6360 1908
rect 6568 1892 6584 1908
rect 6648 1892 6664 1908
rect 6808 1892 6824 1908
rect 6888 1892 6904 1908
rect 888 1872 904 1888
rect 1848 1872 1864 1888
rect 2456 1872 2472 1888
rect 4152 1872 4168 1888
rect 4696 1872 4712 1888
rect 1320 1852 1336 1868
rect 1688 1852 1704 1868
rect 1912 1852 1928 1868
rect 4520 1852 4536 1868
rect 4568 1852 4584 1868
rect 6584 1872 6600 1888
rect 6792 1872 6808 1888
rect 6952 1852 6968 1868
rect 1224 1832 1240 1848
rect 1800 1832 1816 1848
rect 3784 1832 3800 1848
rect 5512 1832 5528 1848
rect 296 1812 312 1828
rect 2136 1812 2152 1828
rect 1768 1792 1784 1808
rect 2120 1792 2136 1808
rect 2158 1802 2186 1818
rect 2392 1812 2408 1828
rect 2872 1792 2888 1808
rect 3432 1792 3448 1808
rect 4206 1802 4234 1818
rect 4568 1812 4584 1828
rect 4824 1792 4840 1808
rect 5288 1792 5304 1808
rect 5640 1792 5656 1808
rect 6200 1792 6216 1808
rect 6238 1802 6266 1818
rect 2360 1752 2376 1768
rect 4504 1772 4520 1788
rect 4744 1772 4760 1788
rect 5352 1772 5368 1788
rect 5400 1772 5416 1788
rect 5608 1772 5624 1788
rect 5624 1772 5640 1788
rect 6056 1772 6072 1788
rect 6280 1772 6296 1788
rect 7240 1772 7256 1788
rect 4792 1752 4808 1768
rect 5384 1752 5400 1768
rect 5736 1752 5752 1768
rect 6296 1752 6312 1768
rect 7304 1752 7320 1768
rect 616 1732 632 1748
rect 744 1732 760 1748
rect 2360 1732 2376 1748
rect 2520 1732 2536 1748
rect 2888 1732 2904 1748
rect 4584 1732 4600 1748
rect 4984 1732 5000 1748
rect 5320 1732 5336 1748
rect 5368 1732 5384 1748
rect 6440 1732 6456 1748
rect 6456 1732 6472 1748
rect 6760 1732 6776 1748
rect 7416 1732 7432 1748
rect 616 1712 632 1728
rect 1592 1712 1608 1728
rect 1784 1712 1800 1728
rect 280 1692 296 1708
rect 3464 1692 3480 1708
rect 3928 1712 3944 1728
rect 4904 1712 4920 1728
rect 5112 1712 5128 1728
rect 5416 1712 5432 1728
rect 5448 1712 5464 1728
rect 5816 1712 5832 1728
rect 6376 1712 6392 1728
rect 6392 1712 6408 1728
rect 7368 1712 7384 1728
rect 3928 1692 3944 1708
rect 4664 1692 4680 1708
rect 4712 1692 4728 1708
rect 5192 1692 5208 1708
rect 5304 1692 5320 1708
rect 7000 1692 7016 1708
rect 808 1672 824 1688
rect 4648 1672 4664 1688
rect 4824 1672 4840 1688
rect 5000 1672 5016 1688
rect 5064 1672 5080 1688
rect 6376 1672 6392 1688
rect 4696 1652 4712 1668
rect 2744 1632 2760 1648
rect 5656 1632 5672 1648
rect 7064 1632 7080 1648
rect 1118 1602 1146 1618
rect 3166 1602 3194 1618
rect 4728 1612 4744 1628
rect 5214 1602 5242 1618
rect 6408 1592 6424 1608
rect 2248 1572 2264 1588
rect 4136 1572 4152 1588
rect 4616 1572 4632 1588
rect 5864 1572 5880 1588
rect 4536 1552 4552 1568
rect 5896 1552 5912 1568
rect 7096 1552 7112 1568
rect 4248 1532 4264 1548
rect 4280 1532 4296 1548
rect 5016 1532 5032 1548
rect 5528 1532 5544 1548
rect 1176 1512 1192 1528
rect 1544 1512 1560 1528
rect 1992 1512 2024 1528
rect 4120 1512 4136 1528
rect 4616 1512 4632 1528
rect 5080 1512 5096 1528
rect 6200 1512 6216 1528
rect 7336 1512 7352 1528
rect 2136 1492 2152 1508
rect 3256 1492 3272 1508
rect 4072 1492 4088 1508
rect 4104 1492 4120 1508
rect 4872 1492 4888 1508
rect 5816 1492 5832 1508
rect 6056 1492 6072 1508
rect 6808 1492 6824 1508
rect 6904 1492 6920 1508
rect 7256 1492 7272 1508
rect 616 1472 632 1488
rect 648 1472 664 1488
rect 3960 1472 3976 1488
rect 4456 1472 4472 1488
rect 4728 1472 4744 1488
rect 4792 1472 4808 1488
rect 5928 1472 5944 1488
rect 4296 1452 4312 1468
rect 5176 1452 5192 1468
rect 7288 1452 7304 1468
rect 7368 1452 7384 1468
rect 2056 1432 2072 1448
rect 3896 1432 3912 1448
rect 4360 1432 4376 1448
rect 6712 1432 6728 1448
rect 824 1412 840 1428
rect 1976 1412 1992 1428
rect 1848 1392 1864 1408
rect 2158 1402 2186 1418
rect 3896 1412 3912 1428
rect 4206 1402 4234 1418
rect 4920 1412 4936 1428
rect 4792 1392 4808 1408
rect 4856 1392 4872 1408
rect 5736 1392 5752 1408
rect 6238 1402 6266 1418
rect 4024 1372 4040 1388
rect 5832 1372 5848 1388
rect 7224 1372 7240 1388
rect 1032 1352 1048 1368
rect 2840 1352 2856 1368
rect 2888 1352 2904 1368
rect 3576 1352 3592 1368
rect 4728 1352 4744 1368
rect 6456 1352 6472 1368
rect 952 1332 968 1348
rect 2808 1332 2824 1348
rect 2824 1332 2840 1348
rect 328 1312 344 1328
rect 648 1312 664 1328
rect 1704 1312 1720 1328
rect 3912 1332 3928 1348
rect 4136 1332 4152 1348
rect 4504 1332 4520 1348
rect 4600 1332 4616 1348
rect 6968 1332 6984 1348
rect 3048 1312 3080 1328
rect 3496 1312 3512 1328
rect 3928 1312 3944 1328
rect 3992 1312 4008 1328
rect 5352 1312 5368 1328
rect 6984 1312 7000 1328
rect 1224 1292 1240 1308
rect 2840 1292 2856 1308
rect 2920 1272 2936 1288
rect 2952 1272 2968 1288
rect 4120 1292 4136 1308
rect 4296 1292 4312 1308
rect 4472 1292 4488 1308
rect 3960 1272 3976 1288
rect 4344 1272 4360 1288
rect 7048 1272 7064 1288
rect 7400 1272 7416 1288
rect 4536 1252 4552 1268
rect 4616 1252 4632 1268
rect 4248 1232 4264 1248
rect 5736 1232 5752 1248
rect 6888 1232 6904 1248
rect 1118 1202 1146 1218
rect 1720 1212 1736 1228
rect 3166 1202 3194 1218
rect 4440 1212 4456 1228
rect 4888 1192 4904 1208
rect 5214 1202 5242 1218
rect 6168 1212 6184 1228
rect 6968 1212 6984 1228
rect 5656 1192 5672 1208
rect 6232 1192 6248 1208
rect 2024 1172 2040 1188
rect 3752 1172 3768 1188
rect 1608 1152 1624 1168
rect 1160 1132 1176 1148
rect 1288 1132 1304 1148
rect 2872 1152 2888 1168
rect 4360 1152 4376 1168
rect 4536 1152 4552 1168
rect 5416 1152 5432 1168
rect 6408 1152 6424 1168
rect 4296 1132 4312 1148
rect 6936 1132 6952 1148
rect 6984 1132 7000 1148
rect 1064 1112 1080 1128
rect 2248 1112 2264 1128
rect 4056 1112 4072 1128
rect 4504 1112 4520 1128
rect 4936 1112 4952 1128
rect 5288 1112 5304 1128
rect 5736 1112 5752 1128
rect 6296 1112 6312 1128
rect 6872 1112 6888 1128
rect 7080 1112 7096 1128
rect 7336 1112 7352 1128
rect 1320 1092 1336 1108
rect 2456 1092 2472 1108
rect 4184 1092 4200 1108
rect 4552 1092 4568 1108
rect 5816 1092 5832 1108
rect 5944 1092 5960 1108
rect 6440 1092 6456 1108
rect 7320 1092 7336 1108
rect 7352 1092 7368 1108
rect 616 1072 632 1088
rect 1064 1072 1080 1088
rect 1560 1072 1576 1088
rect 1976 1072 1992 1088
rect 2920 1072 2952 1088
rect 3624 1072 3640 1088
rect 4040 1072 4056 1088
rect 584 1052 600 1068
rect 648 1052 664 1068
rect 920 1052 936 1068
rect 1048 1052 1064 1068
rect 1960 1052 1976 1068
rect 2232 1052 2248 1068
rect 2392 1052 2408 1068
rect 3768 1052 3784 1068
rect 5336 1072 5352 1088
rect 4120 1052 4136 1068
rect 4904 1052 4920 1068
rect 6392 1052 6408 1068
rect 1432 1032 1448 1048
rect 4680 1032 4696 1048
rect 7000 1032 7016 1048
rect 392 992 408 1008
rect 840 992 856 1008
rect 2158 1002 2186 1018
rect 824 972 840 988
rect 1384 972 1400 988
rect 2344 992 2360 1008
rect 2952 992 2968 1008
rect 3592 992 3608 1008
rect 4024 992 4040 1008
rect 4206 1002 4234 1018
rect 6184 1012 6200 1028
rect 2312 972 2328 988
rect 4536 992 4552 1008
rect 6200 992 6216 1008
rect 6238 1002 6266 1018
rect 6280 992 6296 1008
rect 5336 972 5352 988
rect 5368 972 5384 988
rect 6744 972 6760 988
rect 1848 952 1864 968
rect 1288 932 1304 948
rect 1560 932 1576 948
rect 2120 932 2136 948
rect 1032 912 1048 928
rect 1096 912 1112 928
rect 1704 912 1720 928
rect 2856 912 2872 928
rect 4232 952 4248 968
rect 4584 952 4600 968
rect 5192 932 5208 948
rect 6920 972 6936 988
rect 7112 972 7128 988
rect 7224 972 7240 988
rect 6888 932 6904 948
rect 3736 912 3752 928
rect 4760 912 4776 928
rect 4936 912 4952 928
rect 6088 912 6104 928
rect 6200 912 6216 928
rect 6520 912 6536 928
rect 6984 912 7000 928
rect 7096 912 7112 928
rect 7208 912 7224 928
rect 280 892 296 908
rect 600 892 616 908
rect 1288 892 1304 908
rect 1560 892 1576 908
rect 2392 892 2408 908
rect 2744 892 2760 908
rect 3480 892 3496 908
rect 3592 892 3608 908
rect 3976 892 3992 908
rect 4424 892 4440 908
rect 4552 892 4568 908
rect 4712 892 4728 908
rect 4824 892 4840 908
rect 4872 892 4888 908
rect 5576 892 5592 908
rect 2328 872 2344 888
rect 3528 872 3544 888
rect 3624 872 3640 888
rect 4248 872 4264 888
rect 4456 872 4472 888
rect 4568 872 4584 888
rect 4728 872 4744 888
rect 6744 872 6760 888
rect 1640 852 1656 868
rect 2216 852 2232 868
rect 3720 852 3736 868
rect 3736 852 3752 868
rect 3976 852 3992 868
rect 4248 852 4264 868
rect 4440 852 4456 868
rect 5032 852 5048 868
rect 5464 852 5480 868
rect 5976 852 5992 868
rect 920 832 936 848
rect 1118 802 1146 818
rect 3144 812 3160 828
rect 3166 802 3194 818
rect 3752 792 3768 808
rect 5214 802 5242 818
rect 5256 792 5272 808
rect 3896 772 3912 788
rect 5160 772 5176 788
rect 440 752 456 768
rect 3912 752 3928 768
rect 3992 752 4008 768
rect 5112 752 5128 768
rect 2008 732 2024 748
rect 4328 732 4344 748
rect 5032 732 5048 748
rect 6968 732 6984 748
rect 1592 712 1608 728
rect 4232 712 4248 728
rect 2024 692 2040 708
rect 3464 692 3480 708
rect 3736 692 3752 708
rect 3992 692 4008 708
rect 5592 692 5608 708
rect 7112 692 7128 708
rect 616 672 632 688
rect 6904 652 6920 668
rect 7208 652 7224 668
rect 3720 632 3736 648
rect 600 612 616 628
rect 1976 612 1992 628
rect 2158 602 2186 618
rect 4206 602 4234 618
rect 4680 592 4696 608
rect 5448 592 5464 608
rect 6238 602 6266 618
rect 6808 612 6824 628
rect 6920 612 6936 628
rect 584 572 600 588
rect 3864 572 3880 588
rect 744 552 760 568
rect 952 552 968 568
rect 616 532 632 548
rect 2056 532 2072 548
rect 3416 552 3432 568
rect 3464 552 3480 568
rect 4312 572 4328 588
rect 5336 572 5352 588
rect 6376 552 6392 568
rect 6184 532 6200 548
rect 744 512 760 528
rect 1304 512 1320 528
rect 2328 512 2344 528
rect 4520 512 4536 528
rect 6088 512 6104 528
rect 6744 512 6760 528
rect 648 492 664 508
rect 2136 492 2152 508
rect 3864 492 3880 508
rect 1432 472 1448 488
rect 5768 472 5784 488
rect 6872 452 6888 468
rect 4248 432 4264 448
rect 1118 402 1146 418
rect 3166 402 3194 418
rect 4600 412 4616 428
rect 5214 402 5242 418
rect 5768 412 5784 428
rect 440 372 456 388
rect 1400 372 1416 388
rect 824 352 840 368
rect 3672 352 3688 368
rect 1096 332 1112 348
rect 5176 332 5192 348
rect 6440 332 6456 348
rect 3416 312 3432 328
rect 5016 312 5032 328
rect 5176 312 5192 328
rect 4168 292 4184 308
rect 4888 292 4904 308
rect 5128 292 5144 308
rect 6440 292 6456 308
rect 296 272 312 288
rect 5816 272 5832 288
rect 6312 272 6328 288
rect 7320 272 7336 288
rect 2936 232 2952 248
rect 6920 232 6936 248
rect 2158 202 2186 218
rect 3592 212 3608 228
rect 4206 202 4234 218
rect 4248 192 4264 208
rect 6238 202 6266 218
rect 7128 172 7144 188
rect 7144 172 7160 188
rect 7272 172 7288 188
rect 4248 152 4264 168
rect 1400 132 1416 148
rect 4616 132 4632 148
rect 7160 132 7176 148
rect 7224 132 7240 148
rect 4328 112 4344 128
rect 5032 112 5048 128
rect 5080 112 5096 128
rect 5112 112 5128 128
rect 7192 112 7208 128
rect 7240 112 7256 128
rect 1544 92 1560 108
rect 3592 92 3608 108
rect 4520 92 4536 108
rect 5112 52 5128 68
rect 1118 2 1146 18
rect 3166 2 3194 18
rect 4024 12 4040 28
rect 4856 12 4872 28
rect 4920 12 4936 28
rect 5112 12 5144 28
rect 5214 2 5242 18
rect 5304 12 5320 28
rect 5320 12 5336 28
<< metal4 >>
rect 2186 5406 2192 5414
rect 4234 5406 4240 5414
rect 13 4288 19 4592
rect 29 4068 35 5332
rect 29 3108 35 4052
rect 397 3868 403 4092
rect 509 3888 515 4932
rect 605 4048 611 4512
rect 765 4308 771 5292
rect 1146 5206 1152 5214
rect 813 4928 819 5052
rect 877 4208 883 4892
rect 1245 4828 1251 5172
rect 1437 4908 1443 5052
rect 1885 4968 1891 5052
rect 1146 4806 1152 4814
rect 893 4528 899 4652
rect 1021 4608 1027 4672
rect 893 4188 899 4512
rect 253 3088 259 3472
rect 381 3248 387 3692
rect 205 2728 211 3052
rect 301 2688 307 2992
rect 13 2588 19 2652
rect 381 2528 387 2972
rect 749 2888 755 4112
rect 909 3888 915 4272
rect 1005 4168 1011 4292
rect 1021 4288 1027 4592
rect 1146 4406 1152 4414
rect 1005 4144 1011 4152
rect 1004 4136 1012 4144
rect 1148 4123 1156 4124
rect 1144 4117 1156 4123
rect 1148 4116 1156 4117
rect 925 3908 931 4092
rect 1005 3568 1011 4012
rect 1146 4006 1152 4014
rect 781 2788 787 3552
rect 829 2868 835 3512
rect 604 2783 612 2784
rect 604 2777 616 2783
rect 604 2776 612 2777
rect 333 2128 339 2392
rect 285 908 291 1692
rect 301 288 307 1812
rect 333 1328 339 2112
rect 397 1008 403 2632
rect 413 2168 419 2532
rect 621 1748 627 2092
rect 621 1488 627 1712
rect 653 1488 659 2512
rect 749 1748 755 2152
rect 877 2104 883 2712
rect 1021 2328 1027 3692
rect 1069 2328 1075 3912
rect 1165 3748 1171 3872
rect 1146 3606 1152 3614
rect 876 2096 884 2104
rect 813 1688 819 1932
rect 1021 1928 1027 2312
rect 1069 2048 1075 2312
rect 621 1088 627 1472
rect 653 1328 659 1472
rect 445 388 451 752
rect 589 588 595 1052
rect 605 628 611 892
rect 621 688 627 1072
rect 621 548 627 672
rect 653 508 659 1052
rect 829 988 835 1412
rect 844 1036 852 1044
rect 845 1008 851 1036
rect 749 528 755 552
rect 829 368 835 972
rect 925 848 931 1052
rect 957 568 963 1332
rect 1037 928 1043 1352
rect 1069 1128 1075 2032
rect 1085 2008 1091 3212
rect 1146 3206 1152 3214
rect 1146 2806 1152 2814
rect 1165 2508 1171 3732
rect 1181 2788 1187 4292
rect 1261 4208 1267 4412
rect 1293 4388 1299 4752
rect 1308 4696 1316 4704
rect 1309 4668 1315 4696
rect 1341 4528 1347 4692
rect 1325 4504 1331 4512
rect 1324 4496 1332 4504
rect 1357 4408 1363 4692
rect 1372 4636 1380 4644
rect 1373 4608 1379 4636
rect 1389 4628 1395 4692
rect 1261 3808 1267 4192
rect 1146 2406 1152 2414
rect 1181 2128 1187 2772
rect 1229 2288 1235 3372
rect 1245 2664 1251 2672
rect 1244 2656 1252 2664
rect 1213 2264 1219 2272
rect 1212 2256 1220 2264
rect 1293 2128 1299 3332
rect 1357 3008 1363 4252
rect 1437 3728 1443 4892
rect 1484 4663 1492 4664
rect 1480 4657 1492 4663
rect 1484 4656 1492 4657
rect 1468 4516 1476 4524
rect 1469 4508 1475 4516
rect 1357 2948 1363 2992
rect 1437 2448 1443 3532
rect 1146 2006 1152 2014
rect 1085 1904 1091 1952
rect 1084 1896 1092 1904
rect 1146 1606 1152 1614
rect 1181 1528 1187 2112
rect 1229 1308 1235 1832
rect 1146 1206 1152 1214
rect 1165 1084 1171 1132
rect 1293 1124 1299 1132
rect 1292 1116 1300 1124
rect 1164 1076 1172 1084
rect 1069 1044 1075 1072
rect 1068 1036 1076 1044
rect 1101 348 1107 912
rect 1293 908 1299 932
rect 1146 806 1152 814
rect 1309 528 1315 2112
rect 1469 1928 1475 3512
rect 1485 2788 1491 4492
rect 1501 2108 1507 3712
rect 1549 3648 1555 4412
rect 1581 4328 1587 4712
rect 1596 4516 1604 4524
rect 1597 4508 1603 4516
rect 1709 3768 1715 4512
rect 1821 4484 1827 4492
rect 1820 4476 1828 4484
rect 1725 4208 1731 4232
rect 1741 4208 1747 4252
rect 1821 4144 1827 4332
rect 1869 4228 1875 4352
rect 1965 4308 1971 4992
rect 2013 4768 2019 5012
rect 2186 5006 2192 5014
rect 2541 4828 2547 5132
rect 2556 4716 2564 4724
rect 2557 4688 2563 4716
rect 1981 4644 1987 4652
rect 1980 4636 1988 4644
rect 2444 4636 2452 4644
rect 2186 4606 2192 4614
rect 2076 4583 2084 4584
rect 2076 4577 2088 4583
rect 2076 4576 2084 4577
rect 2172 4576 2180 4584
rect 2061 4564 2067 4572
rect 2060 4556 2068 4564
rect 2173 4548 2179 4576
rect 2204 4536 2212 4544
rect 2205 4508 2211 4536
rect 2381 4484 2387 4492
rect 2380 4476 2388 4484
rect 2348 4436 2356 4444
rect 2077 4328 2083 4432
rect 2186 4206 2192 4214
rect 1820 4136 1828 4144
rect 1821 4128 1827 4136
rect 1965 3788 1971 3912
rect 2204 3863 2212 3864
rect 2200 3857 2212 3863
rect 2204 3856 2212 3857
rect 2186 3806 2192 3814
rect 1549 2048 1555 3512
rect 1596 2263 1604 2264
rect 1592 2257 1604 2263
rect 1596 2256 1604 2257
rect 1613 2128 1619 3692
rect 1645 2328 1651 2532
rect 1709 2168 1715 3752
rect 1741 2688 1747 3672
rect 1757 2988 1763 3432
rect 2093 3288 2099 3792
rect 2186 3406 2192 3414
rect 2253 3328 2259 4372
rect 2333 3548 2339 4392
rect 2349 4308 2355 4436
rect 2365 4148 2371 4272
rect 2349 3904 2355 3912
rect 2348 3896 2356 3904
rect 2365 3328 2371 4012
rect 2381 3928 2387 4476
rect 2365 3188 2371 3312
rect 2186 3006 2192 3014
rect 1757 2728 1763 2972
rect 2044 2836 2052 2844
rect 2045 2788 2051 2836
rect 2060 2763 2068 2764
rect 2056 2757 2068 2763
rect 2060 2756 2068 2757
rect 2092 2743 2100 2744
rect 2092 2737 2104 2743
rect 2092 2736 2100 2737
rect 1900 2723 1908 2724
rect 1896 2717 1908 2723
rect 1900 2716 1908 2717
rect 2109 2704 2115 2712
rect 2108 2696 2116 2704
rect 1836 2676 1844 2684
rect 1709 1948 1715 2152
rect 1676 1903 1684 1904
rect 1672 1897 1684 1903
rect 1676 1896 1684 1897
rect 1325 1108 1331 1852
rect 1437 488 1443 1032
rect 1146 406 1152 414
rect 1405 148 1411 372
rect 1549 108 1555 1512
rect 1580 1083 1588 1084
rect 1576 1077 1588 1083
rect 1580 1076 1588 1077
rect 1565 908 1571 932
rect 1597 728 1603 1712
rect 1709 1328 1715 1932
rect 1613 1104 1619 1152
rect 1612 1096 1620 1104
rect 1709 928 1715 1312
rect 1725 1228 1731 2232
rect 1773 1808 1779 2412
rect 1789 1728 1795 2492
rect 1837 2208 1843 2676
rect 1853 1888 1859 2112
rect 1916 1876 1924 1884
rect 1853 1408 1859 1872
rect 1917 1868 1923 1876
rect 1997 1528 2003 2672
rect 2268 2636 2276 2644
rect 2186 2606 2192 2614
rect 2269 2608 2275 2636
rect 2186 2206 2192 2214
rect 2092 2123 2100 2124
rect 2088 2117 2100 2123
rect 2092 2116 2100 2117
rect 2093 2088 2099 2116
rect 2125 1684 2131 1792
rect 2141 1784 2147 1812
rect 2186 1806 2192 1814
rect 2140 1776 2148 1784
rect 2365 1768 2371 3172
rect 2381 2728 2387 3912
rect 2445 3888 2451 4636
rect 2573 4148 2579 4672
rect 2589 4644 2595 4652
rect 2588 4636 2596 4644
rect 2492 4123 2500 4124
rect 2488 4117 2500 4123
rect 2492 4116 2500 4117
rect 2637 3968 2643 4112
rect 2797 4068 2803 4972
rect 3101 4868 3107 5312
rect 4509 5288 4515 5412
rect 3194 5206 3200 5214
rect 3117 4748 3123 5072
rect 3101 4704 3107 4712
rect 3100 4696 3108 4704
rect 3036 4143 3044 4144
rect 3036 4137 3048 4143
rect 3036 4136 3044 4137
rect 2445 3488 2451 3692
rect 2445 3028 2451 3472
rect 2509 3464 2515 3912
rect 2749 3904 2755 3932
rect 2748 3896 2756 3904
rect 2589 3748 2595 3872
rect 2797 3748 2803 4052
rect 2508 3456 2516 3464
rect 2604 3103 2612 3104
rect 2604 3097 2616 3103
rect 2604 3096 2612 3097
rect 2781 2708 2787 3712
rect 2797 3088 2803 3732
rect 2893 3128 2899 3772
rect 2893 3108 2899 3112
rect 2812 3096 2820 3104
rect 2813 3088 2819 3096
rect 2461 1864 2467 1872
rect 2460 1856 2468 1864
rect 2396 1836 2404 1844
rect 2397 1828 2403 1836
rect 2348 1743 2356 1744
rect 2348 1737 2360 1743
rect 2348 1736 2356 1737
rect 2124 1676 2132 1684
rect 1853 968 1859 1392
rect 1981 1088 1987 1412
rect 1981 628 1987 1072
rect 2013 748 2019 1512
rect 2029 708 2035 1172
rect 2061 548 2067 1432
rect 2125 904 2131 932
rect 2124 896 2132 904
rect 2141 508 2147 1492
rect 2186 1406 2192 1414
rect 2253 1128 2259 1572
rect 2236 1116 2244 1124
rect 2237 1068 2243 1116
rect 2476 1103 2484 1104
rect 2472 1097 2484 1103
rect 2476 1096 2484 1097
rect 2186 1006 2192 1014
rect 2349 984 2355 992
rect 2348 976 2356 984
rect 2220 936 2228 944
rect 2221 868 2227 936
rect 2317 924 2323 972
rect 2316 916 2324 924
rect 2397 908 2403 1052
rect 2749 908 2755 1632
rect 2829 1348 2835 2772
rect 2845 2128 2851 2912
rect 2909 2528 2915 4112
rect 2941 3488 2947 4112
rect 2973 3508 2979 3952
rect 3101 3888 3107 4632
rect 3133 4128 3139 4892
rect 3194 4806 3200 4814
rect 3194 4406 3200 4414
rect 3194 4006 3200 4014
rect 3133 3564 3139 3612
rect 3194 3606 3200 3614
rect 3132 3556 3140 3564
rect 3149 3544 3155 3592
rect 3148 3536 3156 3544
rect 2973 3284 2979 3292
rect 2972 3276 2980 3284
rect 3194 3206 3200 3214
rect 3213 2848 3219 5052
rect 3244 4696 3252 4704
rect 3245 4668 3251 4696
rect 3261 4664 3267 4732
rect 3260 4656 3268 4664
rect 3341 4068 3347 4692
rect 3357 4684 3363 4732
rect 3388 4723 3396 4724
rect 3384 4717 3396 4723
rect 3388 4716 3396 4717
rect 3356 4676 3364 4684
rect 3405 4228 3411 4832
rect 3453 3728 3459 4452
rect 3341 2868 3347 3372
rect 3373 3328 3379 3472
rect 3389 3348 3395 3532
rect 3517 3528 3523 4292
rect 3468 3516 3476 3524
rect 3469 3508 3475 3516
rect 3484 3343 3492 3344
rect 3484 3337 3496 3343
rect 3484 3336 3492 3337
rect 3436 3283 3444 3284
rect 3432 3277 3444 3283
rect 3436 3276 3444 3277
rect 3517 3048 3523 3512
rect 3194 2806 3200 2814
rect 2861 928 2867 2112
rect 2877 1168 2883 1792
rect 2893 1724 2899 1732
rect 2892 1716 2900 1724
rect 2893 1344 2899 1352
rect 2892 1336 2900 1344
rect 3069 1328 3075 2612
rect 3421 2524 3427 2532
rect 3420 2516 3428 2524
rect 3194 2406 3200 2414
rect 3420 2116 3428 2124
rect 3421 2088 3427 2116
rect 3194 2006 3200 2014
rect 3437 1808 3443 2512
rect 3469 2288 3475 2572
rect 3194 1606 3200 1614
rect 2924 1116 2932 1124
rect 2925 1088 2931 1116
rect 2186 606 2192 614
rect 2333 564 2339 872
rect 2332 556 2340 564
rect 2333 528 2339 556
rect 2941 248 2947 1072
rect 2957 1008 2963 1272
rect 3194 1206 3200 1214
rect 3148 876 3156 884
rect 3149 828 3155 876
rect 3194 806 3200 814
rect 3469 708 3475 1692
rect 3484 916 3492 924
rect 3485 908 3491 916
rect 3533 888 3539 5172
rect 3596 4736 3604 4744
rect 3628 4743 3636 4744
rect 3628 4737 3640 4743
rect 3628 4736 3636 4737
rect 3597 4728 3603 4736
rect 3580 4716 3588 4724
rect 3581 4688 3587 4716
rect 3612 4323 3620 4324
rect 3608 4317 3620 4323
rect 3612 4316 3620 4317
rect 3612 4256 3620 4264
rect 3613 4208 3619 4256
rect 3629 4068 3635 4672
rect 3693 4668 3699 5092
rect 3837 4908 3843 4992
rect 3709 4564 3715 4712
rect 3708 4556 3716 4564
rect 3708 4503 3716 4504
rect 3704 4497 3716 4503
rect 3708 4496 3716 4497
rect 3612 3476 3620 3484
rect 3613 3468 3619 3476
rect 3661 3008 3667 4392
rect 3693 3828 3699 4152
rect 3725 3808 3731 4692
rect 3853 4308 3859 4772
rect 3885 4488 3891 5092
rect 3741 3924 3747 4032
rect 3740 3916 3748 3924
rect 3837 3888 3843 4112
rect 3709 3348 3715 3652
rect 3709 3304 3715 3332
rect 3725 3308 3731 3332
rect 3708 3296 3716 3304
rect 3661 2568 3667 2992
rect 3693 2924 3699 2952
rect 3692 2916 3700 2924
rect 3709 2888 3715 3296
rect 3756 3303 3764 3304
rect 3752 3297 3764 3303
rect 3756 3296 3764 3297
rect 3773 3128 3779 3452
rect 3964 3403 3972 3404
rect 3960 3397 3972 3403
rect 3964 3396 3972 3397
rect 3917 3308 3923 3332
rect 3981 3268 3987 5092
rect 4092 5076 4100 5084
rect 4093 4948 4099 5076
rect 4108 4523 4116 4524
rect 4108 4517 4120 4523
rect 4108 4516 4116 4517
rect 4013 4248 4019 4492
rect 4076 4323 4084 4324
rect 4076 4317 4088 4323
rect 4076 4316 4084 4317
rect 4045 4304 4051 4312
rect 4044 4296 4052 4304
rect 4109 4068 4115 4192
rect 4044 3523 4052 3524
rect 4040 3517 4052 3523
rect 4044 3516 4052 3517
rect 4077 3128 4083 3452
rect 3869 2944 3875 2952
rect 3868 2936 3876 2944
rect 4125 2908 4131 4292
rect 4189 3208 4195 5032
rect 4234 5006 4240 5014
rect 4301 4748 4307 5092
rect 4253 4724 4259 4732
rect 4220 4723 4228 4724
rect 4216 4717 4228 4723
rect 4220 4716 4228 4717
rect 4252 4716 4260 4724
rect 4234 4606 4240 4614
rect 4234 4206 4240 4214
rect 4253 3888 4259 4692
rect 4269 4144 4275 4212
rect 4268 4136 4276 4144
rect 4317 3908 4323 4372
rect 4234 3806 4240 3814
rect 4317 3728 4323 3892
rect 4349 3628 4355 4872
rect 4429 4704 4435 4712
rect 4428 4696 4436 4704
rect 4461 4648 4467 4732
rect 4413 4608 4419 4632
rect 4444 4283 4452 4284
rect 4440 4277 4452 4283
rect 4444 4276 4452 4277
rect 4477 4168 4483 4912
rect 4541 4808 4547 5412
rect 4573 5088 4579 5152
rect 4413 3988 4419 4092
rect 4461 4008 4467 4032
rect 4525 3988 4531 4692
rect 4413 3648 4419 3972
rect 4509 3904 4515 3912
rect 4508 3896 4516 3904
rect 4301 3528 4307 3552
rect 4525 3508 4531 3932
rect 4541 3828 4547 3972
rect 4573 3808 4579 5072
rect 4701 4924 4707 4932
rect 4700 4916 4708 4924
rect 4589 3728 4595 4332
rect 4620 3923 4628 3924
rect 4616 3917 4628 3923
rect 4620 3916 4628 3917
rect 4701 3748 4707 4092
rect 4733 3888 4739 5412
rect 4797 5088 4803 5392
rect 4797 4548 4803 5072
rect 4813 4908 4819 5412
rect 4829 4908 4835 5112
rect 4764 4523 4772 4524
rect 4764 4517 4776 4523
rect 4764 4516 4772 4517
rect 4941 4508 4947 5412
rect 4812 4316 4820 4324
rect 4813 4248 4819 4316
rect 4668 3556 4676 3564
rect 4620 3536 4628 3544
rect 4621 3528 4627 3536
rect 4669 3528 4675 3556
rect 4284 3456 4292 3464
rect 4285 3448 4291 3456
rect 4234 3406 4240 3414
rect 4252 3376 4260 3384
rect 4253 3368 4259 3376
rect 4189 2928 4195 3132
rect 4234 3006 4240 3014
rect 4365 2724 4371 2732
rect 4364 2716 4372 2724
rect 4444 2696 4452 2704
rect 4333 2684 4339 2692
rect 4445 2688 4451 2696
rect 4332 2676 4340 2684
rect 4234 2606 4240 2614
rect 3596 2536 3604 2544
rect 3597 2528 3603 2536
rect 3997 1908 4003 2312
rect 4234 2206 4240 2214
rect 3789 1704 3795 1832
rect 3788 1696 3796 1704
rect 3901 1428 3907 1432
rect 3597 908 3603 992
rect 3629 888 3635 1072
rect 3741 868 3747 912
rect 3725 648 3731 852
rect 3757 808 3763 1172
rect 3901 788 3907 1412
rect 3917 768 3923 1332
rect 3933 1328 3939 1692
rect 3965 1288 3971 1472
rect 4029 1388 4035 1912
rect 4109 1508 4115 1972
rect 4253 1908 4259 1932
rect 4156 1896 4164 1904
rect 4157 1888 4163 1896
rect 4234 1806 4240 1814
rect 4092 1503 4100 1504
rect 4088 1497 4100 1503
rect 4092 1496 4100 1497
rect 3981 868 3987 892
rect 3997 768 4003 1312
rect 4125 1308 4131 1512
rect 4141 1348 4147 1572
rect 4285 1548 4291 1912
rect 4234 1406 4240 1414
rect 4253 1248 4259 1532
rect 4300 1476 4308 1484
rect 4301 1468 4307 1476
rect 4301 1284 4307 1292
rect 4300 1276 4308 1284
rect 4301 1124 4307 1132
rect 4076 1123 4084 1124
rect 4072 1117 4084 1123
rect 4076 1116 4084 1117
rect 4300 1116 4308 1124
rect 4172 1103 4180 1104
rect 4172 1097 4184 1103
rect 4172 1096 4180 1097
rect 4140 1063 4148 1064
rect 4136 1057 4148 1063
rect 4140 1056 4148 1057
rect 4234 1006 4240 1014
rect 3740 716 3748 724
rect 3741 708 3747 716
rect 3997 708 4003 752
rect 3452 563 3460 564
rect 3452 557 3464 563
rect 3452 556 3460 557
rect 3194 406 3200 414
rect 3421 328 3427 552
rect 3869 508 3875 572
rect 3677 304 3683 352
rect 3676 296 3684 304
rect 2186 206 2192 214
rect 3597 108 3603 212
rect 4029 28 4035 992
rect 4253 868 4259 872
rect 4234 606 4240 614
rect 4253 448 4259 852
rect 4317 588 4323 2652
rect 4429 2528 4435 2552
rect 4460 2536 4468 2544
rect 4461 2528 4467 2536
rect 4509 2088 4515 2452
rect 4557 2248 4563 3192
rect 4604 2703 4612 2704
rect 4600 2697 4612 2703
rect 4604 2696 4612 2697
rect 4653 2488 4659 3332
rect 4669 2508 4675 2832
rect 4685 2744 4691 3592
rect 4701 3348 4707 3732
rect 4716 3543 4724 3544
rect 4716 3537 4728 3543
rect 4716 3536 4724 3537
rect 4684 2736 4692 2744
rect 4653 2308 4659 2472
rect 4509 1904 4515 1972
rect 4476 1903 4484 1904
rect 4472 1897 4484 1903
rect 4476 1896 4484 1897
rect 4508 1896 4516 1904
rect 4476 1483 4484 1484
rect 4472 1477 4484 1483
rect 4476 1476 4484 1477
rect 4332 1283 4340 1284
rect 4332 1277 4344 1283
rect 4332 1276 4340 1277
rect 4365 1168 4371 1432
rect 4509 1348 4515 1772
rect 4492 1303 4500 1304
rect 4488 1297 4500 1303
rect 4492 1296 4500 1297
rect 4445 924 4451 1212
rect 4509 1128 4515 1332
rect 4460 976 4468 984
rect 4444 916 4452 924
rect 4429 864 4435 892
rect 4461 888 4467 976
rect 4428 856 4436 864
rect 4188 303 4196 304
rect 4184 297 4196 303
rect 4188 296 4196 297
rect 4234 206 4240 214
rect 4253 168 4259 192
rect 4333 128 4339 732
rect 4525 528 4531 1852
rect 4541 1568 4547 1932
rect 4573 1828 4579 1852
rect 4604 1743 4612 1744
rect 4600 1737 4612 1743
rect 4604 1736 4612 1737
rect 4621 1588 4627 2292
rect 4685 2288 4691 2736
rect 4701 2688 4707 3332
rect 4636 1903 4644 1904
rect 4636 1897 4648 1903
rect 4636 1896 4644 1897
rect 4701 1888 4707 2672
rect 4717 2548 4723 3312
rect 4733 3308 4739 3492
rect 4749 2988 4755 3292
rect 4797 3108 4803 3772
rect 4813 3488 4819 3752
rect 4829 3608 4835 4432
rect 5020 4343 5028 4344
rect 5020 4337 5032 4343
rect 5020 4336 5028 4337
rect 4845 3988 4851 4092
rect 4893 4088 4899 4272
rect 4989 4264 4995 4312
rect 4988 4256 4996 4264
rect 4845 3908 4851 3972
rect 4860 3936 4868 3944
rect 4861 3908 4867 3936
rect 4733 2648 4739 2672
rect 4749 2668 4755 2972
rect 4797 2924 4803 2932
rect 4796 2916 4804 2924
rect 4717 2088 4723 2532
rect 4652 1716 4660 1724
rect 4653 1688 4659 1716
rect 4684 1703 4692 1704
rect 4680 1697 4692 1703
rect 4684 1696 4692 1697
rect 4701 1668 4707 1872
rect 4716 1776 4724 1784
rect 4717 1708 4723 1776
rect 4733 1628 4739 2632
rect 4749 1788 4755 2652
rect 4781 2528 4787 2792
rect 4813 2708 4819 3192
rect 4813 2228 4819 2692
rect 4845 2448 4851 3892
rect 4877 3288 4883 3892
rect 4893 3808 4899 3832
rect 4940 2923 4948 2924
rect 4936 2917 4948 2923
rect 4940 2916 4948 2917
rect 4973 2308 4979 3672
rect 5005 3068 5011 4252
rect 5069 3948 5075 5372
rect 5242 5206 5248 5214
rect 5325 4908 5331 5412
rect 5085 4228 5091 4832
rect 5242 4806 5248 4814
rect 5261 4568 5267 4812
rect 5242 4406 5248 4414
rect 5325 4288 5331 4892
rect 4621 1528 4627 1572
rect 4797 1488 4803 1752
rect 4829 1688 4835 1792
rect 4877 1508 4883 2272
rect 4909 1728 4915 1892
rect 4972 1743 4980 1744
rect 4972 1737 4984 1743
rect 4972 1736 4980 1737
rect 5020 1683 5028 1684
rect 5016 1677 5028 1683
rect 5020 1676 5028 1677
rect 4733 1368 4739 1472
rect 4797 1408 4803 1472
rect 4541 1008 4547 1152
rect 4540 903 4548 904
rect 4540 897 4552 903
rect 4540 896 4548 897
rect 4572 896 4580 904
rect 4573 888 4579 896
rect 4525 108 4531 512
rect 4605 428 4611 1332
rect 4621 148 4627 1252
rect 4685 608 4691 1032
rect 4716 916 4724 924
rect 4717 908 4723 916
rect 4733 888 4739 1352
rect 4748 923 4756 924
rect 4748 917 4760 923
rect 4748 916 4756 917
rect 4829 884 4835 892
rect 4828 876 4836 884
rect 4861 28 4867 1392
rect 4876 936 4884 944
rect 4877 908 4883 936
rect 4893 308 4899 1192
rect 4908 1076 4916 1084
rect 4909 1068 4915 1076
rect 4925 28 4931 1412
rect 4956 1123 4964 1124
rect 4952 1117 4964 1123
rect 4956 1116 4964 1117
rect 5021 328 5027 1532
rect 5037 868 5043 3492
rect 5181 3488 5187 4092
rect 5242 4006 5248 4014
rect 5242 3606 5248 3614
rect 5357 3468 5363 5392
rect 5373 3628 5379 5412
rect 6266 5406 6272 5414
rect 5453 4948 5459 5312
rect 5388 4736 5396 4744
rect 5389 4628 5395 4736
rect 5405 4148 5411 4732
rect 5068 3376 5076 3384
rect 5069 3364 5075 3376
rect 5405 3368 5411 3892
rect 5068 3363 5076 3364
rect 5068 3357 5080 3363
rect 5068 3356 5076 3357
rect 5228 3243 5236 3244
rect 5228 3237 5240 3243
rect 5228 3236 5236 3237
rect 5197 3188 5203 3212
rect 5242 3206 5248 3214
rect 5117 1728 5123 2932
rect 5052 1683 5060 1684
rect 5052 1677 5064 1683
rect 5052 1676 5060 1677
rect 5037 128 5043 732
rect 5085 128 5091 1512
rect 5117 128 5123 752
rect 5133 308 5139 3172
rect 5261 2988 5267 3072
rect 5242 2806 5248 2814
rect 5165 2644 5171 2772
rect 5228 2676 5236 2684
rect 5229 2668 5235 2676
rect 5164 2636 5172 2644
rect 5405 2608 5411 2872
rect 5242 2406 5248 2414
rect 5165 788 5171 2112
rect 5181 2008 5187 2112
rect 5242 2006 5248 2014
rect 5181 348 5187 1452
rect 5197 948 5203 1692
rect 5242 1606 5248 1614
rect 5242 1206 5248 1214
rect 5242 806 5248 814
rect 5261 808 5267 2552
rect 5308 2096 5316 2104
rect 5309 1904 5315 2096
rect 5308 1903 5316 1904
rect 5308 1897 5320 1903
rect 5308 1896 5316 1897
rect 5293 1128 5299 1792
rect 5242 406 5248 414
rect 5181 328 5187 332
rect 5117 28 5123 52
rect 5133 28 5139 292
rect 5309 28 5315 1692
rect 5325 28 5331 1732
rect 5341 1088 5347 2292
rect 5357 1328 5363 1772
rect 5389 1768 5395 2592
rect 5421 2108 5427 4912
rect 5437 3328 5443 4072
rect 5437 3208 5443 3312
rect 5453 2784 5459 4932
rect 5468 4703 5476 4704
rect 5468 4697 5480 4703
rect 5468 4696 5476 4697
rect 5468 4676 5476 4684
rect 5469 4588 5475 4676
rect 5501 4348 5507 4852
rect 5628 4656 5636 4664
rect 5629 4588 5635 4656
rect 5596 4583 5604 4584
rect 5596 4577 5608 4583
rect 5596 4576 5604 4577
rect 5869 4528 5875 4732
rect 5980 4716 5988 4724
rect 5981 4648 5987 4716
rect 5740 4483 5748 4484
rect 5740 4477 5752 4483
rect 5740 4476 5748 4477
rect 5517 4308 5523 4392
rect 5789 4308 5795 4372
rect 6013 4368 6019 5112
rect 6044 5083 6052 5084
rect 6040 5077 6052 5083
rect 6044 5076 6052 5077
rect 6045 4328 6051 4932
rect 5932 4296 5940 4304
rect 5517 4148 5523 4292
rect 5485 3744 5491 3752
rect 5484 3736 5492 3744
rect 5501 3588 5507 4112
rect 5789 4068 5795 4292
rect 5933 4288 5939 4296
rect 6045 4288 6051 4312
rect 5517 3508 5523 3892
rect 5613 3748 5619 4052
rect 5469 2924 5475 3092
rect 5468 2916 5476 2924
rect 5452 2776 5460 2784
rect 5405 1724 5411 1772
rect 5453 1728 5459 2776
rect 5485 2548 5491 3452
rect 5404 1716 5412 1724
rect 5421 1168 5427 1712
rect 5341 588 5347 972
rect 5469 868 5475 2512
rect 5485 1988 5491 2532
rect 5517 1848 5523 2672
rect 5581 2508 5587 2612
rect 5533 1548 5539 2332
rect 5549 1908 5555 2192
rect 5564 2143 5572 2144
rect 5564 2137 5576 2143
rect 5564 2136 5572 2137
rect 5581 908 5587 1892
rect 5597 708 5603 3512
rect 5613 2688 5619 3732
rect 5789 3548 5795 4052
rect 5821 3568 5827 3832
rect 5772 3536 5780 3544
rect 5773 3528 5779 3536
rect 5869 3348 5875 3372
rect 5901 3368 5907 3712
rect 5837 3268 5843 3312
rect 5852 3236 5860 3244
rect 5853 3148 5859 3236
rect 5613 1788 5619 2332
rect 5645 2308 5651 2932
rect 5693 2764 5699 2852
rect 5692 2756 5700 2764
rect 5660 2723 5668 2724
rect 5660 2717 5672 2723
rect 5660 2716 5668 2717
rect 5693 2704 5699 2756
rect 5757 2724 5763 2792
rect 5756 2716 5764 2724
rect 5692 2696 5700 2704
rect 5789 2648 5795 2832
rect 5853 2708 5859 3032
rect 5869 2708 5875 3332
rect 5901 2928 5907 3352
rect 5917 3248 5923 4092
rect 5933 2844 5939 4272
rect 6061 4148 6067 4532
rect 6092 4336 6100 4344
rect 6093 4188 6099 4336
rect 6125 3768 6131 5152
rect 6141 4348 6147 4472
rect 6141 3868 6147 4332
rect 6157 3508 6163 5332
rect 6205 4548 6211 5352
rect 6266 5006 6272 5014
rect 6205 4528 6211 4532
rect 6205 4268 6211 4292
rect 6173 3608 6179 3972
rect 5949 3008 5955 3412
rect 5949 2928 5955 2992
rect 5932 2836 5940 2844
rect 5629 1788 5635 2112
rect 5645 1808 5651 2012
rect 5869 1968 5875 2692
rect 5900 2683 5908 2684
rect 5900 2677 5912 2683
rect 5900 2676 5908 2677
rect 5661 1208 5667 1632
rect 5741 1408 5747 1752
rect 5821 1508 5827 1712
rect 5869 1588 5875 1952
rect 5901 1568 5907 2372
rect 5933 1488 5939 2836
rect 6013 2304 6019 2772
rect 6125 2308 6131 2572
rect 6012 2303 6020 2304
rect 6012 2297 6024 2303
rect 6012 2296 6020 2297
rect 5965 2048 5971 2272
rect 5741 1248 5747 1392
rect 5837 1284 5843 1372
rect 5836 1276 5844 1284
rect 5741 1128 5747 1232
rect 5949 1108 5955 1892
rect 6061 1508 6067 1772
rect 6173 1228 6179 3592
rect 6189 2968 6195 4112
rect 6221 4028 6227 4932
rect 6509 4928 6515 5112
rect 6266 4606 6272 4614
rect 6285 4584 6291 4592
rect 6284 4576 6292 4584
rect 6348 4476 6356 4484
rect 6349 4428 6355 4476
rect 6266 4206 6272 4214
rect 6280 4157 6291 4163
rect 6285 4148 6291 4157
rect 6365 4028 6371 4332
rect 6413 4208 6419 4572
rect 6621 4568 6627 4772
rect 6524 4516 6532 4524
rect 6525 4508 6531 4516
rect 6621 4504 6627 4512
rect 6620 4496 6628 4504
rect 6653 4348 6659 4872
rect 6669 4548 6675 5372
rect 7212 5363 7220 5364
rect 7212 5357 7224 5363
rect 7212 5356 7220 5357
rect 6797 4728 6803 5052
rect 6845 4868 6851 5312
rect 6716 4696 6724 4704
rect 6717 4688 6723 4696
rect 6669 4508 6675 4532
rect 6845 4528 6851 4852
rect 6732 4503 6740 4504
rect 6728 4497 6740 4503
rect 6732 4496 6740 4497
rect 6266 3806 6272 3814
rect 6365 3468 6371 4012
rect 6266 3406 6272 3414
rect 6413 3408 6419 4192
rect 6429 3488 6435 4272
rect 6589 4108 6595 4132
rect 6765 4088 6771 4452
rect 6605 3988 6611 4012
rect 6637 3808 6643 4032
rect 6925 3948 6931 4332
rect 6973 4168 6979 5032
rect 7005 4708 7011 4852
rect 7037 4668 7043 4892
rect 6861 3828 6867 3932
rect 6557 3528 6563 3532
rect 6253 3364 6259 3372
rect 6252 3356 6260 3364
rect 6332 3323 6340 3324
rect 6332 3317 6344 3323
rect 6332 3316 6340 3317
rect 6205 2788 6211 3192
rect 6557 3048 6563 3512
rect 6266 3006 6272 3014
rect 6205 1808 6211 2772
rect 6252 2736 6260 2744
rect 6253 2728 6259 2736
rect 6493 2664 6499 2712
rect 6540 2703 6548 2704
rect 6536 2697 6548 2703
rect 6540 2696 6548 2697
rect 6492 2656 6500 2664
rect 6266 2606 6272 2614
rect 6266 2206 6272 2214
rect 6266 1806 6272 1814
rect 6205 1528 6211 1792
rect 6285 1684 6291 1772
rect 6284 1676 6292 1684
rect 6266 1406 6272 1414
rect 6236 1256 6244 1264
rect 6237 1208 6243 1256
rect 6301 1128 6307 1752
rect 5453 564 5459 592
rect 5452 556 5460 564
rect 5773 428 5779 472
rect 5821 288 5827 1092
rect 6093 528 6099 912
rect 6189 548 6195 1012
rect 6266 1006 6272 1014
rect 6205 928 6211 992
rect 6285 904 6291 992
rect 6284 896 6292 904
rect 6266 606 6272 614
rect 6317 288 6323 2632
rect 6493 2328 6499 2656
rect 6509 2188 6515 2572
rect 6332 1956 6340 1964
rect 6333 1928 6339 1956
rect 6349 1908 6355 2112
rect 6381 1688 6387 1712
rect 6381 568 6387 1672
rect 6397 1068 6403 1712
rect 6413 1168 6419 1592
rect 6445 1108 6451 1732
rect 6461 1368 6467 1732
rect 6525 928 6531 2432
rect 6573 2144 6579 3232
rect 6572 2136 6580 2144
rect 6573 1908 6579 2136
rect 6589 1888 6595 2912
rect 6637 2528 6643 2972
rect 6653 1908 6659 2952
rect 6701 2328 6707 3712
rect 6717 3128 6723 3392
rect 6748 3316 6756 3324
rect 6749 3268 6755 3316
rect 6765 3128 6771 3612
rect 6861 3508 6867 3812
rect 6925 3468 6931 3932
rect 6957 3528 6963 4012
rect 6989 3468 6995 4132
rect 6717 1448 6723 2512
rect 6749 2468 6755 2912
rect 6765 1748 6771 3112
rect 6797 2148 6803 2632
rect 6797 1888 6803 2132
rect 6813 1908 6819 2252
rect 6893 2128 6899 2532
rect 6972 2503 6980 2504
rect 6968 2497 6980 2503
rect 6972 2496 6980 2497
rect 6972 2476 6980 2484
rect 6893 1908 6899 2112
rect 6813 1508 6819 1892
rect 6957 1868 6963 2292
rect 6940 1716 6948 1724
rect 6732 983 6740 984
rect 6732 977 6744 983
rect 6732 976 6740 977
rect 6749 528 6755 872
rect 6813 628 6819 1492
rect 6877 468 6883 1112
rect 6893 948 6899 1232
rect 6909 668 6915 1492
rect 6941 1148 6947 1716
rect 6973 1348 6979 2476
rect 6989 1328 6995 2792
rect 7005 1724 7011 4392
rect 7037 4268 7043 4652
rect 7021 2708 7027 3212
rect 7053 3128 7059 3392
rect 7037 2168 7043 2332
rect 7053 2308 7059 2512
rect 7037 1948 7043 2152
rect 7004 1716 7012 1724
rect 6940 983 6948 984
rect 6936 977 6948 983
rect 6940 976 6948 977
rect 6973 748 6979 1212
rect 6989 928 6995 1132
rect 7005 1048 7011 1692
rect 7053 1288 7059 1952
rect 7069 1648 7075 5332
rect 7085 4128 7091 4292
rect 7085 3908 7091 4112
rect 7085 3328 7091 3892
rect 7085 2488 7091 2752
rect 7085 1128 7091 2412
rect 7101 2288 7107 5312
rect 7117 2484 7123 5332
rect 7116 2476 7124 2484
rect 7101 928 7107 1552
rect 7117 708 7123 972
rect 6445 308 6451 332
rect 6925 248 6931 612
rect 6266 206 6272 214
rect 7133 188 7139 4532
rect 7149 2528 7155 5292
rect 7149 2304 7155 2352
rect 7148 2296 7156 2304
rect 7149 164 7155 172
rect 7148 156 7156 164
rect 7165 148 7171 4472
rect 7181 4364 7187 4572
rect 7180 4356 7188 4364
rect 7181 2744 7187 4332
rect 7180 2736 7188 2744
rect 7181 1948 7187 2712
rect 7197 128 7203 5112
rect 7213 2328 7219 4432
rect 7229 2488 7235 4512
rect 7244 2556 7252 2564
rect 7213 943 7219 2132
rect 7245 1803 7251 2556
rect 7229 1797 7251 1803
rect 7229 1388 7235 1797
rect 7228 996 7236 1004
rect 7229 988 7235 996
rect 7213 937 7235 943
rect 7213 668 7219 912
rect 7229 148 7235 937
rect 7245 128 7251 1772
rect 7261 1508 7267 2872
rect 7277 2564 7283 4492
rect 7293 3484 7299 5312
rect 7292 3476 7300 3484
rect 7276 2556 7284 2564
rect 7293 2148 7299 2692
rect 7292 2116 7300 2124
rect 7277 188 7283 1912
rect 7293 1468 7299 2116
rect 7309 1768 7315 5232
rect 7325 1108 7331 4332
rect 7341 2908 7347 3052
rect 7357 2804 7363 5132
rect 7373 3708 7379 4052
rect 7372 3476 7380 3484
rect 7356 2796 7364 2804
rect 7357 2308 7363 2772
rect 7341 1928 7347 2112
rect 7341 1128 7347 1512
rect 7357 1108 7363 2292
rect 7373 1728 7379 3476
rect 7389 2408 7395 3612
rect 7384 1457 7395 1463
rect 7405 1288 7411 3752
rect 7421 1748 7427 3832
rect 7437 2648 7443 2692
rect 7325 288 7331 1092
rect 1146 6 1152 14
rect 3194 6 3200 14
rect 5242 6 5248 14
use OAI21X1  OAI21X1_72
timestamp 1515870181
transform -1 0 72 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_80
timestamp 1515870181
transform -1 0 120 0 -1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_56
timestamp 1515870181
transform 1 0 120 0 -1 5410
box 0 0 192 200
use MUX2X1  MUX2X1_24
timestamp 1515870181
transform -1 0 408 0 -1 5410
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_199
timestamp 1515870181
transform 1 0 408 0 -1 5410
box 0 0 192 200
use BUFX4  BUFX4_77
timestamp 1515870181
transform -1 0 664 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_216
timestamp 1515870181
transform -1 0 856 0 -1 5410
box 0 0 192 200
use NAND2X1  NAND2X1_202
timestamp 1515870181
transform 1 0 856 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_216
timestamp 1515870181
transform -1 0 968 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_196
timestamp 1515870181
transform 1 0 968 0 -1 5410
box 0 0 192 200
use FILL  FILL_26_0_0
timestamp 1515870181
transform 1 0 1160 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_0_1
timestamp 1515870181
transform 1 0 1176 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_10
timestamp 1515870181
transform 1 0 1192 0 -1 5410
box 0 0 96 200
use NAND2X1  NAND2X1_181
timestamp 1515870181
transform 1 0 1288 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_196
timestamp 1515870181
transform -1 0 1400 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_58
timestamp 1515870181
transform 1 0 1400 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_52
timestamp 1515870181
transform -1 0 1512 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_68
timestamp 1515870181
transform -1 0 1704 0 -1 5410
box 0 0 192 200
use BUFX4  BUFX4_63
timestamp 1515870181
transform 1 0 1704 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_72
timestamp 1515870181
transform 1 0 1768 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_56
timestamp 1515870181
transform 1 0 1960 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_62
timestamp 1515870181
transform -1 0 2072 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_1_0
timestamp 1515870181
transform 1 0 2072 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_1_1
timestamp 1515870181
transform 1 0 2088 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_69
timestamp 1515870181
transform 1 0 2104 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_200
timestamp 1515870181
transform 1 0 2296 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_185
timestamp 1515870181
transform -1 0 2408 0 -1 5410
box 0 0 48 200
use MUX2X1  MUX2X1_22
timestamp 1515870181
transform -1 0 2504 0 -1 5410
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_200
timestamp 1515870181
transform -1 0 2696 0 -1 5410
box 0 0 192 200
use BUFX4  BUFX4_31
timestamp 1515870181
transform -1 0 2760 0 -1 5410
box 0 0 64 200
use BUFX4  BUFX4_125
timestamp 1515870181
transform -1 0 2824 0 -1 5410
box 0 0 64 200
use BUFX4  BUFX4_126
timestamp 1515870181
transform -1 0 2888 0 -1 5410
box 0 0 64 200
use BUFX2  BUFX2_21
timestamp 1515870181
transform -1 0 2936 0 -1 5410
box 0 0 48 200
use INVX8  INVX8_4
timestamp 1515870181
transform -1 0 3016 0 -1 5410
box 0 0 80 200
use BUFX2  BUFX2_20
timestamp 1515870181
transform 1 0 3016 0 -1 5410
box 0 0 48 200
use BUFX2  BUFX2_5
timestamp 1515870181
transform -1 0 3112 0 -1 5410
box 0 0 48 200
use BUFX2  BUFX2_4
timestamp 1515870181
transform -1 0 3160 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_2_0
timestamp 1515870181
transform -1 0 3176 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_2_1
timestamp 1515870181
transform -1 0 3192 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_100
timestamp 1515870181
transform -1 0 3384 0 -1 5410
box 0 0 192 200
use INVX1  INVX1_24
timestamp 1515870181
transform 1 0 3384 0 -1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_501
timestamp 1515870181
transform 1 0 3416 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_440
timestamp 1515870181
transform -1 0 3528 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_505
timestamp 1515870181
transform -1 0 3592 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_444
timestamp 1515870181
transform -1 0 3640 0 -1 5410
box 0 0 48 200
use INVX1  INVX1_44
timestamp 1515870181
transform -1 0 3672 0 -1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_104
timestamp 1515870181
transform -1 0 3864 0 -1 5410
box 0 0 192 200
use INVX8  INVX8_8
timestamp 1515870181
transform -1 0 3944 0 -1 5410
box 0 0 80 200
use BUFX4  BUFX4_74
timestamp 1515870181
transform -1 0 4008 0 -1 5410
box 0 0 64 200
use BUFX2  BUFX2_8
timestamp 1515870181
transform -1 0 4056 0 -1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_108
timestamp 1515870181
transform 1 0 4056 0 -1 5410
box 0 0 192 200
use FILL  FILL_26_3_0
timestamp 1515870181
transform 1 0 4248 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_3_1
timestamp 1515870181
transform 1 0 4264 0 -1 5410
box 0 0 16 200
use INVX1  INVX1_64
timestamp 1515870181
transform 1 0 4280 0 -1 5410
box 0 0 32 200
use BUFX2  BUFX2_24
timestamp 1515870181
transform 1 0 4312 0 -1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_266
timestamp 1515870181
transform -1 0 4552 0 -1 5410
box 0 0 192 200
use INVX2  INVX2_11
timestamp 1515870181
transform 1 0 4552 0 -1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_251
timestamp 1515870181
transform -1 0 4648 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_237
timestamp 1515870181
transform -1 0 4696 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_235
timestamp 1515870181
transform 1 0 4696 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_251
timestamp 1515870181
transform 1 0 4744 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_265
timestamp 1515870181
transform -1 0 4856 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_312
timestamp 1515870181
transform 1 0 4856 0 -1 5410
box 0 0 192 200
use INVX2  INVX2_25
timestamp 1515870181
transform 1 0 5048 0 -1 5410
box 0 0 32 200
use BUFX4  BUFX4_90
timestamp 1515870181
transform 1 0 5080 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_249
timestamp 1515870181
transform -1 0 5208 0 -1 5410
box 0 0 64 200
use FILL  FILL_26_4_0
timestamp 1515870181
transform 1 0 5208 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_4_1
timestamp 1515870181
transform 1 0 5224 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_264
timestamp 1515870181
transform 1 0 5240 0 -1 5410
box 0 0 192 200
use INVX2  INVX2_9
timestamp 1515870181
transform 1 0 5432 0 -1 5410
box 0 0 32 200
use BUFX4  BUFX4_29
timestamp 1515870181
transform 1 0 5464 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_231
timestamp 1515870181
transform 1 0 5528 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_247
timestamp 1515870181
transform 1 0 5576 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_261
timestamp 1515870181
transform -1 0 5688 0 -1 5410
box 0 0 64 200
use INVX2  INVX2_21
timestamp 1515870181
transform -1 0 5720 0 -1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_308
timestamp 1515870181
transform -1 0 5912 0 -1 5410
box 0 0 192 200
use NAND2X1  NAND2X1_255
timestamp 1515870181
transform 1 0 5912 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_269
timestamp 1515870181
transform -1 0 6024 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_248
timestamp 1515870181
transform 1 0 6024 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_262
timestamp 1515870181
transform -1 0 6136 0 -1 5410
box 0 0 64 200
use INVX2  INVX2_29
timestamp 1515870181
transform -1 0 6168 0 -1 5410
box 0 0 32 200
use FILL  FILL_26_5_0
timestamp 1515870181
transform -1 0 6184 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_5_1
timestamp 1515870181
transform -1 0 6200 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_316
timestamp 1515870181
transform -1 0 6392 0 -1 5410
box 0 0 192 200
use INVX2  INVX2_22
timestamp 1515870181
transform -1 0 6424 0 -1 5410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_309
timestamp 1515870181
transform -1 0 6616 0 -1 5410
box 0 0 192 200
use BUFX4  BUFX4_93
timestamp 1515870181
transform 1 0 6616 0 -1 5410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_335
timestamp 1515870181
transform -1 0 6872 0 -1 5410
box 0 0 192 200
use AOI21X1  AOI21X1_15
timestamp 1515870181
transform 1 0 6872 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_24
timestamp 1515870181
transform 1 0 6936 0 -1 5410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_286
timestamp 1515870181
transform 1 0 6984 0 -1 5410
box 0 0 192 200
use NOR3X1  NOR3X1_27
timestamp 1515870181
transform 1 0 7176 0 -1 5410
box 0 0 128 200
use NOR2X1  NOR2X1_57
timestamp 1515870181
transform -1 0 7352 0 -1 5410
box 0 0 48 200
use BUFX4  BUFX4_219
timestamp 1515870181
transform 1 0 7352 0 -1 5410
box 0 0 64 200
use FILL  FILL_27_1
timestamp 1515870181
transform -1 0 7432 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_212
timestamp 1515870181
transform -1 0 200 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_71
timestamp 1515870181
transform 1 0 200 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_55
timestamp 1515870181
transform 1 0 392 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_61
timestamp 1515870181
transform -1 0 504 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_199
timestamp 1515870181
transform 1 0 504 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_184
timestamp 1515870181
transform -1 0 616 0 1 5010
box 0 0 48 200
use MUX2X1  MUX2X1_19
timestamp 1515870181
transform 1 0 616 0 1 5010
box 0 0 96 200
use OAI21X1  OAI21X1_207
timestamp 1515870181
transform 1 0 712 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_192
timestamp 1515870181
transform -1 0 824 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_207
timestamp 1515870181
transform 1 0 824 0 1 5010
box 0 0 192 200
use BUFX4  BUFX4_96
timestamp 1515870181
transform -1 0 1080 0 1 5010
box 0 0 64 200
use FILL  FILL_25_0_0
timestamp 1515870181
transform 1 0 1080 0 1 5010
box 0 0 16 200
use FILL  FILL_25_0_1
timestamp 1515870181
transform 1 0 1096 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_180
timestamp 1515870181
transform 1 0 1112 0 1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_164
timestamp 1515870181
transform 1 0 1304 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_180
timestamp 1515870181
transform -1 0 1416 0 1 5010
box 0 0 64 200
use BUFX4  BUFX4_207
timestamp 1515870181
transform 1 0 1416 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_191
timestamp 1515870181
transform -1 0 1672 0 1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_175
timestamp 1515870181
transform 1 0 1672 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_191
timestamp 1515870181
transform -1 0 1784 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_181
timestamp 1515870181
transform 1 0 1784 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_165
timestamp 1515870181
transform -1 0 1896 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_181
timestamp 1515870181
transform 1 0 1896 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_37
timestamp 1515870181
transform 1 0 2088 0 1 5010
box 0 0 64 200
use FILL  FILL_25_1_0
timestamp 1515870181
transform 1 0 2152 0 1 5010
box 0 0 16 200
use FILL  FILL_25_1_1
timestamp 1515870181
transform 1 0 2168 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1515870181
transform 1 0 2184 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_53
timestamp 1515870181
transform 1 0 2376 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_184
timestamp 1515870181
transform 1 0 2440 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_168
timestamp 1515870181
transform -1 0 2552 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_182
timestamp 1515870181
transform 1 0 2552 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_197
timestamp 1515870181
transform -1 0 2664 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_184
timestamp 1515870181
transform 1 0 2664 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_40
timestamp 1515870181
transform 1 0 2856 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1515870181
transform 1 0 2920 0 1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_293
timestamp 1515870181
transform 1 0 3112 0 1 5010
box 0 0 48 200
use FILL  FILL_25_2_0
timestamp 1515870181
transform -1 0 3176 0 1 5010
box 0 0 16 200
use FILL  FILL_25_2_1
timestamp 1515870181
transform -1 0 3192 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_20
timestamp 1515870181
transform -1 0 3384 0 1 5010
box 0 0 192 200
use BUFX4  BUFX4_30
timestamp 1515870181
transform 1 0 3384 0 1 5010
box 0 0 64 200
use BUFX2  BUFX2_23
timestamp 1515870181
transform 1 0 3448 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_85
timestamp 1515870181
transform -1 0 3688 0 1 5010
box 0 0 192 200
use BUFX2  BUFX2_15
timestamp 1515870181
transform 1 0 3688 0 1 5010
box 0 0 48 200
use BUFX4  BUFX4_306
timestamp 1515870181
transform 1 0 3736 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_319
timestamp 1515870181
transform -1 0 3848 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_7
timestamp 1515870181
transform -1 0 3896 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_28
timestamp 1515870181
transform -1 0 3944 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_19
timestamp 1515870181
transform 1 0 3944 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_111
timestamp 1515870181
transform 1 0 3992 0 1 5010
box 0 0 192 200
use INVX1  INVX1_79
timestamp 1515870181
transform 1 0 4184 0 1 5010
box 0 0 32 200
use FILL  FILL_25_3_0
timestamp 1515870181
transform 1 0 4216 0 1 5010
box 0 0 16 200
use FILL  FILL_25_3_1
timestamp 1515870181
transform 1 0 4232 0 1 5010
box 0 0 16 200
use BUFX4  BUFX4_124
timestamp 1515870181
transform 1 0 4248 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_509
timestamp 1515870181
transform 1 0 4312 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_512
timestamp 1515870181
transform 1 0 4376 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_451
timestamp 1515870181
transform -1 0 4488 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_448
timestamp 1515870181
transform -1 0 4536 0 1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_106
timestamp 1515870181
transform -1 0 4728 0 1 5010
box 0 0 192 200
use BUFX4  BUFX4_71
timestamp 1515870181
transform -1 0 4792 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_250
timestamp 1515870181
transform 1 0 4792 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_253
timestamp 1515870181
transform 1 0 4840 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_258
timestamp 1515870181
transform 1 0 4888 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_272
timestamp 1515870181
transform -1 0 5000 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_319
timestamp 1515870181
transform 1 0 5000 0 1 5010
box 0 0 192 200
use INVX2  INVX2_32
timestamp 1515870181
transform 1 0 5192 0 1 5010
box 0 0 32 200
use FILL  FILL_25_4_0
timestamp 1515870181
transform -1 0 5240 0 1 5010
box 0 0 16 200
use FILL  FILL_25_4_1
timestamp 1515870181
transform -1 0 5256 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_303
timestamp 1515870181
transform -1 0 5448 0 1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_72
timestamp 1515870181
transform 1 0 5448 0 1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_63
timestamp 1515870181
transform -1 0 5560 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_245
timestamp 1515870181
transform -1 0 5624 0 1 5010
box 0 0 64 200
use INVX2  INVX2_5
timestamp 1515870181
transform -1 0 5656 0 1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_260
timestamp 1515870181
transform 1 0 5656 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_292
timestamp 1515870181
transform -1 0 6040 0 1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_232
timestamp 1515870181
transform 1 0 6040 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_246
timestamp 1515870181
transform -1 0 6152 0 1 5010
box 0 0 64 200
use INVX2  INVX2_6
timestamp 1515870181
transform -1 0 6184 0 1 5010
box 0 0 32 200
use FILL  FILL_25_5_0
timestamp 1515870181
transform -1 0 6200 0 1 5010
box 0 0 16 200
use FILL  FILL_25_5_1
timestamp 1515870181
transform -1 0 6216 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_261
timestamp 1515870181
transform -1 0 6408 0 1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_65
timestamp 1515870181
transform 1 0 6408 0 1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_56
timestamp 1515870181
transform -1 0 6520 0 1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_296
timestamp 1515870181
transform 1 0 6520 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_280
timestamp 1515870181
transform -1 0 6904 0 1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_324
timestamp 1515870181
transform -1 0 7096 0 1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_13
timestamp 1515870181
transform 1 0 7096 0 1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_4
timestamp 1515870181
transform -1 0 7208 0 1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_29
timestamp 1515870181
transform 1 0 7208 0 1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_20
timestamp 1515870181
transform -1 0 7320 0 1 5010
box 0 0 64 200
use AOI21X1  AOI21X1_8
timestamp 1515870181
transform 1 0 7320 0 1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_17
timestamp 1515870181
transform -1 0 7432 0 1 5010
box 0 0 48 200
use MUX2X1  MUX2X1_12
timestamp 1515870181
transform -1 0 104 0 -1 5010
box 0 0 96 200
use NAND2X1  NAND2X1_198
timestamp 1515870181
transform 1 0 104 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_212
timestamp 1515870181
transform -1 0 216 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_55
timestamp 1515870181
transform 1 0 216 0 -1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_79
timestamp 1515870181
transform 1 0 408 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_71
timestamp 1515870181
transform -1 0 520 0 -1 5010
box 0 0 64 200
use BUFX4  BUFX4_33
timestamp 1515870181
transform -1 0 584 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_223
timestamp 1515870181
transform 1 0 584 0 -1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_223
timestamp 1515870181
transform 1 0 776 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_209
timestamp 1515870181
transform 1 0 840 0 -1 5010
box 0 0 48 200
use BUFX4  BUFX4_208
timestamp 1515870181
transform -1 0 952 0 -1 5010
box 0 0 64 200
use MUX2X1  MUX2X1_43
timestamp 1515870181
transform 1 0 952 0 -1 5010
box 0 0 96 200
use FILL  FILL_24_0_0
timestamp 1515870181
transform 1 0 1048 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_0_1
timestamp 1515870181
transform 1 0 1064 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1515870181
transform 1 0 1080 0 -1 5010
box 0 0 192 200
use MUX2X1  MUX2X1_11
timestamp 1515870181
transform 1 0 1272 0 -1 5010
box 0 0 96 200
use NAND2X1  NAND2X1_41
timestamp 1515870181
transform 1 0 1368 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_36
timestamp 1515870181
transform -1 0 1480 0 -1 5010
box 0 0 64 200
use MUX2X1  MUX2X1_44
timestamp 1515870181
transform -1 0 1576 0 -1 5010
box 0 0 96 200
use OAI21X1  OAI21X1_69
timestamp 1515870181
transform -1 0 1640 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_77
timestamp 1515870181
transform -1 0 1688 0 -1 5010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_53
timestamp 1515870181
transform 1 0 1688 0 -1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_213
timestamp 1515870181
transform 1 0 1880 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_199
timestamp 1515870181
transform -1 0 1992 0 -1 5010
box 0 0 48 200
use MUX2X1  MUX2X1_15
timestamp 1515870181
transform -1 0 2088 0 -1 5010
box 0 0 96 200
use FILL  FILL_24_1_0
timestamp 1515870181
transform -1 0 2104 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_1_1
timestamp 1515870181
transform -1 0 2120 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_213
timestamp 1515870181
transform -1 0 2312 0 -1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_42
timestamp 1515870181
transform -1 0 2360 0 -1 5010
box 0 0 48 200
use MUX2X1  MUX2X1_14
timestamp 1515870181
transform 1 0 2360 0 -1 5010
box 0 0 96 200
use NAND2X1  NAND2X1_59
timestamp 1515870181
transform -1 0 2504 0 -1 5010
box 0 0 48 200
use MUX2X1  MUX2X1_13
timestamp 1515870181
transform -1 0 2600 0 -1 5010
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_197
timestamp 1515870181
transform -1 0 2792 0 -1 5010
box 0 0 192 200
use MUX2X1  MUX2X1_23
timestamp 1515870181
transform 1 0 2792 0 -1 5010
box 0 0 96 200
use NAND2X1  NAND2X1_45
timestamp 1515870181
transform -1 0 2936 0 -1 5010
box 0 0 48 200
use BUFX4  BUFX4_145
timestamp 1515870181
transform -1 0 3000 0 -1 5010
box 0 0 64 200
use BUFX4  BUFX4_146
timestamp 1515870181
transform 1 0 3000 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_20
timestamp 1515870181
transform 1 0 3064 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_23
timestamp 1515870181
transform -1 0 3176 0 -1 5010
box 0 0 48 200
use FILL  FILL_24_2_0
timestamp 1515870181
transform 1 0 3176 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_2_1
timestamp 1515870181
transform 1 0 3192 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_84
timestamp 1515870181
transform 1 0 3208 0 -1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_424
timestamp 1515870181
transform 1 0 3400 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_485
timestamp 1515870181
transform -1 0 3512 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_299
timestamp 1515870181
transform -1 0 3560 0 -1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_425
timestamp 1515870181
transform 1 0 3560 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_486
timestamp 1515870181
transform -1 0 3672 0 -1 5010
box 0 0 64 200
use BUFX2  BUFX2_31
timestamp 1515870181
transform 1 0 3672 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_502
timestamp 1515870181
transform 1 0 3720 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_441
timestamp 1515870181
transform -1 0 3832 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_341
timestamp 1515870181
transform -1 0 3896 0 -1 5010
box 0 0 64 200
use INVX8  INVX8_5
timestamp 1515870181
transform 1 0 3896 0 -1 5010
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_344
timestamp 1515870181
transform -1 0 4168 0 -1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_100
timestamp 1515870181
transform 1 0 4168 0 -1 5010
box 0 0 48 200
use FILL  FILL_24_3_0
timestamp 1515870181
transform -1 0 4232 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_3_1
timestamp 1515870181
transform -1 0 4248 0 -1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_120
timestamp 1515870181
transform -1 0 4312 0 -1 5010
box 0 0 64 200
use BUFX4  BUFX4_305
timestamp 1515870181
transform 1 0 4312 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_446
timestamp 1515870181
transform 1 0 4376 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_507
timestamp 1515870181
transform -1 0 4488 0 -1 5010
box 0 0 64 200
use INVX1  INVX1_54
timestamp 1515870181
transform -1 0 4520 0 -1 5010
box 0 0 32 200
use INVX8  INVX8_15
timestamp 1515870181
transform 1 0 4520 0 -1 5010
box 0 0 80 200
use DFFPOSX1  DFFPOSX1_311
timestamp 1515870181
transform -1 0 4792 0 -1 5010
box 0 0 192 200
use INVX2  INVX2_24
timestamp 1515870181
transform 1 0 4792 0 -1 5010
box 0 0 32 200
use OAI21X1  OAI21X1_264
timestamp 1515870181
transform -1 0 4888 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_242
timestamp 1515870181
transform 1 0 4888 0 -1 5010
box 0 0 48 200
use BUFX4  BUFX4_26
timestamp 1515870181
transform -1 0 5000 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_267
timestamp 1515870181
transform -1 0 5064 0 -1 5010
box 0 0 64 200
use INVX2  INVX2_27
timestamp 1515870181
transform -1 0 5096 0 -1 5010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_314
timestamp 1515870181
transform -1 0 5288 0 -1 5010
box 0 0 192 200
use FILL  FILL_24_4_0
timestamp 1515870181
transform 1 0 5288 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_4_1
timestamp 1515870181
transform 1 0 5304 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_249
timestamp 1515870181
transform 1 0 5320 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_263
timestamp 1515870181
transform -1 0 5432 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_310
timestamp 1515870181
transform 1 0 5432 0 -1 5010
box 0 0 192 200
use INVX2  INVX2_23
timestamp 1515870181
transform 1 0 5624 0 -1 5010
box 0 0 32 200
use BUFX4  BUFX4_87
timestamp 1515870181
transform 1 0 5656 0 -1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_61
timestamp 1515870181
transform 1 0 5720 0 -1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_52
timestamp 1515870181
transform -1 0 5832 0 -1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_45
timestamp 1515870181
transform 1 0 5832 0 -1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_36
timestamp 1515870181
transform -1 0 5944 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_276
timestamp 1515870181
transform -1 0 6136 0 -1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_56
timestamp 1515870181
transform 1 0 6136 0 -1 5010
box 0 0 48 200
use AOI21X1  AOI21X1_47
timestamp 1515870181
transform -1 0 6248 0 -1 5010
box 0 0 64 200
use FILL  FILL_24_5_0
timestamp 1515870181
transform -1 0 6264 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_5_1
timestamp 1515870181
transform -1 0 6280 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_287
timestamp 1515870181
transform -1 0 6472 0 -1 5010
box 0 0 192 200
use AOI21X1  AOI21X1_40
timestamp 1515870181
transform 1 0 6472 0 -1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_49
timestamp 1515870181
transform -1 0 6584 0 -1 5010
box 0 0 48 200
use NAND3X1  NAND3X1_77
timestamp 1515870181
transform -1 0 6648 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_76
timestamp 1515870181
transform -1 0 6712 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_236
timestamp 1515870181
transform -1 0 6776 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_34
timestamp 1515870181
transform -1 0 6840 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_36
timestamp 1515870181
transform -1 0 6904 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_194
timestamp 1515870181
transform -1 0 6968 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_196
timestamp 1515870181
transform -1 0 7032 0 -1 5010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_244
timestamp 1515870181
transform -1 0 7224 0 -1 5010
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_328
timestamp 1515870181
transform 1 0 7224 0 -1 5010
box 0 0 192 200
use FILL  FILL_25_1
timestamp 1515870181
transform -1 0 7432 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_52
timestamp 1515870181
transform -1 0 200 0 1 4610
box 0 0 192 200
use NAND2X1  NAND2X1_76
timestamp 1515870181
transform 1 0 200 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_68
timestamp 1515870181
transform -1 0 312 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_74
timestamp 1515870181
transform 1 0 312 0 1 4610
box 0 0 192 200
use BUFX4  BUFX4_55
timestamp 1515870181
transform -1 0 568 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_58
timestamp 1515870181
transform -1 0 632 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_64
timestamp 1515870181
transform -1 0 680 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_79
timestamp 1515870181
transform 1 0 680 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_63
timestamp 1515870181
transform 1 0 872 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_69
timestamp 1515870181
transform -1 0 984 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_432
timestamp 1515870181
transform -1 0 1048 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_304
timestamp 1515870181
transform -1 0 1112 0 1 4610
box 0 0 64 200
use FILL  FILL_23_0_0
timestamp 1515870181
transform -1 0 1128 0 1 4610
box 0 0 16 200
use FILL  FILL_23_0_1
timestamp 1515870181
transform -1 0 1144 0 1 4610
box 0 0 16 200
use NOR3X1  NOR3X1_8
timestamp 1515870181
transform -1 0 1272 0 1 4610
box 0 0 128 200
use NOR2X1  NOR2X1_89
timestamp 1515870181
transform 1 0 1272 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_90
timestamp 1515870181
transform 1 0 1320 0 1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_4
timestamp 1515870181
transform 1 0 1368 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_140
timestamp 1515870181
transform -1 0 1496 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_52
timestamp 1515870181
transform 1 0 1496 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_47
timestamp 1515870181
transform -1 0 1608 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1515870181
transform -1 0 1800 0 1 4610
box 0 0 192 200
use BUFX4  BUFX4_171
timestamp 1515870181
transform -1 0 1864 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_313
timestamp 1515870181
transform -1 0 1928 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_436
timestamp 1515870181
transform -1 0 1992 0 1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_186
timestamp 1515870181
transform -1 0 2184 0 1 4610
box 0 0 192 200
use FILL  FILL_23_1_0
timestamp 1515870181
transform 1 0 2184 0 1 4610
box 0 0 16 200
use FILL  FILL_23_1_1
timestamp 1515870181
transform 1 0 2200 0 1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_186
timestamp 1515870181
transform 1 0 2216 0 1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_10
timestamp 1515870181
transform -1 0 2408 0 1 4610
box 0 0 128 200
use NOR2X1  NOR2X1_93
timestamp 1515870181
transform 1 0 2408 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_92
timestamp 1515870181
transform -1 0 2504 0 1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_5
timestamp 1515870181
transform 1 0 2504 0 1 4610
box 0 0 80 200
use OAI21X1  OAI21X1_448
timestamp 1515870181
transform 1 0 2584 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_142
timestamp 1515870181
transform 1 0 2648 0 1 4610
box 0 0 48 200
use BUFX4  BUFX4_32
timestamp 1515870181
transform 1 0 2696 0 1 4610
box 0 0 64 200
use OAI22X1  OAI22X1_8
timestamp 1515870181
transform -1 0 2840 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_148
timestamp 1515870181
transform -1 0 2888 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_164
timestamp 1515870181
transform 1 0 2888 0 1 4610
box 0 0 192 200
use INVX1  INVX1_26
timestamp 1515870181
transform 1 0 3080 0 1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_308
timestamp 1515870181
transform 1 0 3112 0 1 4610
box 0 0 64 200
use FILL  FILL_23_2_0
timestamp 1515870181
transform 1 0 3176 0 1 4610
box 0 0 16 200
use FILL  FILL_23_2_1
timestamp 1515870181
transform 1 0 3192 0 1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_211
timestamp 1515870181
transform 1 0 3208 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_292
timestamp 1515870181
transform 1 0 3272 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_41
timestamp 1515870181
transform 1 0 3320 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_51
timestamp 1515870181
transform 1 0 3384 0 1 4610
box 0 0 64 200
use INVX1  INVX1_30
timestamp 1515870181
transform 1 0 3448 0 1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_315
timestamp 1515870181
transform 1 0 3480 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_291
timestamp 1515870181
transform -1 0 3592 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_201
timestamp 1515870181
transform 1 0 3592 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_298
timestamp 1515870181
transform 1 0 3656 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_151
timestamp 1515870181
transform 1 0 3704 0 1 4610
box 0 0 64 200
use INVX1  INVX1_29
timestamp 1515870181
transform -1 0 3800 0 1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_101
timestamp 1515870181
transform -1 0 3992 0 1 4610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_346
timestamp 1515870181
transform 1 0 3992 0 1 4610
box 0 0 192 200
use FILL  FILL_23_3_0
timestamp 1515870181
transform 1 0 4184 0 1 4610
box 0 0 16 200
use FILL  FILL_23_3_1
timestamp 1515870181
transform 1 0 4200 0 1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_241
timestamp 1515870181
transform 1 0 4216 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_347
timestamp 1515870181
transform 1 0 4280 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_368
timestamp 1515870181
transform -1 0 4376 0 1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_333
timestamp 1515870181
transform 1 0 4376 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_81
timestamp 1515870181
transform 1 0 4424 0 1 4610
box 0 0 64 200
use BUFX2  BUFX2_10
timestamp 1515870181
transform -1 0 4536 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_351
timestamp 1515870181
transform -1 0 4728 0 1 4610
box 0 0 192 200
use BUFX4  BUFX4_169
timestamp 1515870181
transform 1 0 4728 0 1 4610
box 0 0 64 200
use BUFX2  BUFX2_6
timestamp 1515870181
transform -1 0 4840 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_256
timestamp 1515870181
transform 1 0 4840 0 1 4610
box 0 0 64 200
use INVX2  INVX2_16
timestamp 1515870181
transform -1 0 4936 0 1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_271
timestamp 1515870181
transform -1 0 5128 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_475
timestamp 1515870181
transform -1 0 5192 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_401
timestamp 1515870181
transform 1 0 5192 0 1 4610
box 0 0 64 200
use FILL  FILL_23_4_0
timestamp 1515870181
transform 1 0 5256 0 1 4610
box 0 0 16 200
use FILL  FILL_23_4_1
timestamp 1515870181
transform 1 0 5272 0 1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_143
timestamp 1515870181
transform 1 0 5288 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_303
timestamp 1515870181
transform 1 0 5352 0 1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_36
timestamp 1515870181
transform 1 0 5416 0 1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_431
timestamp 1515870181
transform 1 0 5544 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_302
timestamp 1515870181
transform 1 0 5608 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_193
timestamp 1515870181
transform -1 0 5736 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_33
timestamp 1515870181
transform 1 0 5736 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_73
timestamp 1515870181
transform -1 0 5864 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_338
timestamp 1515870181
transform -1 0 5928 0 1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_15
timestamp 1515870181
transform 1 0 5928 0 1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_337
timestamp 1515870181
transform 1 0 6056 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_446
timestamp 1515870181
transform 1 0 6120 0 1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_40
timestamp 1515870181
transform 1 0 6184 0 1 4610
box 0 0 128 200
use FILL  FILL_23_5_0
timestamp 1515870181
transform 1 0 6312 0 1 4610
box 0 0 16 200
use FILL  FILL_23_5_1
timestamp 1515870181
transform 1 0 6328 0 1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_447
timestamp 1515870181
transform 1 0 6344 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_233
timestamp 1515870181
transform 1 0 6408 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_72
timestamp 1515870181
transform -1 0 6536 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_232
timestamp 1515870181
transform 1 0 6536 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_75
timestamp 1515870181
transform -1 0 6664 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_74
timestamp 1515870181
transform -1 0 6728 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_237
timestamp 1515870181
transform -1 0 6792 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_235
timestamp 1515870181
transform 1 0 6792 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_37
timestamp 1515870181
transform 1 0 6856 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_234
timestamp 1515870181
transform 1 0 6920 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_197
timestamp 1515870181
transform 1 0 6984 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_35
timestamp 1515870181
transform -1 0 7112 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_195
timestamp 1515870181
transform 1 0 7112 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_33
timestamp 1515870181
transform -1 0 7224 0 1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_248
timestamp 1515870181
transform 1 0 7224 0 1 4610
box 0 0 192 200
use FILL  FILL_24_1
timestamp 1515870181
transform 1 0 7416 0 1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_215
timestamp 1515870181
transform 1 0 8 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_201
timestamp 1515870181
transform -1 0 120 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_215
timestamp 1515870181
transform 1 0 120 0 -1 4610
box 0 0 192 200
use MUX2X1  MUX2X1_21
timestamp 1515870181
transform 1 0 312 0 -1 4610
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_202
timestamp 1515870181
transform 1 0 408 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_202
timestamp 1515870181
transform 1 0 600 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_187
timestamp 1515870181
transform -1 0 712 0 -1 4610
box 0 0 48 200
use MUX2X1  MUX2X1_28
timestamp 1515870181
transform 1 0 712 0 -1 4610
box 0 0 96 200
use MUX2X1  MUX2X1_45
timestamp 1515870181
transform -1 0 904 0 -1 4610
box 0 0 96 200
use NAND2X1  NAND2X1_394
timestamp 1515870181
transform 1 0 904 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_290
timestamp 1515870181
transform 1 0 952 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_416
timestamp 1515870181
transform 1 0 1000 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_367
timestamp 1515870181
transform 1 0 1048 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_403
timestamp 1515870181
transform -1 0 1160 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_0_0
timestamp 1515870181
transform -1 0 1176 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_1
timestamp 1515870181
transform -1 0 1192 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_476
timestamp 1515870181
transform -1 0 1256 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_162
timestamp 1515870181
transform 1 0 1256 0 -1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_15
timestamp 1515870181
transform -1 0 1384 0 -1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_122
timestamp 1515870181
transform 1 0 1384 0 -1 4610
box 0 0 48 200
use BUFX4  BUFX4_174
timestamp 1515870181
transform -1 0 1496 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_123
timestamp 1515870181
transform 1 0 1496 0 -1 4610
box 0 0 48 200
use NOR3X1  NOR3X1_30
timestamp 1515870181
transform 1 0 1544 0 -1 4610
box 0 0 128 200
use NAND2X1  NAND2X1_297
timestamp 1515870181
transform -1 0 1720 0 -1 4610
box 0 0 48 200
use BUFX4  BUFX4_177
timestamp 1515870181
transform 1 0 1720 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_396
timestamp 1515870181
transform 1 0 1784 0 -1 4610
box 0 0 48 200
use BUFX4  BUFX4_99
timestamp 1515870181
transform 1 0 1832 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_10
timestamp 1515870181
transform 1 0 1896 0 -1 4610
box 0 0 192 200
use NAND2X1  NAND2X1_170
timestamp 1515870181
transform 1 0 2088 0 -1 4610
box 0 0 48 200
use FILL  FILL_22_1_0
timestamp 1515870181
transform 1 0 2136 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_1
timestamp 1515870181
transform 1 0 2152 0 -1 4610
box 0 0 16 200
use MUX2X1  MUX2X1_29
timestamp 1515870181
transform 1 0 2168 0 -1 4610
box 0 0 96 200
use NAND2X1  NAND2X1_47
timestamp 1515870181
transform 1 0 2264 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_42
timestamp 1515870181
transform -1 0 2376 0 -1 4610
box 0 0 64 200
use BUFX4  BUFX4_274
timestamp 1515870181
transform -1 0 2440 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_318
timestamp 1515870181
transform 1 0 2440 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_402
timestamp 1515870181
transform 1 0 2488 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_340
timestamp 1515870181
transform -1 0 2600 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_16
timestamp 1515870181
transform -1 0 2728 0 -1 4610
box 0 0 128 200
use NOR2X1  NOR2X1_101
timestamp 1515870181
transform 1 0 2728 0 -1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_102
timestamp 1515870181
transform -1 0 2824 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_164
timestamp 1515870181
transform 1 0 2824 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_147
timestamp 1515870181
transform -1 0 2936 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_133
timestamp 1515870181
transform 1 0 2936 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_114
timestamp 1515870181
transform -1 0 3048 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_133
timestamp 1515870181
transform 1 0 3048 0 -1 4610
box 0 0 192 200
use FILL  FILL_22_2_0
timestamp 1515870181
transform 1 0 3240 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_1
timestamp 1515870181
transform 1 0 3256 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_117
timestamp 1515870181
transform 1 0 3272 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_97
timestamp 1515870181
transform -1 0 3384 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_341
timestamp 1515870181
transform -1 0 3576 0 -1 4610
box 0 0 192 200
use BUFX4  BUFX4_275
timestamp 1515870181
transform 1 0 3576 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_314
timestamp 1515870181
transform 1 0 3640 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_311
timestamp 1515870181
transform 1 0 3704 0 -1 4610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_103
timestamp 1515870181
transform 1 0 3768 0 -1 4610
box 0 0 192 200
use INVX1  INVX1_39
timestamp 1515870181
transform 1 0 3960 0 -1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_122
timestamp 1515870181
transform 1 0 3992 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_504
timestamp 1515870181
transform 1 0 4056 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_102
timestamp 1515870181
transform -1 0 4168 0 -1 4610
box 0 0 48 200
use INVX8  INVX8_10
timestamp 1515870181
transform -1 0 4248 0 -1 4610
box 0 0 80 200
use FILL  FILL_22_3_0
timestamp 1515870181
transform 1 0 4248 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_3_1
timestamp 1515870181
transform 1 0 4264 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_404
timestamp 1515870181
transform 1 0 4280 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_359
timestamp 1515870181
transform 1 0 4344 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_443
timestamp 1515870181
transform -1 0 4456 0 -1 4610
box 0 0 48 200
use BUFX2  BUFX2_26
timestamp 1515870181
transform -1 0 4504 0 -1 4610
box 0 0 48 200
use INVX8  INVX8_7
timestamp 1515870181
transform -1 0 4584 0 -1 4610
box 0 0 80 200
use NAND2X1  NAND2X1_107
timestamp 1515870181
transform 1 0 4584 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_127
timestamp 1515870181
transform -1 0 4696 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_47
timestamp 1515870181
transform -1 0 4824 0 -1 4610
box 0 0 128 200
use NAND2X1  NAND2X1_234
timestamp 1515870181
transform 1 0 4824 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_474
timestamp 1515870181
transform -1 0 4936 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_400
timestamp 1515870181
transform 1 0 4936 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_29
timestamp 1515870181
transform 1 0 5000 0 -1 4610
box 0 0 128 200
use NAND3X1  NAND3X1_302
timestamp 1515870181
transform -1 0 5192 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_142
timestamp 1515870181
transform 1 0 5192 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_4_0
timestamp 1515870181
transform -1 0 5272 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_4_1
timestamp 1515870181
transform -1 0 5288 0 -1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_192
timestamp 1515870181
transform -1 0 5352 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_32
timestamp 1515870181
transform -1 0 5416 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_430
timestamp 1515870181
transform -1 0 5480 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_301
timestamp 1515870181
transform -1 0 5544 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_7
timestamp 1515870181
transform 1 0 5544 0 -1 4610
box 0 0 128 200
use NOR3X1  NOR3X1_37
timestamp 1515870181
transform -1 0 5800 0 -1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_434
timestamp 1515870181
transform 1 0 5800 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_310
timestamp 1515870181
transform 1 0 5864 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_9
timestamp 1515870181
transform 1 0 5928 0 -1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_311
timestamp 1515870181
transform 1 0 6056 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_43
timestamp 1515870181
transform -1 0 6184 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_435
timestamp 1515870181
transform -1 0 6248 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_5_0
timestamp 1515870181
transform 1 0 6248 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_5_1
timestamp 1515870181
transform 1 0 6264 0 -1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_203
timestamp 1515870181
transform 1 0 6280 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_147
timestamp 1515870181
transform -1 0 6408 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_146
timestamp 1515870181
transform -1 0 6472 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_145
timestamp 1515870181
transform -1 0 6536 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_144
timestamp 1515870181
transform -1 0 6600 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_306
timestamp 1515870181
transform -1 0 6664 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_307
timestamp 1515870181
transform -1 0 6728 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_305
timestamp 1515870181
transform 1 0 6728 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_304
timestamp 1515870181
transform 1 0 6792 0 -1 4610
box 0 0 64 200
use AOI21X1  AOI21X1_31
timestamp 1515870181
transform 1 0 6856 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_40
timestamp 1515870181
transform -1 0 6968 0 -1 4610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_255
timestamp 1515870181
transform -1 0 7160 0 -1 4610
box 0 0 192 200
use INVX2  INVX2_31
timestamp 1515870181
transform -1 0 7192 0 -1 4610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_322
timestamp 1515870181
transform 1 0 7192 0 -1 4610
box 0 0 192 200
use INVX2  INVX2_15
timestamp 1515870181
transform -1 0 7416 0 -1 4610
box 0 0 32 200
use FILL  FILL_23_1
timestamp 1515870181
transform -1 0 7432 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_231
timestamp 1515870181
transform 1 0 8 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_218
timestamp 1515870181
transform -1 0 120 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_231
timestamp 1515870181
transform 1 0 120 0 1 4210
box 0 0 192 200
use INVX1  INVX1_23
timestamp 1515870181
transform -1 0 344 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_303
timestamp 1515870181
transform 1 0 344 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_63
timestamp 1515870181
transform 1 0 408 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_79
timestamp 1515870181
transform 1 0 600 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_87
timestamp 1515870181
transform -1 0 712 0 1 4210
box 0 0 48 200
use BUFX4  BUFX4_76
timestamp 1515870181
transform -1 0 776 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_320
timestamp 1515870181
transform -1 0 840 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_444
timestamp 1515870181
transform 1 0 840 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_311
timestamp 1515870181
transform 1 0 904 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_331
timestamp 1515870181
transform -1 0 1016 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_146
timestamp 1515870181
transform 1 0 1016 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_167
timestamp 1515870181
transform 1 0 1064 0 1 4210
box 0 0 48 200
use FILL  FILL_21_0_0
timestamp 1515870181
transform 1 0 1112 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_1
timestamp 1515870181
transform 1 0 1128 0 1 4210
box 0 0 16 200
use MUX2X1  MUX2X1_20
timestamp 1515870181
transform 1 0 1144 0 1 4210
box 0 0 96 200
use OAI22X1  OAI22X1_7
timestamp 1515870181
transform 1 0 1240 0 1 4210
box 0 0 80 200
use NOR2X1  NOR2X1_99
timestamp 1515870181
transform 1 0 1320 0 1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_98
timestamp 1515870181
transform 1 0 1368 0 1 4210
box 0 0 48 200
use NOR3X1  NOR3X1_14
timestamp 1515870181
transform 1 0 1416 0 1 4210
box 0 0 128 200
use BUFX4  BUFX4_159
timestamp 1515870181
transform 1 0 1544 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_160
timestamp 1515870181
transform 1 0 1608 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_60
timestamp 1515870181
transform -1 0 1720 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_70
timestamp 1515870181
transform -1 0 1912 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_54
timestamp 1515870181
transform -1 0 1976 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_60
timestamp 1515870181
transform 1 0 1976 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_170
timestamp 1515870181
transform -1 0 2104 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_293
timestamp 1515870181
transform -1 0 2168 0 1 4210
box 0 0 64 200
use FILL  FILL_21_1_0
timestamp 1515870181
transform -1 0 2184 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_1
timestamp 1515870181
transform -1 0 2200 0 1 4210
box 0 0 16 200
use OAI22X1  OAI22X1_10
timestamp 1515870181
transform -1 0 2280 0 1 4210
box 0 0 80 200
use NOR2X1  NOR2X1_108
timestamp 1515870181
transform 1 0 2280 0 1 4210
box 0 0 48 200
use BUFX4  BUFX4_294
timestamp 1515870181
transform 1 0 2328 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_170
timestamp 1515870181
transform 1 0 2392 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_170
timestamp 1515870181
transform 1 0 2584 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_167
timestamp 1515870181
transform 1 0 2648 0 1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_132
timestamp 1515870181
transform 1 0 2840 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_113
timestamp 1515870181
transform 1 0 3032 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_132
timestamp 1515870181
transform -1 0 3144 0 1 4210
box 0 0 64 200
use INVX1  INVX1_25
timestamp 1515870181
transform 1 0 3144 0 1 4210
box 0 0 32 200
use FILL  FILL_21_2_0
timestamp 1515870181
transform 1 0 3176 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_1
timestamp 1515870181
transform 1 0 3192 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_306
timestamp 1515870181
transform 1 0 3208 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_138
timestamp 1515870181
transform 1 0 3272 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_138
timestamp 1515870181
transform 1 0 3464 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_119
timestamp 1515870181
transform -1 0 3576 0 1 4210
box 0 0 48 200
use INVX1  INVX1_55
timestamp 1515870181
transform 1 0 3576 0 1 4210
box 0 0 32 200
use NAND3X1  NAND3X1_71
timestamp 1515870181
transform 1 0 3608 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_305
timestamp 1515870181
transform -1 0 3736 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_116
timestamp 1515870181
transform 1 0 3736 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_96
timestamp 1515870181
transform -1 0 3848 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_340
timestamp 1515870181
transform -1 0 4040 0 1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_231
timestamp 1515870181
transform 1 0 4040 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_491
timestamp 1515870181
transform 1 0 4104 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_430
timestamp 1515870181
transform -1 0 4216 0 1 4210
box 0 0 48 200
use FILL  FILL_21_3_0
timestamp 1515870181
transform 1 0 4216 0 1 4210
box 0 0 16 200
use FILL  FILL_21_3_1
timestamp 1515870181
transform 1 0 4232 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_90
timestamp 1515870181
transform 1 0 4248 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_360
timestamp 1515870181
transform 1 0 4440 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_334
timestamp 1515870181
transform -1 0 4552 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_102
timestamp 1515870181
transform -1 0 4744 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_305
timestamp 1515870181
transform 1 0 4744 0 1 4210
box 0 0 48 200
use INVX1  INVX1_34
timestamp 1515870181
transform 1 0 4792 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_503
timestamp 1515870181
transform 1 0 4824 0 1 4210
box 0 0 64 200
use BUFX2  BUFX2_22
timestamp 1515870181
transform 1 0 4888 0 1 4210
box 0 0 48 200
use NAND2X1  NAND2X1_442
timestamp 1515870181
transform -1 0 4984 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_221
timestamp 1515870181
transform 1 0 4984 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_248
timestamp 1515870181
transform -1 0 5112 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_263
timestamp 1515870181
transform 1 0 5112 0 1 4210
box 0 0 192 200
use FILL  FILL_21_4_0
timestamp 1515870181
transform 1 0 5304 0 1 4210
box 0 0 16 200
use FILL  FILL_21_4_1
timestamp 1515870181
transform 1 0 5320 0 1 4210
box 0 0 16 200
use INVX2  INVX2_8
timestamp 1515870181
transform 1 0 5336 0 1 4210
box 0 0 32 200
use BUFX4  BUFX4_225
timestamp 1515870181
transform -1 0 5432 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_443
timestamp 1515870181
transform 1 0 5432 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_223
timestamp 1515870181
transform 1 0 5496 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_147
timestamp 1515870181
transform 1 0 5560 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_295
timestamp 1515870181
transform -1 0 5816 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_233
timestamp 1515870181
transform 1 0 5816 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_53
timestamp 1515870181
transform -1 0 5928 0 1 4210
box 0 0 64 200
use BUFX4  BUFX4_228
timestamp 1515870181
transform 1 0 5928 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_213
timestamp 1515870181
transform 1 0 5992 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_320
timestamp 1515870181
transform -1 0 6120 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_202
timestamp 1515870181
transform 1 0 6120 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_42
timestamp 1515870181
transform 1 0 6184 0 1 4210
box 0 0 64 200
use FILL  FILL_21_5_0
timestamp 1515870181
transform -1 0 6264 0 1 4210
box 0 0 16 200
use FILL  FILL_21_5_1
timestamp 1515870181
transform -1 0 6280 0 1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_439
timestamp 1515870181
transform -1 0 6344 0 1 4210
box 0 0 64 200
use AOI21X1  AOI21X1_53
timestamp 1515870181
transform 1 0 6344 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_62
timestamp 1515870181
transform 1 0 6408 0 1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_293
timestamp 1515870181
transform -1 0 6648 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_382
timestamp 1515870181
transform -1 0 6696 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_46
timestamp 1515870181
transform -1 0 6760 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_47
timestamp 1515870181
transform -1 0 6824 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_44
timestamp 1515870181
transform -1 0 6888 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_45
timestamp 1515870181
transform -1 0 6952 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_204
timestamp 1515870181
transform -1 0 7016 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_207
timestamp 1515870181
transform 1 0 7016 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_206
timestamp 1515870181
transform -1 0 7144 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_205
timestamp 1515870181
transform -1 0 7208 0 1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_325
timestamp 1515870181
transform -1 0 7400 0 1 4210
box 0 0 192 200
use FILL  FILL_22_1
timestamp 1515870181
transform 1 0 7400 0 1 4210
box 0 0 16 200
use FILL  FILL_22_2
timestamp 1515870181
transform 1 0 7416 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_232
timestamp 1515870181
transform 1 0 8 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_232
timestamp 1515870181
transform 1 0 200 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_219
timestamp 1515870181
transform -1 0 312 0 -1 4210
box 0 0 48 200
use INVX1  INVX1_43
timestamp 1515870181
transform 1 0 312 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_339
timestamp 1515870181
transform 1 0 344 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_289
timestamp 1515870181
transform -1 0 456 0 -1 4210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_228
timestamp 1515870181
transform -1 0 648 0 -1 4210
box 0 0 192 200
use BUFX4  BUFX4_68
timestamp 1515870181
transform -1 0 712 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_269
timestamp 1515870181
transform -1 0 776 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_51
timestamp 1515870181
transform 1 0 776 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_38
timestamp 1515870181
transform 1 0 840 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_330
timestamp 1515870181
transform 1 0 872 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_400
timestamp 1515870181
transform 1 0 936 0 -1 4210
box 0 0 48 200
use BUFX4  BUFX4_270
timestamp 1515870181
transform 1 0 984 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_358
timestamp 1515870181
transform 1 0 1048 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_0_0
timestamp 1515870181
transform -1 0 1128 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_1
timestamp 1515870181
transform -1 0 1144 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_183
timestamp 1515870181
transform -1 0 1208 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_183
timestamp 1515870181
transform -1 0 1400 0 -1 4210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1515870181
transform 1 0 1400 0 -1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_44
timestamp 1515870181
transform 1 0 1592 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_39
timestamp 1515870181
transform -1 0 1704 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_200
timestamp 1515870181
transform -1 0 1768 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_321
timestamp 1515870181
transform -1 0 1832 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_279
timestamp 1515870181
transform 1 0 1832 0 -1 4210
box 0 0 64 200
use MUX2X1  MUX2X1_16
timestamp 1515870181
transform -1 0 1992 0 -1 4210
box 0 0 96 200
use BUFX4  BUFX4_5
timestamp 1515870181
transform -1 0 2056 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_183
timestamp 1515870181
transform 1 0 2056 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_198
timestamp 1515870181
transform -1 0 2168 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_1_0
timestamp 1515870181
transform -1 0 2184 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_1
timestamp 1515870181
transform -1 0 2200 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_198
timestamp 1515870181
transform -1 0 2392 0 -1 4210
box 0 0 192 200
use NOR2X1  NOR2X1_107
timestamp 1515870181
transform 1 0 2392 0 -1 4210
box 0 0 48 200
use NOR3X1  NOR3X1_20
timestamp 1515870181
transform 1 0 2440 0 -1 4210
box 0 0 128 200
use INVX1  INVX1_56
timestamp 1515870181
transform -1 0 2600 0 -1 4210
box 0 0 32 200
use NAND2X1  NAND2X1_153
timestamp 1515870181
transform 1 0 2600 0 -1 4210
box 0 0 48 200
use OAI22X1  OAI22X1_6
timestamp 1515870181
transform 1 0 2648 0 -1 4210
box 0 0 80 200
use NOR2X1  NOR2X1_144
timestamp 1515870181
transform -1 0 2776 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_167
timestamp 1515870181
transform 1 0 2776 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_150
timestamp 1515870181
transform -1 0 2888 0 -1 4210
box 0 0 48 200
use BUFX4  BUFX4_143
timestamp 1515870181
transform 1 0 2888 0 -1 4210
box 0 0 64 200
use INVX1  INVX1_41
timestamp 1515870181
transform 1 0 2952 0 -1 4210
box 0 0 32 200
use BUFX4  BUFX4_319
timestamp 1515870181
transform -1 0 3048 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_172
timestamp 1515870181
transform 1 0 3048 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_2_0
timestamp 1515870181
transform 1 0 3112 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_1
timestamp 1515870181
transform 1 0 3128 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_31
timestamp 1515870181
transform 1 0 3144 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_31
timestamp 1515870181
transform 1 0 3336 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_34
timestamp 1515870181
transform 1 0 3400 0 -1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_94
timestamp 1515870181
transform -1 0 3496 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_48
timestamp 1515870181
transform -1 0 3560 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_316
timestamp 1515870181
transform -1 0 3624 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_38
timestamp 1515870181
transform 1 0 3624 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_100
timestamp 1515870181
transform 1 0 3688 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_198
timestamp 1515870181
transform -1 0 3800 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_143
timestamp 1515870181
transform 1 0 3800 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_437
timestamp 1515870181
transform 1 0 3848 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_208
timestamp 1515870181
transform 1 0 3912 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_334
timestamp 1515870181
transform -1 0 4040 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_147
timestamp 1515870181
transform 1 0 4040 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_445
timestamp 1515870181
transform -1 0 4152 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_309
timestamp 1515870181
transform -1 0 4216 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_3_0
timestamp 1515870181
transform -1 0 4232 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_3_1
timestamp 1515870181
transform -1 0 4248 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_312
timestamp 1515870181
transform -1 0 4296 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_332
timestamp 1515870181
transform -1 0 4360 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_98
timestamp 1515870181
transform -1 0 4424 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_258
timestamp 1515870181
transform -1 0 4488 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_457
timestamp 1515870181
transform -1 0 4552 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_361
timestamp 1515870181
transform -1 0 4616 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_312
timestamp 1515870181
transform -1 0 4680 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_343
timestamp 1515870181
transform -1 0 4872 0 -1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_99
timestamp 1515870181
transform 1 0 4872 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_119
timestamp 1515870181
transform -1 0 4984 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_318
timestamp 1515870181
transform 1 0 4984 0 -1 4210
box 0 0 64 200
use INVX8  INVX8_6
timestamp 1515870181
transform 1 0 5048 0 -1 4210
box 0 0 80 200
use BUFX4  BUFX4_6
timestamp 1515870181
transform -1 0 5192 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_328
timestamp 1515870181
transform 1 0 5192 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_4_0
timestamp 1515870181
transform 1 0 5256 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_4_1
timestamp 1515870181
transform 1 0 5272 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_329
timestamp 1515870181
transform 1 0 5288 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_63
timestamp 1515870181
transform -1 0 5416 0 -1 4210
box 0 0 64 200
use NOR3X1  NOR3X1_39
timestamp 1515870181
transform -1 0 5544 0 -1 4210
box 0 0 128 200
use OAI21X1  OAI21X1_442
timestamp 1515870181
transform 1 0 5544 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_222
timestamp 1515870181
transform 1 0 5608 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_64
timestamp 1515870181
transform 1 0 5672 0 -1 4210
box 0 0 48 200
use AOI21X1  AOI21X1_55
timestamp 1515870181
transform -1 0 5784 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_20
timestamp 1515870181
transform -1 0 5848 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_218
timestamp 1515870181
transform -1 0 5912 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_21
timestamp 1515870181
transform 1 0 5912 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_182
timestamp 1515870181
transform -1 0 6040 0 -1 4210
box 0 0 64 200
use NOR3X1  NOR3X1_11
timestamp 1515870181
transform 1 0 6040 0 -1 4210
box 0 0 128 200
use OAI21X1  OAI21X1_247
timestamp 1515870181
transform -1 0 6232 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_5_0
timestamp 1515870181
transform 1 0 6232 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_5_1
timestamp 1515870181
transform 1 0 6248 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_319
timestamp 1515870181
transform 1 0 6264 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_52
timestamp 1515870181
transform 1 0 6328 0 -1 4210
box 0 0 64 200
use NOR3X1  NOR3X1_38
timestamp 1515870181
transform 1 0 6392 0 -1 4210
box 0 0 128 200
use OAI21X1  OAI21X1_438
timestamp 1515870181
transform 1 0 6520 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_212
timestamp 1515870181
transform 1 0 6584 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_186
timestamp 1515870181
transform 1 0 6648 0 -1 4210
box 0 0 64 200
use INVX2  INVX2_7
timestamp 1515870181
transform -1 0 6744 0 -1 4210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_262
timestamp 1515870181
transform -1 0 6936 0 -1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_55
timestamp 1515870181
transform -1 0 7000 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_215
timestamp 1515870181
transform 1 0 7000 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_297
timestamp 1515870181
transform -1 0 7128 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_80
timestamp 1515870181
transform 1 0 7128 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_107
timestamp 1515870181
transform 1 0 7192 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_14
timestamp 1515870181
transform 1 0 7256 0 -1 4210
box 0 0 48 200
use AOI21X1  AOI21X1_5
timestamp 1515870181
transform -1 0 7368 0 -1 4210
box 0 0 64 200
use BUFX4  BUFX4_290
timestamp 1515870181
transform 1 0 7368 0 -1 4210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_230
timestamp 1515870181
transform 1 0 8 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_230
timestamp 1515870181
transform -1 0 264 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_217
timestamp 1515870181
transform -1 0 312 0 1 3810
box 0 0 48 200
use INVX1  INVX1_33
timestamp 1515870181
transform 1 0 312 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_321
timestamp 1515870181
transform 1 0 344 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_215
timestamp 1515870181
transform 1 0 408 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_228
timestamp 1515870181
transform -1 0 520 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_220
timestamp 1515870181
transform 1 0 520 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_206
timestamp 1515870181
transform -1 0 632 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_76
timestamp 1515870181
transform 1 0 632 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_220
timestamp 1515870181
transform 1 0 696 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_406
timestamp 1515870181
transform 1 0 888 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_456
timestamp 1515870181
transform -1 0 1000 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_70
timestamp 1515870181
transform 1 0 1000 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_78
timestamp 1515870181
transform -1 0 1112 0 1 3810
box 0 0 48 200
use FILL  FILL_19_0_0
timestamp 1515870181
transform 1 0 1112 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_1
timestamp 1515870181
transform 1 0 1128 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_54
timestamp 1515870181
transform 1 0 1144 0 1 3810
box 0 0 192 200
use MUX2X1  MUX2X1_18
timestamp 1515870181
transform -1 0 1432 0 1 3810
box 0 0 96 200
use NAND2X1  NAND2X1_200
timestamp 1515870181
transform 1 0 1432 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_214
timestamp 1515870181
transform -1 0 1544 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_214
timestamp 1515870181
transform -1 0 1736 0 1 3810
box 0 0 192 200
use BUFX4  BUFX4_197
timestamp 1515870181
transform 1 0 1736 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_203
timestamp 1515870181
transform -1 0 1864 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_166
timestamp 1515870181
transform -1 0 1912 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_38
timestamp 1515870181
transform 1 0 1912 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1515870181
transform 1 0 1976 0 1 3810
box 0 0 192 200
use FILL  FILL_19_1_0
timestamp 1515870181
transform 1 0 2168 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_1
timestamp 1515870181
transform 1 0 2184 0 1 3810
box 0 0 16 200
use NOR2X1  NOR2X1_152
timestamp 1515870181
transform 1 0 2200 0 1 3810
box 0 0 48 200
use MUX2X1  MUX2X1_17
timestamp 1515870181
transform 1 0 2248 0 1 3810
box 0 0 96 200
use NAND2X1  NAND2X1_398
timestamp 1515870181
transform 1 0 2344 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_440
timestamp 1515870181
transform -1 0 2456 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_304
timestamp 1515870181
transform 1 0 2456 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_322
timestamp 1515870181
transform -1 0 2568 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_96
timestamp 1515870181
transform -1 0 2616 0 1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_95
timestamp 1515870181
transform -1 0 2664 0 1 3810
box 0 0 48 200
use NOR3X1  NOR3X1_12
timestamp 1515870181
transform 1 0 2664 0 1 3810
box 0 0 128 200
use NAND2X1  NAND2X1_151
timestamp 1515870181
transform 1 0 2792 0 1 3810
box 0 0 48 200
use BUFX4  BUFX4_144
timestamp 1515870181
transform -1 0 2904 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_165
timestamp 1515870181
transform 1 0 2904 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_165
timestamp 1515870181
transform 1 0 3096 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_148
timestamp 1515870181
transform -1 0 3208 0 1 3810
box 0 0 48 200
use FILL  FILL_19_2_0
timestamp 1515870181
transform 1 0 3208 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_1
timestamp 1515870181
transform 1 0 3224 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_370
timestamp 1515870181
transform 1 0 3240 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_87
timestamp 1515870181
transform 1 0 3288 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_313
timestamp 1515870181
transform -1 0 3528 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_333
timestamp 1515870181
transform -1 0 3592 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_91
timestamp 1515870181
transform 1 0 3592 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_307
timestamp 1515870181
transform -1 0 3704 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_141
timestamp 1515870181
transform 1 0 3704 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_433
timestamp 1515870181
transform -1 0 3816 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_228
timestamp 1515870181
transform -1 0 3880 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_68
timestamp 1515870181
transform -1 0 3944 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_163
timestamp 1515870181
transform 1 0 3944 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_124
timestamp 1515870181
transform 1 0 3992 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_104
timestamp 1515870181
transform -1 0 4104 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_348
timestamp 1515870181
transform 1 0 4104 0 1 3810
box 0 0 192 200
use FILL  FILL_19_3_0
timestamp 1515870181
transform 1 0 4296 0 1 3810
box 0 0 16 200
use FILL  FILL_19_3_1
timestamp 1515870181
transform 1 0 4312 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_477
timestamp 1515870181
transform 1 0 4328 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_377
timestamp 1515870181
transform -1 0 4456 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_153
timestamp 1515870181
transform 1 0 4456 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_261
timestamp 1515870181
transform 1 0 4504 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_109
timestamp 1515870181
transform 1 0 4568 0 1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_101
timestamp 1515870181
transform 1 0 4616 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_98
timestamp 1515870181
transform -1 0 4728 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_323
timestamp 1515870181
transform 1 0 4728 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_118
timestamp 1515870181
transform -1 0 4856 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_61
timestamp 1515870181
transform 1 0 4856 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_342
timestamp 1515870181
transform -1 0 5112 0 1 3810
box 0 0 192 200
use NOR3X1  NOR3X1_13
timestamp 1515870181
transform -1 0 5240 0 1 3810
box 0 0 128 200
use FILL  FILL_19_4_0
timestamp 1515870181
transform 1 0 5240 0 1 3810
box 0 0 16 200
use FILL  FILL_19_4_1
timestamp 1515870181
transform 1 0 5256 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_356
timestamp 1515870181
transform 1 0 5272 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_93
timestamp 1515870181
transform 1 0 5336 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_62
timestamp 1515870181
transform -1 0 5464 0 1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_19
timestamp 1515870181
transform 1 0 5464 0 1 3810
box 0 0 128 200
use DFFPOSX1  DFFPOSX1_279
timestamp 1515870181
transform -1 0 5784 0 1 3810
box 0 0 192 200
use AOI21X1  AOI21X1_54
timestamp 1515870181
transform 1 0 5784 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_63
timestamp 1515870181
transform -1 0 5896 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_277
timestamp 1515870181
transform 1 0 5896 0 1 3810
box 0 0 192 200
use AOI21X1  AOI21X1_37
timestamp 1515870181
transform 1 0 6088 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_46
timestamp 1515870181
transform 1 0 6152 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_38
timestamp 1515870181
transform 1 0 6200 0 1 3810
box 0 0 64 200
use FILL  FILL_19_5_0
timestamp 1515870181
transform -1 0 6280 0 1 3810
box 0 0 16 200
use FILL  FILL_19_5_1
timestamp 1515870181
transform -1 0 6296 0 1 3810
box 0 0 16 200
use NOR2X1  NOR2X1_47
timestamp 1515870181
transform -1 0 6344 0 1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_278
timestamp 1515870181
transform 1 0 6344 0 1 3810
box 0 0 192 200
use BUFX4  BUFX4_298
timestamp 1515870181
transform 1 0 6536 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_262
timestamp 1515870181
transform 1 0 6600 0 1 3810
box 0 0 48 200
use BUFX4  BUFX4_260
timestamp 1515870181
transform -1 0 6712 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_56
timestamp 1515870181
transform -1 0 6776 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_57
timestamp 1515870181
transform -1 0 6840 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_54
timestamp 1515870181
transform -1 0 6904 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_214
timestamp 1515870181
transform -1 0 6968 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_217
timestamp 1515870181
transform 1 0 6968 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_216
timestamp 1515870181
transform 1 0 7032 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_15
timestamp 1515870181
transform 1 0 7096 0 1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_6
timestamp 1515870181
transform -1 0 7208 0 1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_246
timestamp 1515870181
transform -1 0 7400 0 1 3810
box 0 0 192 200
use FILL  FILL_20_1
timestamp 1515870181
transform 1 0 7400 0 1 3810
box 0 0 16 200
use FILL  FILL_20_2
timestamp 1515870181
transform 1 0 7416 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_38
timestamp 1515870181
transform -1 0 200 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_92
timestamp 1515870181
transform -1 0 264 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_88
timestamp 1515870181
transform -1 0 328 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_303
timestamp 1515870181
transform -1 0 376 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_317
timestamp 1515870181
transform -1 0 424 0 -1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_36
timestamp 1515870181
transform -1 0 616 0 -1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_60
timestamp 1515870181
transform 1 0 616 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_74
timestamp 1515870181
transform -1 0 872 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_84
timestamp 1515870181
transform -1 0 920 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_310
timestamp 1515870181
transform -1 0 968 0 -1 3810
box 0 0 48 200
use MUX2X1  MUX2X1_36
timestamp 1515870181
transform 1 0 968 0 -1 3810
box 0 0 96 200
use NAND2X1  NAND2X1_332
timestamp 1515870181
transform 1 0 1064 0 -1 3810
box 0 0 48 200
use FILL  FILL_18_0_0
timestamp 1515870181
transform 1 0 1112 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_1
timestamp 1515870181
transform 1 0 1128 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_464
timestamp 1515870181
transform 1 0 1144 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_410
timestamp 1515870181
transform -1 0 1256 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_346
timestamp 1515870181
transform 1 0 1256 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_376
timestamp 1515870181
transform -1 0 1368 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_178
timestamp 1515870181
transform -1 0 1432 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_209
timestamp 1515870181
transform -1 0 1496 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_156
timestamp 1515870181
transform 1 0 1496 0 -1 3810
box 0 0 48 200
use OAI22X1  OAI22X1_12
timestamp 1515870181
transform 1 0 1544 0 -1 3810
box 0 0 80 200
use NOR2X1  NOR2X1_114
timestamp 1515870181
transform 1 0 1624 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_113
timestamp 1515870181
transform 1 0 1672 0 -1 3810
box 0 0 48 200
use NOR3X1  NOR3X1_24
timestamp 1515870181
transform 1 0 1720 0 -1 3810
box 0 0 128 200
use OAI21X1  OAI21X1_182
timestamp 1515870181
transform 1 0 1848 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_182
timestamp 1515870181
transform 1 0 1912 0 -1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_43
timestamp 1515870181
transform -1 0 2152 0 -1 3810
box 0 0 48 200
use FILL  FILL_18_1_0
timestamp 1515870181
transform 1 0 2152 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_1
timestamp 1515870181
transform 1 0 2168 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_26
timestamp 1515870181
transform 1 0 2184 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_26
timestamp 1515870181
transform 1 0 2376 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_29
timestamp 1515870181
transform -1 0 2488 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_335
timestamp 1515870181
transform -1 0 2536 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_362
timestamp 1515870181
transform -1 0 2600 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_168
timestamp 1515870181
transform 1 0 2600 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_168
timestamp 1515870181
transform 1 0 2792 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_175
timestamp 1515870181
transform 1 0 2856 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_175
timestamp 1515870181
transform -1 0 3112 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_158
timestamp 1515870181
transform -1 0 3160 0 -1 3810
box 0 0 48 200
use INVX1  INVX1_81
timestamp 1515870181
transform 1 0 3160 0 -1 3810
box 0 0 32 200
use FILL  FILL_18_2_0
timestamp 1515870181
transform 1 0 3192 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_1
timestamp 1515870181
transform 1 0 3208 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_407
timestamp 1515870181
transform 1 0 3224 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_31
timestamp 1515870181
transform 1 0 3288 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_488
timestamp 1515870181
transform 1 0 3320 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_427
timestamp 1515870181
transform -1 0 3432 0 -1 3810
box 0 0 48 200
use BUFX4  BUFX4_179
timestamp 1515870181
transform 1 0 3432 0 -1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_39
timestamp 1515870181
transform -1 0 3560 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_295
timestamp 1515870181
transform 1 0 3560 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_199
timestamp 1515870181
transform -1 0 3672 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_395
timestamp 1515870181
transform 1 0 3672 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_149
timestamp 1515870181
transform -1 0 3784 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_372
timestamp 1515870181
transform 1 0 3784 0 -1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_124
timestamp 1515870181
transform 1 0 3832 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_309
timestamp 1515870181
transform -1 0 3944 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_417
timestamp 1515870181
transform 1 0 3944 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_316
timestamp 1515870181
transform -1 0 4040 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_401
timestamp 1515870181
transform 1 0 4040 0 -1 3810
box 0 0 48 200
use BUFX4  BUFX4_38
timestamp 1515870181
transform -1 0 4152 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_406
timestamp 1515870181
transform 1 0 4152 0 -1 3810
box 0 0 64 200
use FILL  FILL_18_3_0
timestamp 1515870181
transform -1 0 4232 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_1
timestamp 1515870181
transform -1 0 4248 0 -1 3810
box 0 0 16 200
use NAND3X1  NAND3X1_99
timestamp 1515870181
transform -1 0 4312 0 -1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_259
timestamp 1515870181
transform -1 0 4376 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_337
timestamp 1515870181
transform 1 0 4376 0 -1 3810
box 0 0 48 200
use NAND2X1  NAND2X1_407
timestamp 1515870181
transform 1 0 4424 0 -1 3810
box 0 0 48 200
use BUFX4  BUFX4_104
timestamp 1515870181
transform -1 0 4536 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_149
timestamp 1515870181
transform 1 0 4536 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_449
timestamp 1515870181
transform 1 0 4584 0 -1 3810
box 0 0 64 200
use BUFX2  BUFX2_12
timestamp 1515870181
transform 1 0 4648 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_343
timestamp 1515870181
transform 1 0 4696 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_103
timestamp 1515870181
transform -1 0 4808 0 -1 3810
box 0 0 48 200
use INVX8  INVX8_12
timestamp 1515870181
transform -1 0 4888 0 -1 3810
box 0 0 80 200
use BUFX4  BUFX4_117
timestamp 1515870181
transform -1 0 4952 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_201
timestamp 1515870181
transform -1 0 5016 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_95
timestamp 1515870181
transform 1 0 5016 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_298
timestamp 1515870181
transform 1 0 5080 0 -1 3810
box 0 0 192 200
use FILL  FILL_18_4_0
timestamp 1515870181
transform 1 0 5272 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_4_1
timestamp 1515870181
transform 1 0 5288 0 -1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_58
timestamp 1515870181
transform 1 0 5304 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_67
timestamp 1515870181
transform 1 0 5368 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_253
timestamp 1515870181
transform 1 0 5416 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_455
timestamp 1515870181
transform -1 0 5544 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_355
timestamp 1515870181
transform 1 0 5544 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_454
timestamp 1515870181
transform 1 0 5608 0 -1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_42
timestamp 1515870181
transform 1 0 5672 0 -1 3810
box 0 0 128 200
use AOI21X1  AOI21X1_39
timestamp 1515870181
transform 1 0 5800 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_48
timestamp 1515870181
transform 1 0 5864 0 -1 3810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_294
timestamp 1515870181
transform 1 0 5912 0 -1 3810
box 0 0 192 200
use BUFX4  BUFX4_18
timestamp 1515870181
transform -1 0 6168 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_262
timestamp 1515870181
transform 1 0 6168 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_239
timestamp 1515870181
transform 1 0 6232 0 -1 3810
box 0 0 48 200
use FILL  FILL_18_5_0
timestamp 1515870181
transform -1 0 6296 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_5_1
timestamp 1515870181
transform -1 0 6312 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_248
timestamp 1515870181
transform -1 0 6376 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_253
timestamp 1515870181
transform -1 0 6440 0 -1 3810
box 0 0 64 200
use INVX2  INVX2_13
timestamp 1515870181
transform -1 0 6472 0 -1 3810
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_268
timestamp 1515870181
transform -1 0 6664 0 -1 3810
box 0 0 192 200
use BUFX4  BUFX4_217
timestamp 1515870181
transform -1 0 6728 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_15
timestamp 1515870181
transform 1 0 6728 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_118
timestamp 1515870181
transform -1 0 6856 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_30
timestamp 1515870181
transform -1 0 6904 0 -1 3810
box 0 0 48 200
use AOI21X1  AOI21X1_21
timestamp 1515870181
transform -1 0 6968 0 -1 3810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_245
timestamp 1515870181
transform -1 0 7160 0 -1 3810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_326
timestamp 1515870181
transform -1 0 7352 0 -1 3810
box 0 0 192 200
use AOI21X1  AOI21X1_22
timestamp 1515870181
transform 1 0 7352 0 -1 3810
box 0 0 64 200
use FILL  FILL_19_1
timestamp 1515870181
transform -1 0 7432 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_91
timestamp 1515870181
transform 1 0 8 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_103
timestamp 1515870181
transform 1 0 72 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_87
timestamp 1515870181
transform 1 0 136 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_104
timestamp 1515870181
transform -1 0 264 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_345
timestamp 1515870181
transform -1 0 312 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_236
timestamp 1515870181
transform 1 0 312 0 1 3410
box 0 0 192 200
use INVX1  INVX1_63
timestamp 1515870181
transform 1 0 504 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_375
timestamp 1515870181
transform 1 0 536 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_58
timestamp 1515870181
transform -1 0 792 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_82
timestamp 1515870181
transform 1 0 792 0 1 3410
box 0 0 48 200
use MUX2X1  MUX2X1_30
timestamp 1515870181
transform -1 0 936 0 1 3410
box 0 0 96 200
use OAI21X1  OAI21X1_312
timestamp 1515870181
transform -1 0 1000 0 1 3410
box 0 0 64 200
use INVX1  INVX1_28
timestamp 1515870181
transform -1 0 1032 0 1 3410
box 0 0 32 200
use MUX2X1  MUX2X1_34
timestamp 1515870181
transform -1 0 1128 0 1 3410
box 0 0 96 200
use FILL  FILL_17_0_0
timestamp 1515870181
transform -1 0 1144 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_1
timestamp 1515870181
transform -1 0 1160 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_204
timestamp 1515870181
transform -1 0 1352 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_189
timestamp 1515870181
transform 1 0 1352 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_204
timestamp 1515870181
transform -1 0 1464 0 1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_35
timestamp 1515870181
transform 1 0 1464 0 1 3410
box 0 0 96 200
use NAND2X1  NAND2X1_172
timestamp 1515870181
transform 1 0 1560 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_188
timestamp 1515870181
transform -1 0 1672 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_188
timestamp 1515870181
transform -1 0 1864 0 1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_116
timestamp 1515870181
transform 1 0 1864 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_4
timestamp 1515870181
transform 1 0 2056 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_6
timestamp 1515870181
transform -1 0 2168 0 1 3410
box 0 0 48 200
use FILL  FILL_17_1_0
timestamp 1515870181
transform -1 0 2184 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_1
timestamp 1515870181
transform -1 0 2200 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_295
timestamp 1515870181
transform -1 0 2264 0 1 3410
box 0 0 64 200
use INVX1  INVX1_27
timestamp 1515870181
transform 1 0 2264 0 1 3410
box 0 0 32 200
use NAND2X1  NAND2X1_294
timestamp 1515870181
transform -1 0 2344 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_309
timestamp 1515870181
transform 1 0 2344 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_119
timestamp 1515870181
transform 1 0 2408 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_7
timestamp 1515870181
transform -1 0 2664 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_23
timestamp 1515870181
transform 1 0 2664 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_23
timestamp 1515870181
transform 1 0 2728 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_314
timestamp 1515870181
transform -1 0 2968 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_335
timestamp 1515870181
transform 1 0 2968 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_143
timestamp 1515870181
transform -1 0 3224 0 1 3410
box 0 0 192 200
use FILL  FILL_17_2_0
timestamp 1515870181
transform 1 0 3224 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_1
timestamp 1515870181
transform 1 0 3240 0 1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_143
timestamp 1515870181
transform 1 0 3256 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_264
timestamp 1515870181
transform -1 0 3368 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_266
timestamp 1515870181
transform 1 0 3368 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_135
timestamp 1515870181
transform 1 0 3416 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_116
timestamp 1515870181
transform -1 0 3528 0 1 3410
box 0 0 48 200
use INVX1  INVX1_40
timestamp 1515870181
transform 1 0 3528 0 1 3410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_135
timestamp 1515870181
transform 1 0 3560 0 1 3410
box 0 0 192 200
use NAND3X1  NAND3X1_200
timestamp 1515870181
transform 1 0 3752 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_40
timestamp 1515870181
transform 1 0 3816 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_150
timestamp 1515870181
transform 1 0 3880 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_310
timestamp 1515870181
transform 1 0 3944 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_229
timestamp 1515870181
transform -1 0 4072 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_69
timestamp 1515870181
transform 1 0 4072 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_230
timestamp 1515870181
transform 1 0 4136 0 1 3410
box 0 0 64 200
use FILL  FILL_17_3_0
timestamp 1515870181
transform 1 0 4200 0 1 3410
box 0 0 16 200
use FILL  FILL_17_3_1
timestamp 1515870181
transform 1 0 4216 0 1 3410
box 0 0 16 200
use NAND3X1  NAND3X1_70
timestamp 1515870181
transform 1 0 4232 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_148
timestamp 1515870181
transform -1 0 4360 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_308
timestamp 1515870181
transform 1 0 4360 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_100
timestamp 1515870181
transform 1 0 4424 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_260
timestamp 1515870181
transform 1 0 4488 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_264
timestamp 1515870181
transform 1 0 4552 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_121
timestamp 1515870181
transform 1 0 4616 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_281
timestamp 1515870181
transform 1 0 4680 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_157
timestamp 1515870181
transform 1 0 4744 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_465
timestamp 1515870181
transform 1 0 4792 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_278
timestamp 1515870181
transform 1 0 4856 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_238
timestamp 1515870181
transform 1 0 4920 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_78
timestamp 1515870181
transform 1 0 4984 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_151
timestamp 1515870181
transform -1 0 5112 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_307
timestamp 1515870181
transform -1 0 5176 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_296
timestamp 1515870181
transform 1 0 5176 0 1 3410
box 0 0 64 200
use FILL  FILL_17_4_0
timestamp 1515870181
transform -1 0 5256 0 1 3410
box 0 0 16 200
use FILL  FILL_17_4_1
timestamp 1515870181
transform -1 0 5272 0 1 3410
box 0 0 16 200
use INVX1  INVX1_5
timestamp 1515870181
transform -1 0 5304 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_76
timestamp 1515870181
transform -1 0 5352 0 1 3410
box 0 0 48 200
use INVX1  INVX1_6
timestamp 1515870181
transform 1 0 5352 0 1 3410
box 0 0 32 200
use NOR2X1  NOR2X1_77
timestamp 1515870181
transform -1 0 5432 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_327
timestamp 1515870181
transform 1 0 5432 0 1 3410
box 0 0 192 200
use NAND3X1  NAND3X1_226
timestamp 1515870181
transform 1 0 5624 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_227
timestamp 1515870181
transform 1 0 5688 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_225
timestamp 1515870181
transform 1 0 5752 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_92
timestamp 1515870181
transform -1 0 5880 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_252
timestamp 1515870181
transform 1 0 5880 0 1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_282
timestamp 1515870181
transform -1 0 6136 0 1 3410
box 0 0 192 200
use BUFX4  BUFX4_113
timestamp 1515870181
transform -1 0 6200 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_149
timestamp 1515870181
transform 1 0 6200 0 1 3410
box 0 0 64 200
use FILL  FILL_17_5_0
timestamp 1515870181
transform -1 0 6280 0 1 3410
box 0 0 16 200
use FILL  FILL_17_5_1
timestamp 1515870181
transform -1 0 6296 0 1 3410
box 0 0 16 200
use NAND3X1  NAND3X1_273
timestamp 1515870181
transform -1 0 6360 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_463
timestamp 1515870181
transform -1 0 6424 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_251
timestamp 1515870181
transform -1 0 6488 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_374
timestamp 1515870181
transform 1 0 6488 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_113
timestamp 1515870181
transform 1 0 6552 0 1 3410
box 0 0 64 200
use NOR3X1  NOR3X1_23
timestamp 1515870181
transform 1 0 6616 0 1 3410
box 0 0 128 200
use NAND2X1  NAND2X1_263
timestamp 1515870181
transform 1 0 6744 0 1 3410
box 0 0 48 200
use BUFX4  BUFX4_148
timestamp 1515870181
transform 1 0 6792 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_114
timestamp 1515870181
transform -1 0 6920 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_117
timestamp 1515870181
transform 1 0 6920 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_116
timestamp 1515870181
transform -1 0 7048 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_115
timestamp 1515870181
transform -1 0 7112 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_78
timestamp 1515870181
transform -1 0 7160 0 1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_332
timestamp 1515870181
transform 1 0 7160 0 1 3410
box 0 0 192 200
use BUFX4  BUFX4_289
timestamp 1515870181
transform 1 0 7352 0 1 3410
box 0 0 64 200
use FILL  FILL_18_1
timestamp 1515870181
transform 1 0 7416 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_40
timestamp 1515870181
transform 1 0 8 0 -1 3410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_44
timestamp 1515870181
transform -1 0 392 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_236
timestamp 1515870181
transform 1 0 392 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_223
timestamp 1515870181
transform -1 0 504 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_39
timestamp 1515870181
transform 1 0 504 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_94
timestamp 1515870181
transform -1 0 760 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_402
timestamp 1515870181
transform 1 0 760 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_296
timestamp 1515870181
transform -1 0 872 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_76
timestamp 1515870181
transform 1 0 872 0 -1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_66
timestamp 1515870181
transform 1 0 1064 0 -1 3410
box 0 0 48 200
use FILL  FILL_16_0_0
timestamp 1515870181
transform -1 0 1128 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_1
timestamp 1515870181
transform -1 0 1144 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_60
timestamp 1515870181
transform -1 0 1208 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_278
timestamp 1515870181
transform -1 0 1272 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_79
timestamp 1515870181
transform -1 0 1336 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_78
timestamp 1515870181
transform -1 0 1400 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_180
timestamp 1515870181
transform 1 0 1400 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_151
timestamp 1515870181
transform 1 0 1464 0 -1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_133
timestamp 1515870181
transform 1 0 1656 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_151
timestamp 1515870181
transform -1 0 1768 0 -1 3410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_148
timestamp 1515870181
transform 1 0 1768 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_148
timestamp 1515870181
transform -1 0 2024 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_130
timestamp 1515870181
transform -1 0 2072 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_98
timestamp 1515870181
transform 1 0 2072 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_42
timestamp 1515870181
transform 1 0 2136 0 -1 3410
box 0 0 32 200
use FILL  FILL_16_1_0
timestamp 1515870181
transform -1 0 2184 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_1
timestamp 1515870181
transform -1 0 2200 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_281
timestamp 1515870181
transform -1 0 2264 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_204
timestamp 1515870181
transform 1 0 2264 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_6
timestamp 1515870181
transform 1 0 2328 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_2
timestamp 1515870181
transform 1 0 2392 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_336
timestamp 1515870181
transform 1 0 2456 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_315
timestamp 1515870181
transform 1 0 2520 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_9
timestamp 1515870181
transform 1 0 2568 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_75
timestamp 1515870181
transform 1 0 2616 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_300
timestamp 1515870181
transform 1 0 2680 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_26
timestamp 1515870181
transform -1 0 2776 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_46
timestamp 1515870181
transform 1 0 2776 0 -1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_405
timestamp 1515870181
transform -1 0 2872 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_80
timestamp 1515870181
transform -1 0 2904 0 -1 3410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_159
timestamp 1515870181
transform 1 0 2904 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_408
timestamp 1515870181
transform -1 0 3160 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_82
timestamp 1515870181
transform -1 0 3192 0 -1 3410
box 0 0 32 200
use FILL  FILL_16_2_0
timestamp 1515870181
transform 1 0 3192 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_1
timestamp 1515870181
transform 1 0 3208 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_141
timestamp 1515870181
transform 1 0 3224 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_159
timestamp 1515870181
transform -1 0 3336 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_124
timestamp 1515870181
transform 1 0 3336 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_317
timestamp 1515870181
transform 1 0 3384 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_265
timestamp 1515870181
transform -1 0 3496 0 -1 3410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_92
timestamp 1515870181
transform 1 0 3496 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_493
timestamp 1515870181
transform 1 0 3688 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_432
timestamp 1515870181
transform -1 0 3800 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_397
timestamp 1515870181
transform -1 0 3848 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_302
timestamp 1515870181
transform -1 0 3896 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_49
timestamp 1515870181
transform 1 0 3896 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_209
timestamp 1515870181
transform 1 0 3960 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_348
timestamp 1515870181
transform -1 0 4072 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_378
timestamp 1515870181
transform 1 0 4072 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_40
timestamp 1515870181
transform 1 0 4136 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_3_0
timestamp 1515870181
transform -1 0 4216 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_3_1
timestamp 1515870181
transform -1 0 4232 0 -1 3410
box 0 0 16 200
use INVX1  INVX1_7
timestamp 1515870181
transform -1 0 4264 0 -1 3410
box 0 0 32 200
use BUFX4  BUFX4_134
timestamp 1515870181
transform -1 0 4328 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_351
timestamp 1515870181
transform 1 0 4328 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_132
timestamp 1515870181
transform 1 0 4376 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_411
timestamp 1515870181
transform 1 0 4440 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_19
timestamp 1515870181
transform -1 0 4552 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_133
timestamp 1515870181
transform -1 0 4616 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_403
timestamp 1515870181
transform -1 0 4664 0 -1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_115
timestamp 1515870181
transform 1 0 4664 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_379
timestamp 1515870181
transform 1 0 4712 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_323
timestamp 1515870181
transform 1 0 4776 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_118
timestamp 1515870181
transform 1 0 4824 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_269
timestamp 1515870181
transform -1 0 4936 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_39
timestamp 1515870181
transform 1 0 4936 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_181
timestamp 1515870181
transform 1 0 5000 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_81
timestamp 1515870181
transform -1 0 5112 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_4
timestamp 1515870181
transform -1 0 5176 0 -1 3410
box 0 0 64 200
use INVX8  INVX8_17
timestamp 1515870181
transform 1 0 5176 0 -1 3410
box 0 0 80 200
use FILL  FILL_16_4_0
timestamp 1515870181
transform -1 0 5272 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_4_1
timestamp 1515870181
transform -1 0 5288 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_261
timestamp 1515870181
transform -1 0 5336 0 -1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_75
timestamp 1515870181
transform 1 0 5336 0 -1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_260
timestamp 1515870181
transform 1 0 5384 0 -1 3410
box 0 0 48 200
use AOI21X1  AOI21X1_7
timestamp 1515870181
transform 1 0 5432 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_16
timestamp 1515870181
transform -1 0 5544 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_67
timestamp 1515870181
transform -1 0 5608 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_66
timestamp 1515870181
transform 1 0 5608 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_65
timestamp 1515870181
transform -1 0 5736 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_97
timestamp 1515870181
transform -1 0 5800 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_257
timestamp 1515870181
transform -1 0 5864 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_95
timestamp 1515870181
transform -1 0 5928 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_255
timestamp 1515870181
transform 1 0 5928 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_51
timestamp 1515870181
transform 1 0 5992 0 -1 3410
box 0 0 48 200
use AOI21X1  AOI21X1_42
timestamp 1515870181
transform -1 0 6104 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_214
timestamp 1515870181
transform -1 0 6168 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_185
timestamp 1515870181
transform 1 0 6168 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_5_0
timestamp 1515870181
transform -1 0 6248 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_5_1
timestamp 1515870181
transform -1 0 6264 0 -1 3410
box 0 0 16 200
use NOR3X1  NOR3X1_44
timestamp 1515870181
transform -1 0 6392 0 -1 3410
box 0 0 128 200
use OAI21X1  OAI21X1_462
timestamp 1515870181
transform 1 0 6392 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_272
timestamp 1515870181
transform -1 0 6520 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_112
timestamp 1515870181
transform -1 0 6584 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_373
timestamp 1515870181
transform -1 0 6648 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_7
timestamp 1515870181
transform -1 0 6712 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_74
timestamp 1515870181
transform 1 0 6712 0 -1 3410
box 0 0 48 200
use INVX1  INVX1_4
timestamp 1515870181
transform -1 0 6792 0 -1 3410
box 0 0 32 200
use BUFX4  BUFX4_313
timestamp 1515870181
transform 1 0 6792 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_230
timestamp 1515870181
transform 1 0 6856 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_274
timestamp 1515870181
transform -1 0 6984 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_302
timestamp 1515870181
transform 1 0 6984 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_277
timestamp 1515870181
transform 1 0 7048 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_275
timestamp 1515870181
transform -1 0 7176 0 -1 3410
box 0 0 64 200
use AOI21X1  AOI21X1_12
timestamp 1515870181
transform 1 0 7176 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_21
timestamp 1515870181
transform -1 0 7288 0 -1 3410
box 0 0 48 200
use BUFX4  BUFX4_231
timestamp 1515870181
transform -1 0 7352 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_234
timestamp 1515870181
transform 1 0 7352 0 -1 3410
box 0 0 64 200
use FILL  FILL_17_1
timestamp 1515870181
transform -1 0 7432 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_96
timestamp 1515870181
transform 1 0 8 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_95
timestamp 1515870181
transform 1 0 72 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_44
timestamp 1515870181
transform -1 0 200 0 1 3010
box 0 0 64 200
use INVX1  INVX1_78
timestamp 1515870181
transform 1 0 200 0 1 3010
box 0 0 32 200
use BUFX4  BUFX4_45
timestamp 1515870181
transform 1 0 232 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_37
timestamp 1515870181
transform 1 0 296 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_90
timestamp 1515870181
transform 1 0 488 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_89
timestamp 1515870181
transform -1 0 616 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_93
timestamp 1515870181
transform 1 0 616 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_218
timestamp 1515870181
transform 1 0 680 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_204
timestamp 1515870181
transform -1 0 792 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_218
timestamp 1515870181
transform 1 0 792 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_229
timestamp 1515870181
transform 1 0 984 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_216
timestamp 1515870181
transform -1 0 1096 0 1 3010
box 0 0 48 200
use FILL  FILL_15_0_0
timestamp 1515870181
transform -1 0 1112 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_1
timestamp 1515870181
transform -1 0 1128 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_229
timestamp 1515870181
transform -1 0 1320 0 1 3010
box 0 0 192 200
use BUFX4  BUFX4_64
timestamp 1515870181
transform -1 0 1384 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1515870181
transform 1 0 1384 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_49
timestamp 1515870181
transform 1 0 1576 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_44
timestamp 1515870181
transform -1 0 1688 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_156
timestamp 1515870181
transform 1 0 1688 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_156
timestamp 1515870181
transform 1 0 1752 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_138
timestamp 1515870181
transform -1 0 1992 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_363
timestamp 1515870181
transform 1 0 1992 0 1 3010
box 0 0 64 200
use INVX1  INVX1_67
timestamp 1515870181
transform 1 0 2056 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_381
timestamp 1515870181
transform 1 0 2088 0 1 3010
box 0 0 64 200
use FILL  FILL_15_1_0
timestamp 1515870181
transform -1 0 2168 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_1
timestamp 1515870181
transform -1 0 2184 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_7
timestamp 1515870181
transform -1 0 2232 0 1 3010
box 0 0 48 200
use BUFX4  BUFX4_84
timestamp 1515870181
transform -1 0 2296 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_118
timestamp 1515870181
transform 1 0 2296 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_8
timestamp 1515870181
transform -1 0 2536 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_21
timestamp 1515870181
transform 1 0 2536 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_24
timestamp 1515870181
transform -1 0 2792 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_24
timestamp 1515870181
transform 1 0 2792 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_21
timestamp 1515870181
transform -1 0 2904 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_308
timestamp 1515870181
transform -1 0 2952 0 1 3010
box 0 0 48 200
use BUFX4  BUFX4_106
timestamp 1515870181
transform 1 0 2952 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_344
timestamp 1515870181
transform 1 0 3016 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_149
timestamp 1515870181
transform 1 0 3080 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_131
timestamp 1515870181
transform 1 0 3144 0 1 3010
box 0 0 48 200
use FILL  FILL_15_2_0
timestamp 1515870181
transform 1 0 3192 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_1
timestamp 1515870181
transform 1 0 3208 0 1 3010
box 0 0 16 200
use INVX1  INVX1_32
timestamp 1515870181
transform 1 0 3224 0 1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_301
timestamp 1515870181
transform -1 0 3304 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_318
timestamp 1515870181
transform 1 0 3304 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_22
timestamp 1515870181
transform 1 0 3368 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_25
timestamp 1515870181
transform -1 0 3480 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_22
timestamp 1515870181
transform 1 0 3480 0 1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_307
timestamp 1515870181
transform -1 0 3720 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_210
timestamp 1515870181
transform -1 0 3784 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_50
timestamp 1515870181
transform 1 0 3784 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_202
timestamp 1515870181
transform 1 0 3848 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_140
timestamp 1515870181
transform 1 0 3912 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_121
timestamp 1515870181
transform -1 0 4024 0 1 3010
box 0 0 48 200
use INVX1  INVX1_65
timestamp 1515870181
transform 1 0 4024 0 1 3010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_140
timestamp 1515870181
transform -1 0 4248 0 1 3010
box 0 0 192 200
use FILL  FILL_15_3_0
timestamp 1515870181
transform 1 0 4248 0 1 3010
box 0 0 16 200
use FILL  FILL_15_3_1
timestamp 1515870181
transform 1 0 4264 0 1 3010
box 0 0 16 200
use NAND3X1  NAND3X1_119
timestamp 1515870181
transform 1 0 4280 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_120
timestamp 1515870181
transform -1 0 4408 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_279
timestamp 1515870181
transform 1 0 4408 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_280
timestamp 1515870181
transform 1 0 4472 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_315
timestamp 1515870181
transform -1 0 4600 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_240
timestamp 1515870181
transform 1 0 4600 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_239
timestamp 1515870181
transform 1 0 4664 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_79
timestamp 1515870181
transform 1 0 4728 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_80
timestamp 1515870181
transform 1 0 4792 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_97
timestamp 1515870181
transform 1 0 4856 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_325
timestamp 1515870181
transform 1 0 4904 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_58
timestamp 1515870181
transform 1 0 4968 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_257
timestamp 1515870181
transform -1 0 5096 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_154
timestamp 1515870181
transform -1 0 5160 0 1 3010
box 0 0 64 200
use FILL  FILL_15_4_0
timestamp 1515870181
transform 1 0 5160 0 1 3010
box 0 0 16 200
use FILL  FILL_15_4_1
timestamp 1515870181
transform 1 0 5176 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_330
timestamp 1515870181
transform 1 0 5192 0 1 3010
box 0 0 192 200
use AOI21X1  AOI21X1_10
timestamp 1515870181
transform 1 0 5384 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_19
timestamp 1515870181
transform -1 0 5496 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_96
timestamp 1515870181
transform -1 0 5560 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_64
timestamp 1515870181
transform -1 0 5624 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_256
timestamp 1515870181
transform 1 0 5624 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_224
timestamp 1515870181
transform 1 0 5688 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_94
timestamp 1515870181
transform -1 0 5816 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_254
timestamp 1515870181
transform -1 0 5880 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_23
timestamp 1515870181
transform 1 0 5880 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_32
timestamp 1515870181
transform -1 0 5992 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_247
timestamp 1515870181
transform -1 0 6184 0 1 3010
box 0 0 192 200
use NOR2X1  NOR2X1_35
timestamp 1515870181
transform -1 0 6232 0 1 3010
box 0 0 48 200
use FILL  FILL_15_5_0
timestamp 1515870181
transform 1 0 6232 0 1 3010
box 0 0 16 200
use FILL  FILL_15_5_1
timestamp 1515870181
transform 1 0 6248 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_108
timestamp 1515870181
transform 1 0 6264 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_26
timestamp 1515870181
transform -1 0 6392 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_250
timestamp 1515870181
transform 1 0 6392 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_300
timestamp 1515870181
transform -1 0 6648 0 1 3010
box 0 0 192 200
use BUFX4  BUFX4_254
timestamp 1515870181
transform 1 0 6648 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_119
timestamp 1515870181
transform -1 0 6776 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_28
timestamp 1515870181
transform 1 0 6776 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_37
timestamp 1515870181
transform -1 0 6888 0 1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_252
timestamp 1515870181
transform 1 0 6888 0 1 3010
box 0 0 192 200
use NAND3X1  NAND3X1_276
timestamp 1515870181
transform 1 0 7080 0 1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_256
timestamp 1515870181
transform 1 0 7144 0 1 3010
box 0 0 192 200
use AOI21X1  AOI21X1_32
timestamp 1515870181
transform -1 0 7400 0 1 3010
box 0 0 64 200
use FILL  FILL_16_1
timestamp 1515870181
transform 1 0 7400 0 1 3010
box 0 0 16 200
use FILL  FILL_16_2
timestamp 1515870181
transform 1 0 7416 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_237
timestamp 1515870181
transform -1 0 72 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_130
timestamp 1515870181
transform -1 0 136 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_42
timestamp 1515870181
transform -1 0 200 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_234
timestamp 1515870181
transform 1 0 200 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_221
timestamp 1515870181
transform -1 0 312 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_234
timestamp 1515870181
transform 1 0 312 0 -1 3010
box 0 0 192 200
use INVX1  INVX1_53
timestamp 1515870181
transform 1 0 504 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_357
timestamp 1515870181
transform 1 0 536 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_129
timestamp 1515870181
transform 1 0 600 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_109
timestamp 1515870181
transform 1 0 664 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_110
timestamp 1515870181
transform -1 0 792 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_366
timestamp 1515870181
transform -1 0 840 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_47
timestamp 1515870181
transform -1 0 1032 0 -1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_12
timestamp 1515870181
transform 1 0 1032 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_10
timestamp 1515870181
transform -1 0 1144 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_0_0
timestamp 1515870181
transform 1 0 1144 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_1
timestamp 1515870181
transform 1 0 1160 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_122
timestamp 1515870181
transform 1 0 1176 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_15
timestamp 1515870181
transform 1 0 1368 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_17
timestamp 1515870181
transform -1 0 1480 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_336
timestamp 1515870181
transform -1 0 1528 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_173
timestamp 1515870181
transform 1 0 1528 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_12
timestamp 1515870181
transform 1 0 1592 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_14
timestamp 1515870181
transform -1 0 1704 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_124
timestamp 1515870181
transform 1 0 1704 0 -1 3010
box 0 0 192 200
use BUFX4  BUFX4_11
timestamp 1515870181
transform -1 0 1960 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_350
timestamp 1515870181
transform -1 0 2008 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_46
timestamp 1515870181
transform -1 0 2072 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_5
timestamp 1515870181
transform 1 0 2072 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_1_0
timestamp 1515870181
transform 1 0 2136 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_1
timestamp 1515870181
transform 1 0 2152 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_117
timestamp 1515870181
transform 1 0 2168 0 -1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_371
timestamp 1515870181
transform -1 0 2408 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_164
timestamp 1515870181
transform -1 0 2472 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_47
timestamp 1515870181
transform -1 0 2536 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_24
timestamp 1515870181
transform 1 0 2536 0 -1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_27
timestamp 1515870181
transform -1 0 2776 0 -1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_369
timestamp 1515870181
transform -1 0 2824 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_166
timestamp 1515870181
transform 1 0 2824 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_321
timestamp 1515870181
transform -1 0 2936 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_10
timestamp 1515870181
transform 1 0 2936 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_149
timestamp 1515870181
transform 1 0 3000 0 -1 3010
box 0 0 192 200
use FILL  FILL_14_2_0
timestamp 1515870181
transform -1 0 3208 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_1
timestamp 1515870181
transform -1 0 3224 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_132
timestamp 1515870181
transform -1 0 3272 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_150
timestamp 1515870181
transform -1 0 3336 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_150
timestamp 1515870181
transform 1 0 3336 0 -1 3010
box 0 0 192 200
use BUFX4  BUFX4_239
timestamp 1515870181
transform -1 0 3592 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_37
timestamp 1515870181
transform 1 0 3592 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_327
timestamp 1515870181
transform 1 0 3624 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_326
timestamp 1515870181
transform -1 0 3752 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_242
timestamp 1515870181
transform 1 0 3752 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_285
timestamp 1515870181
transform -1 0 3880 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_487
timestamp 1515870181
transform 1 0 3880 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_426
timestamp 1515870181
transform -1 0 3992 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_86
timestamp 1515870181
transform 1 0 3992 0 -1 3010
box 0 0 192 200
use FILL  FILL_14_3_0
timestamp 1515870181
transform 1 0 4184 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_3_1
timestamp 1515870181
transform 1 0 4200 0 -1 3010
box 0 0 16 200
use OAI21X1  OAI21X1_134
timestamp 1515870181
transform 1 0 4216 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_115
timestamp 1515870181
transform -1 0 4328 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_134
timestamp 1515870181
transform 1 0 4328 0 -1 3010
box 0 0 192 200
use NAND2X1  NAND2X1_306
timestamp 1515870181
transform -1 0 4568 0 -1 3010
box 0 0 48 200
use INVX1  INVX1_35
timestamp 1515870181
transform 1 0 4568 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_324
timestamp 1515870181
transform 1 0 4600 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_59
timestamp 1515870181
transform -1 0 4728 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_309
timestamp 1515870181
transform 1 0 4728 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_60
timestamp 1515870181
transform 1 0 4776 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_219
timestamp 1515870181
transform -1 0 4904 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_220
timestamp 1515870181
transform -1 0 4968 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_399
timestamp 1515870181
transform 1 0 4968 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_145
timestamp 1515870181
transform 1 0 5016 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_441
timestamp 1515870181
transform 1 0 5064 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_218
timestamp 1515870181
transform 1 0 5128 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_4_0
timestamp 1515870181
transform 1 0 5192 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_4_1
timestamp 1515870181
transform 1 0 5208 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_323
timestamp 1515870181
transform 1 0 5224 0 -1 3010
box 0 0 192 200
use NAND3X1  NAND3X1_23
timestamp 1515870181
transform 1 0 5416 0 -1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1515870181
transform 1 0 5480 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_12
timestamp 1515870181
transform -1 0 5592 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_221
timestamp 1515870181
transform -1 0 5656 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_26
timestamp 1515870181
transform -1 0 5720 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_186
timestamp 1515870181
transform 1 0 5720 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_24
timestamp 1515870181
transform 1 0 5784 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_182
timestamp 1515870181
transform -1 0 5912 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_22
timestamp 1515870181
transform 1 0 5912 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_301
timestamp 1515870181
transform -1 0 6040 0 -1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_35
timestamp 1515870181
transform 1 0 6040 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_44
timestamp 1515870181
transform 1 0 6104 0 -1 3010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_275
timestamp 1515870181
transform -1 0 6344 0 -1 3010
box 0 0 192 200
use FILL  FILL_14_5_0
timestamp 1515870181
transform -1 0 6360 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_5_1
timestamp 1515870181
transform -1 0 6376 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_250
timestamp 1515870181
transform -1 0 6568 0 -1 3010
box 0 0 192 200
use AOI21X1  AOI21X1_60
timestamp 1515870181
transform 1 0 6568 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_69
timestamp 1515870181
transform 1 0 6632 0 -1 3010
box 0 0 48 200
use BUFX4  BUFX4_22
timestamp 1515870181
transform 1 0 6680 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_263
timestamp 1515870181
transform 1 0 6744 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_53
timestamp 1515870181
transform 1 0 6808 0 -1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_44
timestamp 1515870181
transform -1 0 6920 0 -1 3010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_284
timestamp 1515870181
transform 1 0 6920 0 -1 3010
box 0 0 192 200
use NAND3X1  NAND3X1_317
timestamp 1515870181
transform 1 0 7112 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_316
timestamp 1515870181
transform -1 0 7240 0 -1 3010
box 0 0 64 200
use BUFX4  BUFX4_229
timestamp 1515870181
transform -1 0 7304 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_25
timestamp 1515870181
transform 1 0 7304 0 -1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_16
timestamp 1515870181
transform -1 0 7416 0 -1 3010
box 0 0 64 200
use FILL  FILL_15_1
timestamp 1515870181
transform -1 0 7432 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_239
timestamp 1515870181
transform -1 0 200 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_226
timestamp 1515870181
transform 1 0 200 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_239
timestamp 1515870181
transform -1 0 312 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_238
timestamp 1515870181
transform 1 0 312 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_211
timestamp 1515870181
transform 1 0 376 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_89
timestamp 1515870181
transform -1 0 472 0 1 2610
box 0 0 48 200
use INVX4  INVX4_1
timestamp 1515870181
transform -1 0 520 0 1 2610
box 0 0 48 200
use INVX1  INVX1_3
timestamp 1515870181
transform -1 0 552 0 1 2610
box 0 0 32 200
use AND2X2  AND2X2_6
timestamp 1515870181
transform 1 0 552 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_1
timestamp 1515870181
transform -1 0 680 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_5
timestamp 1515870181
transform -1 0 728 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_194
timestamp 1515870181
transform -1 0 776 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_72
timestamp 1515870181
transform -1 0 824 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_5
timestamp 1515870181
transform 1 0 824 0 1 2610
box 0 0 64 200
use INVX2  INVX2_1
timestamp 1515870181
transform 1 0 888 0 1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_177
timestamp 1515870181
transform 1 0 920 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_4
timestamp 1515870181
transform -1 0 1016 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_3
timestamp 1515870181
transform -1 0 1064 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_7
timestamp 1515870181
transform 1 0 1064 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_54
timestamp 1515870181
transform 1 0 1112 0 1 2610
box 0 0 48 200
use FILL  FILL_13_0_0
timestamp 1515870181
transform 1 0 1160 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_1
timestamp 1515870181
transform 1 0 1176 0 1 2610
box 0 0 16 200
use AND2X2  AND2X2_4
timestamp 1515870181
transform 1 0 1192 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_127
timestamp 1515870181
transform 1 0 1256 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_160
timestamp 1515870181
transform 1 0 1448 0 1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_154
timestamp 1515870181
transform 1 0 1496 0 1 2610
box 0 0 192 200
use BUFX4  BUFX4_196
timestamp 1515870181
transform -1 0 1752 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_154
timestamp 1515870181
transform 1 0 1752 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_136
timestamp 1515870181
transform -1 0 1864 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_37
timestamp 1515870181
transform 1 0 1864 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_3
timestamp 1515870181
transform 1 0 1912 0 1 2610
box 0 0 64 200
use INVX1  INVX1_57
timestamp 1515870181
transform 1 0 1976 0 1 2610
box 0 0 32 200
use AND2X2  AND2X2_2
timestamp 1515870181
transform 1 0 2008 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_92
timestamp 1515870181
transform 1 0 2072 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_9
timestamp 1515870181
transform 1 0 2120 0 1 2610
box 0 0 64 200
use FILL  FILL_13_1_0
timestamp 1515870181
transform -1 0 2200 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_1
timestamp 1515870181
transform -1 0 2216 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_165
timestamp 1515870181
transform -1 0 2280 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_28
timestamp 1515870181
transform 1 0 2280 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_31
timestamp 1515870181
transform 1 0 2472 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_28
timestamp 1515870181
transform -1 0 2584 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_139
timestamp 1515870181
transform 1 0 2584 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_172
timestamp 1515870181
transform -1 0 2840 0 1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_172
timestamp 1515870181
transform 1 0 2840 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_155
timestamp 1515870181
transform 1 0 2904 0 1 2610
box 0 0 48 200
use INVX1  INVX1_66
timestamp 1515870181
transform 1 0 2952 0 1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_349
timestamp 1515870181
transform -1 0 3032 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_380
timestamp 1515870181
transform 1 0 3032 0 1 2610
box 0 0 64 200
use FILL  FILL_13_2_0
timestamp 1515870181
transform 1 0 3096 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_1
timestamp 1515870181
transform 1 0 3112 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_120
timestamp 1515870181
transform 1 0 3128 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_10
timestamp 1515870181
transform 1 0 3320 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_8
timestamp 1515870181
transform -1 0 3432 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_322
timestamp 1515870181
transform -1 0 3480 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_345
timestamp 1515870181
transform 1 0 3480 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_188
timestamp 1515870181
transform 1 0 3544 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_166
timestamp 1515870181
transform 1 0 3608 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_149
timestamp 1515870181
transform -1 0 3720 0 1 2610
box 0 0 48 200
use INVX1  INVX1_36
timestamp 1515870181
transform 1 0 3720 0 1 2610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_166
timestamp 1515870181
transform -1 0 3944 0 1 2610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_131
timestamp 1515870181
transform 1 0 3944 0 1 2610
box 0 0 192 200
use INVX1  INVX1_20
timestamp 1515870181
transform 1 0 4136 0 1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_297
timestamp 1515870181
transform 1 0 4168 0 1 2610
box 0 0 64 200
use FILL  FILL_13_3_0
timestamp 1515870181
transform 1 0 4232 0 1 2610
box 0 0 16 200
use FILL  FILL_13_3_1
timestamp 1515870181
transform 1 0 4248 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_127
timestamp 1515870181
transform 1 0 4264 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_31
timestamp 1515870181
transform 1 0 4328 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_88
timestamp 1515870181
transform 1 0 4392 0 1 2610
box 0 0 48 200
use BUFX4  BUFX4_102
timestamp 1515870181
transform -1 0 4504 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_298
timestamp 1515870181
transform 1 0 4504 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_28
timestamp 1515870181
transform -1 0 4632 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_188
timestamp 1515870181
transform -1 0 4696 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_429
timestamp 1515870181
transform -1 0 4760 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_139
timestamp 1515870181
transform -1 0 4808 0 1 2610
box 0 0 48 200
use BUFX4  BUFX4_316
timestamp 1515870181
transform 1 0 4808 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_191
timestamp 1515870181
transform 1 0 4872 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_88
timestamp 1515870181
transform 1 0 4936 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_253
timestamp 1515870181
transform -1 0 5064 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_91
timestamp 1515870181
transform 1 0 5064 0 1 2610
box 0 0 64 200
use NOR3X1  NOR3X1_5
timestamp 1515870181
transform -1 0 5256 0 1 2610
box 0 0 128 200
use FILL  FILL_13_4_0
timestamp 1515870181
transform 1 0 5256 0 1 2610
box 0 0 16 200
use FILL  FILL_13_4_1
timestamp 1515870181
transform 1 0 5272 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_293
timestamp 1515870181
transform 1 0 5288 0 1 2610
box 0 0 64 200
use NOR3X1  NOR3X1_35
timestamp 1515870181
transform -1 0 5480 0 1 2610
box 0 0 128 200
use NAND3X1  NAND3X1_184
timestamp 1515870181
transform -1 0 5544 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_187
timestamp 1515870181
transform 1 0 5544 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_426
timestamp 1515870181
transform 1 0 5608 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_288
timestamp 1515870181
transform 1 0 5672 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_27
timestamp 1515870181
transform -1 0 5800 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_61
timestamp 1515870181
transform 1 0 5800 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_292
timestamp 1515870181
transform 1 0 5864 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_25
timestamp 1515870181
transform -1 0 5992 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_185
timestamp 1515870181
transform 1 0 5992 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_8
timestamp 1515870181
transform -1 0 6120 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_383
timestamp 1515870181
transform 1 0 6120 0 1 2610
box 0 0 48 200
use INVX1  INVX1_88
timestamp 1515870181
transform 1 0 6168 0 1 2610
box 0 0 32 200
use NOR2X1  NOR2X1_128
timestamp 1515870181
transform -1 0 6248 0 1 2610
box 0 0 48 200
use FILL  FILL_13_5_0
timestamp 1515870181
transform -1 0 6264 0 1 2610
box 0 0 16 200
use FILL  FILL_13_5_1
timestamp 1515870181
transform -1 0 6280 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_299
timestamp 1515870181
transform -1 0 6344 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_253
timestamp 1515870181
transform 1 0 6344 0 1 2610
box 0 0 192 200
use BUFX4  BUFX4_292
timestamp 1515870181
transform 1 0 6536 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_232
timestamp 1515870181
transform -1 0 6664 0 1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_249
timestamp 1515870181
transform 1 0 6664 0 1 2610
box 0 0 192 200
use BUFX4  BUFX4_291
timestamp 1515870181
transform -1 0 6920 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_300
timestamp 1515870181
transform 1 0 6920 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_233
timestamp 1515870181
transform 1 0 6984 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_314
timestamp 1515870181
transform -1 0 7112 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_315
timestamp 1515870181
transform 1 0 7112 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_132
timestamp 1515870181
transform 1 0 7176 0 1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_336
timestamp 1515870181
transform -1 0 7416 0 1 2610
box 0 0 192 200
use FILL  FILL_14_1
timestamp 1515870181
transform 1 0 7416 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_241
timestamp 1515870181
transform 1 0 8 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_9
timestamp 1515870181
transform -1 0 120 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_1
timestamp 1515870181
transform 1 0 120 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_90
timestamp 1515870181
transform 1 0 184 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_6
timestamp 1515870181
transform -1 0 280 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_99
timestamp 1515870181
transform 1 0 280 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_100
timestamp 1515870181
transform -1 0 408 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_42
timestamp 1515870181
transform 1 0 408 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_331
timestamp 1515870181
transform -1 0 648 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_71
timestamp 1515870181
transform 1 0 648 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_271
timestamp 1515870181
transform 1 0 696 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_54
timestamp 1515870181
transform -1 0 824 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_1
timestamp 1515870181
transform 1 0 824 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_36
timestamp 1515870181
transform 1 0 856 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_2
timestamp 1515870181
transform -1 0 936 0 -1 2610
box 0 0 32 200
use NAND2X1  NAND2X1_1
timestamp 1515870181
transform 1 0 936 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_91
timestamp 1515870181
transform 1 0 984 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_1
timestamp 1515870181
transform 1 0 1032 0 -1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_2
timestamp 1515870181
transform -1 0 1128 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_0_0
timestamp 1515870181
transform -1 0 1144 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_1
timestamp 1515870181
transform -1 0 1160 0 -1 2610
box 0 0 16 200
use NOR2X1  NOR2X1_8
timestamp 1515870181
transform -1 0 1208 0 -1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_179
timestamp 1515870181
transform 1 0 1208 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_179
timestamp 1515870181
transform 1 0 1400 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_163
timestamp 1515870181
transform -1 0 1512 0 -1 2610
box 0 0 48 200
use MUX2X1  MUX2X1_8
timestamp 1515870181
transform 1 0 1512 0 -1 2610
box 0 0 96 200
use BUFX4  BUFX4_176
timestamp 1515870181
transform 1 0 1608 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_175
timestamp 1515870181
transform 1 0 1672 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_143
timestamp 1515870181
transform 1 0 1736 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_189
timestamp 1515870181
transform 1 0 1784 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_173
timestamp 1515870181
transform -1 0 1896 0 -1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_189
timestamp 1515870181
transform -1 0 2088 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_2
timestamp 1515870181
transform 1 0 2088 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_126
timestamp 1515870181
transform -1 0 2184 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_1_0
timestamp 1515870181
transform 1 0 2184 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_1
timestamp 1515870181
transform 1 0 2200 0 -1 2610
box 0 0 16 200
use AND2X2  AND2X2_1
timestamp 1515870181
transform 1 0 2216 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_19
timestamp 1515870181
transform -1 0 2328 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_109
timestamp 1515870181
transform 1 0 2328 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_420
timestamp 1515870181
transform 1 0 2376 0 -1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_95
timestamp 1515870181
transform 1 0 2424 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_496
timestamp 1515870181
transform 1 0 2616 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_435
timestamp 1515870181
transform -1 0 2728 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_9
timestamp 1515870181
transform -1 0 2792 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_191
timestamp 1515870181
transform 1 0 2792 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_163
timestamp 1515870181
transform 1 0 2856 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_163
timestamp 1515870181
transform 1 0 3048 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_146
timestamp 1515870181
transform -1 0 3160 0 -1 2610
box 0 0 48 200
use INVX1  INVX1_21
timestamp 1515870181
transform 1 0 3160 0 -1 2610
box 0 0 32 200
use FILL  FILL_12_2_0
timestamp 1515870181
transform -1 0 3208 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_1
timestamp 1515870181
transform -1 0 3224 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_286
timestamp 1515870181
transform -1 0 3272 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_299
timestamp 1515870181
transform 1 0 3272 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_48
timestamp 1515870181
transform 1 0 3336 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_140
timestamp 1515870181
transform -1 0 3464 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_47
timestamp 1515870181
transform 1 0 3464 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_300
timestamp 1515870181
transform 1 0 3496 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_187
timestamp 1515870181
transform 1 0 3560 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_283
timestamp 1515870181
transform -1 0 3688 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_484
timestamp 1515870181
transform 1 0 3688 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_423
timestamp 1515870181
transform -1 0 3800 0 -1 2610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_83
timestamp 1515870181
transform 1 0 3800 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_131
timestamp 1515870181
transform 1 0 3992 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_112
timestamp 1515870181
transform -1 0 4104 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_241
timestamp 1515870181
transform 1 0 4104 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_285
timestamp 1515870181
transform -1 0 4216 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_3_0
timestamp 1515870181
transform 1 0 4216 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_3_1
timestamp 1515870181
transform 1 0 4232 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_34
timestamp 1515870181
transform 1 0 4248 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_29
timestamp 1515870181
transform -1 0 4376 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_288
timestamp 1515870181
transform 1 0 4376 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_30
timestamp 1515870181
transform -1 0 4488 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_190
timestamp 1515870181
transform -1 0 4552 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_393
timestamp 1515870181
transform -1 0 4600 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_189
timestamp 1515870181
transform -1 0 4664 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_17
timestamp 1515870181
transform -1 0 4728 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_349
timestamp 1515870181
transform 1 0 4728 0 -1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_105
timestamp 1515870181
transform 1 0 4920 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_125
timestamp 1515870181
transform -1 0 5032 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_243
timestamp 1515870181
transform 1 0 5032 0 -1 2610
box 0 0 192 200
use FILL  FILL_12_4_0
timestamp 1515870181
transform 1 0 5224 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_4_1
timestamp 1515870181
transform 1 0 5240 0 -1 2610
box 0 0 16 200
use AOI21X1  AOI21X1_19
timestamp 1515870181
transform 1 0 5256 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_28
timestamp 1515870181
transform 1 0 5320 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_183
timestamp 1515870181
transform -1 0 5432 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_427
timestamp 1515870181
transform -1 0 5496 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_265
timestamp 1515870181
transform -1 0 5560 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_267
timestamp 1515870181
transform -1 0 5624 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_264
timestamp 1515870181
transform -1 0 5688 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_36
timestamp 1515870181
transform -1 0 5736 0 -1 2610
box 0 0 48 200
use AOI21X1  AOI21X1_27
timestamp 1515870181
transform -1 0 5800 0 -1 2610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_251
timestamp 1515870181
transform 1 0 5800 0 -1 2610
box 0 0 192 200
use NAND3X1  NAND3X1_104
timestamp 1515870181
transform 1 0 5992 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_107
timestamp 1515870181
transform 1 0 6056 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_106
timestamp 1515870181
transform 1 0 6120 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_105
timestamp 1515870181
transform 1 0 6184 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_5_0
timestamp 1515870181
transform -1 0 6264 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_5_1
timestamp 1515870181
transform -1 0 6280 0 -1 2610
box 0 0 16 200
use NAND3X1  NAND3X1_124
timestamp 1515870181
transform -1 0 6344 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_29
timestamp 1515870181
transform 1 0 6344 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_38
timestamp 1515870181
transform -1 0 6456 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_284
timestamp 1515870181
transform 1 0 6456 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_125
timestamp 1515870181
transform -1 0 6584 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_285
timestamp 1515870181
transform 1 0 6584 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_256
timestamp 1515870181
transform 1 0 6648 0 -1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_25
timestamp 1515870181
transform 1 0 6712 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_34
timestamp 1515870181
transform -1 0 6824 0 -1 2610
box 0 0 48 200
use BUFX4  BUFX4_152
timestamp 1515870181
transform 1 0 6824 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1515870181
transform -1 0 6952 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_165
timestamp 1515870181
transform 1 0 6952 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_177
timestamp 1515870181
transform 1 0 7016 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_175
timestamp 1515870181
transform -1 0 7144 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_15
timestamp 1515870181
transform 1 0 7144 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_156
timestamp 1515870181
transform -1 0 7272 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_154
timestamp 1515870181
transform -1 0 7336 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_157
timestamp 1515870181
transform 1 0 7336 0 -1 2610
box 0 0 64 200
use FILL  FILL_13_1
timestamp 1515870181
transform -1 0 7416 0 -1 2610
box 0 0 16 200
use FILL  FILL_13_2
timestamp 1515870181
transform -1 0 7432 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_227
timestamp 1515870181
transform -1 0 200 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_214
timestamp 1515870181
transform 1 0 200 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_227
timestamp 1515870181
transform -1 0 312 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_236
timestamp 1515870181
transform 1 0 312 0 1 2210
box 0 0 64 200
use INVX1  INVX1_18
timestamp 1515870181
transform 1 0 376 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_294
timestamp 1515870181
transform 1 0 408 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_211
timestamp 1515870181
transform 1 0 472 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_197
timestamp 1515870181
transform 1 0 664 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_211
timestamp 1515870181
transform -1 0 776 0 1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_9
timestamp 1515870181
transform 1 0 776 0 1 2210
box 0 0 96 200
use NAND2X1  NAND2X1_207
timestamp 1515870181
transform 1 0 872 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_221
timestamp 1515870181
transform -1 0 984 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_283
timestamp 1515870181
transform 1 0 984 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_392
timestamp 1515870181
transform 1 0 1032 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_428
timestamp 1515870181
transform -1 0 1144 0 1 2210
box 0 0 64 200
use FILL  FILL_11_0_0
timestamp 1515870181
transform -1 0 1160 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1515870181
transform -1 0 1176 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_295
timestamp 1515870181
transform -1 0 1240 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1515870181
transform 1 0 1240 0 1 2210
box 0 0 192 200
use NOR2X1  NOR2X1_87
timestamp 1515870181
transform -1 0 1480 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_40
timestamp 1515870181
transform 1 0 1480 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_35
timestamp 1515870181
transform -1 0 1592 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_138
timestamp 1515870181
transform 1 0 1592 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_161
timestamp 1515870181
transform -1 0 1688 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_177
timestamp 1515870181
transform -1 0 1880 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_177
timestamp 1515870181
transform -1 0 1944 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_38
timestamp 1515870181
transform 1 0 1944 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_33
timestamp 1515870181
transform -1 0 2056 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_19
timestamp 1515870181
transform 1 0 2056 0 1 2210
box 0 0 192 200
use FILL  FILL_11_1_0
timestamp 1515870181
transform 1 0 2248 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1515870181
transform 1 0 2264 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_19
timestamp 1515870181
transform 1 0 2280 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_22
timestamp 1515870181
transform -1 0 2392 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_29
timestamp 1515870181
transform 1 0 2392 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_32
timestamp 1515870181
transform 1 0 2584 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_29
timestamp 1515870181
transform -1 0 2696 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_81
timestamp 1515870181
transform 1 0 2696 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_421
timestamp 1515870181
transform 1 0 2888 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_482
timestamp 1515870181
transform -1 0 3000 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_494
timestamp 1515870181
transform 1 0 3000 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_433
timestamp 1515870181
transform -1 0 3112 0 1 2210
box 0 0 48 200
use FILL  FILL_11_2_0
timestamp 1515870181
transform -1 0 3128 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1515870181
transform -1 0 3144 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_93
timestamp 1515870181
transform -1 0 3336 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_5
timestamp 1515870181
transform 1 0 3336 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_3
timestamp 1515870181
transform -1 0 3448 0 1 2210
box 0 0 64 200
use INVX1  INVX1_22
timestamp 1515870181
transform 1 0 3448 0 1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_271
timestamp 1515870181
transform -1 0 3528 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_113
timestamp 1515870181
transform 1 0 3528 0 1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_273
timestamp 1515870181
transform 1 0 3720 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_3
timestamp 1515870181
transform 1 0 3768 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_1
timestamp 1515870181
transform -1 0 3880 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_161
timestamp 1515870181
transform 1 0 3880 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_144
timestamp 1515870181
transform -1 0 3992 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_161
timestamp 1515870181
transform -1 0 4184 0 1 2210
box 0 0 192 200
use FILL  FILL_11_3_0
timestamp 1515870181
transform 1 0 4184 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_1
timestamp 1515870181
transform 1 0 4200 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_129
timestamp 1515870181
transform 1 0 4216 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_110
timestamp 1515870181
transform -1 0 4328 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_129
timestamp 1515870181
transform -1 0 4520 0 1 2210
box 0 0 192 200
use BUFX4  BUFX4_255
timestamp 1515870181
transform -1 0 4584 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_259
timestamp 1515870181
transform -1 0 4648 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_310
timestamp 1515870181
transform -1 0 4712 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_138
timestamp 1515870181
transform 1 0 4712 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_133
timestamp 1515870181
transform -1 0 4824 0 1 2210
box 0 0 48 200
use INVX8  INVX8_18
timestamp 1515870181
transform 1 0 4824 0 1 2210
box 0 0 80 200
use BUFX4  BUFX4_153
timestamp 1515870181
transform -1 0 4968 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_115
timestamp 1515870181
transform 1 0 4968 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_291
timestamp 1515870181
transform 1 0 5032 0 1 2210
box 0 0 192 200
use FILL  FILL_11_4_0
timestamp 1515870181
transform 1 0 5224 0 1 2210
box 0 0 16 200
use FILL  FILL_11_4_1
timestamp 1515870181
transform 1 0 5240 0 1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_51
timestamp 1515870181
transform 1 0 5256 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_60
timestamp 1515870181
transform 1 0 5320 0 1 2210
box 0 0 48 200
use AOI21X1  AOI21X1_11
timestamp 1515870181
transform 1 0 5368 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_20
timestamp 1515870181
transform -1 0 5480 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_282
timestamp 1515870181
transform 1 0 5480 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_266
timestamp 1515870181
transform -1 0 5608 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_54
timestamp 1515870181
transform 1 0 5608 0 1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_333
timestamp 1515870181
transform 1 0 5656 0 1 2210
box 0 0 192 200
use AOI21X1  AOI21X1_13
timestamp 1515870181
transform 1 0 5848 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_22
timestamp 1515870181
transform 1 0 5912 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_222
timestamp 1515870181
transform -1 0 6024 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_150
timestamp 1515870181
transform -1 0 6088 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_286
timestamp 1515870181
transform -1 0 6152 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_126
timestamp 1515870181
transform 1 0 6152 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_127
timestamp 1515870181
transform -1 0 6280 0 1 2210
box 0 0 64 200
use FILL  FILL_11_5_0
timestamp 1515870181
transform -1 0 6296 0 1 2210
box 0 0 16 200
use FILL  FILL_11_5_1
timestamp 1515870181
transform -1 0 6312 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_258
timestamp 1515870181
transform -1 0 6376 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_287
timestamp 1515870181
transform -1 0 6440 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_252
timestamp 1515870181
transform -1 0 6504 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_314
timestamp 1515870181
transform 1 0 6504 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_249
timestamp 1515870181
transform 1 0 6568 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_4
timestamp 1515870181
transform 1 0 6632 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_7
timestamp 1515870181
transform 1 0 6696 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_6
timestamp 1515870181
transform -1 0 6824 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_14
timestamp 1515870181
transform -1 0 6888 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_17
timestamp 1515870181
transform 1 0 6888 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_174
timestamp 1515870181
transform 1 0 6952 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_176
timestamp 1515870181
transform -1 0 7080 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_16
timestamp 1515870181
transform 1 0 7080 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_223
timestamp 1515870181
transform 1 0 7144 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_2
timestamp 1515870181
transform 1 0 7208 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_11
timestamp 1515870181
transform 1 0 7272 0 1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_41
timestamp 1515870181
transform 1 0 7320 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_220
timestamp 1515870181
transform -1 0 7432 0 1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_35
timestamp 1515870181
transform -1 0 200 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_86
timestamp 1515870181
transform 1 0 200 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_85
timestamp 1515870181
transform -1 0 328 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_131
timestamp 1515870181
transform 1 0 328 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_282
timestamp 1515870181
transform -1 0 440 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_51
timestamp 1515870181
transform 1 0 440 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_67
timestamp 1515870181
transform 1 0 632 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_75
timestamp 1515870181
transform -1 0 744 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_85
timestamp 1515870181
transform -1 0 792 0 -1 2210
box 0 0 48 200
use MUX2X1  MUX2X1_39
timestamp 1515870181
transform -1 0 888 0 -1 2210
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_221
timestamp 1515870181
transform -1 0 1080 0 -1 2210
box 0 0 192 200
use BUFX4  BUFX4_162
timestamp 1515870181
transform -1 0 1144 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_0_0
timestamp 1515870181
transform 1 0 1144 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1515870181
transform 1 0 1160 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_206
timestamp 1515870181
transform 1 0 1176 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_287
timestamp 1515870181
transform -1 0 1304 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_210
timestamp 1515870181
transform -1 0 1368 0 -1 2210
box 0 0 64 200
use NOR3X1  NOR3X1_6
timestamp 1515870181
transform -1 0 1496 0 -1 2210
box 0 0 128 200
use NOR2X1  NOR2X1_86
timestamp 1515870181
transform -1 0 1544 0 -1 2210
box 0 0 48 200
use OAI22X1  OAI22X1_3
timestamp 1515870181
transform 1 0 1544 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_205
timestamp 1515870181
transform 1 0 1624 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_268
timestamp 1515870181
transform 1 0 1688 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_2
timestamp 1515870181
transform 1 0 1752 0 -1 2210
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1515870181
transform -1 0 2040 0 -1 2210
box 0 0 192 200
use BUFX4  BUFX4_213
timestamp 1515870181
transform -1 0 2104 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_38
timestamp 1515870181
transform 1 0 2104 0 -1 2210
box 0 0 96 200
use FILL  FILL_10_1_0
timestamp 1515870181
transform 1 0 2200 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1515870181
transform 1 0 2216 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_45
timestamp 1515870181
transform 1 0 2232 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_50
timestamp 1515870181
transform -1 0 2344 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1515870181
transform -1 0 2536 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_147
timestamp 1515870181
transform -1 0 2728 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_147
timestamp 1515870181
transform -1 0 2792 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_129
timestamp 1515870181
transform 1 0 2792 0 -1 2210
box 0 0 48 200
use BUFX4  BUFX4_167
timestamp 1515870181
transform 1 0 2840 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_212
timestamp 1515870181
transform -1 0 2968 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_115
timestamp 1515870181
transform 1 0 2968 0 -1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_355
timestamp 1515870181
transform -1 0 3208 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_2_0
timestamp 1515870181
transform 1 0 3208 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1515870181
transform 1 0 3224 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_287
timestamp 1515870181
transform 1 0 3240 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_152
timestamp 1515870181
transform 1 0 3288 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_134
timestamp 1515870181
transform -1 0 3400 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_152
timestamp 1515870181
transform -1 0 3592 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_17
timestamp 1515870181
transform 1 0 3592 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_20
timestamp 1515870181
transform -1 0 3704 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_17
timestamp 1515870181
transform 1 0 3704 0 -1 2210
box 0 0 192 200
use NAND2X1  NAND2X1_272
timestamp 1515870181
transform -1 0 3944 0 -1 2210
box 0 0 48 200
use INVX1  INVX1_11
timestamp 1515870181
transform 1 0 3944 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_281
timestamp 1515870181
transform 1 0 3976 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_58
timestamp 1515870181
transform -1 0 4104 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_279
timestamp 1515870181
transform -1 0 4168 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_10
timestamp 1515870181
transform -1 0 4200 0 -1 2210
box 0 0 32 200
use FILL  FILL_10_3_0
timestamp 1515870181
transform -1 0 4216 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_3_1
timestamp 1515870181
transform -1 0 4232 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_317
timestamp 1515870181
transform -1 0 4296 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_169
timestamp 1515870181
transform -1 0 4360 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1515870181
transform -1 0 4424 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1515870181
transform -1 0 4488 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_168
timestamp 1515870181
transform -1 0 4552 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_91
timestamp 1515870181
transform -1 0 4584 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_113
timestamp 1515870181
transform 1 0 4584 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_337
timestamp 1515870181
transform 1 0 4648 0 -1 2210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_285
timestamp 1515870181
transform 1 0 4840 0 -1 2210
box 0 0 192 200
use BUFX4  BUFX4_265
timestamp 1515870181
transform 1 0 5032 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_211
timestamp 1515870181
transform 1 0 5096 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_4_0
timestamp 1515870181
transform 1 0 5160 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_4_1
timestamp 1515870181
transform 1 0 5176 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_331
timestamp 1515870181
transform 1 0 5192 0 -1 2210
box 0 0 192 200
use BUFX4  BUFX4_59
timestamp 1515870181
transform 1 0 5384 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_45
timestamp 1515870181
transform 1 0 5448 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_216
timestamp 1515870181
transform -1 0 5576 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_122
timestamp 1515870181
transform 1 0 5576 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_9
timestamp 1515870181
transform 1 0 5640 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_18
timestamp 1515870181
transform -1 0 5752 0 -1 2210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_329
timestamp 1515870181
transform 1 0 5752 0 -1 2210
box 0 0 192 200
use NAND3X1  NAND3X1_87
timestamp 1515870181
transform -1 0 6008 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_86
timestamp 1515870181
transform 1 0 6008 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_84
timestamp 1515870181
transform -1 0 6136 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_246
timestamp 1515870181
transform 1 0 6136 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_244
timestamp 1515870181
transform 1 0 6200 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_5_0
timestamp 1515870181
transform 1 0 6264 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_5_1
timestamp 1515870181
transform 1 0 6280 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_241
timestamp 1515870181
transform 1 0 6296 0 -1 2210
box 0 0 192 200
use AOI21X1  AOI21X1_17
timestamp 1515870181
transform 1 0 6488 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_26
timestamp 1515870181
transform -1 0 6600 0 -1 2210
box 0 0 48 200
use BUFX4  BUFX4_16
timestamp 1515870181
transform 1 0 6600 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_164
timestamp 1515870181
transform 1 0 6664 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_167
timestamp 1515870181
transform 1 0 6728 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_166
timestamp 1515870181
transform 1 0 6792 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_294
timestamp 1515870181
transform -1 0 6920 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_134
timestamp 1515870181
transform -1 0 6984 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_136
timestamp 1515870181
transform -1 0 7048 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_137
timestamp 1515870181
transform 1 0 7048 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_135
timestamp 1515870181
transform -1 0 7176 0 -1 2210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_321
timestamp 1515870181
transform -1 0 7368 0 -1 2210
box 0 0 192 200
use AOI21X1  AOI21X1_1
timestamp 1515870181
transform 1 0 7368 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_235
timestamp 1515870181
transform -1 0 72 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_3
timestamp 1515870181
transform -1 0 168 0 1 1810
box 0 0 96 200
use NAND2X1  NAND2X1_73
timestamp 1515870181
transform 1 0 168 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_212
timestamp 1515870181
transform 1 0 216 0 1 1810
box 0 0 48 200
use INVX1  INVX1_8
timestamp 1515870181
transform 1 0 264 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_276
timestamp 1515870181
transform 1 0 296 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_45
timestamp 1515870181
transform 1 0 360 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_77
timestamp 1515870181
transform 1 0 552 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_61
timestamp 1515870181
transform 1 0 616 0 1 1810
box 0 0 192 200
use NAND2X1  NAND2X1_387
timestamp 1515870181
transform 1 0 808 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_420
timestamp 1515870181
transform -1 0 920 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_268
timestamp 1515870181
transform 1 0 920 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_277
timestamp 1515870181
transform -1 0 1032 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_67
timestamp 1515870181
transform -1 0 1080 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_385
timestamp 1515870181
transform 1 0 1080 0 1 1810
box 0 0 64 200
use FILL  FILL_9_0_0
timestamp 1515870181
transform -1 0 1160 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1515870181
transform -1 0 1176 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_353
timestamp 1515870181
transform -1 0 1224 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_412
timestamp 1515870181
transform 1 0 1224 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_468
timestamp 1515870181
transform -1 0 1336 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_37
timestamp 1515870181
transform -1 0 1432 0 1 1810
box 0 0 96 200
use NAND2X1  NAND2X1_190
timestamp 1515870181
transform 1 0 1432 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_205
timestamp 1515870181
transform -1 0 1544 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_267
timestamp 1515870181
transform -1 0 1608 0 1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_2
timestamp 1515870181
transform -1 0 1736 0 1 1810
box 0 0 128 200
use NOR2X1  NOR2X1_80
timestamp 1515870181
transform -1 0 1784 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_79
timestamp 1515870181
transform -1 0 1832 0 1 1810
box 0 0 48 200
use OAI22X1  OAI22X1_1
timestamp 1515870181
transform 1 0 1832 0 1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_134
timestamp 1515870181
transform 1 0 1912 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_193
timestamp 1515870181
transform 1 0 1960 0 1 1810
box 0 0 192 200
use FILL  FILL_9_1_0
timestamp 1515870181
transform 1 0 2152 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1515870181
transform 1 0 2168 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_178
timestamp 1515870181
transform 1 0 2184 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_193
timestamp 1515870181
transform -1 0 2296 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_7
timestamp 1515870181
transform -1 0 2392 0 1 1810
box 0 0 96 200
use NOR2X1  NOR2X1_158
timestamp 1515870181
transform 1 0 2392 0 1 1810
box 0 0 48 200
use OAI22X1  OAI22X1_13
timestamp 1515870181
transform -1 0 2520 0 1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_117
timestamp 1515870181
transform 1 0 2520 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_116
timestamp 1515870181
transform 1 0 2568 0 1 1810
box 0 0 48 200
use NOR3X1  NOR3X1_26
timestamp 1515870181
transform 1 0 2616 0 1 1810
box 0 0 128 200
use NAND2X1  NAND2X1_356
timestamp 1515870181
transform -1 0 2792 0 1 1810
box 0 0 48 200
use BUFX4  BUFX4_83
timestamp 1515870181
transform -1 0 2856 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_286
timestamp 1515870181
transform -1 0 2920 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_8
timestamp 1515870181
transform 1 0 2920 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_62
timestamp 1515870181
transform 1 0 2984 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_266
timestamp 1515870181
transform 1 0 3048 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_57
timestamp 1515870181
transform -1 0 3176 0 1 1810
box 0 0 64 200
use FILL  FILL_9_2_0
timestamp 1515870181
transform 1 0 3176 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1515870181
transform 1 0 3192 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_176
timestamp 1515870181
transform 1 0 3208 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_145
timestamp 1515870181
transform 1 0 3400 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_127
timestamp 1515870181
transform -1 0 3512 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_145
timestamp 1515870181
transform 1 0 3512 0 1 1810
box 0 0 192 200
use INVX1  INVX1_12
timestamp 1515870181
transform 1 0 3704 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_282
timestamp 1515870181
transform 1 0 3736 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_387
timestamp 1515870181
transform -1 0 3864 0 1 1810
box 0 0 64 200
use INVX1  INVX1_70
timestamp 1515870181
transform -1 0 3896 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_122
timestamp 1515870181
transform 1 0 3896 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_386
timestamp 1515870181
transform -1 0 3992 0 1 1810
box 0 0 48 200
use BUFX4  BUFX4_243
timestamp 1515870181
transform 1 0 3992 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_36
timestamp 1515870181
transform -1 0 4120 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_261
timestamp 1515870181
transform -1 0 4184 0 1 1810
box 0 0 64 200
use FILL  FILL_9_3_0
timestamp 1515870181
transform -1 0 4200 0 1 1810
box 0 0 16 200
use FILL  FILL_9_3_1
timestamp 1515870181
transform -1 0 4216 0 1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_128
timestamp 1515870181
transform -1 0 4280 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_118
timestamp 1515870181
transform 1 0 4280 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_388
timestamp 1515870181
transform -1 0 4392 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_274
timestamp 1515870181
transform 1 0 4392 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_10
timestamp 1515870181
transform -1 0 4504 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_14
timestamp 1515870181
transform -1 0 4568 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_170
timestamp 1515870181
transform -1 0 4632 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_389
timestamp 1515870181
transform 1 0 4632 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_82
timestamp 1515870181
transform 1 0 4680 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_280
timestamp 1515870181
transform -1 0 4792 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_93
timestamp 1515870181
transform 1 0 4792 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_421
timestamp 1515870181
transform -1 0 4904 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_386
timestamp 1515870181
transform 1 0 4904 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_278
timestamp 1515870181
transform 1 0 4968 0 1 1810
box 0 0 64 200
use INVX8  INVX8_13
timestamp 1515870181
transform -1 0 5112 0 1 1810
box 0 0 80 200
use INVX1  INVX1_90
timestamp 1515870181
transform 1 0 5112 0 1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_131
timestamp 1515870181
transform -1 0 5192 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_130
timestamp 1515870181
transform 1 0 5192 0 1 1810
box 0 0 48 200
use FILL  FILL_9_4_0
timestamp 1515870181
transform -1 0 5256 0 1 1810
box 0 0 16 200
use FILL  FILL_9_4_1
timestamp 1515870181
transform -1 0 5272 0 1 1810
box 0 0 16 200
use INVX1  INVX1_89
timestamp 1515870181
transform -1 0 5304 0 1 1810
box 0 0 32 200
use BUFX4  BUFX4_23
timestamp 1515870181
transform 1 0 5304 0 1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_25
timestamp 1515870181
transform -1 0 5496 0 1 1810
box 0 0 128 200
use OAI21X1  OAI21X1_466
timestamp 1515870181
transform -1 0 5560 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_382
timestamp 1515870181
transform 1 0 5560 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_301
timestamp 1515870181
transform -1 0 5816 0 1 1810
box 0 0 192 200
use NOR2X1  NOR2X1_70
timestamp 1515870181
transform 1 0 5816 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_61
timestamp 1515870181
transform -1 0 5928 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_49
timestamp 1515870181
transform 1 0 5928 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_58
timestamp 1515870181
transform -1 0 6040 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_85
timestamp 1515870181
transform -1 0 6104 0 1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1515870181
transform -1 0 6232 0 1 1810
box 0 0 128 200
use FILL  FILL_9_5_0
timestamp 1515870181
transform 1 0 6232 0 1 1810
box 0 0 16 200
use FILL  FILL_9_5_1
timestamp 1515870181
transform 1 0 6248 0 1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_247
timestamp 1515870181
transform 1 0 6264 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_245
timestamp 1515870181
transform 1 0 6328 0 1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_33
timestamp 1515870181
transform 1 0 6392 0 1 1810
box 0 0 128 200
use BUFX4  BUFX4_215
timestamp 1515870181
transform -1 0 6584 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_33
timestamp 1515870181
transform -1 0 6648 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_24
timestamp 1515870181
transform 1 0 6648 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_27
timestamp 1515870181
transform -1 0 6760 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_18
timestamp 1515870181
transform -1 0 6824 0 1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_242
timestamp 1515870181
transform 1 0 6824 0 1 1810
box 0 0 192 200
use NAND3X1  NAND3X1_296
timestamp 1515870181
transform -1 0 7080 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_297
timestamp 1515870181
transform 1 0 7080 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_295
timestamp 1515870181
transform 1 0 7144 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_14
timestamp 1515870181
transform 1 0 7208 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_23
timestamp 1515870181
transform 1 0 7272 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_155
timestamp 1515870181
transform 1 0 7320 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_10
timestamp 1515870181
transform -1 0 7432 0 1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_49
timestamp 1515870181
transform -1 0 200 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_65
timestamp 1515870181
transform -1 0 264 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_225
timestamp 1515870181
transform -1 0 328 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_267
timestamp 1515870181
transform -1 0 376 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_225
timestamp 1515870181
transform -1 0 568 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_81
timestamp 1515870181
transform -1 0 632 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_105
timestamp 1515870181
transform 1 0 632 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_106
timestamp 1515870181
transform -1 0 760 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_89
timestamp 1515870181
transform -1 0 824 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_352
timestamp 1515870181
transform -1 0 872 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_384
timestamp 1515870181
transform 1 0 872 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_61
timestamp 1515870181
transform 1 0 936 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_77
timestamp 1515870181
transform 1 0 1000 0 -1 1810
box 0 0 192 200
use FILL  FILL_8_0_0
timestamp 1515870181
transform 1 0 1192 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1515870181
transform 1 0 1208 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_173
timestamp 1515870181
transform 1 0 1224 0 -1 1810
box 0 0 192 200
use NAND2X1  NAND2X1_156
timestamp 1515870181
transform 1 0 1416 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_173
timestamp 1515870181
transform -1 0 1528 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_205
timestamp 1515870181
transform 1 0 1528 0 -1 1810
box 0 0 192 200
use BUFX4  BUFX4_141
timestamp 1515870181
transform -1 0 1784 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_192
timestamp 1515870181
transform -1 0 1976 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_192
timestamp 1515870181
transform 1 0 1976 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_176
timestamp 1515870181
transform -1 0 2088 0 -1 1810
box 0 0 48 200
use MUX2X1  MUX2X1_1
timestamp 1515870181
transform -1 0 2184 0 -1 1810
box 0 0 96 200
use FILL  FILL_8_1_0
timestamp 1515870181
transform -1 0 2200 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1515870181
transform -1 0 2216 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_56
timestamp 1515870181
transform -1 0 2280 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_67
timestamp 1515870181
transform 1 0 2280 0 -1 1810
box 0 0 192 200
use INVX1  INVX1_71
timestamp 1515870181
transform 1 0 2472 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_57
timestamp 1515870181
transform 1 0 2504 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_51
timestamp 1515870181
transform -1 0 2616 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_195
timestamp 1515870181
transform 1 0 2616 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_180
timestamp 1515870181
transform -1 0 2728 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_389
timestamp 1515870181
transform 1 0 2728 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_195
timestamp 1515870181
transform -1 0 2984 0 -1 1810
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_32
timestamp 1515870181
transform 1 0 2984 0 -1 1810
box 0 0 192 200
use FILL  FILL_8_2_0
timestamp 1515870181
transform 1 0 3176 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1515870181
transform 1 0 3192 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_35
timestamp 1515870181
transform 1 0 3208 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_32
timestamp 1515870181
transform -1 0 3320 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_176
timestamp 1515870181
transform 1 0 3320 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_159
timestamp 1515870181
transform -1 0 3432 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_142
timestamp 1515870181
transform 1 0 3432 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_86
timestamp 1515870181
transform 1 0 3496 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_377
timestamp 1515870181
transform -1 0 3576 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_416
timestamp 1515870181
transform 1 0 3576 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_141
timestamp 1515870181
transform 1 0 3640 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_141
timestamp 1515870181
transform 1 0 3704 0 -1 1810
box 0 0 192 200
use BUFX4  BUFX4_240
timestamp 1515870181
transform -1 0 3960 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_284
timestamp 1515870181
transform -1 0 4024 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_384
timestamp 1515870181
transform 1 0 4024 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_129
timestamp 1515870181
transform -1 0 4136 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_358
timestamp 1515870181
transform 1 0 4136 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_3_0
timestamp 1515870181
transform 1 0 4184 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_3_1
timestamp 1515870181
transform 1 0 4200 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_319
timestamp 1515870181
transform 1 0 4216 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_289
timestamp 1515870181
transform -1 0 4344 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_413
timestamp 1515870181
transform 1 0 4344 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_288
timestamp 1515870181
transform -1 0 4456 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_469
timestamp 1515870181
transform -1 0 4520 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_159
timestamp 1515870181
transform -1 0 4568 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_385
timestamp 1515870181
transform -1 0 4616 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_291
timestamp 1515870181
transform 1 0 4616 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_131
timestamp 1515870181
transform 1 0 4680 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_11
timestamp 1515870181
transform 1 0 4744 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_135
timestamp 1515870181
transform 1 0 4808 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_114
timestamp 1515870181
transform -1 0 4920 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_354
timestamp 1515870181
transform 1 0 4920 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_388
timestamp 1515870181
transform 1 0 4968 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_171
timestamp 1515870181
transform 1 0 5016 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_510
timestamp 1515870181
transform 1 0 5080 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_449
timestamp 1515870181
transform -1 0 5192 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_270
timestamp 1515870181
transform -1 0 5240 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_4_0
timestamp 1515870181
transform -1 0 5256 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_4_1
timestamp 1515870181
transform -1 0 5272 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_381
timestamp 1515870181
transform -1 0 5320 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_129
timestamp 1515870181
transform -1 0 5368 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_28
timestamp 1515870181
transform -1 0 5432 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_380
timestamp 1515870181
transform 1 0 5432 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_383
timestamp 1515870181
transform 1 0 5480 0 -1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_45
timestamp 1515870181
transform 1 0 5544 0 -1 1810
box 0 0 128 200
use OAI21X1  OAI21X1_467
timestamp 1515870181
transform 1 0 5672 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_123
timestamp 1515870181
transform 1 0 5736 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_283
timestamp 1515870181
transform 1 0 5800 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_289
timestamp 1515870181
transform 1 0 5864 0 -1 1810
box 0 0 192 200
use NAND3X1  NAND3X1_3
timestamp 1515870181
transform -1 0 6120 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_183
timestamp 1515870181
transform 1 0 6120 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_275
timestamp 1515870181
transform -1 0 6248 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_5_0
timestamp 1515870181
transform 1 0 6248 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_5_1
timestamp 1515870181
transform 1 0 6264 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_163
timestamp 1515870181
transform 1 0 6280 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_419
timestamp 1515870181
transform -1 0 6408 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_418
timestamp 1515870181
transform 1 0 6408 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_274
timestamp 1515870181
transform 1 0 6472 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_42
timestamp 1515870181
transform -1 0 6584 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_13
timestamp 1515870181
transform -1 0 6648 0 -1 1810
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_273
timestamp 1515870181
transform -1 0 6840 0 -1 1810
box 0 0 192 200
use BUFX4  BUFX4_116
timestamp 1515870181
transform 1 0 6840 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_39
timestamp 1515870181
transform 1 0 6904 0 -1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_30
timestamp 1515870181
transform -1 0 7016 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_73
timestamp 1515870181
transform -1 0 7064 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_254
timestamp 1515870181
transform -1 0 7256 0 -1 1810
box 0 0 192 200
use AOI21X1  AOI21X1_46
timestamp 1515870181
transform 1 0 7256 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_132
timestamp 1515870181
transform -1 0 7384 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_55
timestamp 1515870181
transform -1 0 7432 0 -1 1810
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_209
timestamp 1515870181
transform -1 0 200 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_195
timestamp 1515870181
transform 1 0 200 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_209
timestamp 1515870181
transform -1 0 312 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_33
timestamp 1515870181
transform -1 0 504 0 1 1410
box 0 0 192 200
use BUFX4  BUFX4_52
timestamp 1515870181
transform -1 0 568 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_82
timestamp 1515870181
transform -1 0 632 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_222
timestamp 1515870181
transform 1 0 632 0 1 1410
box 0 0 192 200
use BUFX4  BUFX4_53
timestamp 1515870181
transform 1 0 824 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_86
timestamp 1515870181
transform 1 0 888 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_273
timestamp 1515870181
transform 1 0 952 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_64
timestamp 1515870181
transform 1 0 1016 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_70
timestamp 1515870181
transform -1 0 1128 0 1 1410
box 0 0 48 200
use FILL  FILL_7_0_0
timestamp 1515870181
transform -1 0 1144 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1515870181
transform -1 0 1160 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_154
timestamp 1515870181
transform -1 0 1208 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_80
timestamp 1515870181
transform 1 0 1208 0 1 1410
box 0 0 192 200
use BUFX4  BUFX4_163
timestamp 1515870181
transform 1 0 1400 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_105
timestamp 1515870181
transform 1 0 1464 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_193
timestamp 1515870181
transform 1 0 1528 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_208
timestamp 1515870181
transform -1 0 1640 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_208
timestamp 1515870181
transform -1 0 1832 0 1 1410
box 0 0 192 200
use MUX2X1  MUX2X1_47
timestamp 1515870181
transform 1 0 1832 0 1 1410
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1515870181
transform -1 0 2120 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_53
timestamp 1515870181
transform 1 0 2120 0 1 1410
box 0 0 48 200
use FILL  FILL_7_1_0
timestamp 1515870181
transform -1 0 2184 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1515870181
transform -1 0 2200 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_48
timestamp 1515870181
transform -1 0 2264 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_198
timestamp 1515870181
transform 1 0 2264 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_146
timestamp 1515870181
transform 1 0 2328 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_128
timestamp 1515870181
transform -1 0 2440 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_161
timestamp 1515870181
transform 1 0 2440 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_244
timestamp 1515870181
transform 1 0 2504 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_157
timestamp 1515870181
transform -1 0 2760 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_157
timestamp 1515870181
transform 1 0 2760 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_139
timestamp 1515870181
transform -1 0 2872 0 1 1410
box 0 0 48 200
use INVX1  INVX1_72
timestamp 1515870181
transform 1 0 2872 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_390
timestamp 1515870181
transform 1 0 2904 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_357
timestamp 1515870181
transform -1 0 3016 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_125
timestamp 1515870181
transform -1 0 3208 0 1 1410
box 0 0 192 200
use FILL  FILL_7_2_0
timestamp 1515870181
transform 1 0 3208 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1515870181
transform 1 0 3224 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_15
timestamp 1515870181
transform 1 0 3240 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_13
timestamp 1515870181
transform -1 0 3352 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_160
timestamp 1515870181
transform 1 0 3352 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_142
timestamp 1515870181
transform -1 0 3464 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_160
timestamp 1515870181
transform 1 0 3464 0 1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_144
timestamp 1515870181
transform 1 0 3656 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_144
timestamp 1515870181
transform -1 0 3912 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_125
timestamp 1515870181
transform -1 0 3960 0 1 1410
box 0 0 48 200
use INVX1  INVX1_85
timestamp 1515870181
transform 1 0 3960 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_414
timestamp 1515870181
transform 1 0 3992 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_37
timestamp 1515870181
transform -1 0 4120 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_130
timestamp 1515870181
transform -1 0 4184 0 1 1410
box 0 0 64 200
use FILL  FILL_7_3_0
timestamp 1515870181
transform 1 0 4184 0 1 1410
box 0 0 16 200
use FILL  FILL_7_3_1
timestamp 1515870181
transform 1 0 4200 0 1 1410
box 0 0 16 200
use NAND3X1  NAND3X1_159
timestamp 1515870181
transform 1 0 4216 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_290
timestamp 1515870181
transform 1 0 4280 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_136
timestamp 1515870181
transform -1 0 4408 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_160
timestamp 1515870181
transform -1 0 4472 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_379
timestamp 1515870181
transform 1 0 4472 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_127
timestamp 1515870181
transform 1 0 4520 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_137
timestamp 1515870181
transform -1 0 4632 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_158
timestamp 1515870181
transform -1 0 4696 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_415
timestamp 1515870181
transform -1 0 4760 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_327
timestamp 1515870181
transform -1 0 4808 0 1 1410
box 0 0 48 200
use BUFX4  BUFX4_35
timestamp 1515870181
transform -1 0 4872 0 1 1410
box 0 0 64 200
use BUFX2  BUFX2_29
timestamp 1515870181
transform -1 0 4920 0 1 1410
box 0 0 48 200
use BUFX2  BUFX2_17
timestamp 1515870181
transform -1 0 4968 0 1 1410
box 0 0 48 200
use INVX1  INVX1_69
timestamp 1515870181
transform 1 0 4968 0 1 1410
box 0 0 32 200
use BUFX4  BUFX4_135
timestamp 1515870181
transform -1 0 5064 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_308
timestamp 1515870181
transform 1 0 5064 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_296
timestamp 1515870181
transform -1 0 5192 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_311
timestamp 1515870181
transform 1 0 5192 0 1 1410
box 0 0 64 200
use FILL  FILL_7_4_0
timestamp 1515870181
transform -1 0 5272 0 1 1410
box 0 0 16 200
use FILL  FILL_7_4_1
timestamp 1515870181
transform -1 0 5288 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_339
timestamp 1515870181
transform -1 0 5480 0 1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_95
timestamp 1515870181
transform 1 0 5480 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_115
timestamp 1515870181
transform -1 0 5592 0 1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_43
timestamp 1515870181
transform 1 0 5592 0 1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_458
timestamp 1515870181
transform 1 0 5720 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_262
timestamp 1515870181
transform -1 0 5848 0 1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_21
timestamp 1515870181
transform 1 0 5848 0 1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_364
timestamp 1515870181
transform 1 0 5976 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_102
timestamp 1515870181
transform 1 0 6040 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_283
timestamp 1515870181
transform -1 0 6296 0 1 1410
box 0 0 192 200
use FILL  FILL_7_5_0
timestamp 1515870181
transform -1 0 6312 0 1 1410
box 0 0 16 200
use FILL  FILL_7_5_1
timestamp 1515870181
transform -1 0 6328 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_281
timestamp 1515870181
transform -1 0 6520 0 1 1410
box 0 0 192 200
use NAND3X1  NAND3X1_2
timestamp 1515870181
transform -1 0 6584 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_162
timestamp 1515870181
transform 1 0 6584 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_184
timestamp 1515870181
transform 1 0 6648 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_43
timestamp 1515870181
transform -1 0 6760 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_34
timestamp 1515870181
transform -1 0 6824 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_274
timestamp 1515870181
transform -1 0 7016 0 1 1410
box 0 0 192 200
use BUFX4  BUFX4_247
timestamp 1515870181
transform 1 0 7016 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_64
timestamp 1515870181
transform -1 0 7144 0 1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_304
timestamp 1515870181
transform -1 0 7336 0 1 1410
box 0 0 192 200
use AOI21X1  AOI21X1_48
timestamp 1515870181
transform 1 0 7336 0 1 1410
box 0 0 64 200
use FILL  FILL_8_1
timestamp 1515870181
transform 1 0 7400 0 1 1410
box 0 0 16 200
use FILL  FILL_8_2
timestamp 1515870181
transform 1 0 7416 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_62
timestamp 1515870181
transform 1 0 8 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_78
timestamp 1515870181
transform 1 0 200 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_86
timestamp 1515870181
transform -1 0 312 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_128
timestamp 1515870181
transform -1 0 376 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_83
timestamp 1515870181
transform 1 0 376 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_75
timestamp 1515870181
transform -1 0 488 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_222
timestamp 1515870181
transform 1 0 488 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_208
timestamp 1515870181
transform -1 0 600 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_272
timestamp 1515870181
transform -1 0 664 0 -1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_42
timestamp 1515870181
transform -1 0 760 0 -1 1410
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_210
timestamp 1515870181
transform 1 0 760 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_210
timestamp 1515870181
transform 1 0 952 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_196
timestamp 1515870181
transform -1 0 1064 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_171
timestamp 1515870181
transform 1 0 1064 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_0_0
timestamp 1515870181
transform 1 0 1128 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1515870181
transform 1 0 1144 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_171
timestamp 1515870181
transform 1 0 1160 0 -1 1410
box 0 0 192 200
use MUX2X1  MUX2X1_46
timestamp 1515870181
transform -1 0 1448 0 -1 1410
box 0 0 96 200
use OAI21X1  OAI21X1_49
timestamp 1515870181
transform 1 0 1448 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_55
timestamp 1515870181
transform -1 0 1560 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_61
timestamp 1515870181
transform 1 0 1560 0 -1 1410
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_65
timestamp 1515870181
transform -1 0 1784 0 -1 1410
box 0 0 192 200
use NOR2X1  NOR2X1_125
timestamp 1515870181
transform -1 0 1832 0 -1 1410
box 0 0 48 200
use OAI22X1  OAI22X1_16
timestamp 1515870181
transform -1 0 1912 0 -1 1410
box 0 0 80 200
use NOR2X1  NOR2X1_126
timestamp 1515870181
transform -1 0 1960 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_164
timestamp 1515870181
transform -1 0 2008 0 -1 1410
box 0 0 48 200
use NOR3X1  NOR3X1_32
timestamp 1515870181
transform 1 0 2008 0 -1 1410
box 0 0 128 200
use FILL  FILL_6_1_0
timestamp 1515870181
transform 1 0 2136 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1515870181
transform 1 0 2152 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_3
timestamp 1515870181
transform 1 0 2168 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_146
timestamp 1515870181
transform 1 0 2232 0 -1 1410
box 0 0 192 200
use INVX1  INVX1_17
timestamp 1515870181
transform 1 0 2424 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_291
timestamp 1515870181
transform 1 0 2456 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_280
timestamp 1515870181
transform 1 0 2520 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_114
timestamp 1515870181
transform -1 0 2760 0 -1 1410
box 0 0 192 200
use BUFX4  BUFX4_70
timestamp 1515870181
transform -1 0 2824 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_49
timestamp 1515870181
transform 1 0 2824 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_371
timestamp 1515870181
transform 1 0 2888 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_4
timestamp 1515870181
transform 1 0 2952 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_2
timestamp 1515870181
transform -1 0 3064 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_189
timestamp 1515870181
transform 1 0 3064 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_378
timestamp 1515870181
transform 1 0 3128 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_2_0
timestamp 1515870181
transform 1 0 3176 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1515870181
transform 1 0 3192 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_497
timestamp 1515870181
transform 1 0 3208 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_436
timestamp 1515870181
transform -1 0 3320 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_96
timestamp 1515870181
transform 1 0 3320 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_417
timestamp 1515870181
transform -1 0 3576 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_87
timestamp 1515870181
transform -1 0 3608 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_376
timestamp 1515870181
transform 1 0 3608 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_190
timestamp 1515870181
transform 1 0 3656 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_109
timestamp 1515870181
transform -1 0 3784 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_20
timestamp 1515870181
transform -1 0 3848 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_269
timestamp 1515870181
transform -1 0 3912 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_180
timestamp 1515870181
transform -1 0 3976 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_320
timestamp 1515870181
transform -1 0 4040 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_318
timestamp 1515870181
transform -1 0 4104 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_419
timestamp 1515870181
transform -1 0 4152 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_165
timestamp 1515870181
transform 1 0 4152 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_3_0
timestamp 1515870181
transform -1 0 4216 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_3_1
timestamp 1515870181
transform -1 0 4232 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_481
timestamp 1515870181
transform -1 0 4296 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_321
timestamp 1515870181
transform 1 0 4296 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_248
timestamp 1515870181
transform -1 0 4424 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_88
timestamp 1515870181
transform -1 0 4488 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_161
timestamp 1515870181
transform 1 0 4488 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_351
timestamp 1515870181
transform -1 0 4616 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_490
timestamp 1515870181
transform 1 0 4616 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_429
timestamp 1515870181
transform -1 0 4728 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_89
timestamp 1515870181
transform -1 0 4920 0 -1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_109
timestamp 1515870181
transform -1 0 5112 0 -1 1410
box 0 0 192 200
use NAND2X1  NAND2X1_284
timestamp 1515870181
transform 1 0 5112 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_4_0
timestamp 1515870181
transform 1 0 5160 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_4_1
timestamp 1515870181
transform 1 0 5176 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_297
timestamp 1515870181
transform 1 0 5192 0 -1 1410
box 0 0 192 200
use NOR2X1  NOR2X1_66
timestamp 1515870181
transform -1 0 5432 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_57
timestamp 1515870181
transform -1 0 5496 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_459
timestamp 1515870181
transform 1 0 5496 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_263
timestamp 1515870181
transform -1 0 5624 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_103
timestamp 1515870181
transform 1 0 5624 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_365
timestamp 1515870181
transform -1 0 5752 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_83
timestamp 1515870181
transform 1 0 5752 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_243
timestamp 1515870181
transform 1 0 5816 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_43
timestamp 1515870181
transform 1 0 5880 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_52
timestamp 1515870181
transform -1 0 5992 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_226
timestamp 1515870181
transform 1 0 5992 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_82
timestamp 1515870181
transform -1 0 6120 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_50
timestamp 1515870181
transform -1 0 6168 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_41
timestamp 1515870181
transform -1 0 6232 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_5_0
timestamp 1515870181
transform 1 0 6232 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_5_1
timestamp 1515870181
transform 1 0 6248 0 -1 1410
box 0 0 16 200
use NAND3X1  NAND3X1_242
timestamp 1515870181
transform 1 0 6264 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_173
timestamp 1515870181
transform -1 0 6392 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_172
timestamp 1515870181
transform -1 0 6456 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_13
timestamp 1515870181
transform -1 0 6520 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_133
timestamp 1515870181
transform -1 0 6584 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_153
timestamp 1515870181
transform -1 0 6648 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_313
timestamp 1515870181
transform -1 0 6712 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_293
timestamp 1515870181
transform -1 0 6776 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_12
timestamp 1515870181
transform 1 0 6776 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_479
timestamp 1515870181
transform -1 0 6904 0 -1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_48
timestamp 1515870181
transform 1 0 6904 0 -1 1410
box 0 0 128 200
use NAND3X1  NAND3X1_152
timestamp 1515870181
transform -1 0 7096 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_312
timestamp 1515870181
transform -1 0 7160 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_292
timestamp 1515870181
transform -1 0 7224 0 -1 1410
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_288
timestamp 1515870181
transform -1 0 7416 0 -1 1410
box 0 0 192 200
use FILL  FILL_7_1
timestamp 1515870181
transform -1 0 7432 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_219
timestamp 1515870181
transform 1 0 8 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_219
timestamp 1515870181
transform 1 0 200 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_205
timestamp 1515870181
transform -1 0 312 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_59
timestamp 1515870181
transform -1 0 504 0 1 1010
box 0 0 192 200
use MUX2X1  MUX2X1_33
timestamp 1515870181
transform 1 0 504 0 1 1010
box 0 0 96 200
use INVX1  INVX1_68
timestamp 1515870181
transform 1 0 600 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_111
timestamp 1515870181
transform 1 0 632 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_48
timestamp 1515870181
transform -1 0 888 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_112
timestamp 1515870181
transform -1 0 952 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_373
timestamp 1515870181
transform -1 0 1000 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_411
timestamp 1515870181
transform -1 0 1064 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_408
timestamp 1515870181
transform 1 0 1064 0 1 1010
box 0 0 48 200
use FILL  FILL_5_0_0
timestamp 1515870181
transform -1 0 1128 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1515870181
transform -1 0 1144 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_460
timestamp 1515870181
transform -1 0 1208 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_414
timestamp 1515870181
transform -1 0 1256 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_360
timestamp 1515870181
transform 1 0 1256 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_276
timestamp 1515870181
transform 1 0 1304 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_390
timestamp 1515870181
transform 1 0 1352 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_339
timestamp 1515870181
transform 1 0 1400 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_404
timestamp 1515870181
transform -1 0 1496 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_325
timestamp 1515870181
transform 1 0 1496 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_367
timestamp 1515870181
transform -1 0 1608 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_169
timestamp 1515870181
transform 1 0 1608 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_152
timestamp 1515870181
transform -1 0 1720 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_169
timestamp 1515870181
transform 1 0 1720 0 1 1010
box 0 0 192 200
use BUFX4  BUFX4_103
timestamp 1515870181
transform -1 0 1976 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_418
timestamp 1515870181
transform 1 0 1976 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_480
timestamp 1515870181
transform -1 0 2088 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_374
timestamp 1515870181
transform 1 0 2088 0 1 1010
box 0 0 48 200
use FILL  FILL_5_1_0
timestamp 1515870181
transform -1 0 2152 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1515870181
transform -1 0 2168 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_412
timestamp 1515870181
transform -1 0 2232 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_154
timestamp 1515870181
transform 1 0 2232 0 1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_11
timestamp 1515870181
transform -1 0 2360 0 1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_111
timestamp 1515870181
transform -1 0 2408 0 1 1010
box 0 0 48 200
use NOR3X1  NOR3X1_22
timestamp 1515870181
transform -1 0 2536 0 1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_110
timestamp 1515870181
transform -1 0 2584 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_69
timestamp 1515870181
transform 1 0 2584 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_25
timestamp 1515870181
transform 1 0 2648 0 1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_28
timestamp 1515870181
transform 1 0 2840 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_25
timestamp 1515870181
transform -1 0 2952 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_328
timestamp 1515870181
transform -1 0 3000 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_128
timestamp 1515870181
transform 1 0 3000 0 1 1010
box 0 0 192 200
use FILL  FILL_5_2_0
timestamp 1515870181
transform 1 0 3192 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1515870181
transform 1 0 3208 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_18
timestamp 1515870181
transform 1 0 3224 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_16
timestamp 1515870181
transform -1 0 3336 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_82
timestamp 1515870181
transform 1 0 3336 0 1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_278
timestamp 1515870181
transform -1 0 3576 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_290
timestamp 1515870181
transform -1 0 3640 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_344
timestamp 1515870181
transform 1 0 3640 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_110
timestamp 1515870181
transform -1 0 3752 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_19
timestamp 1515870181
transform -1 0 3816 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_281
timestamp 1515870181
transform 1 0 3816 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_179
timestamp 1515870181
transform -1 0 3928 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_391
timestamp 1515870181
transform 1 0 3928 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_409
timestamp 1515870181
transform 1 0 3976 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_27
timestamp 1515870181
transform -1 0 4072 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_111
timestamp 1515870181
transform 1 0 4072 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_112
timestamp 1515870181
transform 1 0 4136 0 1 1010
box 0 0 48 200
use FILL  FILL_5_3_0
timestamp 1515870181
transform -1 0 4200 0 1 1010
box 0 0 16 200
use FILL  FILL_5_3_1
timestamp 1515870181
transform -1 0 4216 0 1 1010
box 0 0 16 200
use NAND3X1  NAND3X1_138
timestamp 1515870181
transform -1 0 4280 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_298
timestamp 1515870181
transform 1 0 4280 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_178
timestamp 1515870181
transform -1 0 4408 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_137
timestamp 1515870181
transform 1 0 4408 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_425
timestamp 1515870181
transform -1 0 4520 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_18
timestamp 1515870181
transform 1 0 4520 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_289
timestamp 1515870181
transform -1 0 4648 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_108
timestamp 1515870181
transform -1 0 4712 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_370
timestamp 1515870181
transform -1 0 4776 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_268
timestamp 1515870181
transform -1 0 4840 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_461
timestamp 1515870181
transform -1 0 4904 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_155
timestamp 1515870181
transform 1 0 4904 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_271
timestamp 1515870181
transform 1 0 4952 0 1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_347
timestamp 1515870181
transform -1 0 5208 0 1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_103
timestamp 1515870181
transform 1 0 5208 0 1 1010
box 0 0 48 200
use FILL  FILL_5_4_0
timestamp 1515870181
transform -1 0 5272 0 1 1010
box 0 0 16 200
use FILL  FILL_5_4_1
timestamp 1515870181
transform -1 0 5288 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_123
timestamp 1515870181
transform -1 0 5352 0 1 1010
box 0 0 64 200
use INVX8  INVX8_1
timestamp 1515870181
transform 1 0 5352 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_256
timestamp 1515870181
transform 1 0 5432 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_270
timestamp 1515870181
transform -1 0 5544 0 1 1010
box 0 0 64 200
use INVX2  INVX2_30
timestamp 1515870181
transform -1 0 5576 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_317
timestamp 1515870181
transform -1 0 5768 0 1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_347
timestamp 1515870181
transform -1 0 5832 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_451
timestamp 1515870181
transform -1 0 5896 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_17
timestamp 1515870181
transform 1 0 5896 0 1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_346
timestamp 1515870181
transform 1 0 6024 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_228
timestamp 1515870181
transform 1 0 6088 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_242
timestamp 1515870181
transform -1 0 6200 0 1 1010
box 0 0 64 200
use FILL  FILL_5_5_0
timestamp 1515870181
transform 1 0 6200 0 1 1010
box 0 0 16 200
use FILL  FILL_5_5_1
timestamp 1515870181
transform 1 0 6216 0 1 1010
box 0 0 16 200
use NOR3X1  NOR3X1_41
timestamp 1515870181
transform 1 0 6232 0 1 1010
box 0 0 128 200
use INVX2  INVX2_2
timestamp 1515870181
transform 1 0 6360 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_450
timestamp 1515870181
transform -1 0 6456 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_423
timestamp 1515870181
transform -1 0 6520 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_422
timestamp 1515870181
transform -1 0 6584 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_284
timestamp 1515870181
transform -1 0 6648 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_3
timestamp 1515870181
transform 1 0 6648 0 1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_283
timestamp 1515870181
transform -1 0 6840 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_410
timestamp 1515870181
transform -1 0 6904 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_392
timestamp 1515870181
transform -1 0 6968 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_31
timestamp 1515870181
transform 1 0 6968 0 1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_409
timestamp 1515870181
transform -1 0 7160 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_478
timestamp 1515870181
transform -1 0 7224 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_470
timestamp 1515870181
transform -1 0 7288 0 1 1010
box 0 0 64 200
use INVX2  INVX2_3
timestamp 1515870181
transform -1 0 7320 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_391
timestamp 1515870181
transform 1 0 7320 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_31
timestamp 1515870181
transform -1 0 7432 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_235
timestamp 1515870181
transform 1 0 8 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_235
timestamp 1515870181
transform 1 0 200 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_222
timestamp 1515870181
transform -1 0 312 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_43
timestamp 1515870181
transform -1 0 376 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_41
timestamp 1515870181
transform 1 0 376 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_58
timestamp 1515870181
transform 1 0 440 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_366
timestamp 1515870181
transform 1 0 472 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_348
timestamp 1515870181
transform 1 0 536 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_393
timestamp 1515870181
transform -1 0 664 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_65
timestamp 1515870181
transform -1 0 728 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_57
timestamp 1515870181
transform 1 0 728 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_73
timestamp 1515870181
transform 1 0 920 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_81
timestamp 1515870181
transform -1 0 1032 0 -1 1010
box 0 0 48 200
use MUX2X1  MUX2X1_6
timestamp 1515870181
transform 1 0 1032 0 -1 1010
box 0 0 96 200
use FILL  FILL_4_0_0
timestamp 1515870181
transform 1 0 1128 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1515870181
transform 1 0 1144 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_472
timestamp 1515870181
transform 1 0 1160 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_394
timestamp 1515870181
transform 1 0 1224 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_286
timestamp 1515870181
transform 1 0 1288 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_424
timestamp 1515870181
transform 1 0 1352 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_452
timestamp 1515870181
transform 1 0 1416 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_349
timestamp 1515870181
transform 1 0 1480 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_136
timestamp 1515870181
transform 1 0 1544 0 -1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_2
timestamp 1515870181
transform -1 0 1672 0 -1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_83
timestamp 1515870181
transform 1 0 1672 0 -1 1010
box 0 0 48 200
use NOR3X1  NOR3X1_4
timestamp 1515870181
transform -1 0 1848 0 -1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_84
timestamp 1515870181
transform 1 0 1848 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_121
timestamp 1515870181
transform -1 0 1960 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_150
timestamp 1515870181
transform 1 0 1960 0 -1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_9
timestamp 1515870181
transform -1 0 2088 0 -1 1010
box 0 0 80 200
use NOR3X1  NOR3X1_28
timestamp 1515870181
transform -1 0 2216 0 -1 1010
box 0 0 128 200
use FILL  FILL_4_1_0
timestamp 1515870181
transform -1 0 2232 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1515870181
transform -1 0 2248 0 -1 1010
box 0 0 16 200
use NOR2X1  NOR2X1_119
timestamp 1515870181
transform -1 0 2296 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_120
timestamp 1515870181
transform -1 0 2344 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_160
timestamp 1515870181
transform 1 0 2344 0 -1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_14
timestamp 1515870181
transform -1 0 2472 0 -1 1010
box 0 0 80 200
use MUX2X1  MUX2X1_40
timestamp 1515870181
transform 1 0 2472 0 -1 1010
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_78
timestamp 1515870181
transform -1 0 2760 0 -1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_68
timestamp 1515870181
transform 1 0 2760 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_62
timestamp 1515870181
transform -1 0 2872 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_51
timestamp 1515870181
transform 1 0 2872 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_353
timestamp 1515870181
transform 1 0 2904 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_168
timestamp 1515870181
transform 1 0 2968 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_18
timestamp 1515870181
transform 1 0 3032 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_21
timestamp 1515870181
transform -1 0 3144 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_2_0
timestamp 1515870181
transform 1 0 3144 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1515870181
transform 1 0 3160 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_18
timestamp 1515870181
transform 1 0 3176 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_483
timestamp 1515870181
transform 1 0 3368 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_422
timestamp 1515870181
transform -1 0 3480 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_141
timestamp 1515870181
transform 1 0 3480 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_279
timestamp 1515870181
transform -1 0 3592 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_288
timestamp 1515870181
transform -1 0 3656 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_121
timestamp 1515870181
transform -1 0 3704 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_365
timestamp 1515870181
transform -1 0 3752 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_139
timestamp 1515870181
transform -1 0 3816 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_89
timestamp 1515870181
transform -1 0 3880 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_249
timestamp 1515870181
transform -1 0 3944 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_397
timestamp 1515870181
transform 1 0 3944 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_299
timestamp 1515870181
transform -1 0 4072 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_330
timestamp 1515870181
transform 1 0 4072 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_415
timestamp 1515870181
transform 1 0 4120 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_161
timestamp 1515870181
transform 1 0 4168 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_3_0
timestamp 1515870181
transform 1 0 4216 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_1
timestamp 1515870181
transform 1 0 4232 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_473
timestamp 1515870181
transform 1 0 4248 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_301
timestamp 1515870181
transform 1 0 4312 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_405
timestamp 1515870181
transform 1 0 4376 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_181
timestamp 1515870181
transform 1 0 4424 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_85
timestamp 1515870181
transform 1 0 4488 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_21
timestamp 1515870181
transform 1 0 4536 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_106
timestamp 1515870181
transform 1 0 4600 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_352
timestamp 1515870181
transform -1 0 4712 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_453
timestamp 1515870181
transform -1 0 4776 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_151
timestamp 1515870181
transform -1 0 4824 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_91
timestamp 1515870181
transform 1 0 4824 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_251
timestamp 1515870181
transform 1 0 4888 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_94
timestamp 1515870181
transform -1 0 5016 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_368
timestamp 1515870181
transform 1 0 5016 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_350
timestamp 1515870181
transform 1 0 5080 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_4_0
timestamp 1515870181
transform -1 0 5160 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_4_1
timestamp 1515870181
transform -1 0 5176 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_345
timestamp 1515870181
transform -1 0 5368 0 -1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_101
timestamp 1515870181
transform 1 0 5368 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_121
timestamp 1515870181
transform -1 0 5480 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_193
timestamp 1515870181
transform 1 0 5480 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_120
timestamp 1515870181
transform -1 0 5608 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_68
timestamp 1515870181
transform 1 0 5608 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_59
timestamp 1515870181
transform -1 0 5720 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_72
timestamp 1515870181
transform 1 0 5720 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_266
timestamp 1515870181
transform 1 0 5784 0 -1 1010
box 0 0 64 200
use INVX2  INVX2_26
timestamp 1515870181
transform -1 0 5880 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_313
timestamp 1515870181
transform -1 0 6072 0 -1 1010
box 0 0 192 200
use BUFX4  BUFX4_25
timestamp 1515870181
transform 1 0 6072 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_257
timestamp 1515870181
transform 1 0 6136 0 -1 1010
box 0 0 192 200
use FILL  FILL_4_5_0
timestamp 1515870181
transform -1 0 6344 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_5_1
timestamp 1515870181
transform -1 0 6360 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_254
timestamp 1515870181
transform -1 0 6424 0 -1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_34
timestamp 1515870181
transform -1 0 6552 0 -1 1010
box 0 0 128 200
use DFFPOSX1  DFFPOSX1_302
timestamp 1515870181
transform 1 0 6552 0 -1 1010
box 0 0 192 200
use BUFX4  BUFX4_101
timestamp 1515870181
transform 1 0 6744 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_112
timestamp 1515870181
transform 1 0 6808 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_62
timestamp 1515870181
transform 1 0 6872 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_71
timestamp 1515870181
transform 1 0 6936 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_471
timestamp 1515870181
transform 1 0 6984 0 -1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_46
timestamp 1515870181
transform 1 0 7048 0 -1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_271
timestamp 1515870181
transform -1 0 7240 0 -1 1010
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_318
timestamp 1515870181
transform -1 0 7432 0 -1 1010
box 0 0 192 200
use OAI21X1  OAI21X1_238
timestamp 1515870181
transform -1 0 72 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_238
timestamp 1515870181
transform 1 0 72 0 1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_41
timestamp 1515870181
transform 1 0 264 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_98
timestamp 1515870181
transform 1 0 456 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_97
timestamp 1515870181
transform -1 0 584 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_324
timestamp 1515870181
transform -1 0 632 0 1 610
box 0 0 48 200
use INVX1  INVX1_73
timestamp 1515870181
transform 1 0 632 0 1 610
box 0 0 32 200
use BUFX4  BUFX4_92
timestamp 1515870181
transform -1 0 728 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_240
timestamp 1515870181
transform 1 0 728 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_240
timestamp 1515870181
transform 1 0 920 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_227
timestamp 1515870181
transform -1 0 1032 0 1 610
box 0 0 48 200
use INVX1  INVX1_83
timestamp 1515870181
transform 1 0 1032 0 1 610
box 0 0 32 200
use MUX2X1  MUX2X1_27
timestamp 1515870181
transform 1 0 1064 0 1 610
box 0 0 96 200
use FILL  FILL_3_0_0
timestamp 1515870181
transform 1 0 1160 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1515870181
transform 1 0 1176 0 1 610
box 0 0 16 200
use OAI21X1  OAI21X1_224
timestamp 1515870181
transform 1 0 1192 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_210
timestamp 1515870181
transform -1 0 1304 0 1 610
box 0 0 48 200
use MUX2X1  MUX2X1_48
timestamp 1515870181
transform 1 0 1304 0 1 610
box 0 0 96 200
use OAI21X1  OAI21X1_80
timestamp 1515870181
transform 1 0 1400 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_88
timestamp 1515870181
transform -1 0 1512 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_178
timestamp 1515870181
transform 1 0 1512 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_162
timestamp 1515870181
transform -1 0 1624 0 1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_178
timestamp 1515870181
transform 1 0 1624 0 1 610
box 0 0 192 200
use MUX2X1  MUX2X1_5
timestamp 1515870181
transform 1 0 1816 0 1 610
box 0 0 96 200
use BUFX4  BUFX4_246
timestamp 1515870181
transform -1 0 1976 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_199
timestamp 1515870181
transform 1 0 1976 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_104
timestamp 1515870181
transform 1 0 2040 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_105
timestamp 1515870181
transform 1 0 2088 0 1 610
box 0 0 48 200
use FILL  FILL_3_1_0
timestamp 1515870181
transform 1 0 2136 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1515870181
transform 1 0 2152 0 1 610
box 0 0 16 200
use NOR3X1  NOR3X1_18
timestamp 1515870181
transform 1 0 2168 0 1 610
box 0 0 128 200
use OAI21X1  OAI21X1_187
timestamp 1515870181
transform 1 0 2296 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_171
timestamp 1515870181
transform -1 0 2408 0 1 610
box 0 0 48 200
use MUX2X1  MUX2X1_32
timestamp 1515870181
transform -1 0 2504 0 1 610
box 0 0 96 200
use NAND2X1  NAND2X1_191
timestamp 1515870181
transform 1 0 2504 0 1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_187
timestamp 1515870181
transform -1 0 2744 0 1 610
box 0 0 192 200
use NAND2X1  NAND2X1_188
timestamp 1515870181
transform -1 0 2792 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_59
timestamp 1515870181
transform 1 0 2792 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_65
timestamp 1515870181
transform -1 0 2904 0 1 610
box 0 0 48 200
use MUX2X1  MUX2X1_31
timestamp 1515870181
transform 1 0 2904 0 1 610
box 0 0 96 200
use BUFX4  BUFX4_12
timestamp 1515870181
transform 1 0 3000 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_75
timestamp 1515870181
transform -1 0 3256 0 1 610
box 0 0 192 200
use FILL  FILL_3_2_0
timestamp 1515870181
transform 1 0 3256 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1515870181
transform 1 0 3272 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_50
timestamp 1515870181
transform 1 0 3288 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_162
timestamp 1515870181
transform 1 0 3352 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_162
timestamp 1515870181
transform 1 0 3544 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_145
timestamp 1515870181
transform -1 0 3656 0 1 610
box 0 0 48 200
use INVX1  INVX1_16
timestamp 1515870181
transform 1 0 3656 0 1 610
box 0 0 32 200
use INVX1  INVX1_15
timestamp 1515870181
transform -1 0 3720 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_130
timestamp 1515870181
transform 1 0 3720 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_111
timestamp 1515870181
transform 1 0 3784 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_140
timestamp 1515870181
transform 1 0 3832 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_120
timestamp 1515870181
transform -1 0 3944 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_270
timestamp 1515870181
transform -1 0 4008 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_245
timestamp 1515870181
transform -1 0 4072 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_90
timestamp 1515870181
transform -1 0 4136 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_300
timestamp 1515870181
transform 1 0 4136 0 1 610
box 0 0 64 200
use FILL  FILL_3_3_0
timestamp 1515870181
transform -1 0 4216 0 1 610
box 0 0 16 200
use FILL  FILL_3_3_1
timestamp 1515870181
transform -1 0 4232 0 1 610
box 0 0 16 200
use NAND3X1  NAND3X1_250
timestamp 1515870181
transform -1 0 4296 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_157
timestamp 1515870181
transform 1 0 4296 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_174
timestamp 1515870181
transform -1 0 4408 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_174
timestamp 1515870181
transform -1 0 4600 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_495
timestamp 1515870181
transform 1 0 4600 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_434
timestamp 1515870181
transform -1 0 4712 0 1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_94
timestamp 1515870181
transform -1 0 4904 0 1 610
box 0 0 192 200
use BUFX2  BUFX2_18
timestamp 1515870181
transform 1 0 4904 0 1 610
box 0 0 48 200
use INVX1  INVX1_45
timestamp 1515870181
transform 1 0 4952 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_489
timestamp 1515870181
transform 1 0 4984 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_428
timestamp 1515870181
transform -1 0 5096 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_342
timestamp 1515870181
transform 1 0 5096 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_320
timestamp 1515870181
transform -1 0 5208 0 1 610
box 0 0 48 200
use FILL  FILL_3_4_0
timestamp 1515870181
transform -1 0 5224 0 1 610
box 0 0 16 200
use FILL  FILL_3_4_1
timestamp 1515870181
transform -1 0 5240 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_88
timestamp 1515870181
transform -1 0 5432 0 1 610
box 0 0 192 200
use INVX8  INVX8_3
timestamp 1515870181
transform 1 0 5432 0 1 610
box 0 0 80 200
use INVX1  INVX1_59
timestamp 1515870181
transform 1 0 5512 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_340
timestamp 1515870181
transform 1 0 5544 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_303
timestamp 1515870181
transform 1 0 5592 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_447
timestamp 1515870181
transform -1 0 5704 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_304
timestamp 1515870181
transform 1 0 5704 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_299
timestamp 1515870181
transform -1 0 5960 0 1 610
box 0 0 192 200
use INVX2  INVX2_20
timestamp 1515870181
transform -1 0 5992 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_260
timestamp 1515870181
transform 1 0 5992 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_27
timestamp 1515870181
transform 1 0 6056 0 1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_307
timestamp 1515870181
transform -1 0 6312 0 1 610
box 0 0 192 200
use FILL  FILL_3_5_0
timestamp 1515870181
transform 1 0 6312 0 1 610
box 0 0 16 200
use FILL  FILL_3_5_1
timestamp 1515870181
transform 1 0 6328 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_240
timestamp 1515870181
transform 1 0 6344 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_250
timestamp 1515870181
transform -1 0 6456 0 1 610
box 0 0 64 200
use INVX2  INVX2_14
timestamp 1515870181
transform -1 0 6488 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_269
timestamp 1515870181
transform -1 0 6680 0 1 610
box 0 0 192 200
use INVX2  INVX2_10
timestamp 1515870181
transform -1 0 6712 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_265
timestamp 1515870181
transform 1 0 6712 0 1 610
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_290
timestamp 1515870181
transform -1 0 7096 0 1 610
box 0 0 192 200
use NOR2X1  NOR2X1_59
timestamp 1515870181
transform 1 0 7096 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_50
timestamp 1515870181
transform -1 0 7208 0 1 610
box 0 0 64 200
use INVX2  INVX2_17
timestamp 1515870181
transform -1 0 7240 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_258
timestamp 1515870181
transform 1 0 7240 0 1 610
box 0 0 192 200
use NAND2X1  NAND2X1_225
timestamp 1515870181
transform -1 0 56 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_108
timestamp 1515870181
transform 1 0 56 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_107
timestamp 1515870181
transform -1 0 184 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_43
timestamp 1515870181
transform 1 0 184 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_102
timestamp 1515870181
transform 1 0 376 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_101
timestamp 1515870181
transform -1 0 504 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_338
timestamp 1515870181
transform -1 0 552 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_359
timestamp 1515870181
transform -1 0 600 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_83
timestamp 1515870181
transform -1 0 664 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_84
timestamp 1515870181
transform -1 0 728 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_217
timestamp 1515870181
transform 1 0 728 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_203
timestamp 1515870181
transform 1 0 920 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_217
timestamp 1515870181
transform 1 0 968 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_224
timestamp 1515870181
transform 1 0 1032 0 -1 610
box 0 0 192 200
use FILL  FILL_2_0_0
timestamp 1515870181
transform -1 0 1240 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1515870181
transform -1 0 1256 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_276
timestamp 1515870181
transform -1 0 1320 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_64
timestamp 1515870181
transform 1 0 1320 0 -1 610
box 0 0 192 200
use BUFX4  BUFX4_157
timestamp 1515870181
transform -1 0 1576 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1515870181
transform 1 0 1576 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_34
timestamp 1515870181
transform 1 0 1768 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_39
timestamp 1515870181
transform 1 0 1832 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1515870181
transform 1 0 1880 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_43
timestamp 1515870181
transform -1 0 2136 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_48
timestamp 1515870181
transform -1 0 2184 0 -1 610
box 0 0 48 200
use FILL  FILL_2_1_0
timestamp 1515870181
transform -1 0 2200 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1515870181
transform -1 0 2216 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_67
timestamp 1515870181
transform -1 0 2280 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_123
timestamp 1515870181
transform -1 0 2344 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_206
timestamp 1515870181
transform -1 0 2536 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_206
timestamp 1515870181
transform -1 0 2600 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_203
timestamp 1515870181
transform 1 0 2600 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_203
timestamp 1515870181
transform 1 0 2664 0 -1 610
box 0 0 192 200
use BUFX4  BUFX4_109
timestamp 1515870181
transform -1 0 2920 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_110
timestamp 1515870181
transform -1 0 2984 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_342
timestamp 1515870181
transform 1 0 2984 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_277
timestamp 1515870181
transform -1 0 3096 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_82
timestamp 1515870181
transform -1 0 3160 0 -1 610
box 0 0 64 200
use FILL  FILL_2_2_0
timestamp 1515870181
transform 1 0 3160 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1515870181
transform 1 0 3176 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_282
timestamp 1515870181
transform 1 0 3192 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_73
timestamp 1515870181
transform 1 0 3256 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_156
timestamp 1515870181
transform 1 0 3320 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_194
timestamp 1515870181
transform -1 0 3448 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_122
timestamp 1515870181
transform 1 0 3448 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_130
timestamp 1515870181
transform 1 0 3512 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_492
timestamp 1515870181
transform 1 0 3704 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_431
timestamp 1515870181
transform -1 0 3816 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_139
timestamp 1515870181
transform 1 0 3816 0 -1 610
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_139
timestamp 1515870181
transform 1 0 3880 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_341
timestamp 1515870181
transform -1 0 4120 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_398
timestamp 1515870181
transform -1 0 4184 0 -1 610
box 0 0 64 200
use INVX1  INVX1_76
timestamp 1515870181
transform -1 0 4216 0 -1 610
box 0 0 32 200
use FILL  FILL_2_3_0
timestamp 1515870181
transform -1 0 4232 0 -1 610
box 0 0 16 200
use FILL  FILL_2_3_1
timestamp 1515870181
transform -1 0 4248 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_111
timestamp 1515870181
transform -1 0 4312 0 -1 610
box 0 0 64 200
use INVX1  INVX1_60
timestamp 1515870181
transform 1 0 4312 0 -1 610
box 0 0 32 200
use BUFX2  BUFX2_16
timestamp 1515870181
transform 1 0 4344 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_369
timestamp 1515870181
transform -1 0 4456 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_396
timestamp 1515870181
transform 1 0 4456 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_362
timestamp 1515870181
transform 1 0 4520 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_136
timestamp 1515870181
transform 1 0 4568 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_117
timestamp 1515870181
transform -1 0 4680 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_136
timestamp 1515870181
transform 1 0 4680 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_361
timestamp 1515870181
transform 1 0 4872 0 -1 610
box 0 0 48 200
use BUFX2  BUFX2_25
timestamp 1515870181
transform 1 0 4920 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_97
timestamp 1515870181
transform 1 0 4968 0 -1 610
box 0 0 192 200
use INVX1  INVX1_9
timestamp 1515870181
transform 1 0 5160 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_498
timestamp 1515870181
transform 1 0 5192 0 -1 610
box 0 0 64 200
use FILL  FILL_2_4_0
timestamp 1515870181
transform -1 0 5272 0 -1 610
box 0 0 16 200
use FILL  FILL_2_4_1
timestamp 1515870181
transform -1 0 5288 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_437
timestamp 1515870181
transform -1 0 5336 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_326
timestamp 1515870181
transform 1 0 5336 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_439
timestamp 1515870181
transform 1 0 5384 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_107
timestamp 1515870181
transform -1 0 5624 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_508
timestamp 1515870181
transform 1 0 5624 0 -1 610
box 0 0 64 200
use INVX8  INVX8_11
timestamp 1515870181
transform 1 0 5688 0 -1 610
box 0 0 80 200
use INVX1  INVX1_74
timestamp 1515870181
transform -1 0 5800 0 -1 610
box 0 0 32 200
use NAND2X1  NAND2X1_252
timestamp 1515870181
transform 1 0 5800 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_110
timestamp 1515870181
transform -1 0 6040 0 -1 610
box 0 0 192 200
use NAND2X1  NAND2X1_246
timestamp 1515870181
transform -1 0 6088 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_244
timestamp 1515870181
transform 1 0 6088 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_511
timestamp 1515870181
transform 1 0 6136 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_450
timestamp 1515870181
transform -1 0 6248 0 -1 610
box 0 0 48 200
use FILL  FILL_2_5_0
timestamp 1515870181
transform 1 0 6248 0 -1 610
box 0 0 16 200
use FILL  FILL_2_5_1
timestamp 1515870181
transform 1 0 6264 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_236
timestamp 1515870181
transform 1 0 6280 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_258
timestamp 1515870181
transform -1 0 6392 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_227
timestamp 1515870181
transform -1 0 6456 0 -1 610
box 0 0 64 200
use INVX2  INVX2_18
timestamp 1515870181
transform -1 0 6488 0 -1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_305
timestamp 1515870181
transform -1 0 6680 0 -1 610
box 0 0 192 200
use BUFX4  BUFX4_224
timestamp 1515870181
transform 1 0 6680 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_97
timestamp 1515870181
transform 1 0 6744 0 -1 610
box 0 0 64 200
use INVX8  INVX8_14
timestamp 1515870181
transform 1 0 6808 0 -1 610
box 0 0 80 200
use INVX8  INVX8_16
timestamp 1515870181
transform -1 0 6968 0 -1 610
box 0 0 80 200
use NAND2X1  NAND2X1_243
timestamp 1515870181
transform 1 0 6968 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_243
timestamp 1515870181
transform -1 0 7080 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_257
timestamp 1515870181
transform -1 0 7144 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_257
timestamp 1515870181
transform 1 0 7144 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_272
timestamp 1515870181
transform -1 0 7384 0 -1 610
box 0 0 192 200
use BUFX2  BUFX2_3
timestamp 1515870181
transform 1 0 7384 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_237
timestamp 1515870181
transform 1 0 8 0 1 210
box 0 0 192 200
use NAND2X1  NAND2X1_224
timestamp 1515870181
transform 1 0 200 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_237
timestamp 1515870181
transform -1 0 312 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_220
timestamp 1515870181
transform -1 0 360 0 1 210
box 0 0 48 200
use INVX1  INVX1_48
timestamp 1515870181
transform 1 0 360 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_34
timestamp 1515870181
transform 1 0 392 0 1 210
box 0 0 192 200
use NAND2X1  NAND2X1_275
timestamp 1515870181
transform 1 0 584 0 1 210
box 0 0 48 200
use INVX1  INVX1_13
timestamp 1515870181
transform 1 0 632 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_285
timestamp 1515870181
transform 1 0 664 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_74
timestamp 1515870181
transform 1 0 728 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_66
timestamp 1515870181
transform -1 0 840 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_50
timestamp 1515870181
transform 1 0 840 0 1 210
box 0 0 192 200
use BUFX4  BUFX4_85
timestamp 1515870181
transform 1 0 1032 0 1 210
box 0 0 64 200
use FILL  FILL_1_0_0
timestamp 1515870181
transform 1 0 1096 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1515870181
transform 1 0 1112 0 1 210
box 0 0 16 200
use MUX2X1  MUX2X1_4
timestamp 1515870181
transform 1 0 1128 0 1 210
box 0 0 96 200
use NAND2X1  NAND2X1_56
timestamp 1515870181
transform 1 0 1224 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_73
timestamp 1515870181
transform -1 0 1464 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_57
timestamp 1515870181
transform 1 0 1464 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_63
timestamp 1515870181
transform -1 0 1576 0 1 210
box 0 0 48 200
use MUX2X1  MUX2X1_25
timestamp 1515870181
transform -1 0 1672 0 1 210
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1515870181
transform 1 0 1672 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_41
timestamp 1515870181
transform 1 0 1864 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_46
timestamp 1515870181
transform -1 0 1976 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_1
timestamp 1515870181
transform -1 0 2040 0 1 210
box 0 0 64 200
use MUX2X1  MUX2X1_26
timestamp 1515870181
transform -1 0 2136 0 1 210
box 0 0 96 200
use FILL  FILL_1_1_0
timestamp 1515870181
transform 1 0 2136 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1515870181
transform 1 0 2152 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_14
timestamp 1515870181
transform 1 0 2168 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_46
timestamp 1515870181
transform 1 0 2360 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_51
timestamp 1515870181
transform -1 0 2472 0 1 210
box 0 0 48 200
use MUX2X1  MUX2X1_41
timestamp 1515870181
transform -1 0 2568 0 1 210
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_126
timestamp 1515870181
transform 1 0 2568 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_14
timestamp 1515870181
transform 1 0 2760 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_16
timestamp 1515870181
transform -1 0 2872 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_364
timestamp 1515870181
transform -1 0 2920 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_399
timestamp 1515870181
transform 1 0 2920 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_27
timestamp 1515870181
transform -1 0 3176 0 1 210
box 0 0 192 200
use FILL  FILL_1_2_0
timestamp 1515870181
transform 1 0 3176 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1515870181
transform 1 0 3192 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_30
timestamp 1515870181
transform 1 0 3208 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_27
timestamp 1515870181
transform -1 0 3320 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_11
timestamp 1515870181
transform 1 0 3320 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_13
timestamp 1515870181
transform -1 0 3432 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_123
timestamp 1515870181
transform 1 0 3432 0 1 210
box 0 0 192 200
use NAND2X1  NAND2X1_135
timestamp 1515870181
transform -1 0 3672 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_329
timestamp 1515870181
transform -1 0 3720 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_343
timestamp 1515870181
transform 1 0 3720 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_372
timestamp 1515870181
transform -1 0 3832 0 1 210
box 0 0 64 200
use INVX1  INVX1_52
timestamp 1515870181
transform 1 0 3832 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_354
timestamp 1515870181
transform 1 0 3864 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_91
timestamp 1515870181
transform 1 0 3928 0 1 210
box 0 0 192 200
use NAND2X1  NAND2X1_363
timestamp 1515870181
transform -1 0 4168 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_30
timestamp 1515870181
transform 1 0 4168 0 1 210
box 0 0 64 200
use FILL  FILL_1_3_0
timestamp 1515870181
transform 1 0 4232 0 1 210
box 0 0 16 200
use FILL  FILL_1_3_1
timestamp 1515870181
transform 1 0 4248 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_33
timestamp 1515870181
transform 1 0 4264 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_128
timestamp 1515870181
transform 1 0 4312 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_108
timestamp 1515870181
transform -1 0 4424 0 1 210
box 0 0 48 200
use INVX1  INVX1_75
timestamp 1515870181
transform 1 0 4424 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_352
timestamp 1515870181
transform 1 0 4456 0 1 210
box 0 0 192 200
use BUFX4  BUFX4_280
timestamp 1515870181
transform 1 0 4648 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_413
timestamp 1515870181
transform -1 0 4776 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_2
timestamp 1515870181
transform 1 0 4776 0 1 210
box 0 0 48 200
use INVX1  INVX1_50
timestamp 1515870181
transform -1 0 4856 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_395
timestamp 1515870181
transform 1 0 4856 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_32
timestamp 1515870181
transform 1 0 4920 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_66
timestamp 1515870181
transform -1 0 5032 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_13
timestamp 1515870181
transform 1 0 5032 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_7
timestamp 1515870181
transform -1 0 5144 0 1 210
box 0 0 64 200
use INVX1  INVX1_19
timestamp 1515870181
transform -1 0 5176 0 1 210
box 0 0 32 200
use FILL  FILL_1_4_0
timestamp 1515870181
transform -1 0 5192 0 1 210
box 0 0 16 200
use FILL  FILL_1_4_1
timestamp 1515870181
transform -1 0 5208 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_99
timestamp 1515870181
transform -1 0 5400 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_500
timestamp 1515870181
transform -1 0 5464 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_94
timestamp 1515870181
transform -1 0 5512 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_287
timestamp 1515870181
transform 1 0 5512 0 1 210
box 0 0 64 200
use INVX1  INVX1_49
timestamp 1515870181
transform -1 0 5608 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_506
timestamp 1515870181
transform 1 0 5608 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_445
timestamp 1515870181
transform 1 0 5672 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_105
timestamp 1515870181
transform -1 0 5912 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_268
timestamp 1515870181
transform 1 0 5912 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_254
timestamp 1515870181
transform -1 0 6024 0 1 210
box 0 0 48 200
use INVX2  INVX2_28
timestamp 1515870181
transform -1 0 6056 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_315
timestamp 1515870181
transform -1 0 6248 0 1 210
box 0 0 192 200
use FILL  FILL_1_5_0
timestamp 1515870181
transform 1 0 6248 0 1 210
box 0 0 16 200
use FILL  FILL_1_5_1
timestamp 1515870181
transform 1 0 6264 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_238
timestamp 1515870181
transform 1 0 6280 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_244
timestamp 1515870181
transform 1 0 6328 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_230
timestamp 1515870181
transform -1 0 6440 0 1 210
box 0 0 48 200
use INVX2  INVX2_4
timestamp 1515870181
transform -1 0 6472 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_259
timestamp 1515870181
transform 1 0 6472 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_252
timestamp 1515870181
transform -1 0 6728 0 1 210
box 0 0 64 200
use INVX2  INVX2_12
timestamp 1515870181
transform -1 0 6760 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_267
timestamp 1515870181
transform -1 0 6952 0 1 210
box 0 0 192 200
use NAND2X1  NAND2X1_229
timestamp 1515870181
transform 1 0 6952 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_273
timestamp 1515870181
transform -1 0 7064 0 1 210
box 0 0 64 200
use INVX2  INVX2_33
timestamp 1515870181
transform -1 0 7096 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_320
timestamp 1515870181
transform -1 0 7288 0 1 210
box 0 0 192 200
use NAND2X1  NAND2X1_241
timestamp 1515870181
transform 1 0 7288 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_255
timestamp 1515870181
transform -1 0 7400 0 1 210
box 0 0 64 200
use FILL  FILL_2_1
timestamp 1515870181
transform 1 0 7400 0 1 210
box 0 0 16 200
use FILL  FILL_2_2
timestamp 1515870181
transform 1 0 7416 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_46
timestamp 1515870181
transform 1 0 8 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_233
timestamp 1515870181
transform 1 0 200 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_233
timestamp 1515870181
transform -1 0 456 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_226
timestamp 1515870181
transform -1 0 648 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_213
timestamp 1515870181
transform 1 0 648 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_226
timestamp 1515870181
transform -1 0 760 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_194
timestamp 1515870181
transform 1 0 760 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_194
timestamp 1515870181
transform 1 0 952 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_179
timestamp 1515870181
transform 1 0 1016 0 -1 210
box 0 0 48 200
use FILL  FILL_0_0_0
timestamp 1515870181
transform -1 0 1080 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1515870181
transform -1 0 1096 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_66
timestamp 1515870181
transform -1 0 1288 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_50
timestamp 1515870181
transform -1 0 1352 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_158
timestamp 1515870181
transform -1 0 1416 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_192
timestamp 1515870181
transform -1 0 1480 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_201
timestamp 1515870181
transform 1 0 1480 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_186
timestamp 1515870181
transform -1 0 1592 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_201
timestamp 1515870181
transform -1 0 1784 0 -1 210
box 0 0 192 200
use BUFX4  BUFX4_195
timestamp 1515870181
transform -1 0 1848 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_185
timestamp 1515870181
transform 1 0 1848 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_185
timestamp 1515870181
transform 1 0 1912 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_169
timestamp 1515870181
transform 1 0 2104 0 -1 210
box 0 0 48 200
use FILL  FILL_0_1_0
timestamp 1515870181
transform -1 0 2168 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1515870181
transform -1 0 2184 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_174
timestamp 1515870181
transform -1 0 2232 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_190
timestamp 1515870181
transform -1 0 2296 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_190
timestamp 1515870181
transform -1 0 2488 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_158
timestamp 1515870181
transform 1 0 2488 0 -1 210
box 0 0 192 200
use INVX1  INVX1_77
timestamp 1515870181
transform 1 0 2680 0 -1 210
box 0 0 32 200
use NAND2X1  NAND2X1_140
timestamp 1515870181
transform 1 0 2712 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_158
timestamp 1515870181
transform -1 0 2824 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_121
timestamp 1515870181
transform 1 0 2824 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_9
timestamp 1515870181
transform 1 0 3016 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_11
timestamp 1515870181
transform -1 0 3128 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_155
timestamp 1515870181
transform 1 0 3128 0 -1 210
box 0 0 64 200
use FILL  FILL_0_2_0
timestamp 1515870181
transform -1 0 3208 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1515870181
transform -1 0 3224 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_137
timestamp 1515870181
transform -1 0 3272 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_155
timestamp 1515870181
transform 1 0 3272 0 -1 210
box 0 0 192 200
use INVX1  INVX1_62
timestamp 1515870181
transform 1 0 3464 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_30
timestamp 1515870181
transform 1 0 3496 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_153
timestamp 1515870181
transform 1 0 3544 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_153
timestamp 1515870181
transform 1 0 3608 0 -1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_30
timestamp 1515870181
transform 1 0 3800 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_106
timestamp 1515870181
transform 1 0 3992 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_126
timestamp 1515870181
transform -1 0 4104 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_350
timestamp 1515870181
transform -1 0 4296 0 -1 210
box 0 0 192 200
use FILL  FILL_0_3_0
timestamp 1515870181
transform 1 0 4296 0 -1 210
box 0 0 16 200
use FILL  FILL_0_3_1
timestamp 1515870181
transform 1 0 4312 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_14
timestamp 1515870181
transform 1 0 4328 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_142
timestamp 1515870181
transform 1 0 4376 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_123
timestamp 1515870181
transform 1 0 4440 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_142
timestamp 1515870181
transform -1 0 4680 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_375
timestamp 1515870181
transform 1 0 4680 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_137
timestamp 1515870181
transform 1 0 4728 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_118
timestamp 1515870181
transform -1 0 4840 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_137
timestamp 1515870181
transform -1 0 5032 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_11
timestamp 1515870181
transform 1 0 5032 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_1
timestamp 1515870181
transform 1 0 5080 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_9
timestamp 1515870181
transform 1 0 5128 0 -1 210
box 0 0 48 200
use FILL  FILL_0_4_0
timestamp 1515870181
transform -1 0 5192 0 -1 210
box 0 0 16 200
use FILL  FILL_0_4_1
timestamp 1515870181
transform -1 0 5208 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_338
timestamp 1515870181
transform -1 0 5400 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_114
timestamp 1515870181
transform -1 0 5464 0 -1 210
box 0 0 64 200
use INVX8  INVX8_9
timestamp 1515870181
transform -1 0 5544 0 -1 210
box 0 0 80 200
use NAND2X1  NAND2X1_277
timestamp 1515870181
transform 1 0 5544 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_155
timestamp 1515870181
transform -1 0 5656 0 -1 210
box 0 0 64 200
use INVX8  INVX8_2
timestamp 1515870181
transform -1 0 5736 0 -1 210
box 0 0 80 200
use NAND2X1  NAND2X1_438
timestamp 1515870181
transform 1 0 5736 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_499
timestamp 1515870181
transform -1 0 5848 0 -1 210
box 0 0 64 200
use INVX1  INVX1_14
timestamp 1515870181
transform -1 0 5880 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_98
timestamp 1515870181
transform -1 0 6072 0 -1 210
box 0 0 192 200
use BUFX4  BUFX4_100
timestamp 1515870181
transform -1 0 6136 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_513
timestamp 1515870181
transform -1 0 6200 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_452
timestamp 1515870181
transform -1 0 6248 0 -1 210
box 0 0 48 200
use FILL  FILL_0_5_0
timestamp 1515870181
transform -1 0 6264 0 -1 210
box 0 0 16 200
use FILL  FILL_0_5_1
timestamp 1515870181
transform -1 0 6280 0 -1 210
box 0 0 16 200
use INVX1  INVX1_84
timestamp 1515870181
transform -1 0 6312 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_112
timestamp 1515870181
transform -1 0 6504 0 -1 210
box 0 0 192 200
use BUFX4  BUFX4_81
timestamp 1515870181
transform 1 0 6504 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_245
timestamp 1515870181
transform 1 0 6568 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_259
timestamp 1515870181
transform -1 0 6680 0 -1 210
box 0 0 64 200
use INVX2  INVX2_19
timestamp 1515870181
transform -1 0 6712 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_306
timestamp 1515870181
transform -1 0 6904 0 -1 210
box 0 0 192 200
use NAND2X1  NAND2X1_259
timestamp 1515870181
transform 1 0 6904 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_270
timestamp 1515870181
transform 1 0 6952 0 -1 210
box 0 0 192 200
use AOI21X1  AOI21X1_24
timestamp 1515870181
transform -1 0 7208 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_334
timestamp 1515870181
transform 1 0 7208 0 -1 210
box 0 0 192 200
use FILL  FILL_1_1
timestamp 1515870181
transform -1 0 7416 0 -1 210
box 0 0 16 200
use FILL  FILL_1_2
timestamp 1515870181
transform -1 0 7432 0 -1 210
box 0 0 16 200
<< labels >>
flabel space 1348 42 1356 136 6 FreeSans 48 0 0 0 vdd
port 0 nsew
flabel space 2388 42 2396 136 6 FreeSans 48 0 0 0 gnd
port 1 nsew
flabel metal2 5408 -40 5408 -40 7 FreeSans 48 270 0 0 REG_D<0>
port 2 nsew
flabel metal2 6576 -40 6576 -40 7 FreeSans 48 270 0 0 REG_D<1>
port 3 nsew
flabel metal2 6432 -40 6432 -40 7 FreeSans 48 270 0 0 REG_D<2>
port 4 nsew
flabel metal2 3520 5460 3520 5460 3 FreeSans 48 90 0 0 REG_D<3>
port 5 nsew
flabel metal2 6032 5460 6032 5460 3 FreeSans 48 90 0 0 REG_D<4>
port 6 nsew
flabel metal2 5328 5460 5328 5460 3 FreeSans 48 90 0 0 REG_D<5>
port 7 nsew
flabel metal2 4848 5460 4848 5460 3 FreeSans 48 90 0 0 REG_D<6>
port 8 nsew
flabel metal2 3632 5460 3632 5460 3 FreeSans 48 90 0 0 REG_D<7>
port 9 nsew
flabel metal2 5536 -40 5536 -40 7 FreeSans 48 270 0 0 REG_D<8>
port 10 nsew
flabel metal2 4688 5460 4688 5460 3 FreeSans 48 90 0 0 REG_D<9>
port 11 nsew
flabel metal2 6016 -40 6016 -40 7 FreeSans 48 270 0 0 REG_D<10>
port 12 nsew
flabel metal2 5920 5460 5920 5460 3 FreeSans 48 90 0 0 REG_D<11>
port 13 nsew
flabel metal2 6352 -40 6352 -40 7 FreeSans 48 270 0 0 REG_D<12>
port 14 nsew
flabel metal3 7488 320 7488 320 3 FreeSans 48 0 0 0 REG_D<13>
port 15 nsew
flabel metal2 4512 5460 4512 5460 3 FreeSans 48 90 0 0 REG_D<14>
port 16 nsew
flabel metal2 6272 -40 6272 -40 7 FreeSans 48 270 0 0 REG_D<15>
port 17 nsew
flabel metal2 5328 -40 5328 -40 7 FreeSans 48 270 0 0 REG_RF1<0>
port 18 nsew
flabel metal2 5360 -40 5360 -40 7 FreeSans 48 270 0 0 REG_RF1<1>
port 19 nsew
flabel metal3 7488 2700 7488 2700 3 FreeSans 48 0 0 0 REG_RF1<2>
port 20 nsew
flabel metal3 7488 2660 7488 2660 3 FreeSans 48 0 0 0 REG_RF1<3>
port 21 nsew
flabel metal2 5440 5460 5440 5460 3 FreeSans 48 90 0 0 REG_RF2<0>
port 22 nsew
flabel metal2 5376 5460 5376 5460 3 FreeSans 48 90 0 0 REG_RF2<1>
port 23 nsew
flabel metal3 7488 3520 7488 3520 3 FreeSans 48 0 0 0 REG_RF2<2>
port 24 nsew
flabel metal3 7488 3560 7488 3560 3 FreeSans 48 0 0 0 REG_RF2<3>
port 25 nsew
flabel metal3 -48 2660 -48 2660 7 FreeSans 48 0 0 0 REG_RFD<0>
port 26 nsew
flabel metal3 -48 2560 -48 2560 7 FreeSans 48 0 0 0 REG_RFD<1>
port 27 nsew
flabel metal3 -48 2520 -48 2520 7 FreeSans 48 0 0 0 REG_RFD<2>
port 28 nsew
flabel metal3 -48 2600 -48 2600 7 FreeSans 48 0 0 0 REG_RFD<3>
port 29 nsew
flabel metal3 7488 2500 7488 2500 3 FreeSans 48 0 0 0 REG_R1<0>
port 30 nsew
flabel metal3 7488 2580 7488 2580 3 FreeSans 48 0 0 0 REG_R1<1>
port 31 nsew
flabel metal3 7488 2740 7488 2740 3 FreeSans 48 0 0 0 REG_R1<2>
port 32 nsew
flabel metal3 7488 4720 7488 4720 3 FreeSans 48 0 0 0 REG_R1<3>
port 33 nsew
flabel metal3 7488 4320 7488 4320 3 FreeSans 48 0 0 0 REG_R1<4>
port 34 nsew
flabel metal3 7488 4100 7488 4100 3 FreeSans 48 0 0 0 REG_R1<5>
port 35 nsew
flabel metal3 7488 3600 7488 3600 3 FreeSans 48 0 0 0 REG_R1<6>
port 36 nsew
flabel metal2 6800 5460 6800 5460 3 FreeSans 48 90 0 0 REG_R1<7>
port 37 nsew
flabel metal3 7488 1960 7488 1960 3 FreeSans 48 0 0 0 REG_R1<8>
port 38 nsew
flabel metal3 7488 3300 7488 3300 3 FreeSans 48 0 0 0 REG_R1<9>
port 39 nsew
flabel metal3 7488 2540 7488 2540 3 FreeSans 48 0 0 0 REG_R1<10>
port 40 nsew
flabel metal3 7488 3340 7488 3340 3 FreeSans 48 0 0 0 REG_R1<11>
port 41 nsew
flabel metal3 7488 2620 7488 2620 3 FreeSans 48 0 0 0 REG_R1<12>
port 42 nsew
flabel metal3 7488 2100 7488 2100 3 FreeSans 48 0 0 0 REG_R1<13>
port 43 nsew
flabel metal3 7488 4500 7488 4500 3 FreeSans 48 0 0 0 REG_R1<14>
port 44 nsew
flabel metal3 7488 1920 7488 1920 3 FreeSans 48 0 0 0 REG_R1<15>
port 45 nsew
flabel metal3 -48 2480 -48 2480 7 FreeSans 48 0 0 0 REG_Write
port 46 nsew
flabel metal2 4656 -40 4656 -40 7 FreeSans 48 270 0 0 REG_Interrupt_flag
port 47 nsew
flabel metal2 5248 -40 5248 -40 7 FreeSans 48 270 0 0 clk
port 48 nsew
flabel space -48 120 -48 120 7 FreeSans 48 0 0 0 rst
port 49 nsew
flabel metal2 5168 -40 5168 -40 7 FreeSans 48 270 0 0 REG_A<0>
port 50 nsew
flabel metal2 4816 -40 4816 -40 7 FreeSans 48 270 0 0 REG_A<1>
port 51 nsew
flabel metal3 7488 520 7488 520 3 FreeSans 48 0 0 0 REG_A<2>
port 52 nsew
flabel metal2 3168 5460 3168 5460 3 FreeSans 48 90 0 0 REG_A<3>
port 53 nsew
flabel metal2 3136 5460 3136 5460 3 FreeSans 48 90 0 0 REG_A<4>
port 54 nsew
flabel metal2 4800 5460 4800 5460 3 FreeSans 48 90 0 0 REG_A<5>
port 55 nsew
flabel metal2 3856 5460 3856 5460 3 FreeSans 48 90 0 0 REG_A<6>
port 56 nsew
flabel metal2 4032 5460 4032 5460 3 FreeSans 48 90 0 0 REG_A<7>
port 57 nsew
flabel metal2 5280 -40 5280 -40 7 FreeSans 48 270 0 0 REG_A<8>
port 58 nsew
flabel metal2 4544 5460 4544 5460 3 FreeSans 48 90 0 0 REG_A<9>
port 59 nsew
flabel metal2 5200 -40 5200 -40 7 FreeSans 48 270 0 0 REG_A<10>
port 60 nsew
flabel metal2 4736 5460 4736 5460 3 FreeSans 48 90 0 0 REG_A<11>
port 61 nsew
flabel metal2 5120 -40 5120 -40 7 FreeSans 48 270 0 0 REG_A<12>
port 62 nsew
flabel metal2 4368 -40 4368 -40 7 FreeSans 48 270 0 0 REG_A<13>
port 63 nsew
flabel metal2 3760 5460 3760 5460 3 FreeSans 48 90 0 0 REG_A<14>
port 64 nsew
flabel metal2 4416 -40 4416 -40 7 FreeSans 48 270 0 0 REG_A<15>
port 65 nsew
flabel metal2 4928 -40 4928 -40 7 FreeSans 48 270 0 0 REG_B<0>
port 66 nsew
flabel metal2 4976 -40 4976 -40 7 FreeSans 48 270 0 0 REG_B<1>
port 67 nsew
flabel metal2 3984 5460 3984 5460 3 FreeSans 48 90 0 0 REG_B<2>
port 68 nsew
flabel metal2 3088 5460 3088 5460 3 FreeSans 48 90 0 0 REG_B<3>
port 69 nsew
flabel metal2 2896 5460 2896 5460 3 FreeSans 48 90 0 0 REG_B<4>
port 70 nsew
flabel metal2 4944 5460 4944 5460 3 FreeSans 48 90 0 0 REG_B<5>
port 71 nsew
flabel metal2 3472 5460 3472 5460 3 FreeSans 48 90 0 0 REG_B<6>
port 72 nsew
flabel metal2 4352 5460 4352 5460 3 FreeSans 48 90 0 0 REG_B<7>
port 73 nsew
flabel metal2 5008 -40 5008 -40 7 FreeSans 48 270 0 0 REG_B<8>
port 74 nsew
flabel metal2 4464 5460 4464 5460 3 FreeSans 48 90 0 0 REG_B<9>
port 75 nsew
flabel metal2 4032 -40 4032 -40 7 FreeSans 48 270 0 0 REG_B<10>
port 76 nsew
flabel metal2 3936 5460 3936 5460 3 FreeSans 48 90 0 0 REG_B<11>
port 77 nsew
flabel metal2 4864 -40 4864 -40 7 FreeSans 48 270 0 0 REG_B<12>
port 78 nsew
flabel metal2 3536 -40 3536 -40 7 FreeSans 48 270 0 0 REG_B<13>
port 79 nsew
flabel metal2 3712 5460 3712 5460 3 FreeSans 48 90 0 0 REG_B<14>
port 80 nsew
flabel metal2 5056 -40 5056 -40 7 FreeSans 48 270 0 0 REG_B<15>
port 81 nsew
<< end >>
