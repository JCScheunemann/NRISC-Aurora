module NRISC_IData ( gnd, vdd, IDATA_CORE_addr, IDATA_PROG_write, IDATA_PROG_addr, IDATA_PROG_data, clk, rst, IDATA_CORE_out);

input gnd, vdd;
input IDATA_PROG_write;
input clk;
input rst;
input [15:0] IDATA_CORE_addr;
input [9:0] IDATA_PROG_addr;
input [15:0] IDATA_PROG_data;
output [15:0] IDATA_CORE_out;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf15) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf14) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf13) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf12) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf11) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf10) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf9) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf7) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf6) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf5) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf4) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf3) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf2) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf1) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .Y(_3393__hier0_bF_buf0) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf250), .Y(clk_bF_buf250_bF_buf3) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf250), .Y(clk_bF_buf250_bF_buf2) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf250), .Y(clk_bF_buf250_bF_buf1) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf250), .Y(clk_bF_buf250_bF_buf0) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf251), .Y(clk_bF_buf251_bF_buf3) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf251), .Y(clk_bF_buf251_bF_buf2) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf251), .Y(clk_bF_buf251_bF_buf1) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf251), .Y(clk_bF_buf251_bF_buf0) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf252), .Y(clk_bF_buf252_bF_buf3) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf252), .Y(clk_bF_buf252_bF_buf2) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf252), .Y(clk_bF_buf252_bF_buf1) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf252), .Y(clk_bF_buf252_bF_buf0) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf253), .Y(clk_bF_buf253_bF_buf3) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf253), .Y(clk_bF_buf253_bF_buf2) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf253), .Y(clk_bF_buf253_bF_buf1) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf253), .Y(clk_bF_buf253_bF_buf0) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf254), .Y(clk_bF_buf254_bF_buf3) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf254), .Y(clk_bF_buf254_bF_buf2) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf254), .Y(clk_bF_buf254_bF_buf1) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf254), .Y(clk_bF_buf254_bF_buf0) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf255), .Y(clk_bF_buf255_bF_buf3) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf255), .Y(clk_bF_buf255_bF_buf2) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf255), .Y(clk_bF_buf255_bF_buf1) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf255), .Y(clk_bF_buf255_bF_buf0) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf8) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf7) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf6) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf5) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf4) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf3) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf2) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf1) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .Y(_3313__hier0_bF_buf0) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf240), .Y(clk_bF_buf240_bF_buf3) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf240), .Y(clk_bF_buf240_bF_buf2) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf240), .Y(clk_bF_buf240_bF_buf1) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf240), .Y(clk_bF_buf240_bF_buf0) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf241), .Y(clk_bF_buf241_bF_buf3) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf241), .Y(clk_bF_buf241_bF_buf2) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf241), .Y(clk_bF_buf241_bF_buf1) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf241), .Y(clk_bF_buf241_bF_buf0) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf242), .Y(clk_bF_buf242_bF_buf3) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf242), .Y(clk_bF_buf242_bF_buf2) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf242), .Y(clk_bF_buf242_bF_buf1) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf242), .Y(clk_bF_buf242_bF_buf0) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf243), .Y(clk_bF_buf243_bF_buf3) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf243), .Y(clk_bF_buf243_bF_buf2) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf243), .Y(clk_bF_buf243_bF_buf1) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf243), .Y(clk_bF_buf243_bF_buf0) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf244), .Y(clk_bF_buf244_bF_buf3) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf244), .Y(clk_bF_buf244_bF_buf2) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf244), .Y(clk_bF_buf244_bF_buf1) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf244), .Y(clk_bF_buf244_bF_buf0) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf245), .Y(clk_bF_buf245_bF_buf3) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf245), .Y(clk_bF_buf245_bF_buf2) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf245), .Y(clk_bF_buf245_bF_buf1) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf245), .Y(clk_bF_buf245_bF_buf0) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf246), .Y(clk_bF_buf246_bF_buf3) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf246), .Y(clk_bF_buf246_bF_buf2) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf246), .Y(clk_bF_buf246_bF_buf1) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf246), .Y(clk_bF_buf246_bF_buf0) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf247), .Y(clk_bF_buf247_bF_buf3) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf247), .Y(clk_bF_buf247_bF_buf2) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf247), .Y(clk_bF_buf247_bF_buf1) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf247), .Y(clk_bF_buf247_bF_buf0) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf248), .Y(clk_bF_buf248_bF_buf3) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf248), .Y(clk_bF_buf248_bF_buf2) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf248), .Y(clk_bF_buf248_bF_buf1) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf248), .Y(clk_bF_buf248_bF_buf0) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf249), .Y(clk_bF_buf249_bF_buf3) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf249), .Y(clk_bF_buf249_bF_buf2) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf249), .Y(clk_bF_buf249_bF_buf1) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(clk_bF_buf249), .Y(clk_bF_buf249_bF_buf0) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf13), .Y(_14882__bF_buf13_bF_buf3) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf13), .Y(_14882__bF_buf13_bF_buf2) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf13), .Y(_14882__bF_buf13_bF_buf1) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf13), .Y(_14882__bF_buf13_bF_buf0) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14), .Y(_14882__bF_buf14_bF_buf3) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14), .Y(_14882__bF_buf14_bF_buf2) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14), .Y(_14882__bF_buf14_bF_buf1) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14), .Y(_14882__bF_buf14_bF_buf0) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf15), .Y(_14882__bF_buf15_bF_buf3) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf15), .Y(_14882__bF_buf15_bF_buf2) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf15), .Y(_14882__bF_buf15_bF_buf1) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf15), .Y(_14882__bF_buf15_bF_buf0) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf6) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf5) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf4) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf3) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf2) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf1) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .Y(_3306__bF_buf0) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_15120_), .Y(_15120__bF_buf3) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(_15120_), .Y(_15120__bF_buf2) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(_15120_), .Y(_15120__bF_buf1) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(_15120_), .Y(_15120__bF_buf0) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .Y(_8476__bF_buf3) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .Y(_8476__bF_buf2) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .Y(_8476__bF_buf1) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(_8476_), .Y(_8476__bF_buf0) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(_8820_), .Y(_8820__bF_buf3) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(_8820_), .Y(_8820__bF_buf2) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(_8820_), .Y(_8820__bF_buf1) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(_8820_), .Y(_8820__bF_buf0) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(_15575_), .Y(_15575__bF_buf3) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(_15575_), .Y(_15575__bF_buf2) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(_15575_), .Y(_15575__bF_buf1) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(_15575_), .Y(_15575__bF_buf0) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf3) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf2) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf1) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .Y(_2497__bF_buf0) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .Y(_3952__bF_buf3) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .Y(_3952__bF_buf2) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .Y(_3952__bF_buf1) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .Y(_3952__bF_buf0) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_14978_), .Y(_14978__bF_buf4) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_14978_), .Y(_14978__bF_buf3) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(_14978_), .Y(_14978__bF_buf2) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(_14978_), .Y(_14978__bF_buf1) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(_14978_), .Y(_14978__bF_buf0) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf13) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf12) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf11) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf10) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf9) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf8) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf7) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf6) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf5) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf4) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf3) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf2) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf1) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(_14902_), .Y(_14902__bF_buf0) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .Y(_2418__bF_buf3) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .Y(_2418__bF_buf2) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .Y(_2418__bF_buf1) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .Y(_2418__bF_buf0) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_8279_), .Y(_8279__bF_buf3) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_8279_), .Y(_8279__bF_buf2) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_8279_), .Y(_8279__bF_buf1) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_8279_), .Y(_8279__bF_buf0) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf13) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf12) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf11) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf10) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf9) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf8) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf7) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf6) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf5) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf4) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf3) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf2) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf1) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_15055_), .Y(_15055__bF_buf0) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[14]), .Y(IDATA_PROG_data_14_bF_buf4) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[14]), .Y(IDATA_PROG_data_14_bF_buf3) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[14]), .Y(IDATA_PROG_data_14_bF_buf2) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[14]), .Y(IDATA_PROG_data_14_bF_buf1) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[14]), .Y(IDATA_PROG_data_14_bF_buf0) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[8]), .Y(IDATA_PROG_data_8_bF_buf4) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[8]), .Y(IDATA_PROG_data_8_bF_buf3) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[8]), .Y(IDATA_PROG_data_8_bF_buf2) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[8]), .Y(IDATA_PROG_data_8_bF_buf1) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[8]), .Y(IDATA_PROG_data_8_bF_buf0) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf13) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf12) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf11) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf10) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf9) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf8) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf7) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf6) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf5) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf4) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf3) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf2) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf1) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(_15052_), .Y(_15052__bF_buf0) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(_7259_), .Y(_7259__bF_buf3) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(_7259_), .Y(_7259__bF_buf2) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(_7259_), .Y(_7259__bF_buf1) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(_7259_), .Y(_7259__bF_buf0) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf14) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf13) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf12) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf11) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf10) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf9) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf8) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf7) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf6) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf5) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf4) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf3) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf2) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf1) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_15049_), .Y(_15049__bF_buf0) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .Y(_6912__bF_buf3) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .Y(_6912__bF_buf2) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .Y(_6912__bF_buf1) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(_6912_), .Y(_6912__bF_buf0) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[11]), .Y(IDATA_PROG_data_11_bF_buf4) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[11]), .Y(IDATA_PROG_data_11_bF_buf3) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[11]), .Y(IDATA_PROG_data_11_bF_buf2) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[11]), .Y(IDATA_PROG_data_11_bF_buf1) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[11]), .Y(IDATA_PROG_data_11_bF_buf0) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[5]), .Y(IDATA_PROG_data_5_bF_buf4) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[5]), .Y(IDATA_PROG_data_5_bF_buf3) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[5]), .Y(IDATA_PROG_data_5_bF_buf2) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[5]), .Y(IDATA_PROG_data_5_bF_buf1) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[5]), .Y(IDATA_PROG_data_5_bF_buf0) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(_15011_), .Y(_15011__bF_buf3) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(_15011_), .Y(_15011__bF_buf2) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(_15011_), .Y(_15011__bF_buf1) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(_15011_), .Y(_15011__bF_buf0) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf8) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf7) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf6) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf5) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf4) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf3) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf2) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf1) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write), .Y(IDATA_PROG_write_bF_buf0) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .Y(_1815__bF_buf3) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .Y(_1815__bF_buf2) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .Y(_1815__bF_buf1) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .Y(_1815__bF_buf0) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .Y(_2065__bF_buf3) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .Y(_2065__bF_buf2) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .Y(_2065__bF_buf1) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .Y(_2065__bF_buf0) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .Y(_4763__bF_buf3) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .Y(_4763__bF_buf2) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .Y(_4763__bF_buf1) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_4763_), .Y(_4763__bF_buf0) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[2]), .Y(IDATA_PROG_data_2_bF_buf3) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[2]), .Y(IDATA_PROG_data_2_bF_buf2) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[2]), .Y(IDATA_PROG_data_2_bF_buf1) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[2]), .Y(IDATA_PROG_data_2_bF_buf0) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(_8364_), .Y(_8364__bF_buf3) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(_8364_), .Y(_8364__bF_buf2) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(_8364_), .Y(_8364__bF_buf1) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(_8364_), .Y(_8364__bF_buf0) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(_1812_), .Y(_1812__bF_buf3) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(_1812_), .Y(_1812__bF_buf2) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_1812_), .Y(_1812__bF_buf1) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_1812_), .Y(_1812__bF_buf0) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf255) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf254) );
BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf253) );
BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf252) );
BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf251) );
BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf250) );
BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf249) );
BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf248) );
BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf247) );
BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf246) );
BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf245) );
BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf244) );
BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf243) );
BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf242) );
BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf241) );
BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf240) );
BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf239) );
BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf238) );
BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf237) );
BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf236) );
BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf235) );
BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf234) );
BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf233) );
BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf232) );
BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf231) );
BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf230) );
BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf229) );
BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf228) );
BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf227) );
BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf226) );
BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf225) );
BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf224) );
BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf223) );
BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf222) );
BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf221) );
BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf220) );
BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf219) );
BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf218) );
BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf217) );
BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf216) );
BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf215) );
BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf214) );
BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf213) );
BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf212) );
BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf211) );
BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf210) );
BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf209) );
BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf208) );
BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf207) );
BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf206) );
BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf205) );
BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf204) );
BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf203) );
BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf202) );
BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf201) );
BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf200) );
BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf199) );
BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf198) );
BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf197) );
BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf196) );
BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf195) );
BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf194) );
BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf193) );
BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf192) );
BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf191) );
BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf190) );
BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf189) );
BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf188) );
BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf187) );
BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf186) );
BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf185) );
BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf184) );
BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf183) );
BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf182) );
BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf181) );
BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf180) );
BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf179) );
BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf178) );
BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf177) );
BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf176) );
BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf175) );
BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf174) );
BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf173) );
BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf172) );
BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf171) );
BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf170) );
BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf169) );
BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf168) );
BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf167) );
BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf166) );
BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf165) );
BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf164) );
BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf163) );
BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf162) );
BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf161) );
BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf160) );
BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf159) );
BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf158) );
BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf157) );
BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf156) );
BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf155) );
BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf154) );
BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf153) );
BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf152) );
BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf151) );
BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf150) );
BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf149) );
BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf148) );
BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf147) );
BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf146) );
BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf145) );
BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf144) );
BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf143) );
BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf142) );
BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf141) );
BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf140) );
BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf139) );
BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf138) );
BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf137) );
BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf136) );
BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf135) );
BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf134) );
BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf133) );
BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf132) );
BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf131) );
BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf130) );
BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf129) );
BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf128) );
BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf127) );
BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf126) );
BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf125) );
BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf124) );
BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf123) );
BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf122) );
BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf121) );
BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf120) );
BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf119) );
BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf118) );
BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf117) );
BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf116) );
BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf115) );
BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf114) );
BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf113) );
BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf112) );
BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf111) );
BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf110) );
BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf109) );
BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf108) );
BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf107) );
BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf106) );
BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf105) );
BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf104) );
BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf103) );
BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf102) );
BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf101) );
BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf100) );
BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf99) );
BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf98) );
BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf97) );
BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf96) );
BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf95) );
BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf94) );
BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf93) );
BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf92) );
BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf91) );
BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf90) );
BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf89) );
BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf88) );
BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf87) );
BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf86) );
BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf85) );
BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf84) );
BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf83) );
BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf82) );
BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf81) );
BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf80) );
BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf79) );
BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf78) );
BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf77) );
BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf76) );
BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf75) );
BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf74) );
BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf73) );
BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf72) );
BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf71) );
BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf70) );
BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf69) );
BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf68) );
BUFX4 BUFX4_464 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf67) );
BUFX4 BUFX4_465 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf66) );
BUFX4 BUFX4_466 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf65) );
BUFX4 BUFX4_467 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf64) );
BUFX4 BUFX4_468 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf63) );
BUFX4 BUFX4_469 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf62) );
BUFX4 BUFX4_470 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf61) );
BUFX4 BUFX4_471 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf60) );
BUFX4 BUFX4_472 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf59) );
BUFX4 BUFX4_473 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf58) );
BUFX4 BUFX4_474 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf57) );
BUFX4 BUFX4_475 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf56) );
BUFX4 BUFX4_476 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf55) );
BUFX4 BUFX4_477 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf54) );
BUFX4 BUFX4_478 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf53) );
BUFX4 BUFX4_479 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf52) );
BUFX4 BUFX4_480 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf51) );
BUFX4 BUFX4_481 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf50) );
BUFX4 BUFX4_482 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf49) );
BUFX4 BUFX4_483 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf48) );
BUFX4 BUFX4_484 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf47) );
BUFX4 BUFX4_485 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf46) );
BUFX4 BUFX4_486 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf45) );
BUFX4 BUFX4_487 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf44) );
BUFX4 BUFX4_488 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf43) );
BUFX4 BUFX4_489 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf42) );
BUFX4 BUFX4_490 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf41) );
BUFX4 BUFX4_491 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf40) );
BUFX4 BUFX4_492 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf39) );
BUFX4 BUFX4_493 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf38) );
BUFX4 BUFX4_494 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf37) );
BUFX4 BUFX4_495 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf36) );
BUFX4 BUFX4_496 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf35) );
BUFX4 BUFX4_497 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf34) );
BUFX4 BUFX4_498 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf33) );
BUFX4 BUFX4_499 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf32) );
BUFX4 BUFX4_500 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf31) );
BUFX4 BUFX4_501 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf30) );
BUFX4 BUFX4_502 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf29) );
BUFX4 BUFX4_503 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf28) );
BUFX4 BUFX4_504 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf27) );
BUFX4 BUFX4_505 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf26) );
BUFX4 BUFX4_506 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf25) );
BUFX4 BUFX4_507 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf24) );
BUFX4 BUFX4_508 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf23) );
BUFX4 BUFX4_509 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf22) );
BUFX4 BUFX4_510 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf21) );
BUFX4 BUFX4_511 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf20) );
BUFX4 BUFX4_512 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf19) );
BUFX4 BUFX4_513 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf18) );
BUFX4 BUFX4_514 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf17) );
BUFX4 BUFX4_515 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf16) );
BUFX4 BUFX4_516 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf15), .Y(clk_bF_buf15) );
BUFX4 BUFX4_517 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf14), .Y(clk_bF_buf14) );
BUFX4 BUFX4_518 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf13), .Y(clk_bF_buf13) );
BUFX4 BUFX4_519 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf12), .Y(clk_bF_buf12) );
BUFX4 BUFX4_520 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf11), .Y(clk_bF_buf11) );
BUFX4 BUFX4_521 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf10), .Y(clk_bF_buf10) );
BUFX4 BUFX4_522 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf9), .Y(clk_bF_buf9) );
BUFX4 BUFX4_523 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf8) );
BUFX4 BUFX4_524 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf7) );
BUFX4 BUFX4_525 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf6) );
BUFX4 BUFX4_526 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf5) );
BUFX4 BUFX4_527 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf4) );
BUFX4 BUFX4_528 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf3) );
BUFX4 BUFX4_529 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf2) );
BUFX4 BUFX4_530 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf1) );
BUFX4 BUFX4_531 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf0) );
BUFX4 BUFX4_532 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf9) );
BUFX4 BUFX4_533 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf8) );
BUFX4 BUFX4_534 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf7) );
BUFX4 BUFX4_535 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf6) );
BUFX4 BUFX4_536 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf5) );
BUFX4 BUFX4_537 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf4) );
BUFX4 BUFX4_538 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf3) );
BUFX4 BUFX4_539 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf2) );
BUFX4 BUFX4_540 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf1) );
BUFX4 BUFX4_541 ( .gnd(gnd), .vdd(vdd), .A(_7118_), .Y(_7118__bF_buf0) );
BUFX4 BUFX4_542 ( .gnd(gnd), .vdd(vdd), .A(_15005_), .Y(_15005__bF_buf3) );
BUFX4 BUFX4_543 ( .gnd(gnd), .vdd(vdd), .A(_15005_), .Y(_15005__bF_buf2) );
BUFX4 BUFX4_544 ( .gnd(gnd), .vdd(vdd), .A(_15005_), .Y(_15005__bF_buf1) );
BUFX4 BUFX4_545 ( .gnd(gnd), .vdd(vdd), .A(_15005_), .Y(_15005__bF_buf0) );
BUFX4 BUFX4_546 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf7) );
BUFX4 BUFX4_547 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf6) );
BUFX4 BUFX4_548 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf5) );
BUFX4 BUFX4_549 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf4) );
BUFX4 BUFX4_550 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf3) );
BUFX4 BUFX4_551 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf2) );
BUFX4 BUFX4_552 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf1) );
BUFX4 BUFX4_553 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2958__bF_buf0) );
BUFX4 BUFX4_554 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .Y(_1562__bF_buf3) );
BUFX4 BUFX4_555 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .Y(_1562__bF_buf2) );
BUFX4 BUFX4_556 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .Y(_1562__bF_buf1) );
BUFX4 BUFX4_557 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .Y(_1562__bF_buf0) );
BUFX4 BUFX4_558 ( .gnd(gnd), .vdd(vdd), .A(_893_), .Y(_893__bF_buf3) );
BUFX4 BUFX4_559 ( .gnd(gnd), .vdd(vdd), .A(_893_), .Y(_893__bF_buf2) );
BUFX4 BUFX4_560 ( .gnd(gnd), .vdd(vdd), .A(_893_), .Y(_893__bF_buf1) );
BUFX4 BUFX4_561 ( .gnd(gnd), .vdd(vdd), .A(_893_), .Y(_893__bF_buf0) );
BUFX4 BUFX4_562 ( .gnd(gnd), .vdd(vdd), .A(_14963_), .Y(_14963__bF_buf3) );
BUFX4 BUFX4_563 ( .gnd(gnd), .vdd(vdd), .A(_14963_), .Y(_14963__bF_buf2) );
BUFX4 BUFX4_564 ( .gnd(gnd), .vdd(vdd), .A(_14963_), .Y(_14963__bF_buf1) );
BUFX4 BUFX4_565 ( .gnd(gnd), .vdd(vdd), .A(_14963_), .Y(_14963__bF_buf0) );
BUFX4 BUFX4_566 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .Y(_5354__bF_buf3) );
BUFX4 BUFX4_567 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .Y(_5354__bF_buf2) );
BUFX4 BUFX4_568 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .Y(_5354__bF_buf1) );
BUFX4 BUFX4_569 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .Y(_5354__bF_buf0) );
BUFX4 BUFX4_570 ( .gnd(gnd), .vdd(vdd), .A(_1694_), .Y(_1694__bF_buf3) );
BUFX4 BUFX4_571 ( .gnd(gnd), .vdd(vdd), .A(_1694_), .Y(_1694__bF_buf2) );
BUFX4 BUFX4_572 ( .gnd(gnd), .vdd(vdd), .A(_1694_), .Y(_1694__bF_buf1) );
BUFX4 BUFX4_573 ( .gnd(gnd), .vdd(vdd), .A(_1694_), .Y(_1694__bF_buf0) );
BUFX4 BUFX4_574 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .Y(_15175__bF_buf4) );
BUFX4 BUFX4_575 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .Y(_15175__bF_buf3) );
BUFX4 BUFX4_576 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .Y(_15175__bF_buf2) );
BUFX4 BUFX4_577 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .Y(_15175__bF_buf1) );
BUFX4 BUFX4_578 ( .gnd(gnd), .vdd(vdd), .A(_15175_), .Y(_15175__bF_buf0) );
BUFX4 BUFX4_579 ( .gnd(gnd), .vdd(vdd), .A(_14998_), .Y(_14998__bF_buf3) );
BUFX4 BUFX4_580 ( .gnd(gnd), .vdd(vdd), .A(_14998_), .Y(_14998__bF_buf2) );
BUFX4 BUFX4_581 ( .gnd(gnd), .vdd(vdd), .A(_14998_), .Y(_14998__bF_buf1) );
BUFX4 BUFX4_582 ( .gnd(gnd), .vdd(vdd), .A(_14998_), .Y(_14998__bF_buf0) );
BUFX4 BUFX4_583 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .Y(_2573__bF_buf3) );
BUFX4 BUFX4_584 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .Y(_2573__bF_buf2) );
BUFX4 BUFX4_585 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .Y(_2573__bF_buf1) );
BUFX4 BUFX4_586 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .Y(_2573__bF_buf0) );
BUFX4 BUFX4_587 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .Y(_15457__bF_buf3) );
BUFX4 BUFX4_588 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .Y(_15457__bF_buf2) );
BUFX4 BUFX4_589 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .Y(_15457__bF_buf1) );
BUFX4 BUFX4_590 ( .gnd(gnd), .vdd(vdd), .A(_15457_), .Y(_15457__bF_buf0) );
BUFX4 BUFX4_591 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .Y(_5025__bF_buf3) );
BUFX4 BUFX4_592 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .Y(_5025__bF_buf2) );
BUFX4 BUFX4_593 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .Y(_5025__bF_buf1) );
BUFX4 BUFX4_594 ( .gnd(gnd), .vdd(vdd), .A(_5025_), .Y(_5025__bF_buf0) );
BUFX4 BUFX4_595 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .Y(_2532__bF_buf3) );
BUFX4 BUFX4_596 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .Y(_2532__bF_buf2) );
BUFX4 BUFX4_597 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .Y(_2532__bF_buf1) );
BUFX4 BUFX4_598 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .Y(_2532__bF_buf0) );
BUFX4 BUFX4_599 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf69) );
BUFX4 BUFX4_600 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf68) );
BUFX4 BUFX4_601 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf67) );
BUFX4 BUFX4_602 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf66) );
BUFX4 BUFX4_603 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf65) );
BUFX4 BUFX4_604 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf64) );
BUFX4 BUFX4_605 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf63) );
BUFX4 BUFX4_606 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf62) );
BUFX4 BUFX4_607 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf61) );
BUFX4 BUFX4_608 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf60) );
BUFX4 BUFX4_609 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf59) );
BUFX4 BUFX4_610 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf58) );
BUFX4 BUFX4_611 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf57) );
BUFX4 BUFX4_612 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf56) );
BUFX4 BUFX4_613 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf55) );
BUFX4 BUFX4_614 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf54) );
BUFX4 BUFX4_615 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf53) );
BUFX4 BUFX4_616 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf52) );
BUFX4 BUFX4_617 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf51) );
BUFX4 BUFX4_618 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf50) );
BUFX4 BUFX4_619 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf49) );
BUFX4 BUFX4_620 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf48) );
BUFX4 BUFX4_621 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf47) );
BUFX4 BUFX4_622 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf46) );
BUFX4 BUFX4_623 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf45) );
BUFX4 BUFX4_624 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf44) );
BUFX4 BUFX4_625 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf43) );
BUFX4 BUFX4_626 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf42) );
BUFX4 BUFX4_627 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf41) );
BUFX4 BUFX4_628 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf40) );
BUFX4 BUFX4_629 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf39) );
BUFX4 BUFX4_630 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf38) );
BUFX4 BUFX4_631 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf37) );
BUFX4 BUFX4_632 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf36) );
BUFX4 BUFX4_633 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf35) );
BUFX4 BUFX4_634 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf34) );
BUFX4 BUFX4_635 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf33) );
BUFX4 BUFX4_636 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf32) );
BUFX4 BUFX4_637 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf31) );
BUFX4 BUFX4_638 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf30) );
BUFX4 BUFX4_639 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf29) );
BUFX4 BUFX4_640 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf28) );
BUFX4 BUFX4_641 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf27) );
BUFX4 BUFX4_642 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf26) );
BUFX4 BUFX4_643 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf25) );
BUFX4 BUFX4_644 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf24) );
BUFX4 BUFX4_645 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf23) );
BUFX4 BUFX4_646 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf22) );
BUFX4 BUFX4_647 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf21) );
BUFX4 BUFX4_648 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf20) );
BUFX4 BUFX4_649 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf19) );
BUFX4 BUFX4_650 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf18) );
BUFX4 BUFX4_651 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf17) );
BUFX4 BUFX4_652 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf16) );
BUFX4 BUFX4_653 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf15) );
BUFX4 BUFX4_654 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf14) );
BUFX4 BUFX4_655 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf13) );
BUFX4 BUFX4_656 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf12) );
BUFX4 BUFX4_657 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf11) );
BUFX4 BUFX4_658 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf10) );
BUFX4 BUFX4_659 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf9) );
BUFX4 BUFX4_660 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf8) );
BUFX4 BUFX4_661 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf1), .Y(_3393__bF_buf7) );
BUFX4 BUFX4_662 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf0), .Y(_3393__bF_buf6) );
BUFX4 BUFX4_663 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf7), .Y(_3393__bF_buf5) );
BUFX4 BUFX4_664 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf6), .Y(_3393__bF_buf4) );
BUFX4 BUFX4_665 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf5), .Y(_3393__bF_buf3) );
BUFX4 BUFX4_666 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf4), .Y(_3393__bF_buf2) );
BUFX4 BUFX4_667 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf3), .Y(_3393__bF_buf1) );
BUFX4 BUFX4_668 ( .gnd(gnd), .vdd(vdd), .A(_3393__hier0_bF_buf2), .Y(_3393__bF_buf0) );
BUFX4 BUFX4_669 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .Y(_1036__bF_buf3) );
BUFX4 BUFX4_670 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .Y(_1036__bF_buf2) );
BUFX4 BUFX4_671 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .Y(_1036__bF_buf1) );
BUFX4 BUFX4_672 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .Y(_1036__bF_buf0) );
BUFX4 BUFX4_673 ( .gnd(gnd), .vdd(vdd), .A(_14895_), .Y(_14895__bF_buf3) );
BUFX4 BUFX4_674 ( .gnd(gnd), .vdd(vdd), .A(_14895_), .Y(_14895__bF_buf2) );
BUFX4 BUFX4_675 ( .gnd(gnd), .vdd(vdd), .A(_14895_), .Y(_14895__bF_buf1) );
BUFX4 BUFX4_676 ( .gnd(gnd), .vdd(vdd), .A(_14895_), .Y(_14895__bF_buf0) );
BUFX4 BUFX4_677 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf14) );
BUFX4 BUFX4_678 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf13) );
BUFX4 BUFX4_679 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf12) );
BUFX4 BUFX4_680 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf11) );
BUFX4 BUFX4_681 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf10) );
BUFX4 BUFX4_682 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf9) );
BUFX4 BUFX4_683 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf8) );
BUFX4 BUFX4_684 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf7) );
BUFX4 BUFX4_685 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf6) );
BUFX4 BUFX4_686 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf5) );
BUFX4 BUFX4_687 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf4) );
BUFX4 BUFX4_688 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf3) );
BUFX4 BUFX4_689 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf2) );
BUFX4 BUFX4_690 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf1) );
BUFX4 BUFX4_691 ( .gnd(gnd), .vdd(vdd), .A(_14913_), .Y(_14913__bF_buf0) );
BUFX4 BUFX4_692 ( .gnd(gnd), .vdd(vdd), .A(_15031_), .Y(_15031__bF_buf3) );
BUFX4 BUFX4_693 ( .gnd(gnd), .vdd(vdd), .A(_15031_), .Y(_15031__bF_buf2) );
BUFX4 BUFX4_694 ( .gnd(gnd), .vdd(vdd), .A(_15031_), .Y(_15031__bF_buf1) );
BUFX4 BUFX4_695 ( .gnd(gnd), .vdd(vdd), .A(_15031_), .Y(_15031__bF_buf0) );
BUFX4 BUFX4_696 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf6) );
BUFX4 BUFX4_697 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf5) );
BUFX4 BUFX4_698 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf4) );
BUFX4 BUFX4_699 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf3) );
BUFX4 BUFX4_700 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf2) );
BUFX4 BUFX4_701 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf1) );
BUFX4 BUFX4_702 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .Y(_2984__bF_buf0) );
BUFX4 BUFX4_703 ( .gnd(gnd), .vdd(vdd), .A(_15066_), .Y(_15066__bF_buf3) );
BUFX4 BUFX4_704 ( .gnd(gnd), .vdd(vdd), .A(_15066_), .Y(_15066__bF_buf2) );
BUFX4 BUFX4_705 ( .gnd(gnd), .vdd(vdd), .A(_15066_), .Y(_15066__bF_buf1) );
BUFX4 BUFX4_706 ( .gnd(gnd), .vdd(vdd), .A(_15066_), .Y(_15066__bF_buf0) );
BUFX4 BUFX4_707 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .Y(_7655__bF_buf3) );
BUFX4 BUFX4_708 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .Y(_7655__bF_buf2) );
BUFX4 BUFX4_709 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .Y(_7655__bF_buf1) );
BUFX4 BUFX4_710 ( .gnd(gnd), .vdd(vdd), .A(_7655_), .Y(_7655__bF_buf0) );
BUFX4 BUFX4_711 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_361__bF_buf5) );
BUFX4 BUFX4_712 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_361__bF_buf4) );
BUFX4 BUFX4_713 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_361__bF_buf3) );
BUFX4 BUFX4_714 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_361__bF_buf2) );
BUFX4 BUFX4_715 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_361__bF_buf1) );
BUFX4 BUFX4_716 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_361__bF_buf0) );
BUFX4 BUFX4_717 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .Y(_15025__bF_buf4) );
BUFX4 BUFX4_718 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .Y(_15025__bF_buf3) );
BUFX4 BUFX4_719 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .Y(_15025__bF_buf2) );
BUFX4 BUFX4_720 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .Y(_15025__bF_buf1) );
BUFX4 BUFX4_721 ( .gnd(gnd), .vdd(vdd), .A(_15025_), .Y(_15025__bF_buf0) );
BUFX4 BUFX4_722 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .Y(_14886__bF_buf3) );
BUFX4 BUFX4_723 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .Y(_14886__bF_buf2) );
BUFX4 BUFX4_724 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .Y(_14886__bF_buf1) );
BUFX4 BUFX4_725 ( .gnd(gnd), .vdd(vdd), .A(_14886_), .Y(_14886__bF_buf0) );
BUFX4 BUFX4_726 ( .gnd(gnd), .vdd(vdd), .A(_6388_), .Y(_6388__bF_buf3) );
BUFX4 BUFX4_727 ( .gnd(gnd), .vdd(vdd), .A(_6388_), .Y(_6388__bF_buf2) );
BUFX4 BUFX4_728 ( .gnd(gnd), .vdd(vdd), .A(_6388_), .Y(_6388__bF_buf1) );
BUFX4 BUFX4_729 ( .gnd(gnd), .vdd(vdd), .A(_6388_), .Y(_6388__bF_buf0) );
BUFX4 BUFX4_730 ( .gnd(gnd), .vdd(vdd), .A(_14942_), .Y(_14942__bF_buf3) );
BUFX4 BUFX4_731 ( .gnd(gnd), .vdd(vdd), .A(_14942_), .Y(_14942__bF_buf2) );
BUFX4 BUFX4_732 ( .gnd(gnd), .vdd(vdd), .A(_14942_), .Y(_14942__bF_buf1) );
BUFX4 BUFX4_733 ( .gnd(gnd), .vdd(vdd), .A(_14942_), .Y(_14942__bF_buf0) );
BUFX4 BUFX4_734 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .Y(_3989__bF_buf4) );
BUFX4 BUFX4_735 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .Y(_3989__bF_buf3) );
BUFX4 BUFX4_736 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .Y(_3989__bF_buf2) );
BUFX4 BUFX4_737 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .Y(_3989__bF_buf1) );
BUFX4 BUFX4_738 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .Y(_3989__bF_buf0) );
BUFX4 BUFX4_739 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf14) );
BUFX4 BUFX4_740 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf13) );
BUFX4 BUFX4_741 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf12) );
BUFX4 BUFX4_742 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf11) );
BUFX4 BUFX4_743 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf10) );
BUFX4 BUFX4_744 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf9) );
BUFX4 BUFX4_745 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf8) );
BUFX4 BUFX4_746 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf7) );
BUFX4 BUFX4_747 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf6) );
BUFX4 BUFX4_748 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf5) );
BUFX4 BUFX4_749 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf4) );
BUFX4 BUFX4_750 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf3) );
BUFX4 BUFX4_751 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf2) );
BUFX4 BUFX4_752 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf1) );
BUFX4 BUFX4_753 ( .gnd(gnd), .vdd(vdd), .A(_15060_), .Y(_15060__bF_buf0) );
BUFX4 BUFX4_754 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .Y(_5944__bF_buf3) );
BUFX4 BUFX4_755 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .Y(_5944__bF_buf2) );
BUFX4 BUFX4_756 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .Y(_5944__bF_buf1) );
BUFX4 BUFX4_757 ( .gnd(gnd), .vdd(vdd), .A(_5944_), .Y(_5944__bF_buf0) );
BUFX4 BUFX4_758 ( .gnd(gnd), .vdd(vdd), .A(_15019_), .Y(_15019__bF_buf3) );
BUFX4 BUFX4_759 ( .gnd(gnd), .vdd(vdd), .A(_15019_), .Y(_15019__bF_buf2) );
BUFX4 BUFX4_760 ( .gnd(gnd), .vdd(vdd), .A(_15019_), .Y(_15019__bF_buf1) );
BUFX4 BUFX4_761 ( .gnd(gnd), .vdd(vdd), .A(_15019_), .Y(_15019__bF_buf0) );
BUFX4 BUFX4_762 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf7) );
BUFX4 BUFX4_763 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf6) );
BUFX4 BUFX4_764 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf5) );
BUFX4 BUFX4_765 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf4) );
BUFX4 BUFX4_766 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf3) );
BUFX4 BUFX4_767 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf2) );
BUFX4 BUFX4_768 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf1) );
BUFX4 BUFX4_769 ( .gnd(gnd), .vdd(vdd), .A(_678_), .Y(_678__bF_buf0) );
BUFX4 BUFX4_770 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .Y(_14977__bF_buf3) );
BUFX4 BUFX4_771 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .Y(_14977__bF_buf2) );
BUFX4 BUFX4_772 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .Y(_14977__bF_buf1) );
BUFX4 BUFX4_773 ( .gnd(gnd), .vdd(vdd), .A(_14977_), .Y(_14977__bF_buf0) );
BUFX4 BUFX4_774 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf3) );
BUFX4 BUFX4_775 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf2) );
BUFX4 BUFX4_776 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf1) );
BUFX4 BUFX4_777 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .Y(_2552__bF_buf0) );
BUFX4 BUFX4_778 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .Y(_7167__bF_buf3) );
BUFX4 BUFX4_779 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .Y(_7167__bF_buf2) );
BUFX4 BUFX4_780 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .Y(_7167__bF_buf1) );
BUFX4 BUFX4_781 ( .gnd(gnd), .vdd(vdd), .A(_7167_), .Y(_7167__bF_buf0) );
BUFX4 BUFX4_782 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .Y(_14936__bF_buf3) );
BUFX4 BUFX4_783 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .Y(_14936__bF_buf2) );
BUFX4 BUFX4_784 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .Y(_14936__bF_buf1) );
BUFX4 BUFX4_785 ( .gnd(gnd), .vdd(vdd), .A(_14936_), .Y(_14936__bF_buf0) );
BUFX4 BUFX4_786 ( .gnd(gnd), .vdd(vdd), .A(_5459_), .Y(_5459__bF_buf3) );
BUFX4 BUFX4_787 ( .gnd(gnd), .vdd(vdd), .A(_5459_), .Y(_5459__bF_buf2) );
BUFX4 BUFX4_788 ( .gnd(gnd), .vdd(vdd), .A(_5459_), .Y(_5459__bF_buf1) );
BUFX4 BUFX4_789 ( .gnd(gnd), .vdd(vdd), .A(_5459_), .Y(_5459__bF_buf0) );
BUFX4 BUFX4_790 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[13]), .Y(IDATA_PROG_data_13_bF_buf4) );
BUFX4 BUFX4_791 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[13]), .Y(IDATA_PROG_data_13_bF_buf3) );
BUFX4 BUFX4_792 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[13]), .Y(IDATA_PROG_data_13_bF_buf2) );
BUFX4 BUFX4_793 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[13]), .Y(IDATA_PROG_data_13_bF_buf1) );
BUFX4 BUFX4_794 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[13]), .Y(IDATA_PROG_data_13_bF_buf0) );
BUFX4 BUFX4_795 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[7]), .Y(IDATA_PROG_data_7_bF_buf5) );
BUFX4 BUFX4_796 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[7]), .Y(IDATA_PROG_data_7_bF_buf4) );
BUFX4 BUFX4_797 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[7]), .Y(IDATA_PROG_data_7_bF_buf3) );
BUFX4 BUFX4_798 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[7]), .Y(IDATA_PROG_data_7_bF_buf2) );
BUFX4 BUFX4_799 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[7]), .Y(IDATA_PROG_data_7_bF_buf1) );
BUFX4 BUFX4_800 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[7]), .Y(IDATA_PROG_data_7_bF_buf0) );
BUFX4 BUFX4_801 ( .gnd(gnd), .vdd(vdd), .A(_995_), .Y(_995__bF_buf3) );
BUFX4 BUFX4_802 ( .gnd(gnd), .vdd(vdd), .A(_995_), .Y(_995__bF_buf2) );
BUFX4 BUFX4_803 ( .gnd(gnd), .vdd(vdd), .A(_995_), .Y(_995__bF_buf1) );
BUFX4 BUFX4_804 ( .gnd(gnd), .vdd(vdd), .A(_995_), .Y(_995__bF_buf0) );
BUFX4 BUFX4_805 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf8) );
BUFX4 BUFX4_806 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf7) );
BUFX4 BUFX4_807 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf6) );
BUFX4 BUFX4_808 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf5) );
BUFX4 BUFX4_809 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf4) );
BUFX4 BUFX4_810 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf3) );
BUFX4 BUFX4_811 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf2) );
BUFX4 BUFX4_812 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf1) );
BUFX4 BUFX4_813 ( .gnd(gnd), .vdd(vdd), .A(_15183_), .Y(_15183__bF_buf0) );
BUFX4 BUFX4_814 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .Y(_15086__bF_buf4) );
BUFX4 BUFX4_815 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .Y(_15086__bF_buf3) );
BUFX4 BUFX4_816 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .Y(_15086__bF_buf2) );
BUFX4 BUFX4_817 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .Y(_15086__bF_buf1) );
BUFX4 BUFX4_818 ( .gnd(gnd), .vdd(vdd), .A(_15086_), .Y(_15086__bF_buf0) );
BUFX4 BUFX4_819 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[10]), .Y(IDATA_PROG_data_10_bF_buf4) );
BUFX4 BUFX4_820 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[10]), .Y(IDATA_PROG_data_10_bF_buf3) );
BUFX4 BUFX4_821 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[10]), .Y(IDATA_PROG_data_10_bF_buf2) );
BUFX4 BUFX4_822 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[10]), .Y(IDATA_PROG_data_10_bF_buf1) );
BUFX4 BUFX4_823 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[10]), .Y(IDATA_PROG_data_10_bF_buf0) );
BUFX4 BUFX4_824 ( .gnd(gnd), .vdd(vdd), .A(_7123_), .Y(_7123__bF_buf3) );
BUFX4 BUFX4_825 ( .gnd(gnd), .vdd(vdd), .A(_7123_), .Y(_7123__bF_buf2) );
BUFX4 BUFX4_826 ( .gnd(gnd), .vdd(vdd), .A(_7123_), .Y(_7123__bF_buf1) );
BUFX4 BUFX4_827 ( .gnd(gnd), .vdd(vdd), .A(_7123_), .Y(_7123__bF_buf0) );
BUFX4 BUFX4_828 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[4]), .Y(IDATA_PROG_data_4_bF_buf4) );
BUFX4 BUFX4_829 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[4]), .Y(IDATA_PROG_data_4_bF_buf3) );
BUFX4 BUFX4_830 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[4]), .Y(IDATA_PROG_data_4_bF_buf2) );
BUFX4 BUFX4_831 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[4]), .Y(IDATA_PROG_data_4_bF_buf1) );
BUFX4 BUFX4_832 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[4]), .Y(IDATA_PROG_data_4_bF_buf0) );
BUFX4 BUFX4_833 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .Y(_1890__bF_buf3) );
BUFX4 BUFX4_834 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .Y(_1890__bF_buf2) );
BUFX4 BUFX4_835 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .Y(_1890__bF_buf1) );
BUFX4 BUFX4_836 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .Y(_1890__bF_buf0) );
BUFX4 BUFX4_837 ( .gnd(gnd), .vdd(vdd), .A(_14965_), .Y(_14965__bF_buf3) );
BUFX4 BUFX4_838 ( .gnd(gnd), .vdd(vdd), .A(_14965_), .Y(_14965__bF_buf2) );
BUFX4 BUFX4_839 ( .gnd(gnd), .vdd(vdd), .A(_14965_), .Y(_14965__bF_buf1) );
BUFX4 BUFX4_840 ( .gnd(gnd), .vdd(vdd), .A(_14965_), .Y(_14965__bF_buf0) );
BUFX4 BUFX4_841 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .Y(_2387__bF_buf3) );
BUFX4 BUFX4_842 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .Y(_2387__bF_buf2) );
BUFX4 BUFX4_843 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .Y(_2387__bF_buf1) );
BUFX4 BUFX4_844 ( .gnd(gnd), .vdd(vdd), .A(_2387_), .Y(_2387__bF_buf0) );
BUFX4 BUFX4_845 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf9) );
BUFX4 BUFX4_846 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf8) );
BUFX4 BUFX4_847 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf7) );
BUFX4 BUFX4_848 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf6) );
BUFX4 BUFX4_849 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf5) );
BUFX4 BUFX4_850 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf4) );
BUFX4 BUFX4_851 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf3) );
BUFX4 BUFX4_852 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf2) );
BUFX4 BUFX4_853 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf1) );
BUFX4 BUFX4_854 ( .gnd(gnd), .vdd(vdd), .A(_15788_), .Y(_15788__bF_buf0) );
BUFX4 BUFX4_855 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[1]), .Y(IDATA_PROG_data_1_bF_buf4) );
BUFX4 BUFX4_856 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[1]), .Y(IDATA_PROG_data_1_bF_buf3) );
BUFX4 BUFX4_857 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[1]), .Y(IDATA_PROG_data_1_bF_buf2) );
BUFX4 BUFX4_858 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[1]), .Y(IDATA_PROG_data_1_bF_buf1) );
BUFX4 BUFX4_859 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[1]), .Y(IDATA_PROG_data_1_bF_buf0) );
BUFX4 BUFX4_860 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf3) );
BUFX4 BUFX4_861 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf2) );
BUFX4 BUFX4_862 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf1) );
BUFX4 BUFX4_863 ( .gnd(gnd), .vdd(vdd), .A(_913_), .Y(_913__bF_buf0) );
BUFX4 BUFX4_864 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf13) );
BUFX4 BUFX4_865 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf12) );
BUFX4 BUFX4_866 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf11) );
BUFX4 BUFX4_867 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf10) );
BUFX4 BUFX4_868 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf9) );
BUFX4 BUFX4_869 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf8) );
BUFX4 BUFX4_870 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf7) );
BUFX4 BUFX4_871 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf6) );
BUFX4 BUFX4_872 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf5) );
BUFX4 BUFX4_873 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf4) );
BUFX4 BUFX4_874 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf3) );
BUFX4 BUFX4_875 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf2) );
BUFX4 BUFX4_876 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf1) );
BUFX4 BUFX4_877 ( .gnd(gnd), .vdd(vdd), .A(_14924_), .Y(_14924__bF_buf0) );
BUFX4 BUFX4_878 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .Y(_15042__bF_buf3) );
BUFX4 BUFX4_879 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .Y(_15042__bF_buf2) );
BUFX4 BUFX4_880 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .Y(_15042__bF_buf1) );
BUFX4 BUFX4_881 ( .gnd(gnd), .vdd(vdd), .A(_15042_), .Y(_15042__bF_buf0) );
BUFX4 BUFX4_882 ( .gnd(gnd), .vdd(vdd), .A(_948_), .Y(_948__bF_buf4) );
BUFX4 BUFX4_883 ( .gnd(gnd), .vdd(vdd), .A(_948_), .Y(_948__bF_buf3) );
BUFX4 BUFX4_884 ( .gnd(gnd), .vdd(vdd), .A(_948_), .Y(_948__bF_buf2) );
BUFX4 BUFX4_885 ( .gnd(gnd), .vdd(vdd), .A(_948_), .Y(_948__bF_buf1) );
BUFX4 BUFX4_886 ( .gnd(gnd), .vdd(vdd), .A(_948_), .Y(_948__bF_buf0) );
BUFX4 BUFX4_887 ( .gnd(gnd), .vdd(vdd), .A(_15688_), .Y(_15688__bF_buf3) );
BUFX4 BUFX4_888 ( .gnd(gnd), .vdd(vdd), .A(_15688_), .Y(_15688__bF_buf2) );
BUFX4 BUFX4_889 ( .gnd(gnd), .vdd(vdd), .A(_15688_), .Y(_15688__bF_buf1) );
BUFX4 BUFX4_890 ( .gnd(gnd), .vdd(vdd), .A(_15688_), .Y(_15688__bF_buf0) );
BUFX4 BUFX4_891 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf10) );
BUFX4 BUFX4_892 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf9) );
BUFX4 BUFX4_893 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf8) );
BUFX4 BUFX4_894 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf7) );
BUFX4 BUFX4_895 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf6) );
BUFX4 BUFX4_896 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf5) );
BUFX4 BUFX4_897 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf4) );
BUFX4 BUFX4_898 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf3) );
BUFX4 BUFX4_899 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf2) );
BUFX4 BUFX4_900 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf1) );
BUFX4 BUFX4_901 ( .gnd(gnd), .vdd(vdd), .A(_15900_), .Y(_15900__bF_buf0) );
BUFX4 BUFX4_902 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .Y(_1079__bF_buf3) );
BUFX4 BUFX4_903 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .Y(_1079__bF_buf2) );
BUFX4 BUFX4_904 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .Y(_1079__bF_buf1) );
BUFX4 BUFX4_905 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .Y(_1079__bF_buf0) );
BUFX4 BUFX4_906 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .Y(_15515__bF_buf3) );
BUFX4 BUFX4_907 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .Y(_15515__bF_buf2) );
BUFX4 BUFX4_908 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .Y(_15515__bF_buf1) );
BUFX4 BUFX4_909 ( .gnd(gnd), .vdd(vdd), .A(_15515_), .Y(_15515__bF_buf0) );
BUFX4 BUFX4_910 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .Y(_3395__bF_buf3) );
BUFX4 BUFX4_911 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .Y(_3395__bF_buf2) );
BUFX4 BUFX4_912 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .Y(_3395__bF_buf1) );
BUFX4 BUFX4_913 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .Y(_3395__bF_buf0) );
BUFX4 BUFX4_914 ( .gnd(gnd), .vdd(vdd), .A(_15838_), .Y(_15838__bF_buf3) );
BUFX4 BUFX4_915 ( .gnd(gnd), .vdd(vdd), .A(_15838_), .Y(_15838__bF_buf2) );
BUFX4 BUFX4_916 ( .gnd(gnd), .vdd(vdd), .A(_15838_), .Y(_15838__bF_buf1) );
BUFX4 BUFX4_917 ( .gnd(gnd), .vdd(vdd), .A(_15838_), .Y(_15838__bF_buf0) );
BUFX4 BUFX4_918 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf13) );
BUFX4 BUFX4_919 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf12) );
BUFX4 BUFX4_920 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf11) );
BUFX4 BUFX4_921 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf10) );
BUFX4 BUFX4_922 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf9) );
BUFX4 BUFX4_923 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf8) );
BUFX4 BUFX4_924 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf7) );
BUFX4 BUFX4_925 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf6) );
BUFX4 BUFX4_926 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf5) );
BUFX4 BUFX4_927 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf4) );
BUFX4 BUFX4_928 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf3) );
BUFX4 BUFX4_929 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf2) );
BUFX4 BUFX4_930 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf1) );
BUFX4 BUFX4_931 ( .gnd(gnd), .vdd(vdd), .A(_14918_), .Y(_14918__bF_buf0) );
BUFX4 BUFX4_932 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf12) );
BUFX4 BUFX4_933 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf11) );
BUFX4 BUFX4_934 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf10) );
BUFX4 BUFX4_935 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf9) );
BUFX4 BUFX4_936 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf8) );
BUFX4 BUFX4_937 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf7) );
BUFX4 BUFX4_938 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf6) );
BUFX4 BUFX4_939 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf5) );
BUFX4 BUFX4_940 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf4) );
BUFX4 BUFX4_941 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf3) );
BUFX4 BUFX4_942 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf2) );
BUFX4 BUFX4_943 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf1) );
BUFX4 BUFX4_944 ( .gnd(gnd), .vdd(vdd), .A(_15074_), .Y(_15074__bF_buf0) );
BUFX4 BUFX4_945 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .Y(_1229__bF_buf4) );
BUFX4 BUFX4_946 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .Y(_1229__bF_buf3) );
BUFX4 BUFX4_947 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .Y(_1229__bF_buf2) );
BUFX4 BUFX4_948 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .Y(_1229__bF_buf1) );
BUFX4 BUFX4_949 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .Y(_1229__bF_buf0) );
BUFX4 BUFX4_950 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .Y(_7302__bF_buf3) );
BUFX4 BUFX4_951 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .Y(_7302__bF_buf2) );
BUFX4 BUFX4_952 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .Y(_7302__bF_buf1) );
BUFX4 BUFX4_953 ( .gnd(gnd), .vdd(vdd), .A(_7302_), .Y(_7302__bF_buf0) );
BUFX4 BUFX4_954 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf14) );
BUFX4 BUFX4_955 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf13) );
BUFX4 BUFX4_956 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf12) );
BUFX4 BUFX4_957 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf11) );
BUFX4 BUFX4_958 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf10) );
BUFX4 BUFX4_959 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf9) );
BUFX4 BUFX4_960 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf8) );
BUFX4 BUFX4_961 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf7) );
BUFX4 BUFX4_962 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf6) );
BUFX4 BUFX4_963 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf5) );
BUFX4 BUFX4_964 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf4) );
BUFX4 BUFX4_965 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf3) );
BUFX4 BUFX4_966 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf2) );
BUFX4 BUFX4_967 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf1) );
BUFX4 BUFX4_968 ( .gnd(gnd), .vdd(vdd), .A(_14897_), .Y(_14897__bF_buf0) );
BUFX4 BUFX4_969 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .Y(_8125__bF_buf5) );
BUFX4 BUFX4_970 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .Y(_8125__bF_buf4) );
BUFX4 BUFX4_971 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .Y(_8125__bF_buf3) );
BUFX4 BUFX4_972 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .Y(_8125__bF_buf2) );
BUFX4 BUFX4_973 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .Y(_8125__bF_buf1) );
BUFX4 BUFX4_974 ( .gnd(gnd), .vdd(vdd), .A(_8125_), .Y(_8125__bF_buf0) );
BUFX4 BUFX4_975 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .Y(_3354__bF_buf3) );
BUFX4 BUFX4_976 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .Y(_3354__bF_buf2) );
BUFX4 BUFX4_977 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .Y(_3354__bF_buf1) );
BUFX4 BUFX4_978 ( .gnd(gnd), .vdd(vdd), .A(_3354_), .Y(_3354__bF_buf0) );
BUFX4 BUFX4_979 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf4) );
BUFX4 BUFX4_980 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf3) );
BUFX4 BUFX4_981 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf2) );
BUFX4 BUFX4_982 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf1) );
BUFX4 BUFX4_983 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf0) );
BUFX4 BUFX4_984 ( .gnd(gnd), .vdd(vdd), .A(_425_), .Y(_425__bF_buf3) );
BUFX4 BUFX4_985 ( .gnd(gnd), .vdd(vdd), .A(_425_), .Y(_425__bF_buf2) );
BUFX4 BUFX4_986 ( .gnd(gnd), .vdd(vdd), .A(_425_), .Y(_425__bF_buf1) );
BUFX4 BUFX4_987 ( .gnd(gnd), .vdd(vdd), .A(_425_), .Y(_425__bF_buf0) );
BUFX4 BUFX4_988 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf14) );
BUFX4 BUFX4_989 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf13) );
BUFX4 BUFX4_990 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf12) );
BUFX4 BUFX4_991 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf11) );
BUFX4 BUFX4_992 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf10) );
BUFX4 BUFX4_993 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf9) );
BUFX4 BUFX4_994 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf8) );
BUFX4 BUFX4_995 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf7) );
BUFX4 BUFX4_996 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf6) );
BUFX4 BUFX4_997 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf5) );
BUFX4 BUFX4_998 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf4) );
BUFX4 BUFX4_999 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf3) );
BUFX4 BUFX4_1000 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf2) );
BUFX4 BUFX4_1001 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf1) );
BUFX4 BUFX4_1002 ( .gnd(gnd), .vdd(vdd), .A(_14894_), .Y(_14894__bF_buf0) );
BUFX4 BUFX4_1003 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf91) );
BUFX4 BUFX4_1004 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf90) );
BUFX4 BUFX4_1005 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf89) );
BUFX4 BUFX4_1006 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf88) );
BUFX4 BUFX4_1007 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf87) );
BUFX4 BUFX4_1008 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf86) );
BUFX4 BUFX4_1009 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf85) );
BUFX4 BUFX4_1010 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf84) );
BUFX4 BUFX4_1011 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf83) );
BUFX4 BUFX4_1012 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf82) );
BUFX4 BUFX4_1013 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf81) );
BUFX4 BUFX4_1014 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf80) );
BUFX4 BUFX4_1015 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf79) );
BUFX4 BUFX4_1016 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf78) );
BUFX4 BUFX4_1017 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf77) );
BUFX4 BUFX4_1018 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf76) );
BUFX4 BUFX4_1019 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf75) );
BUFX4 BUFX4_1020 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf74) );
BUFX4 BUFX4_1021 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf73) );
BUFX4 BUFX4_1022 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf72) );
BUFX4 BUFX4_1023 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf71) );
BUFX4 BUFX4_1024 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf70) );
BUFX4 BUFX4_1025 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf69) );
BUFX4 BUFX4_1026 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf68) );
BUFX4 BUFX4_1027 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf67) );
BUFX4 BUFX4_1028 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf66) );
BUFX4 BUFX4_1029 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf65) );
BUFX4 BUFX4_1030 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf64) );
BUFX4 BUFX4_1031 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf63) );
BUFX4 BUFX4_1032 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf62) );
BUFX4 BUFX4_1033 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf61) );
BUFX4 BUFX4_1034 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf60) );
BUFX4 BUFX4_1035 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf59) );
BUFX4 BUFX4_1036 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf58) );
BUFX4 BUFX4_1037 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf57) );
BUFX4 BUFX4_1038 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf56) );
BUFX4 BUFX4_1039 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf55) );
BUFX4 BUFX4_1040 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf54) );
BUFX4 BUFX4_1041 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf53) );
BUFX4 BUFX4_1042 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf52) );
BUFX4 BUFX4_1043 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf51) );
BUFX4 BUFX4_1044 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf50) );
BUFX4 BUFX4_1045 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf49) );
BUFX4 BUFX4_1046 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf48) );
BUFX4 BUFX4_1047 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf47) );
BUFX4 BUFX4_1048 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf46) );
BUFX4 BUFX4_1049 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf45) );
BUFX4 BUFX4_1050 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf44) );
BUFX4 BUFX4_1051 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf43) );
BUFX4 BUFX4_1052 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf42) );
BUFX4 BUFX4_1053 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf41) );
BUFX4 BUFX4_1054 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf40) );
BUFX4 BUFX4_1055 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf39) );
BUFX4 BUFX4_1056 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf38) );
BUFX4 BUFX4_1057 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf37) );
BUFX4 BUFX4_1058 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf36) );
BUFX4 BUFX4_1059 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf35) );
BUFX4 BUFX4_1060 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf34) );
BUFX4 BUFX4_1061 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf33) );
BUFX4 BUFX4_1062 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf32) );
BUFX4 BUFX4_1063 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf31) );
BUFX4 BUFX4_1064 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf30) );
BUFX4 BUFX4_1065 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf29) );
BUFX4 BUFX4_1066 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf28) );
BUFX4 BUFX4_1067 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf27) );
BUFX4 BUFX4_1068 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf26) );
BUFX4 BUFX4_1069 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf25) );
BUFX4 BUFX4_1070 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf24) );
BUFX4 BUFX4_1071 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf23) );
BUFX4 BUFX4_1072 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf22) );
BUFX4 BUFX4_1073 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf21) );
BUFX4 BUFX4_1074 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf20) );
BUFX4 BUFX4_1075 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf19) );
BUFX4 BUFX4_1076 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf18) );
BUFX4 BUFX4_1077 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf17) );
BUFX4 BUFX4_1078 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf16) );
BUFX4 BUFX4_1079 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf15) );
BUFX4 BUFX4_1080 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf14) );
BUFX4 BUFX4_1081 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf13) );
BUFX4 BUFX4_1082 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf12) );
BUFX4 BUFX4_1083 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf11) );
BUFX4 BUFX4_1084 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf10) );
BUFX4 BUFX4_1085 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf9) );
BUFX4 BUFX4_1086 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf6), .Y(_3313__bF_buf8) );
BUFX4 BUFX4_1087 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf5), .Y(_3313__bF_buf7) );
BUFX4 BUFX4_1088 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf4), .Y(_3313__bF_buf6) );
BUFX4 BUFX4_1089 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf3), .Y(_3313__bF_buf5) );
BUFX4 BUFX4_1090 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf2), .Y(_3313__bF_buf4) );
BUFX4 BUFX4_1091 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf1), .Y(_3313__bF_buf3) );
BUFX4 BUFX4_1092 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf0), .Y(_3313__bF_buf2) );
BUFX4 BUFX4_1093 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf8), .Y(_3313__bF_buf1) );
BUFX4 BUFX4_1094 ( .gnd(gnd), .vdd(vdd), .A(_3313__hier0_bF_buf7), .Y(_3313__bF_buf0) );
BUFX4 BUFX4_1095 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[3]), .Y(IDATA_PROG_addr_3_bF_buf3) );
BUFX4 BUFX4_1096 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[3]), .Y(IDATA_PROG_addr_3_bF_buf2) );
BUFX4 BUFX4_1097 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[3]), .Y(IDATA_PROG_addr_3_bF_buf1) );
BUFX4 BUFX4_1098 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[3]), .Y(IDATA_PROG_addr_3_bF_buf0) );
BUFX4 BUFX4_1099 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .Y(_7431__bF_buf4) );
BUFX4 BUFX4_1100 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .Y(_7431__bF_buf3) );
BUFX4 BUFX4_1101 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .Y(_7431__bF_buf2) );
BUFX4 BUFX4_1102 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .Y(_7431__bF_buf1) );
BUFX4 BUFX4_1103 ( .gnd(gnd), .vdd(vdd), .A(_7431_), .Y(_7431__bF_buf0) );
BUFX4 BUFX4_1104 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .Y(_2619__bF_buf3) );
BUFX4 BUFX4_1105 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .Y(_2619__bF_buf2) );
BUFX4 BUFX4_1106 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .Y(_2619__bF_buf1) );
BUFX4 BUFX4_1107 ( .gnd(gnd), .vdd(vdd), .A(_2619_), .Y(_2619__bF_buf0) );
BUFX4 BUFX4_1108 ( .gnd(gnd), .vdd(vdd), .A(_974_), .Y(_974__bF_buf3) );
BUFX4 BUFX4_1109 ( .gnd(gnd), .vdd(vdd), .A(_974_), .Y(_974__bF_buf2) );
BUFX4 BUFX4_1110 ( .gnd(gnd), .vdd(vdd), .A(_974_), .Y(_974__bF_buf1) );
BUFX4 BUFX4_1111 ( .gnd(gnd), .vdd(vdd), .A(_974_), .Y(_974__bF_buf0) );
BUFX4 BUFX4_1112 ( .gnd(gnd), .vdd(vdd), .A(_15065_), .Y(_15065__bF_buf3) );
BUFX4 BUFX4_1113 ( .gnd(gnd), .vdd(vdd), .A(_15065_), .Y(_15065__bF_buf2) );
BUFX4 BUFX4_1114 ( .gnd(gnd), .vdd(vdd), .A(_15065_), .Y(_15065__bF_buf1) );
BUFX4 BUFX4_1115 ( .gnd(gnd), .vdd(vdd), .A(_15065_), .Y(_15065__bF_buf0) );
BUFX4 BUFX4_1116 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(_4171__bF_buf4) );
BUFX4 BUFX4_1117 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(_4171__bF_buf3) );
BUFX4 BUFX4_1118 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(_4171__bF_buf2) );
BUFX4 BUFX4_1119 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(_4171__bF_buf1) );
BUFX4 BUFX4_1120 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .Y(_4171__bF_buf0) );
BUFX4 BUFX4_1121 ( .gnd(gnd), .vdd(vdd), .A(_14888_), .Y(_14888__bF_buf3) );
BUFX4 BUFX4_1122 ( .gnd(gnd), .vdd(vdd), .A(_14888_), .Y(_14888__bF_buf2) );
BUFX4 BUFX4_1123 ( .gnd(gnd), .vdd(vdd), .A(_14888_), .Y(_14888__bF_buf1) );
BUFX4 BUFX4_1124 ( .gnd(gnd), .vdd(vdd), .A(_14888_), .Y(_14888__bF_buf0) );
BUFX4 BUFX4_1125 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .Y(_5911__bF_buf3) );
BUFX4 BUFX4_1126 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .Y(_5911__bF_buf2) );
BUFX4 BUFX4_1127 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .Y(_5911__bF_buf1) );
BUFX4 BUFX4_1128 ( .gnd(gnd), .vdd(vdd), .A(_5911_), .Y(_5911__bF_buf0) );
BUFX4 BUFX4_1129 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf13) );
BUFX4 BUFX4_1130 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf12) );
BUFX4 BUFX4_1131 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf11) );
BUFX4 BUFX4_1132 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf10) );
BUFX4 BUFX4_1133 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf9) );
BUFX4 BUFX4_1134 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf8) );
BUFX4 BUFX4_1135 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf7) );
BUFX4 BUFX4_1136 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf6) );
BUFX4 BUFX4_1137 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf5) );
BUFX4 BUFX4_1138 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf4) );
BUFX4 BUFX4_1139 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf3) );
BUFX4 BUFX4_1140 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf2) );
BUFX4 BUFX4_1141 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf1) );
BUFX4 BUFX4_1142 ( .gnd(gnd), .vdd(vdd), .A(_15062_), .Y(_15062__bF_buf0) );
BUFX4 BUFX4_1143 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .Y(_14885__bF_buf3) );
BUFX4 BUFX4_1144 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .Y(_14885__bF_buf2) );
BUFX4 BUFX4_1145 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .Y(_14885__bF_buf1) );
BUFX4 BUFX4_1146 ( .gnd(gnd), .vdd(vdd), .A(_14885_), .Y(_14885__bF_buf0) );
BUFX4 BUFX4_1147 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .Y(_15632__bF_buf3) );
BUFX4 BUFX4_1148 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .Y(_15632__bF_buf2) );
BUFX4 BUFX4_1149 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .Y(_15632__bF_buf1) );
BUFX4 BUFX4_1150 ( .gnd(gnd), .vdd(vdd), .A(_15632_), .Y(_15632__bF_buf0) );
BUFX4 BUFX4_1151 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf13) );
BUFX4 BUFX4_1152 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf12) );
BUFX4 BUFX4_1153 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf11) );
BUFX4 BUFX4_1154 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf10) );
BUFX4 BUFX4_1155 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf9) );
BUFX4 BUFX4_1156 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf8) );
BUFX4 BUFX4_1157 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf7) );
BUFX4 BUFX4_1158 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf6) );
BUFX4 BUFX4_1159 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf5) );
BUFX4 BUFX4_1160 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf4) );
BUFX4 BUFX4_1161 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf3) );
BUFX4 BUFX4_1162 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf2) );
BUFX4 BUFX4_1163 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf1) );
BUFX4 BUFX4_1164 ( .gnd(gnd), .vdd(vdd), .A(_14903_), .Y(_14903__bF_buf0) );
BUFX4 BUFX4_1165 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf15) );
BUFX4 BUFX4_1166 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf14) );
BUFX4 BUFX4_1167 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf13) );
BUFX4 BUFX4_1168 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf12) );
BUFX4 BUFX4_1169 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf11) );
BUFX4 BUFX4_1170 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf10) );
BUFX4 BUFX4_1171 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf9) );
BUFX4 BUFX4_1172 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf8) );
BUFX4 BUFX4_1173 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf7) );
BUFX4 BUFX4_1174 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf6) );
BUFX4 BUFX4_1175 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf5) );
BUFX4 BUFX4_1176 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf4) );
BUFX4 BUFX4_1177 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf3) );
BUFX4 BUFX4_1178 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf2) );
BUFX4 BUFX4_1179 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf1) );
BUFX4 BUFX4_1180 ( .gnd(gnd), .vdd(vdd), .A(_14882_), .Y(_14882__bF_buf0) );
BUFX4 BUFX4_1181 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .Y(_3089__bF_buf3) );
BUFX4 BUFX4_1182 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .Y(_3089__bF_buf2) );
BUFX4 BUFX4_1183 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .Y(_3089__bF_buf1) );
BUFX4 BUFX4_1184 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .Y(_3089__bF_buf0) );
BUFX4 BUFX4_1185 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf3) );
BUFX4 BUFX4_1186 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf2) );
BUFX4 BUFX4_1187 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf1) );
BUFX4 BUFX4_1188 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .Y(_2513__bF_buf0) );
BUFX4 BUFX4_1189 ( .gnd(gnd), .vdd(vdd), .A(_8145_), .Y(_8145__bF_buf3) );
BUFX4 BUFX4_1190 ( .gnd(gnd), .vdd(vdd), .A(_8145_), .Y(_8145__bF_buf2) );
BUFX4 BUFX4_1191 ( .gnd(gnd), .vdd(vdd), .A(_8145_), .Y(_8145__bF_buf1) );
BUFX4 BUFX4_1192 ( .gnd(gnd), .vdd(vdd), .A(_8145_), .Y(_8145__bF_buf0) );
BUFX4 BUFX4_1193 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[15]), .Y(IDATA_PROG_data_15_bF_buf5) );
BUFX4 BUFX4_1194 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[15]), .Y(IDATA_PROG_data_15_bF_buf4) );
BUFX4 BUFX4_1195 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[15]), .Y(IDATA_PROG_data_15_bF_buf3) );
BUFX4 BUFX4_1196 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[15]), .Y(IDATA_PROG_data_15_bF_buf2) );
BUFX4 BUFX4_1197 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[15]), .Y(IDATA_PROG_data_15_bF_buf1) );
BUFX4 BUFX4_1198 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[15]), .Y(IDATA_PROG_data_15_bF_buf0) );
BUFX4 BUFX4_1199 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .Y(_2319__bF_buf4) );
BUFX4 BUFX4_1200 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .Y(_2319__bF_buf3) );
BUFX4 BUFX4_1201 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .Y(_2319__bF_buf2) );
BUFX4 BUFX4_1202 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .Y(_2319__bF_buf1) );
BUFX4 BUFX4_1203 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .Y(_2319__bF_buf0) );
BUFX4 BUFX4_1204 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[9]), .Y(IDATA_PROG_data_9_bF_buf4) );
BUFX4 BUFX4_1205 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[9]), .Y(IDATA_PROG_data_9_bF_buf3) );
BUFX4 BUFX4_1206 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[9]), .Y(IDATA_PROG_data_9_bF_buf2) );
BUFX4 BUFX4_1207 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[9]), .Y(IDATA_PROG_data_9_bF_buf1) );
BUFX4 BUFX4_1208 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[9]), .Y(IDATA_PROG_data_9_bF_buf0) );
BUFX4 BUFX4_1209 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf8) );
BUFX4 BUFX4_1210 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf7) );
BUFX4 BUFX4_1211 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf6) );
BUFX4 BUFX4_1212 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf5) );
BUFX4 BUFX4_1213 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf4) );
BUFX4 BUFX4_1214 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf3) );
BUFX4 BUFX4_1215 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf2) );
BUFX4 BUFX4_1216 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf1) );
BUFX4 BUFX4_1217 ( .gnd(gnd), .vdd(vdd), .A(_15949_), .Y(_15949__bF_buf0) );
BUFX4 BUFX4_1218 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf3) );
BUFX4 BUFX4_1219 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf2) );
BUFX4 BUFX4_1220 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf1) );
BUFX4 BUFX4_1221 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .Y(_5076__bF_buf0) );
BUFX4 BUFX4_1222 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .Y(_2871__bF_buf4) );
BUFX4 BUFX4_1223 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .Y(_2871__bF_buf3) );
BUFX4 BUFX4_1224 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .Y(_2871__bF_buf2) );
BUFX4 BUFX4_1225 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .Y(_2871__bF_buf1) );
BUFX4 BUFX4_1226 ( .gnd(gnd), .vdd(vdd), .A(_2871_), .Y(_2871__bF_buf0) );
BUFX4 BUFX4_1227 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[12]), .Y(IDATA_PROG_data_12_bF_buf4) );
BUFX4 BUFX4_1228 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[12]), .Y(IDATA_PROG_data_12_bF_buf3) );
BUFX4 BUFX4_1229 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[12]), .Y(IDATA_PROG_data_12_bF_buf2) );
BUFX4 BUFX4_1230 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[12]), .Y(IDATA_PROG_data_12_bF_buf1) );
BUFX4 BUFX4_1231 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[12]), .Y(IDATA_PROG_data_12_bF_buf0) );
BUFX4 BUFX4_1232 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[6]), .Y(IDATA_PROG_data_6_bF_buf4) );
BUFX4 BUFX4_1233 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[6]), .Y(IDATA_PROG_data_6_bF_buf3) );
BUFX4 BUFX4_1234 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[6]), .Y(IDATA_PROG_data_6_bF_buf2) );
BUFX4 BUFX4_1235 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[6]), .Y(IDATA_PROG_data_6_bF_buf1) );
BUFX4 BUFX4_1236 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[6]), .Y(IDATA_PROG_data_6_bF_buf0) );
BUFX4 BUFX4_1237 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .Y(_5420__bF_buf3) );
BUFX4 BUFX4_1238 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .Y(_5420__bF_buf2) );
BUFX4 BUFX4_1239 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .Y(_5420__bF_buf1) );
BUFX4 BUFX4_1240 ( .gnd(gnd), .vdd(vdd), .A(_5420_), .Y(_5420__bF_buf0) );
BUFX4 BUFX4_1241 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf14) );
BUFX4 BUFX4_1242 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf13) );
BUFX4 BUFX4_1243 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf12) );
BUFX4 BUFX4_1244 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf11) );
BUFX4 BUFX4_1245 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf10) );
BUFX4 BUFX4_1246 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf9) );
BUFX4 BUFX4_1247 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf8) );
BUFX4 BUFX4_1248 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf7) );
BUFX4 BUFX4_1249 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf6) );
BUFX4 BUFX4_1250 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf5) );
BUFX4 BUFX4_1251 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf4) );
BUFX4 BUFX4_1252 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf3) );
BUFX4 BUFX4_1253 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf2) );
BUFX4 BUFX4_1254 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf1) );
BUFX4 BUFX4_1255 ( .gnd(gnd), .vdd(vdd), .A(_14932_), .Y(_14932__bF_buf0) );
BUFX4 BUFX4_1256 ( .gnd(gnd), .vdd(vdd), .A(_7448_), .Y(_7448__bF_buf3) );
BUFX4 BUFX4_1257 ( .gnd(gnd), .vdd(vdd), .A(_7448_), .Y(_7448__bF_buf2) );
BUFX4 BUFX4_1258 ( .gnd(gnd), .vdd(vdd), .A(_7448_), .Y(_7448__bF_buf1) );
BUFX4 BUFX4_1259 ( .gnd(gnd), .vdd(vdd), .A(_7448_), .Y(_7448__bF_buf0) );
BUFX4 BUFX4_1260 ( .gnd(gnd), .vdd(vdd), .A(_15335_), .Y(_15335__bF_buf3) );
BUFX4 BUFX4_1261 ( .gnd(gnd), .vdd(vdd), .A(_15335_), .Y(_15335__bF_buf2) );
BUFX4 BUFX4_1262 ( .gnd(gnd), .vdd(vdd), .A(_15335_), .Y(_15335__bF_buf1) );
BUFX4 BUFX4_1263 ( .gnd(gnd), .vdd(vdd), .A(_15335_), .Y(_15335__bF_buf0) );
BUFX4 BUFX4_1264 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .Y(_15793__bF_buf5) );
BUFX4 BUFX4_1265 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .Y(_15793__bF_buf4) );
BUFX4 BUFX4_1266 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .Y(_15793__bF_buf3) );
BUFX4 BUFX4_1267 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .Y(_15793__bF_buf2) );
BUFX4 BUFX4_1268 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .Y(_15793__bF_buf1) );
BUFX4 BUFX4_1269 ( .gnd(gnd), .vdd(vdd), .A(_15793_), .Y(_15793__bF_buf0) );
BUFX4 BUFX4_1270 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1528__bF_buf5) );
BUFX4 BUFX4_1271 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1528__bF_buf4) );
BUFX4 BUFX4_1272 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1528__bF_buf3) );
BUFX4 BUFX4_1273 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1528__bF_buf2) );
BUFX4 BUFX4_1274 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1528__bF_buf1) );
BUFX4 BUFX4_1275 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .Y(_1528__bF_buf0) );
BUFX4 BUFX4_1276 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .Y(_2601__bF_buf4) );
BUFX4 BUFX4_1277 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .Y(_2601__bF_buf3) );
BUFX4 BUFX4_1278 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .Y(_2601__bF_buf2) );
BUFX4 BUFX4_1279 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .Y(_2601__bF_buf1) );
BUFX4 BUFX4_1280 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .Y(_2601__bF_buf0) );
BUFX4 BUFX4_1281 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[3]), .Y(IDATA_PROG_data_3_bF_buf4) );
BUFX4 BUFX4_1282 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[3]), .Y(IDATA_PROG_data_3_bF_buf3) );
BUFX4 BUFX4_1283 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[3]), .Y(IDATA_PROG_data_3_bF_buf2) );
BUFX4 BUFX4_1284 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[3]), .Y(IDATA_PROG_data_3_bF_buf1) );
BUFX4 BUFX4_1285 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[3]), .Y(IDATA_PROG_data_3_bF_buf0) );
BUFX4 BUFX4_1286 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_342__bF_buf4) );
BUFX4 BUFX4_1287 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_342__bF_buf3) );
BUFX4 BUFX4_1288 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_342__bF_buf2) );
BUFX4 BUFX4_1289 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_342__bF_buf1) );
BUFX4 BUFX4_1290 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_342__bF_buf0) );
BUFX4 BUFX4_1291 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3039__bF_buf4) );
BUFX4 BUFX4_1292 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3039__bF_buf3) );
BUFX4 BUFX4_1293 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3039__bF_buf2) );
BUFX4 BUFX4_1294 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3039__bF_buf1) );
BUFX4 BUFX4_1295 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .Y(_3039__bF_buf0) );
BUFX4 BUFX4_1296 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .Y(_1525__bF_buf4) );
BUFX4 BUFX4_1297 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .Y(_1525__bF_buf3) );
BUFX4 BUFX4_1298 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .Y(_1525__bF_buf2) );
BUFX4 BUFX4_1299 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .Y(_1525__bF_buf1) );
BUFX4 BUFX4_1300 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .Y(_1525__bF_buf0) );
BUFX4 BUFX4_1301 ( .gnd(gnd), .vdd(vdd), .A(_15006_), .Y(_15006__bF_buf4) );
BUFX4 BUFX4_1302 ( .gnd(gnd), .vdd(vdd), .A(_15006_), .Y(_15006__bF_buf3) );
BUFX4 BUFX4_1303 ( .gnd(gnd), .vdd(vdd), .A(_15006_), .Y(_15006__bF_buf2) );
BUFX4 BUFX4_1304 ( .gnd(gnd), .vdd(vdd), .A(_15006_), .Y(_15006__bF_buf1) );
BUFX4 BUFX4_1305 ( .gnd(gnd), .vdd(vdd), .A(_15006_), .Y(_15006__bF_buf0) );
BUFX4 BUFX4_1306 ( .gnd(gnd), .vdd(vdd), .A(_2063_), .Y(_2063__bF_buf3) );
BUFX4 BUFX4_1307 ( .gnd(gnd), .vdd(vdd), .A(_2063_), .Y(_2063__bF_buf2) );
BUFX4 BUFX4_1308 ( .gnd(gnd), .vdd(vdd), .A(_2063_), .Y(_2063__bF_buf1) );
BUFX4 BUFX4_1309 ( .gnd(gnd), .vdd(vdd), .A(_2063_), .Y(_2063__bF_buf0) );
BUFX4 BUFX4_1310 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf4) );
BUFX4 BUFX4_1311 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf3) );
BUFX4 BUFX4_1312 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf2) );
BUFX4 BUFX4_1313 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf1) );
BUFX4 BUFX4_1314 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .Y(_2959__bF_buf0) );
BUFX4 BUFX4_1315 ( .gnd(gnd), .vdd(vdd), .A(_15235_), .Y(_15235__bF_buf3) );
BUFX4 BUFX4_1316 ( .gnd(gnd), .vdd(vdd), .A(_15235_), .Y(_15235__bF_buf2) );
BUFX4 BUFX4_1317 ( .gnd(gnd), .vdd(vdd), .A(_15235_), .Y(_15235__bF_buf1) );
BUFX4 BUFX4_1318 ( .gnd(gnd), .vdd(vdd), .A(_15235_), .Y(_15235__bF_buf0) );
BUFX4 BUFX4_1319 ( .gnd(gnd), .vdd(vdd), .A(_15367_), .Y(_15367__bF_buf3) );
BUFX4 BUFX4_1320 ( .gnd(gnd), .vdd(vdd), .A(_15367_), .Y(_15367__bF_buf2) );
BUFX4 BUFX4_1321 ( .gnd(gnd), .vdd(vdd), .A(_15367_), .Y(_15367__bF_buf1) );
BUFX4 BUFX4_1322 ( .gnd(gnd), .vdd(vdd), .A(_15367_), .Y(_15367__bF_buf0) );
BUFX4 BUFX4_1323 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[0]), .Y(IDATA_PROG_data_0_bF_buf4) );
BUFX4 BUFX4_1324 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[0]), .Y(IDATA_PROG_data_0_bF_buf3) );
BUFX4 BUFX4_1325 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[0]), .Y(IDATA_PROG_data_0_bF_buf2) );
BUFX4 BUFX4_1326 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[0]), .Y(IDATA_PROG_data_0_bF_buf1) );
BUFX4 BUFX4_1327 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data[0]), .Y(IDATA_PROG_data_0_bF_buf0) );
BUFX4 BUFX4_1328 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .Y(_8782__bF_buf3) );
BUFX4 BUFX4_1329 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .Y(_8782__bF_buf2) );
BUFX4 BUFX4_1330 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .Y(_8782__bF_buf1) );
BUFX4 BUFX4_1331 ( .gnd(gnd), .vdd(vdd), .A(_8782_), .Y(_8782__bF_buf0) );
BUFX4 BUFX4_1332 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf7) );
BUFX4 BUFX4_1333 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf6) );
BUFX4 BUFX4_1334 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf5) );
BUFX4 BUFX4_1335 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf4) );
BUFX4 BUFX4_1336 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf3) );
BUFX4 BUFX4_1337 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf2) );
BUFX4 BUFX4_1338 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf1) );
BUFX4 BUFX4_1339 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .Y(_1810__bF_buf0) );
BUFX4 BUFX4_1340 ( .gnd(gnd), .vdd(vdd), .A(_7213_), .Y(_7213__bF_buf3) );
BUFX4 BUFX4_1341 ( .gnd(gnd), .vdd(vdd), .A(_7213_), .Y(_7213__bF_buf2) );
BUFX4 BUFX4_1342 ( .gnd(gnd), .vdd(vdd), .A(_7213_), .Y(_7213__bF_buf1) );
BUFX4 BUFX4_1343 ( .gnd(gnd), .vdd(vdd), .A(_7213_), .Y(_7213__bF_buf0) );
BUFX4 BUFX4_1344 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .Y(_1942__bF_buf3) );
BUFX4 BUFX4_1345 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .Y(_1942__bF_buf2) );
BUFX4 BUFX4_1346 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .Y(_1942__bF_buf1) );
BUFX4 BUFX4_1347 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .Y(_1942__bF_buf0) );
BUFX4 BUFX4_1348 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .Y(_7345__bF_buf3) );
BUFX4 BUFX4_1349 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .Y(_7345__bF_buf2) );
BUFX4 BUFX4_1350 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .Y(_7345__bF_buf1) );
BUFX4 BUFX4_1351 ( .gnd(gnd), .vdd(vdd), .A(_7345_), .Y(_7345__bF_buf0) );
BUFX4 BUFX4_1352 ( .gnd(gnd), .vdd(vdd), .A(_16111_), .Y(_16111__bF_buf3) );
BUFX4 BUFX4_1353 ( .gnd(gnd), .vdd(vdd), .A(_16111_), .Y(_16111__bF_buf2) );
BUFX4 BUFX4_1354 ( .gnd(gnd), .vdd(vdd), .A(_16111_), .Y(_16111__bF_buf1) );
BUFX4 BUFX4_1355 ( .gnd(gnd), .vdd(vdd), .A(_16111_), .Y(_16111__bF_buf0) );
BUFX4 BUFX4_1356 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf14) );
BUFX4 BUFX4_1357 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf13) );
BUFX4 BUFX4_1358 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf12) );
BUFX4 BUFX4_1359 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf11) );
BUFX4 BUFX4_1360 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf10) );
BUFX4 BUFX4_1361 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf9) );
BUFX4 BUFX4_1362 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf8) );
BUFX4 BUFX4_1363 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf7) );
BUFX4 BUFX4_1364 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf6) );
BUFX4 BUFX4_1365 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf5) );
BUFX4 BUFX4_1366 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf4) );
BUFX4 BUFX4_1367 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf3) );
BUFX4 BUFX4_1368 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf2) );
BUFX4 BUFX4_1369 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf1) );
BUFX4 BUFX4_1370 ( .gnd(gnd), .vdd(vdd), .A(_14899_), .Y(_14899__bF_buf0) );
BUFX4 BUFX4_1371 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf13) );
BUFX4 BUFX4_1372 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf12) );
BUFX4 BUFX4_1373 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf11) );
BUFX4 BUFX4_1374 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf10) );
BUFX4 BUFX4_1375 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf9) );
BUFX4 BUFX4_1376 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf8) );
BUFX4 BUFX4_1377 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf7) );
BUFX4 BUFX4_1378 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf6) );
BUFX4 BUFX4_1379 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf5) );
BUFX4 BUFX4_1380 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf4) );
BUFX4 BUFX4_1381 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf3) );
BUFX4 BUFX4_1382 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf2) );
BUFX4 BUFX4_1383 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf1) );
BUFX4 BUFX4_1384 ( .gnd(gnd), .vdd(vdd), .A(_14920_), .Y(_14920__bF_buf0) );
BUFX4 BUFX4_1385 ( .gnd(gnd), .vdd(vdd), .A(_6842_), .Y(_6842__bF_buf3) );
BUFX4 BUFX4_1386 ( .gnd(gnd), .vdd(vdd), .A(_6842_), .Y(_6842__bF_buf2) );
BUFX4 BUFX4_1387 ( .gnd(gnd), .vdd(vdd), .A(_6842_), .Y(_6842__bF_buf1) );
BUFX4 BUFX4_1388 ( .gnd(gnd), .vdd(vdd), .A(_6842_), .Y(_6842__bF_buf0) );
BUFX4 BUFX4_1389 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .Y(_1040__bF_buf3) );
BUFX4 BUFX4_1390 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .Y(_1040__bF_buf2) );
BUFX4 BUFX4_1391 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .Y(_1040__bF_buf1) );
BUFX4 BUFX4_1392 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .Y(_1040__bF_buf0) );
BUFX4 BUFX4_1393 ( .gnd(gnd), .vdd(vdd), .A(_15170_), .Y(_15170__bF_buf3) );
BUFX4 BUFX4_1394 ( .gnd(gnd), .vdd(vdd), .A(_15170_), .Y(_15170__bF_buf2) );
BUFX4 BUFX4_1395 ( .gnd(gnd), .vdd(vdd), .A(_15170_), .Y(_15170__bF_buf1) );
BUFX4 BUFX4_1396 ( .gnd(gnd), .vdd(vdd), .A(_15170_), .Y(_15170__bF_buf0) );
BUFX4 BUFX4_1397 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .Y(_2339__bF_buf3) );
BUFX4 BUFX4_1398 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .Y(_2339__bF_buf2) );
BUFX4 BUFX4_1399 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .Y(_2339__bF_buf1) );
BUFX4 BUFX4_1400 ( .gnd(gnd), .vdd(vdd), .A(_2339_), .Y(_2339__bF_buf0) );
BUFX4 BUFX4_1401 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .Y(_1266__bF_buf5) );
BUFX4 BUFX4_1402 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .Y(_1266__bF_buf4) );
BUFX4 BUFX4_1403 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .Y(_1266__bF_buf3) );
BUFX4 BUFX4_1404 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .Y(_1266__bF_buf2) );
BUFX4 BUFX4_1405 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .Y(_1266__bF_buf1) );
BUFX4 BUFX4_1406 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .Y(_1266__bF_buf0) );
BUFX4 BUFX4_1407 ( .gnd(gnd), .vdd(vdd), .A(_5384_), .Y(_5384__bF_buf3) );
BUFX4 BUFX4_1408 ( .gnd(gnd), .vdd(vdd), .A(_5384_), .Y(_5384__bF_buf2) );
BUFX4 BUFX4_1409 ( .gnd(gnd), .vdd(vdd), .A(_5384_), .Y(_5384__bF_buf1) );
BUFX4 BUFX4_1410 ( .gnd(gnd), .vdd(vdd), .A(_5384_), .Y(_5384__bF_buf0) );
BUFX4 BUFX4_1411 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .Y(_3353__bF_buf4) );
BUFX4 BUFX4_1412 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .Y(_3353__bF_buf3) );
BUFX4 BUFX4_1413 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .Y(_3353__bF_buf2) );
BUFX4 BUFX4_1414 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .Y(_3353__bF_buf1) );
BUFX4 BUFX4_1415 ( .gnd(gnd), .vdd(vdd), .A(_3353_), .Y(_3353__bF_buf0) );
BUFX4 BUFX4_1416 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf6) );
BUFX4 BUFX4_1417 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf5) );
BUFX4 BUFX4_1418 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf4) );
BUFX4 BUFX4_1419 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf3) );
BUFX4 BUFX4_1420 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf2) );
BUFX4 BUFX4_1421 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf1) );
BUFX4 BUFX4_1422 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3391__bF_buf0) );
BUFX4 BUFX4_1423 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .Y(_15834__bF_buf4) );
BUFX4 BUFX4_1424 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .Y(_15834__bF_buf3) );
BUFX4 BUFX4_1425 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .Y(_15834__bF_buf2) );
BUFX4 BUFX4_1426 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .Y(_15834__bF_buf1) );
BUFX4 BUFX4_1427 ( .gnd(gnd), .vdd(vdd), .A(_15834_), .Y(_15834__bF_buf0) );
BUFX4 BUFX4_1428 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .Y(_2471__bF_buf3) );
BUFX4 BUFX4_1429 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .Y(_2471__bF_buf2) );
BUFX4 BUFX4_1430 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .Y(_2471__bF_buf1) );
BUFX4 BUFX4_1431 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .Y(_2471__bF_buf0) );
BUFX4 BUFX4_1432 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .Y(_2280__bF_buf4) );
BUFX4 BUFX4_1433 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .Y(_2280__bF_buf3) );
BUFX4 BUFX4_1434 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .Y(_2280__bF_buf2) );
BUFX4 BUFX4_1435 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .Y(_2280__bF_buf1) );
BUFX4 BUFX4_1436 ( .gnd(gnd), .vdd(vdd), .A(_2280_), .Y(_2280__bF_buf0) );
BUFX4 BUFX4_1437 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf3) );
BUFX4 BUFX4_1438 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf2) );
BUFX4 BUFX4_1439 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf1) );
BUFX4 BUFX4_1440 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf0) );
BUFX4 BUFX4_1441 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .Y(_14952__bF_buf4) );
BUFX4 BUFX4_1442 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .Y(_14952__bF_buf3) );
BUFX4 BUFX4_1443 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .Y(_14952__bF_buf2) );
BUFX4 BUFX4_1444 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .Y(_14952__bF_buf1) );
BUFX4 BUFX4_1445 ( .gnd(gnd), .vdd(vdd), .A(_14952_), .Y(_14952__bF_buf0) );
BUFX4 BUFX4_1446 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf6) );
BUFX4 BUFX4_1447 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf5) );
BUFX4 BUFX4_1448 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf4) );
BUFX4 BUFX4_1449 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf3) );
BUFX4 BUFX4_1450 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf2) );
BUFX4 BUFX4_1451 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf1) );
BUFX4 BUFX4_1452 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .Y(_1225__bF_buf0) );
BUFX4 BUFX4_1453 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf7) );
BUFX4 BUFX4_1454 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf6) );
BUFX4 BUFX4_1455 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf5) );
BUFX4 BUFX4_1456 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf4) );
BUFX4 BUFX4_1457 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf3) );
BUFX4 BUFX4_1458 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf2) );
BUFX4 BUFX4_1459 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf1) );
BUFX4 BUFX4_1460 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .Y(_2621__bF_buf0) );
BUFX4 BUFX4_1461 ( .gnd(gnd), .vdd(vdd), .A(_2791_), .Y(_2791__bF_buf3) );
BUFX4 BUFX4_1462 ( .gnd(gnd), .vdd(vdd), .A(_2791_), .Y(_2791__bF_buf2) );
BUFX4 BUFX4_1463 ( .gnd(gnd), .vdd(vdd), .A(_2791_), .Y(_2791__bF_buf1) );
BUFX4 BUFX4_1464 ( .gnd(gnd), .vdd(vdd), .A(_2791_), .Y(_2791__bF_buf0) );
BUFX4 BUFX4_1465 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf13) );
BUFX4 BUFX4_1466 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf12) );
BUFX4 BUFX4_1467 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf11) );
BUFX4 BUFX4_1468 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf10) );
BUFX4 BUFX4_1469 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf9) );
BUFX4 BUFX4_1470 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf8) );
BUFX4 BUFX4_1471 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf7) );
BUFX4 BUFX4_1472 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf6) );
BUFX4 BUFX4_1473 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf5) );
BUFX4 BUFX4_1474 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf4) );
BUFX4 BUFX4_1475 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf3) );
BUFX4 BUFX4_1476 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf2) );
BUFX4 BUFX4_1477 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf1) );
BUFX4 BUFX4_1478 ( .gnd(gnd), .vdd(vdd), .A(_14908_), .Y(_14908__bF_buf0) );
BUFX4 BUFX4_1479 ( .gnd(gnd), .vdd(vdd), .A(_14946_), .Y(_14946__bF_buf4) );
BUFX4 BUFX4_1480 ( .gnd(gnd), .vdd(vdd), .A(_14946_), .Y(_14946__bF_buf3) );
BUFX4 BUFX4_1481 ( .gnd(gnd), .vdd(vdd), .A(_14946_), .Y(_14946__bF_buf2) );
BUFX4 BUFX4_1482 ( .gnd(gnd), .vdd(vdd), .A(_14946_), .Y(_14946__bF_buf1) );
BUFX4 BUFX4_1483 ( .gnd(gnd), .vdd(vdd), .A(_14946_), .Y(_14946__bF_buf0) );
BUFX4 BUFX4_1484 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .Y(_14984__bF_buf4) );
BUFX4 BUFX4_1485 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .Y(_14984__bF_buf3) );
BUFX4 BUFX4_1486 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .Y(_14984__bF_buf2) );
BUFX4 BUFX4_1487 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .Y(_14984__bF_buf1) );
BUFX4 BUFX4_1488 ( .gnd(gnd), .vdd(vdd), .A(_14984_), .Y(_14984__bF_buf0) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .Y(_14882_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .B(IDATA_PROG_addr[7]), .Y(_14883_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(IDATA_PROG_addr[4]), .Y(_14884_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14883_), .B(_14884_), .Y(_14885_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf3), .B(IDATA_PROG_addr[2]), .Y(_14886_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(IDATA_PROG_addr[0]), .Y(_14887_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf3), .B(_14887_), .Y(_14888_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf3), .B(_14888__bF_buf3), .Y(_14889_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf15_bF_buf3), .Y(_14890_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(data_255__0_), .Y(_14891_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf14_bF_buf3), .C(_14891_), .Y(_14892_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14890_), .B(IDATA_PROG_data_0_bF_buf4), .C(_14892_), .Y(_14893_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_14893_), .Y(_173__0_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf4), .Y(_14894_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf13_bF_buf3), .B(_14889_), .Y(_14895_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(data_255__1_), .B(_14895__bF_buf3), .Y(_14896_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_14895__bF_buf2), .C(_14896_), .Y(_173__1_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf3), .Y(_14897_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(data_255__2_), .B(_14895__bF_buf1), .Y(_14898_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_14895__bF_buf0), .C(_14898_), .Y(_173__2_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf4), .Y(_14899_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(data_255__3_), .B(_14895__bF_buf3), .Y(_14900_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_14895__bF_buf2), .C(_14900_), .Y(_173__3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(data_255__4_), .Y(_14901_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf4), .Y(_14902_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_14901_), .S(_14895__bF_buf1), .Y(_173__4_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf4), .Y(_14903_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(data_255__5_), .B(_14895__bF_buf0), .Y(_14904_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_14895__bF_buf3), .C(_14904_), .Y(_173__5_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(data_255__6_), .Y(_14905_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf12), .C(_14905_), .Y(_14906_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_14890_), .B(IDATA_PROG_data_6_bF_buf4), .C(_14906_), .Y(_14907_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_14907_), .Y(_173__6_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf5), .Y(_14908_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(data_255__7_), .B(_14895__bF_buf2), .Y(_14909_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_14895__bF_buf1), .C(_14909_), .Y(_173__7_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(data_255__8_), .Y(_14910_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf11), .C(_14910_), .Y(_14911_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14890_), .B(IDATA_PROG_data_8_bF_buf4), .C(_14911_), .Y(_14912_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .Y(_173__8_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf4), .Y(_14913_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(data_255__9_), .B(_14895__bF_buf0), .Y(_14914_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf14), .B(_14895__bF_buf3), .C(_14914_), .Y(_173__9_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(data_255__10_), .Y(_14915_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf10), .C(_14915_), .Y(_14916_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_14890_), .B(IDATA_PROG_data_10_bF_buf4), .C(_14916_), .Y(_14917_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_14917_), .Y(_173__10_) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf4), .Y(_14918_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(data_255__11_), .B(_14895__bF_buf2), .Y(_14919_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_14895__bF_buf1), .C(_14919_), .Y(_173__11_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf4), .Y(_14920_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(data_255__12_), .B(_14895__bF_buf0), .Y(_14921_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_14895__bF_buf3), .C(_14921_), .Y(_173__12_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(data_255__13_), .Y(_14922_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf9), .C(_14922_), .Y(_14923_) );
INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf4), .Y(_14924_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_14895__bF_buf2), .Y(_14925_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_14925_), .B(_14923_), .Y(_173__13_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(data_255__14_), .Y(_14926_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf8), .C(_14926_), .Y(_14927_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_14890_), .B(IDATA_PROG_data_14_bF_buf4), .C(_14927_), .Y(_14928_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_14928_), .Y(_173__14_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(data_255__15_), .Y(_14929_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_14889_), .B(_14882__bF_buf7), .C(_14929_), .Y(_14930_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_14890_), .B(IDATA_PROG_data_15_bF_buf5), .C(_14930_), .Y(_14931_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_14931_), .Y(_173__15_) );
INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf3), .Y(_14932_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(IDATA_PROG_addr[4]), .Y(_14933_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[7]), .Y(_14934_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .B(_14934_), .Y(_14935_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14933_), .B(_14935_), .Y(_14936_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .Y(_14937_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[7]), .B(_14937_), .Y(_14938_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .Y(_14939_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[4]), .B(_14939_), .Y(_14940_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14940_), .Y(_14941_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf2), .B(IDATA_PROG_addr[2]), .Y(_14942_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .B(IDATA_PROG_addr[7]), .Y(_14943_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[4]), .Y(_14944_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(_14944_), .Y(_14945_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_14943_), .B(_14945_), .Y(_14946_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[0]), .Y(_14947_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(_14947_), .Y(_14948_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .Y(_14949_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[0]), .B(_14949_), .Y(_14950_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[2]), .Y(_14951_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf1), .B(_14951_), .Y(_14952_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14950_), .C(_14952__bF_buf4), .Y(_14953_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(IDATA_PROG_addr[0]), .Y(_14954_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(IDATA_PROG_addr[0]), .Y(_14955_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf0), .Y(_14956_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[2]), .B(_14956_), .Y(_14957_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf3), .B(_14954_), .C(_14955_), .D(_14957_), .Y(_14958_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_14953_), .B(_14958_), .Y(_14959_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(_14942__bF_buf3), .C(_14959_), .D(_14946__bF_buf4), .Y(_14960_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf2), .B(_14955_), .Y(_14961_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14950_), .C(_14957_), .Y(_14962_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf3), .B(IDATA_PROG_addr[2]), .Y(_14963_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf3), .B(_14955_), .C(_14957_), .D(_14954_), .Y(_14964_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_14962_), .Y(_14965_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf3), .B(_14961_), .C(_14946__bF_buf3), .Y(_14966_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf3), .B(_14966_), .C(_14960_), .Y(_14967_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(IDATA_PROG_addr[4]), .Y(_14968_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[4]), .B(_14939_), .Y(_14969_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[7]), .B(_14937_), .Y(_14970_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .B(_14968_), .C(_14970_), .Y(_14971_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_14971_), .Y(_14972_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14972_), .B(_14967_), .Y(_14973_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf2), .B(IDATA_PROG_addr[2]), .Y(_14974_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14955_), .C(_14974_), .Y(_14975_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(IDATA_PROG_addr[0]), .Y(_14976_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[2]), .B(_14956_), .Y(_14977_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_14887_), .B(_14974_), .C(_14977__bF_buf3), .D(_14976_), .Y(_14978_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf4), .B(_14975_), .C(_14946__bF_buf2), .Y(_14979_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[0]), .B(_14949_), .Y(_14980_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf1), .B(_14980_), .Y(_14981_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(_14947_), .Y(_14982_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf0), .B(_14982_), .Y(_14983_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_14943_), .B(_14940_), .Y(_14984_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_14983_), .C(_14984__bF_buf4), .Y(_14985_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14976_), .Y(_14986_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf1), .B(_14986_), .C(_14888__bF_buf2), .D(_14984__bF_buf3), .Y(_14987_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14985_), .B(_14987_), .C(_14979_), .Y(_14988_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf1), .B(_14951_), .Y(_14989_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14982_), .C(_14989_), .Y(_14990_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf3), .B(_14976_), .C(_14989_), .D(_14887_), .Y(_14991_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .B(_14990_), .C(_14984__bF_buf2), .Y(_14992_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_14992_), .Y(_14993_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14982_), .C(_14977__bF_buf2), .Y(_14994_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf1), .B(_14994_), .Y(_14995_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_14977__bF_buf1), .B(_14887_), .C(_14976_), .D(_14989_), .Y(_14996_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf0), .B(_14996_), .Y(_14997_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14884_), .B(_14943_), .Y(_14998_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_14939_), .B(_14970_), .C(_14998__bF_buf3), .Y(_14999_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_14999_), .B(_14995_), .C(_14997_), .Y(_15000_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14993_), .B(_15000_), .C(_14988_), .Y(_15001_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .B(IDATA_PROG_addr[7]), .Y(_15002_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_15002_), .B(_14968_), .Y(_15003_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_15003_), .Y(_15004_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(_14944_), .C(_15002_), .Y(_15005_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14939_), .B(IDATA_PROG_addr[4]), .C(_15002_), .Y(_15006_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf4), .B(_14942__bF_buf2), .C(_15005__bF_buf3), .Y(_15007_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_15007_), .B(_15004_), .Y(_15008_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf3), .B(_14975_), .C(_14984__bF_buf4), .Y(_15009_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .B(IDATA_PROG_addr[7]), .Y(_15010_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_14933_), .B(_15010_), .Y(_15011_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_14983_), .C(_15011__bF_buf3), .Y(_15012_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf1), .B(_15011__bF_buf2), .C(_14984__bF_buf3), .D(_14986_), .Y(_15013_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_15012_), .B(_15013_), .C(_15009_), .Y(_15014_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .B(_14990_), .C(_15011__bF_buf1), .Y(_15015_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_14994_), .C(_15011__bF_buf0), .Y(_15016_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_15015_), .B(_15016_), .Y(_15017_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_15017_), .B(_15008_), .C(_15014_), .Y(_15018_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_14935_), .B(_14969_), .Y(_15019_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(_14944_), .Y(_15020_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14935_), .C(_15020_), .Y(_15021_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_14968_), .B(_14942__bF_buf1), .C(_14935_), .Y(_15022_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf3), .B(_15022_), .C(_15021_), .Y(_15023_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_15002_), .B(_14942__bF_buf0), .C(_15020_), .Y(_15024_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14933_), .B(_15002_), .Y(_15025_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_14968_), .B(_14974_), .C(_14935_), .Y(_15026_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf4), .B(_15024_), .C(_15026_), .Y(_15027_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_15023_), .B(_15027_), .Y(_15028_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf2), .B(_14975_), .C(_15011__bF_buf3), .Y(_15029_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf3), .B(_14955_), .Y(_15030_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_14933_), .B(_15010_), .Y(_15031_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_15031__bF_buf3), .Y(_15032_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(_15032_), .Y(_15033_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf0), .B(IDATA_PROG_addr[2]), .Y(_15034_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .Y(_15035_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf2), .B(_14950_), .Y(_15036_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_15036_), .C(_14885__bF_buf2), .Y(_15037_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_15029_), .C(_15037_), .Y(_15038_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_15038_), .B(_15028_), .Y(_15039_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .B(_15039_), .Y(_15040_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_15001_), .C(_15040_), .Y(_15041_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf6), .B(_15041_), .Y(_15042_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(data_254__0_), .B(_15042__bF_buf3), .Y(_15043_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_15042__bF_buf2), .C(_15043_), .Y(_172__0_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(data_254__1_), .B(_15042__bF_buf1), .Y(_15044_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_15042__bF_buf0), .C(_15044_), .Y(_172__1_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(data_254__2_), .Y(_15045_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf13), .B(_15045_), .S(_15042__bF_buf3), .Y(_172__2_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(data_254__3_), .B(_15042__bF_buf2), .Y(_15046_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_15042__bF_buf1), .C(_15046_), .Y(_172__3_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(data_254__4_), .B(_15042__bF_buf0), .Y(_15047_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_15042__bF_buf3), .C(_15047_), .Y(_172__4_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(data_254__5_), .B(_15042__bF_buf2), .Y(_15048_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_15042__bF_buf1), .C(_15048_), .Y(_172__5_) );
INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf3), .Y(_15049_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(data_254__6_), .Y(_15050_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_15050_), .S(_15042__bF_buf0), .Y(_172__6_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(data_254__7_), .B(_15042__bF_buf3), .Y(_15051_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_15042__bF_buf2), .C(_15051_), .Y(_172__7_) );
INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf3), .Y(_15052_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(data_254__8_), .Y(_15053_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_15053_), .S(_15042__bF_buf1), .Y(_172__8_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(data_254__9_), .Y(_15054_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_15054_), .S(_15042__bF_buf0), .Y(_172__9_) );
INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf3), .Y(_15055_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(data_254__10_), .Y(_15056_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_15056_), .S(_15042__bF_buf3), .Y(_172__10_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(data_254__11_), .B(_15042__bF_buf2), .Y(_15057_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_15042__bF_buf1), .C(_15057_), .Y(_172__11_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(data_254__12_), .B(_15042__bF_buf0), .Y(_15058_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_15042__bF_buf3), .C(_15058_), .Y(_172__12_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(data_254__13_), .Y(_15059_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_15059_), .S(_15042__bF_buf2), .Y(_172__13_) );
INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf3), .Y(_15060_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(data_254__14_), .Y(_15061_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf14), .B(_15061_), .S(_15042__bF_buf1), .Y(_172__14_) );
INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf4), .Y(_15062_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(data_254__15_), .Y(_15063_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_15063_), .S(_15042__bF_buf0), .Y(_172__15_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14939_), .B(_14944_), .Y(_15064_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_15064_), .Y(_15065_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14935_), .B(_15020_), .Y(_15066_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_14994_), .C(_14946__bF_buf0), .Y(_15067_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf3), .B(_14974_), .C(_15067_), .Y(_15068_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_14961_), .B(_14946__bF_buf4), .Y(_15069_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf3), .B(_14990_), .Y(_15070_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf2), .B(_14991_), .Y(_15071_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_15069_), .B(_15070_), .C(_15071_), .Y(_15072_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf3), .B(_15072_), .C(_15068_), .Y(_15073_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_14971_), .C(_15001_), .Y(_15074_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_15029_), .Y(_15075_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf1), .B(_14888__bF_buf0), .C(_15032_), .Y(_15076_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14955_), .B(_14963__bF_buf2), .Y(_15077_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf1), .B(_14982_), .C(_15077_), .Y(_15078_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .B(_15035_), .C(_14885__bF_buf0), .Y(_15079_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_15076_), .B(_15079_), .Y(_15080_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_15075_), .B(_15080_), .Y(_15081_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf5), .B(_15023_), .Y(_15082_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_15082_), .Y(_15083_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_15027_), .B(_15083_), .Y(_15084_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .B(_15081_), .C(_15084_), .Y(_15085_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf12), .B(_15085_), .Y(_15086_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_15086__bF_buf4), .Y(_15087_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(data_253__0_), .B(_15086__bF_buf3), .C(_15087_), .Y(_15088_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_15088_), .Y(_171__0_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_15086__bF_buf2), .Y(_15089_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(data_253__1_), .B(_15086__bF_buf1), .C(_15089_), .Y(_15090_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_15090_), .Y(_171__1_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf12), .B(_15086__bF_buf0), .Y(_15091_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(data_253__2_), .B(_15086__bF_buf4), .C(_15091_), .Y(_15092_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_15092_), .Y(_171__2_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_15086__bF_buf3), .Y(_15093_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(data_253__3_), .B(_15086__bF_buf2), .C(_15093_), .Y(_15094_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_15094_), .Y(_171__3_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_15086__bF_buf1), .Y(_15095_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(data_253__4_), .B(_15086__bF_buf0), .C(_15095_), .Y(_15096_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_15096_), .Y(_171__4_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_15086__bF_buf4), .Y(_15097_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(data_253__5_), .B(_15086__bF_buf3), .C(_15097_), .Y(_15098_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_15098_), .Y(_171__5_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_15086__bF_buf2), .Y(_15099_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(data_253__6_), .B(_15086__bF_buf1), .C(_15099_), .Y(_15100_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .Y(_171__6_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_15086__bF_buf0), .Y(_15101_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(data_253__7_), .B(_15086__bF_buf4), .C(_15101_), .Y(_15102_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_15102_), .Y(_171__7_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_15086__bF_buf3), .Y(_15103_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(data_253__8_), .B(_15086__bF_buf2), .C(_15103_), .Y(_15104_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_15104_), .Y(_171__8_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_15086__bF_buf1), .Y(_15105_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(data_253__9_), .B(_15086__bF_buf0), .C(_15105_), .Y(_15106_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_15106_), .Y(_171__9_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_15086__bF_buf4), .Y(_15107_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(data_253__10_), .B(_15086__bF_buf3), .C(_15107_), .Y(_15108_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_15108_), .Y(_171__10_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_15086__bF_buf2), .Y(_15109_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(data_253__11_), .B(_15086__bF_buf1), .C(_15109_), .Y(_15110_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_15110_), .Y(_171__11_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_15086__bF_buf0), .Y(_15111_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(data_253__12_), .B(_15086__bF_buf4), .C(_15111_), .Y(_15112_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_15112_), .Y(_171__12_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_15086__bF_buf3), .Y(_15113_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(data_253__13_), .B(_15086__bF_buf2), .C(_15113_), .Y(_15114_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_15114_), .Y(_171__13_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_15086__bF_buf1), .Y(_15115_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(data_253__14_), .B(_15086__bF_buf0), .C(_15115_), .Y(_15116_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_15116_), .Y(_171__14_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_15086__bF_buf4), .Y(_15117_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(data_253__15_), .B(_15086__bF_buf3), .C(_15117_), .Y(_15118_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_15118_), .Y(_171__15_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(data_252__0_), .Y(_15119_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_15023_), .B(_15027_), .Y(_15120_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_14983_), .C(_14885__bF_buf3), .Y(_15121_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_15029_), .B(_15121_), .C(_15076_), .Y(_15122_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_15034_), .C(IDATA_PROG_write_bF_buf7), .Y(_15123_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_15123_), .B(_15122_), .Y(_15124_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf3), .B(_15124_), .C(_15018_), .Y(_15125_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf11), .B(_15125_), .Y(_15126_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_15119_), .S(_15126_), .Y(_170__0_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(data_252__1_), .Y(_15127_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_15127_), .S(_15126_), .Y(_170__1_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(data_252__2_), .Y(_15128_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf10), .B(_15125_), .C(_15128_), .Y(_15129_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_15126_), .Y(_15130_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_15130_), .B(_15129_), .Y(_170__2_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(data_252__3_), .Y(_15131_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_15131_), .S(_15126_), .Y(_170__3_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(data_252__4_), .Y(_15132_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_15132_), .S(_15126_), .Y(_170__4_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(data_252__5_), .Y(_15133_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_15133_), .S(_15126_), .Y(_170__5_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(data_252__6_), .Y(_15134_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf9), .B(_15125_), .C(_15134_), .Y(_15135_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_15126_), .Y(_15136_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_15136_), .B(_15135_), .Y(_170__6_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(data_252__7_), .Y(_15137_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_15137_), .S(_15126_), .Y(_170__7_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(data_252__8_), .Y(_15138_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf8), .B(_15125_), .C(_15138_), .Y(_15139_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_15126_), .Y(_15140_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_15140_), .B(_15139_), .Y(_170__8_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(data_252__9_), .Y(_15141_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf7), .B(_15125_), .C(_15141_), .Y(_15142_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_15126_), .Y(_15143_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_15143_), .B(_15142_), .Y(_170__9_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(data_252__10_), .Y(_15144_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf6), .B(_15125_), .C(_15144_), .Y(_15145_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_15126_), .Y(_15146_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_15146_), .B(_15145_), .Y(_170__10_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(data_252__11_), .Y(_15147_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_15147_), .S(_15126_), .Y(_170__11_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(data_252__12_), .Y(_15148_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_15148_), .S(_15126_), .Y(_170__12_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(data_252__13_), .Y(_15149_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf5), .B(_15125_), .C(_15149_), .Y(_15150_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_15126_), .Y(_15151_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_15151_), .B(_15150_), .Y(_170__13_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(data_252__14_), .Y(_15152_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf4), .B(_15125_), .C(_15152_), .Y(_15153_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_15126_), .Y(_15154_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_15154_), .B(_15153_), .Y(_170__14_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(data_252__15_), .Y(_15155_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf3), .B(_15125_), .C(_15155_), .Y(_15156_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_15126_), .Y(_15157_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_15157_), .B(_15156_), .Y(_170__15_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(data_251__0_), .Y(_15158_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .Y(_15159_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14955_), .C(_14957_), .Y(_15160_) );
INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .Y(_15161_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf2), .B(_15161_), .C(_15122_), .Y(_15162_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14989_), .C(_15077_), .Y(_15163_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf1), .B(_15163_), .Y(_15164_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf2), .B(_14885__bF_buf0), .C(_14882__bF_buf4), .Y(_15165_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf2), .B(_15165_), .Y(_15166_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_15164_), .B(_15166_), .C(_15162_), .Y(_15167_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_15167_), .B(_15159_), .Y(_15168_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf2), .C(_15158_), .Y(_15169_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[5]), .B(_14944_), .C(_15010_), .Y(_15170_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14887_), .B(_14942__bF_buf2), .C(_14976_), .Y(_15171_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14942__bF_buf1), .C(_14952__bF_buf1), .D(_14955_), .Y(_15172_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_15171_), .B(_15172_), .C(_15170__bF_buf3), .Y(_15173_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf1), .B(_14887_), .C(_14976_), .Y(_15174_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_15010_), .B(_15020_), .Y(_15175_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15175__bF_buf4), .Y(_15176_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf0), .B(_14954_), .Y(_15177_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_15170__bF_buf2), .C(_15175__bF_buf3), .D(_15177_), .Y(_15178_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15176_), .B(_15178_), .C(_15173_), .Y(_15179_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_14958_), .B(_15175__bF_buf2), .C(_14999_), .Y(_15180_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_14994_), .B(_14984__bF_buf2), .C(_15180_), .Y(_15181_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_14992_), .B(_15181_), .C(_15179_), .Y(_15182_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .B(_14972_), .C(_15182_), .Y(_15183_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_15159_), .B(_15167_), .Y(_15184_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_15183__bF_buf8), .C(_15184_), .Y(_15185_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_15169_), .B(_15185_), .Y(_169__0_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(data_251__1_), .Y(_15186_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf1), .C(_15186_), .Y(_15187_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_15183__bF_buf7), .C(_15184_), .Y(_15188_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_15187_), .B(_15188_), .Y(_169__1_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(data_251__2_), .Y(_15189_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf0), .C(_15189_), .Y(_15190_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_15183__bF_buf6), .C(_15184_), .Y(_15191_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_15190_), .B(_15191_), .Y(_169__2_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(data_251__3_), .Y(_15192_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf12), .C(_15192_), .Y(_15193_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_15183__bF_buf5), .C(_15184_), .Y(_15194_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_15193_), .B(_15194_), .Y(_169__3_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(data_251__4_), .Y(_15195_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf11), .C(_15195_), .Y(_15196_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_15183__bF_buf4), .C(_15184_), .Y(_15197_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_15196_), .B(_15197_), .Y(_169__4_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(data_251__5_), .Y(_15198_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf10), .C(_15198_), .Y(_15199_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_15183__bF_buf3), .C(_15184_), .Y(_15200_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_15199_), .B(_15200_), .Y(_169__5_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(data_251__6_), .Y(_15201_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf9), .C(_15201_), .Y(_15202_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_15183__bF_buf2), .C(_15184_), .Y(_15203_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_15202_), .B(_15203_), .Y(_169__6_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(data_251__7_), .Y(_15204_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf8), .C(_15204_), .Y(_15205_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_15183__bF_buf1), .C(_15184_), .Y(_15206_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_15205_), .B(_15206_), .Y(_169__7_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(data_251__8_), .Y(_15207_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf7), .C(_15207_), .Y(_15208_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_15183__bF_buf0), .C(_15184_), .Y(_15209_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_15208_), .B(_15209_), .Y(_169__8_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(data_251__9_), .Y(_15210_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf6), .C(_15210_), .Y(_15211_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_15183__bF_buf8), .C(_15184_), .Y(_15212_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_15211_), .B(_15212_), .Y(_169__9_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(data_251__10_), .Y(_15213_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf5), .C(_15213_), .Y(_15214_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_15183__bF_buf7), .C(_15184_), .Y(_15215_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_15214_), .B(_15215_), .Y(_169__10_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(data_251__11_), .Y(_15216_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf4), .C(_15216_), .Y(_15217_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_15183__bF_buf6), .C(_15184_), .Y(_15218_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_15217_), .B(_15218_), .Y(_169__11_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(data_251__12_), .Y(_15219_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf3), .C(_15219_), .Y(_15220_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_15183__bF_buf5), .C(_15184_), .Y(_15221_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_15220_), .B(_15221_), .Y(_169__12_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(data_251__13_), .Y(_15222_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf2), .C(_15222_), .Y(_15223_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_15183__bF_buf4), .C(_15184_), .Y(_15224_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_15223_), .B(_15224_), .Y(_169__13_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(data_251__14_), .Y(_15225_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf1), .C(_15225_), .Y(_15226_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_15183__bF_buf3), .C(_15184_), .Y(_15227_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_15226_), .B(_15227_), .Y(_169__14_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(data_251__15_), .Y(_15228_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_15168_), .B(_15074__bF_buf0), .C(_15228_), .Y(_15229_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf10), .B(_15183__bF_buf2), .C(_15184_), .Y(_15230_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_15229_), .B(_15230_), .Y(_169__15_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(data_250__0_), .Y(_15231_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_15165_), .B(_15120__bF_buf1), .Y(_15232_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_14964_), .Y(_15233_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_15233_), .B(_15232_), .Y(_15234_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .B(_15162_), .C(_15234_), .Y(_15235_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf3), .B(_15074__bF_buf12), .C(_15231_), .Y(_15236_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf11), .B(_15235__bF_buf2), .Y(_15237_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_15237_), .Y(_15238_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_15238_), .B(_15236_), .Y(_168__0_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(data_250__1_), .Y(_15239_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf1), .B(_15074__bF_buf10), .C(_15239_), .Y(_15240_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_15237_), .Y(_15241_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_15241_), .B(_15240_), .Y(_168__1_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(data_250__2_), .Y(_15242_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf0), .B(_15074__bF_buf9), .C(_15242_), .Y(_15243_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_15237_), .Y(_15244_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_15244_), .B(_15243_), .Y(_168__2_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(data_250__3_), .Y(_15245_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf3), .B(_15074__bF_buf8), .C(_15245_), .Y(_15246_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_15237_), .Y(_15247_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_15247_), .B(_15246_), .Y(_168__3_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(data_250__4_), .Y(_15248_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf2), .B(_15074__bF_buf7), .C(_15248_), .Y(_15249_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_15237_), .Y(_15250_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_15250_), .B(_15249_), .Y(_168__4_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(data_250__5_), .Y(_15251_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf1), .B(_15074__bF_buf6), .C(_15251_), .Y(_15252_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_15237_), .Y(_15253_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_15253_), .B(_15252_), .Y(_168__5_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(data_250__6_), .Y(_15254_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf0), .B(_15074__bF_buf5), .C(_15254_), .Y(_15255_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_15237_), .Y(_15256_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_15256_), .B(_15255_), .Y(_168__6_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(data_250__7_), .Y(_15257_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf3), .B(_15074__bF_buf4), .C(_15257_), .Y(_15258_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_15237_), .Y(_15259_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_15259_), .B(_15258_), .Y(_168__7_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(data_250__8_), .Y(_15260_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf2), .B(_15074__bF_buf3), .C(_15260_), .Y(_15261_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_15237_), .Y(_15262_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_15262_), .B(_15261_), .Y(_168__8_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(data_250__9_), .Y(_15263_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf1), .B(_15074__bF_buf2), .C(_15263_), .Y(_15264_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_15237_), .Y(_15265_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_15265_), .B(_15264_), .Y(_168__9_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(data_250__10_), .Y(_15266_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf0), .B(_15074__bF_buf1), .C(_15266_), .Y(_15267_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_15237_), .Y(_15268_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_15268_), .B(_15267_), .Y(_168__10_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(data_250__11_), .Y(_15269_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf3), .B(_15074__bF_buf0), .C(_15269_), .Y(_15270_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_15237_), .Y(_15271_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_15271_), .B(_15270_), .Y(_168__11_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(data_250__12_), .Y(_15272_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf2), .B(_15074__bF_buf12), .C(_15272_), .Y(_15273_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_15237_), .Y(_15274_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_15274_), .B(_15273_), .Y(_168__12_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(data_250__13_), .Y(_15275_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf1), .B(_15074__bF_buf11), .C(_15275_), .Y(_15276_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_15237_), .Y(_15277_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_15277_), .B(_15276_), .Y(_168__13_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(data_250__14_), .Y(_15278_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf0), .B(_15074__bF_buf10), .C(_15278_), .Y(_15279_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_15237_), .Y(_15280_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_15280_), .B(_15279_), .Y(_168__14_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(data_250__15_), .Y(_15281_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_15235__bF_buf3), .B(_15074__bF_buf9), .C(_15281_), .Y(_15282_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_15237_), .Y(_15283_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_15283_), .B(_15282_), .Y(_168__15_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_14955_), .B(_14957_), .Y(_15284_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14989_), .C(_15284_), .Y(_15285_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf3), .B(_15285_), .C(_15122_), .Y(_15286_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .B(_15286_), .C(_15234_), .Y(_15287_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf8), .B(_15287_), .Y(_15288_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_15288_), .Y(_15289_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(data_249__0_), .B(_15288_), .C(_15289_), .Y(_15290_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_15290_), .Y(_166__0_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_15288_), .Y(_15291_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(data_249__1_), .B(_15288_), .C(_15291_), .Y(_15292_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_15292_), .Y(_166__1_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(data_249__2_), .Y(_15293_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf7), .C(_15293_), .Y(_15294_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_14964_), .C(_15166_), .Y(_15295_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_15286_), .B(_15018_), .Y(_15296_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_15295_), .B(_15296_), .Y(_15297_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_15183__bF_buf1), .C(_15297_), .Y(_15298_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_15298_), .B(_15294_), .Y(_166__2_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_15288_), .Y(_15299_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(data_249__3_), .B(_15288_), .C(_15299_), .Y(_15300_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_15300_), .Y(_166__3_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_15288_), .Y(_15301_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(data_249__4_), .B(_15288_), .C(_15301_), .Y(_15302_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_15302_), .Y(_166__4_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_15288_), .Y(_15303_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(data_249__5_), .B(_15288_), .C(_15303_), .Y(_15304_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_15304_), .Y(_166__5_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(data_249__6_), .Y(_15305_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf6), .C(_15305_), .Y(_15306_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_15183__bF_buf0), .C(_15297_), .Y(_15307_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_15307_), .B(_15306_), .Y(_166__6_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_15288_), .Y(_15308_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(data_249__7_), .B(_15288_), .C(_15308_), .Y(_15309_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_15309_), .Y(_166__7_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(data_249__8_), .Y(_15310_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf5), .C(_15310_), .Y(_15311_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_15183__bF_buf8), .C(_15297_), .Y(_15312_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_15312_), .B(_15311_), .Y(_166__8_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(data_249__9_), .Y(_15313_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf4), .C(_15313_), .Y(_15314_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_15183__bF_buf7), .C(_15297_), .Y(_15315_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_15315_), .B(_15314_), .Y(_166__9_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(data_249__10_), .Y(_15316_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf3), .C(_15316_), .Y(_15317_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_15183__bF_buf6), .C(_15297_), .Y(_15318_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_15318_), .B(_15317_), .Y(_166__10_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_15288_), .Y(_15319_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(data_249__11_), .B(_15288_), .C(_15319_), .Y(_15320_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_15320_), .Y(_166__11_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_15288_), .Y(_15321_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(data_249__12_), .B(_15288_), .C(_15321_), .Y(_15322_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_15322_), .Y(_166__12_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(data_249__13_), .Y(_15323_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf2), .C(_15323_), .Y(_15324_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_15183__bF_buf5), .C(_15297_), .Y(_15325_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_15325_), .B(_15324_), .Y(_166__13_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(data_249__14_), .Y(_15326_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf1), .C(_15326_), .Y(_15327_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_15183__bF_buf4), .C(_15297_), .Y(_15328_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_15328_), .B(_15327_), .Y(_166__14_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(data_249__15_), .Y(_15329_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_15287_), .B(_15074__bF_buf0), .C(_15329_), .Y(_15330_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_15183__bF_buf3), .C(_15297_), .Y(_15331_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_15331_), .B(_15330_), .Y(_166__15_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(data_248__0_), .Y(_15332_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf2), .B(_14965__bF_buf2), .C(_15122_), .Y(_15333_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_15333_), .B(_15166_), .C(_15018_), .Y(_15334_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf12), .B(_15334_), .Y(_15335_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_15332_), .S(_15335__bF_buf3), .Y(_165__0_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(data_248__1_), .Y(_15336_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_15336_), .S(_15335__bF_buf2), .Y(_165__1_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_15335__bF_buf1), .Y(_15337_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(data_248__2_), .B(_15335__bF_buf0), .C(_15337_), .Y(_15338_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_15338_), .Y(_165__2_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(data_248__3_), .Y(_15339_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_15339_), .S(_15335__bF_buf3), .Y(_165__3_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(data_248__4_), .Y(_15340_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_15340_), .S(_15335__bF_buf2), .Y(_165__4_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(data_248__5_), .Y(_15341_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_15341_), .S(_15335__bF_buf1), .Y(_165__5_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_15335__bF_buf0), .Y(_15342_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(data_248__6_), .B(_15335__bF_buf3), .C(_15342_), .Y(_15343_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_15343_), .Y(_165__6_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(data_248__7_), .Y(_15344_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_15344_), .S(_15335__bF_buf2), .Y(_165__7_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_15335__bF_buf1), .Y(_15345_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(data_248__8_), .B(_15335__bF_buf0), .C(_15345_), .Y(_15346_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_15346_), .Y(_165__8_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf7), .B(_15335__bF_buf3), .Y(_15347_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(data_248__9_), .B(_15335__bF_buf2), .C(_15347_), .Y(_15348_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_15348_), .Y(_165__9_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_15335__bF_buf1), .Y(_15349_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(data_248__10_), .B(_15335__bF_buf0), .C(_15349_), .Y(_15350_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_15350_), .Y(_165__10_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(data_248__11_), .Y(_15351_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_15351_), .S(_15335__bF_buf3), .Y(_165__11_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(data_248__12_), .Y(_15352_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_15352_), .S(_15335__bF_buf2), .Y(_165__12_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_15335__bF_buf1), .Y(_15353_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(data_248__13_), .B(_15335__bF_buf0), .C(_15353_), .Y(_15354_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_15354_), .Y(_165__13_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_15335__bF_buf3), .Y(_15355_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(data_248__14_), .B(_15335__bF_buf2), .C(_15355_), .Y(_15356_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_15356_), .Y(_165__14_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_15335__bF_buf1), .Y(_15357_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(data_248__15_), .B(_15335__bF_buf0), .C(_15357_), .Y(_15358_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_15358_), .Y(_165__15_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(data_247__0_), .Y(_15359_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14955_), .C(_14952__bF_buf0), .Y(_15360_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_15360_), .B(_15003_), .C(IDATA_PROG_write_bF_buf6), .Y(_15361_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_15361_), .B(_15028_), .Y(_15362_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14977__bF_buf0), .C(_15284_), .Y(_15363_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf1), .B(_15363_), .Y(_15364_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf1), .B(_15364_), .C(_15122_), .Y(_15365_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_15365_), .B(_15362_), .C(_15018_), .Y(_15366_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf11), .B(_15366_), .Y(_15367_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_15359_), .S(_15367__bF_buf3), .Y(_164__0_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(data_247__1_), .Y(_15368_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_15368_), .S(_15367__bF_buf2), .Y(_164__1_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(data_247__2_), .Y(_15369_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf10), .C(_15369_), .Y(_15370_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_15367__bF_buf1), .Y(_15371_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_15371_), .B(_15370_), .Y(_164__2_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(data_247__3_), .Y(_15372_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_15372_), .S(_15367__bF_buf0), .Y(_164__3_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(data_247__4_), .Y(_15373_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_15373_), .S(_15367__bF_buf3), .Y(_164__4_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(data_247__5_), .Y(_15374_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_15374_), .S(_15367__bF_buf2), .Y(_164__5_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(data_247__6_), .Y(_15375_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf9), .C(_15375_), .Y(_15376_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_15367__bF_buf1), .Y(_15377_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_15377_), .B(_15376_), .Y(_164__6_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(data_247__7_), .Y(_15378_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_15378_), .S(_15367__bF_buf0), .Y(_164__7_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(data_247__8_), .Y(_15379_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf8), .C(_15379_), .Y(_15380_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_15367__bF_buf3), .Y(_15381_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_15381_), .B(_15380_), .Y(_164__8_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(data_247__9_), .Y(_15382_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf7), .C(_15382_), .Y(_15383_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_15367__bF_buf2), .Y(_15384_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_15384_), .B(_15383_), .Y(_164__9_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(data_247__10_), .Y(_15385_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf6), .C(_15385_), .Y(_15386_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_15367__bF_buf1), .Y(_15387_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_15387_), .B(_15386_), .Y(_164__10_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(data_247__11_), .Y(_15388_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_15388_), .S(_15367__bF_buf0), .Y(_164__11_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(data_247__12_), .Y(_15389_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_15389_), .S(_15367__bF_buf3), .Y(_164__12_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(data_247__13_), .Y(_15390_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf5), .C(_15390_), .Y(_15391_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_15367__bF_buf2), .Y(_15392_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_15392_), .B(_15391_), .Y(_164__13_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(data_247__14_), .Y(_15393_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_15366_), .B(_15074__bF_buf4), .C(_15393_), .Y(_15394_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_15367__bF_buf1), .Y(_15395_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_15395_), .B(_15394_), .Y(_164__14_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_15367__bF_buf0), .B(data_247__15_), .Y(_15396_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_15367__bF_buf3), .Y(_15397_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_15396_), .B(_15397_), .Y(_164__15_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(data_246__0_), .Y(_15398_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf0), .B(_15018_), .Y(_15399_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_14958_), .Y(_15400_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_15400_), .B(_15361_), .Y(_15401_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_15401_), .B(_15333_), .Y(_15402_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_15399_), .B(_15402_), .Y(_15403_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf3), .C(_15398_), .Y(_15404_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_15402_), .B(_15399_), .Y(_15405_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_15183__bF_buf2), .C(_15405_), .Y(_15406_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_15404_), .B(_15406_), .Y(_163__0_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(data_246__1_), .Y(_15407_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf2), .C(_15407_), .Y(_15408_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_15183__bF_buf1), .C(_15405_), .Y(_15409_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_15408_), .B(_15409_), .Y(_163__1_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(data_246__2_), .Y(_15410_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf1), .C(_15410_), .Y(_15411_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_15183__bF_buf0), .C(_15405_), .Y(_15412_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_15411_), .B(_15412_), .Y(_163__2_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(data_246__3_), .Y(_15413_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf0), .C(_15413_), .Y(_15414_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_15183__bF_buf8), .C(_15405_), .Y(_15415_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_15414_), .B(_15415_), .Y(_163__3_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(data_246__4_), .Y(_15416_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf12), .C(_15416_), .Y(_15417_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_15183__bF_buf7), .C(_15405_), .Y(_15418_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_15417_), .B(_15418_), .Y(_163__4_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(data_246__5_), .Y(_15419_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf11), .C(_15419_), .Y(_15420_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_15183__bF_buf6), .C(_15405_), .Y(_15421_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_15420_), .B(_15421_), .Y(_163__5_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(data_246__6_), .Y(_15422_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf10), .C(_15422_), .Y(_15423_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_15183__bF_buf5), .C(_15405_), .Y(_15424_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_15423_), .B(_15424_), .Y(_163__6_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(data_246__7_), .Y(_15425_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf9), .C(_15425_), .Y(_15426_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_15183__bF_buf4), .C(_15405_), .Y(_15427_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_15426_), .B(_15427_), .Y(_163__7_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(data_246__8_), .Y(_15428_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf8), .C(_15428_), .Y(_15429_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_15183__bF_buf3), .C(_15405_), .Y(_15430_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_15429_), .B(_15430_), .Y(_163__8_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(data_246__9_), .Y(_15431_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf7), .C(_15431_), .Y(_15432_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_15183__bF_buf2), .C(_15405_), .Y(_15433_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_15432_), .B(_15433_), .Y(_163__9_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(data_246__10_), .Y(_15434_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf6), .C(_15434_), .Y(_15435_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_15183__bF_buf1), .C(_15405_), .Y(_15436_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_15435_), .B(_15436_), .Y(_163__10_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(data_246__11_), .Y(_15437_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf5), .C(_15437_), .Y(_15438_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_15183__bF_buf0), .C(_15405_), .Y(_15439_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_15438_), .B(_15439_), .Y(_163__11_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(data_246__12_), .Y(_15440_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf4), .C(_15440_), .Y(_15441_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_15183__bF_buf8), .C(_15405_), .Y(_15442_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_15441_), .B(_15442_), .Y(_163__12_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(data_246__13_), .Y(_15443_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf3), .C(_15443_), .Y(_15444_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_15183__bF_buf7), .C(_15405_), .Y(_15445_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_15444_), .B(_15445_), .Y(_163__13_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(data_246__14_), .Y(_15446_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf2), .C(_15446_), .Y(_15447_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_15183__bF_buf6), .C(_15405_), .Y(_15448_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_15447_), .B(_15448_), .Y(_163__14_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(data_246__15_), .Y(_15449_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_15403_), .B(_15074__bF_buf1), .C(_15449_), .Y(_15450_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_15183__bF_buf5), .C(_15405_), .Y(_15451_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_15450_), .B(_15451_), .Y(_163__15_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(data_245__0_), .Y(_15452_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_14950_), .B(_14955_), .C(_14952__bF_buf4), .Y(_15453_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_15453_), .B(_15003_), .C(IDATA_PROG_write_bF_buf5), .Y(_15454_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_15400_), .B(_15454_), .Y(_15455_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_15455_), .B(_15120__bF_buf3), .Y(_15456_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_15333_), .B(_15456_), .C(_15018_), .Y(_15457_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf0), .B(_15457__bF_buf3), .C(_15452_), .Y(_15458_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf12), .B(_15457__bF_buf2), .Y(_15459_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_15459_), .Y(_15460_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_15460_), .B(_15458_), .Y(_162__0_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(data_245__1_), .Y(_15461_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf11), .B(_15457__bF_buf1), .C(_15461_), .Y(_15462_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_15459_), .Y(_15463_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_15463_), .B(_15462_), .Y(_162__1_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(data_245__2_), .Y(_15464_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf10), .B(_15457__bF_buf0), .C(_15464_), .Y(_15465_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_15459_), .Y(_15466_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_15466_), .B(_15465_), .Y(_162__2_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(data_245__3_), .Y(_15467_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf9), .B(_15457__bF_buf3), .C(_15467_), .Y(_15468_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_15459_), .Y(_15469_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_15469_), .B(_15468_), .Y(_162__3_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(data_245__4_), .Y(_15470_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf8), .B(_15457__bF_buf2), .C(_15470_), .Y(_15471_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_15459_), .Y(_15472_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_15472_), .B(_15471_), .Y(_162__4_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(data_245__5_), .Y(_15473_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf7), .B(_15457__bF_buf1), .C(_15473_), .Y(_15474_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_15459_), .Y(_15475_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_15475_), .B(_15474_), .Y(_162__5_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(data_245__6_), .Y(_15476_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf6), .B(_15457__bF_buf0), .C(_15476_), .Y(_15477_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_15459_), .Y(_15478_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_15478_), .B(_15477_), .Y(_162__6_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(data_245__7_), .Y(_15479_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf5), .B(_15457__bF_buf3), .C(_15479_), .Y(_15480_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_15459_), .Y(_15481_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_15481_), .B(_15480_), .Y(_162__7_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(data_245__8_), .Y(_15482_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf4), .B(_15457__bF_buf2), .C(_15482_), .Y(_15483_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_15459_), .Y(_15484_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_15484_), .B(_15483_), .Y(_162__8_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(data_245__9_), .Y(_15485_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf3), .B(_15457__bF_buf1), .C(_15485_), .Y(_15486_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_15459_), .Y(_15487_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_15487_), .B(_15486_), .Y(_162__9_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(data_245__10_), .Y(_15488_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf2), .B(_15457__bF_buf0), .C(_15488_), .Y(_15489_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_15459_), .Y(_15490_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_15490_), .B(_15489_), .Y(_162__10_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(data_245__11_), .Y(_15491_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf1), .B(_15457__bF_buf3), .C(_15491_), .Y(_15492_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_15459_), .Y(_15493_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_15493_), .B(_15492_), .Y(_162__11_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(data_245__12_), .Y(_15494_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf0), .B(_15457__bF_buf2), .C(_15494_), .Y(_15495_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_15459_), .Y(_15496_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_15496_), .B(_15495_), .Y(_162__12_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(data_245__13_), .Y(_15497_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf12), .B(_15457__bF_buf1), .C(_15497_), .Y(_15498_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_15459_), .Y(_15499_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_15499_), .B(_15498_), .Y(_162__13_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(data_245__14_), .Y(_15500_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf11), .B(_15457__bF_buf0), .C(_15500_), .Y(_15501_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf5), .B(_15459_), .Y(_15502_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_15502_), .B(_15501_), .Y(_162__14_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(data_245__15_), .Y(_15503_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf10), .B(_15457__bF_buf3), .C(_15503_), .Y(_15504_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_15459_), .Y(_15505_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_15505_), .B(_15504_), .Y(_162__15_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(data_244__0_), .Y(_15506_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_15017_), .B(_15014_), .Y(_15507_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_14994_), .B(_14996_), .Y(_15508_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_14990_), .B(_14991_), .Y(_15509_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_15509_), .B(_15508_), .C(_15003_), .Y(_15510_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_15510_), .B(_15122_), .Y(_15511_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_15004_), .B(_15007_), .Y(_15512_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_15512_), .Y(_15513_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_15513_), .Y(_15514_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_15507_), .B(_15511_), .C(_15514_), .Y(_15515_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf3), .B(_15074__bF_buf9), .C(_15506_), .Y(_15516_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf8), .B(_15515__bF_buf2), .Y(_15517_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_15517_), .Y(_15518_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_15518_), .B(_15516_), .Y(_161__0_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(data_244__1_), .Y(_15519_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf1), .B(_15074__bF_buf7), .C(_15519_), .Y(_15520_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_15517_), .Y(_15521_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_15521_), .B(_15520_), .Y(_161__1_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(data_244__2_), .Y(_15522_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf0), .B(_15074__bF_buf6), .C(_15522_), .Y(_15523_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_15517_), .Y(_15524_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_15524_), .B(_15523_), .Y(_161__2_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(data_244__3_), .Y(_15525_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf3), .B(_15074__bF_buf5), .C(_15525_), .Y(_15526_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_15517_), .Y(_15527_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_15527_), .B(_15526_), .Y(_161__3_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(data_244__4_), .Y(_15528_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf2), .B(_15074__bF_buf4), .C(_15528_), .Y(_15529_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_15517_), .Y(_15530_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_15530_), .B(_15529_), .Y(_161__4_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(data_244__5_), .Y(_15531_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf1), .B(_15074__bF_buf3), .C(_15531_), .Y(_15532_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_15517_), .Y(_15533_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_15533_), .B(_15532_), .Y(_161__5_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(data_244__6_), .Y(_15534_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf0), .B(_15074__bF_buf2), .C(_15534_), .Y(_15535_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_15517_), .Y(_15536_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_15536_), .B(_15535_), .Y(_161__6_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(data_244__7_), .Y(_15537_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf3), .B(_15074__bF_buf1), .C(_15537_), .Y(_15538_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_15517_), .Y(_15539_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_15539_), .B(_15538_), .Y(_161__7_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(data_244__8_), .Y(_15540_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf2), .B(_15074__bF_buf0), .C(_15540_), .Y(_15541_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_15517_), .Y(_15542_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_15542_), .B(_15541_), .Y(_161__8_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(data_244__9_), .Y(_15543_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf1), .B(_15074__bF_buf12), .C(_15543_), .Y(_15544_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_15517_), .Y(_15545_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_15545_), .B(_15544_), .Y(_161__9_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(data_244__10_), .Y(_15546_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf0), .B(_15074__bF_buf11), .C(_15546_), .Y(_15547_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf3), .B(_15517_), .Y(_15548_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_15548_), .B(_15547_), .Y(_161__10_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(data_244__11_), .Y(_15549_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf3), .B(_15074__bF_buf10), .C(_15549_), .Y(_15550_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_15517_), .Y(_15551_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_15551_), .B(_15550_), .Y(_161__11_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(data_244__12_), .Y(_15552_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf2), .B(_15074__bF_buf9), .C(_15552_), .Y(_15553_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_15517_), .Y(_15554_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_15554_), .B(_15553_), .Y(_161__12_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(data_244__13_), .Y(_15555_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf1), .B(_15074__bF_buf8), .C(_15555_), .Y(_15556_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_15517_), .Y(_15557_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_15557_), .B(_15556_), .Y(_161__13_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(data_244__14_), .Y(_15558_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf0), .B(_15074__bF_buf7), .C(_15558_), .Y(_15559_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_15517_), .Y(_15560_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_15560_), .B(_15559_), .Y(_161__14_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(data_244__15_), .Y(_15561_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_15515__bF_buf3), .B(_15074__bF_buf6), .C(_15561_), .Y(_15562_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_15517_), .Y(_15563_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_15563_), .B(_15562_), .Y(_161__15_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .B(_15017_), .Y(_15564_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .Y(_15565_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_15031__bF_buf2), .C(_14889_), .Y(_15566_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf0), .B(_15565_), .C(_15566_), .Y(_15567_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14965__bF_buf0), .C(_14885__bF_buf3), .Y(_15568_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_15029_), .B(_15567_), .C(_15568_), .Y(_15569_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_15569_), .B(_15564_), .Y(_15570_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14955_), .C(_14942__bF_buf0), .Y(_15571_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .Y(_15572_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf2), .B(_15034_), .C(IDATA_PROG_write_bF_buf3), .Y(_15573_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf2), .B(_15572_), .C(_15573_), .Y(_15574_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_14883_), .B(_14945_), .Y(_15575_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf1), .B(_15006__bF_buf3), .S(_14942__bF_buf3), .Y(_15576_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf3), .B(_15575__bF_buf3), .C(_15576_), .Y(_15577_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_15577_), .B(_15574_), .Y(_15578_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_14955_), .B(_14952__bF_buf3), .Y(_15579_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14982_), .C(_15579_), .Y(_15580_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .Y(_15581_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_15581_), .C(_15120__bF_buf2), .Y(_15582_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_15578_), .B(_15582_), .Y(_15583_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_15583_), .B(_15570_), .Y(_15584_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf5), .B(_15584_), .Y(_15585_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_15585_), .Y(_15586_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(data_243__0_), .B(_15585_), .C(_15586_), .Y(_15587_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_15587_), .Y(_160__0_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_15585_), .Y(_15588_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(data_243__1_), .B(_15585_), .C(_15588_), .Y(_15589_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_15589_), .Y(_160__1_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(data_243__2_), .Y(_15590_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf4), .C(_15590_), .Y(_15591_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_15507_), .B(_15511_), .Y(_15592_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_15582_), .B(_15578_), .Y(_15593_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_15593_), .Y(_15594_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_15183__bF_buf4), .C(_15594_), .Y(_15595_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_15591_), .B(_15595_), .Y(_160__2_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_15585_), .Y(_15596_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(data_243__3_), .B(_15585_), .C(_15596_), .Y(_15597_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_15597_), .Y(_160__3_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_15585_), .Y(_15598_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(data_243__4_), .B(_15585_), .C(_15598_), .Y(_15599_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_15599_), .Y(_160__4_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_15585_), .Y(_15600_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(data_243__5_), .B(_15585_), .C(_15600_), .Y(_15601_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_15601_), .Y(_160__5_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(data_243__6_), .Y(_15602_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf3), .C(_15602_), .Y(_15603_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_15183__bF_buf3), .C(_15594_), .Y(_15604_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_15603_), .B(_15604_), .Y(_160__6_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_15585_), .Y(_15605_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(data_243__7_), .B(_15585_), .C(_15605_), .Y(_15606_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_15606_), .Y(_160__7_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(data_243__8_), .Y(_15607_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf2), .C(_15607_), .Y(_15608_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_15183__bF_buf2), .C(_15594_), .Y(_15609_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_15608_), .B(_15609_), .Y(_160__8_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(data_243__9_), .Y(_15610_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf1), .C(_15610_), .Y(_15611_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_15183__bF_buf1), .C(_15594_), .Y(_15612_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_15611_), .B(_15612_), .Y(_160__9_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(data_243__10_), .Y(_15613_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf0), .C(_15613_), .Y(_15614_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_15183__bF_buf0), .C(_15594_), .Y(_15615_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_15614_), .B(_15615_), .Y(_160__10_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_15585_), .Y(_15616_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(data_243__11_), .B(_15585_), .C(_15616_), .Y(_15617_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_15617_), .Y(_160__11_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_15585_), .Y(_15618_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(data_243__12_), .B(_15585_), .C(_15618_), .Y(_15619_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_15619_), .Y(_160__12_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(data_243__13_), .Y(_15620_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf12), .C(_15620_), .Y(_15621_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_15183__bF_buf8), .C(_15594_), .Y(_15622_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_15621_), .B(_15622_), .Y(_160__13_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(data_243__14_), .Y(_15623_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf11), .C(_15623_), .Y(_15624_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_15183__bF_buf7), .C(_15594_), .Y(_15625_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_15624_), .B(_15625_), .Y(_160__14_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(data_243__15_), .Y(_15626_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_15584_), .B(_15074__bF_buf10), .C(_15626_), .Y(_15627_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf2), .B(_15183__bF_buf6), .C(_15594_), .Y(_15628_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_15627_), .B(_15628_), .Y(_160__15_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(data_242__0_), .Y(_15629_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_15003_), .B(_15172_), .C(_15120__bF_buf1), .Y(_15630_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_15578_), .B(_15630_), .Y(_15631_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_15631_), .B(_15570_), .Y(_15632_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf3), .B(_15074__bF_buf9), .C(_15629_), .Y(_15633_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf8), .B(_15632__bF_buf2), .Y(_15634_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_15634_), .Y(_15635_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_15635_), .B(_15633_), .Y(_159__0_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(data_242__1_), .Y(_15636_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf1), .B(_15074__bF_buf7), .C(_15636_), .Y(_15637_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_15634_), .Y(_15638_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_15638_), .B(_15637_), .Y(_159__1_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(data_242__2_), .Y(_15639_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf0), .B(_15074__bF_buf6), .C(_15639_), .Y(_15640_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_15631_), .Y(_15641_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_15183__bF_buf5), .C(_15641_), .Y(_15642_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_15642_), .B(_15640_), .Y(_159__2_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(data_242__3_), .Y(_15643_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf3), .B(_15074__bF_buf5), .C(_15643_), .Y(_15644_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_15634_), .Y(_15645_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_15645_), .B(_15644_), .Y(_159__3_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(data_242__4_), .Y(_15646_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf2), .B(_15074__bF_buf4), .C(_15646_), .Y(_15647_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_15634_), .Y(_15648_) );
AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_15648_), .B(_15647_), .Y(_159__4_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(data_242__5_), .Y(_15649_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf1), .B(_15074__bF_buf3), .C(_15649_), .Y(_15650_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_15634_), .Y(_15651_) );
AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_15651_), .B(_15650_), .Y(_159__5_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(data_242__6_), .Y(_15652_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf0), .B(_15074__bF_buf2), .C(_15652_), .Y(_15653_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_15183__bF_buf4), .C(_15641_), .Y(_15654_) );
AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_15654_), .B(_15653_), .Y(_159__6_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(data_242__7_), .Y(_15655_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf3), .B(_15074__bF_buf1), .C(_15655_), .Y(_15656_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_15634_), .Y(_15657_) );
AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_15657_), .B(_15656_), .Y(_159__7_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(data_242__8_), .Y(_15658_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf2), .B(_15074__bF_buf0), .C(_15658_), .Y(_15659_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_15183__bF_buf3), .C(_15641_), .Y(_15660_) );
AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_15660_), .B(_15659_), .Y(_159__8_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(data_242__9_), .Y(_15661_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf1), .B(_15074__bF_buf12), .C(_15661_), .Y(_15662_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_15183__bF_buf2), .C(_15641_), .Y(_15663_) );
AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_15663_), .B(_15662_), .Y(_159__9_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(data_242__10_), .Y(_15664_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf0), .B(_15074__bF_buf11), .C(_15664_), .Y(_15665_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_15183__bF_buf1), .C(_15641_), .Y(_15666_) );
AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_15666_), .B(_15665_), .Y(_159__10_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(data_242__11_), .Y(_15667_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf3), .B(_15074__bF_buf10), .C(_15667_), .Y(_15668_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_15634_), .Y(_15669_) );
AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_15669_), .B(_15668_), .Y(_159__11_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(data_242__12_), .Y(_15670_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf2), .B(_15074__bF_buf9), .C(_15670_), .Y(_15671_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_15634_), .Y(_15672_) );
AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_15672_), .B(_15671_), .Y(_159__12_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(data_242__13_), .Y(_15673_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf1), .B(_15074__bF_buf8), .C(_15673_), .Y(_15674_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_15183__bF_buf0), .C(_15641_), .Y(_15675_) );
AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_15675_), .B(_15674_), .Y(_159__13_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(data_242__14_), .Y(_15676_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf0), .B(_15074__bF_buf7), .C(_15676_), .Y(_15677_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_15183__bF_buf8), .C(_15641_), .Y(_15678_) );
AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_15678_), .B(_15677_), .Y(_159__14_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(data_242__15_), .Y(_15679_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_15632__bF_buf3), .B(_15074__bF_buf6), .C(_15679_), .Y(_15680_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_15183__bF_buf7), .C(_15641_), .Y(_15681_) );
AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_15681_), .B(_15680_), .Y(_159__15_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(data_241__0_), .Y(_15682_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf1), .B(_14978__bF_buf1), .Y(_15683_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14982_), .C(_15030_), .Y(_15684_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf0), .B(_15684_), .C(_15573_), .Y(_15685_) );
AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_15685_), .B(_15683_), .Y(_15686_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf0), .B(_15577_), .C(_15686_), .Y(_15687_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_15687_), .Y(_15688_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf3), .B(_15074__bF_buf5), .C(_15682_), .Y(_15689_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf4), .B(_15688__bF_buf2), .Y(_15690_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_15690_), .Y(_15691_) );
AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_15691_), .B(_15689_), .Y(_158__0_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(data_241__1_), .Y(_15692_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf1), .B(_15074__bF_buf3), .C(_15692_), .Y(_15693_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_15690_), .Y(_15694_) );
AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_15694_), .B(_15693_), .Y(_158__1_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(data_241__2_), .Y(_15695_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf0), .B(_15074__bF_buf2), .C(_15695_), .Y(_15696_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_15687_), .B(_15592_), .Y(_15697_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_15183__bF_buf6), .C(_15697_), .Y(_15698_) );
AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_15696_), .B(_15698_), .Y(_158__2_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(data_241__3_), .Y(_15699_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf3), .B(_15074__bF_buf1), .C(_15699_), .Y(_15700_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_15690_), .Y(_15701_) );
AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_15701_), .B(_15700_), .Y(_158__3_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(data_241__4_), .Y(_15702_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf2), .B(_15074__bF_buf0), .C(_15702_), .Y(_15703_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_15690_), .Y(_15704_) );
AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_15704_), .B(_15703_), .Y(_158__4_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(data_241__5_), .Y(_15705_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf1), .B(_15074__bF_buf12), .C(_15705_), .Y(_15706_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_15690_), .Y(_15707_) );
AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_15707_), .B(_15706_), .Y(_158__5_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(data_241__6_), .Y(_15708_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf0), .B(_15074__bF_buf11), .C(_15708_), .Y(_15709_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_15183__bF_buf5), .C(_15697_), .Y(_15710_) );
AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_15709_), .B(_15710_), .Y(_158__6_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(data_241__7_), .Y(_15711_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf3), .B(_15074__bF_buf10), .C(_15711_), .Y(_15712_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_15690_), .Y(_15713_) );
AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_15713_), .B(_15712_), .Y(_158__7_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(data_241__8_), .Y(_15714_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf2), .B(_15074__bF_buf9), .C(_15714_), .Y(_15715_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_15183__bF_buf4), .C(_15697_), .Y(_15716_) );
AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_15715_), .B(_15716_), .Y(_158__8_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(data_241__9_), .Y(_15717_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf1), .B(_15074__bF_buf8), .C(_15717_), .Y(_15718_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_15183__bF_buf3), .C(_15697_), .Y(_15719_) );
AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_15718_), .B(_15719_), .Y(_158__9_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(data_241__10_), .Y(_15720_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf0), .B(_15074__bF_buf7), .C(_15720_), .Y(_15721_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_15183__bF_buf2), .C(_15697_), .Y(_15722_) );
AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_15721_), .B(_15722_), .Y(_158__10_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(data_241__11_), .Y(_15723_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf3), .B(_15074__bF_buf6), .C(_15723_), .Y(_15724_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_15690_), .Y(_15725_) );
AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_15725_), .B(_15724_), .Y(_158__11_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(data_241__12_), .Y(_15726_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf2), .B(_15074__bF_buf5), .C(_15726_), .Y(_15727_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_15690_), .Y(_15728_) );
AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_15728_), .B(_15727_), .Y(_158__12_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(data_241__13_), .Y(_15729_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf1), .B(_15074__bF_buf4), .C(_15729_), .Y(_15730_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_15183__bF_buf1), .C(_15697_), .Y(_15731_) );
AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_15730_), .B(_15731_), .Y(_158__13_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(data_241__14_), .Y(_15732_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf0), .B(_15074__bF_buf3), .C(_15732_), .Y(_15733_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_15183__bF_buf0), .C(_15697_), .Y(_15734_) );
AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_15733_), .B(_15734_), .Y(_158__14_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(data_241__15_), .Y(_15735_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_15688__bF_buf3), .B(_15074__bF_buf2), .C(_15735_), .Y(_15736_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_15183__bF_buf8), .C(_15697_), .Y(_15737_) );
AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_15736_), .B(_15737_), .Y(_158__15_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(data_240__0_), .Y(_15738_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf3), .B(_15074__bF_buf1), .Y(_15739_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf2), .B(_15006__bF_buf2), .Y(_15740_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_15575__bF_buf2), .B(_15740_), .Y(_15741_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf0), .B(_14975_), .C(_14885__bF_buf3), .Y(_15742_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_15741_), .B(_15742_), .C(_15120__bF_buf3), .Y(_15743_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_15743_), .B(_15592_), .Y(_15744_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_15744_), .B(_15739_), .Y(_15745_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_15738_), .B(_14932__bF_buf0), .S(_15745_), .Y(_157__0_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(data_240__1_), .Y(_15746_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_15746_), .B(_14894__bF_buf14), .S(_15745_), .Y(_157__1_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(data_240__2_), .Y(_15747_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_15747_), .B(_14897__bF_buf14), .S(_15745_), .Y(_157__2_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(data_240__3_), .Y(_15748_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_15748_), .B(_14899__bF_buf14), .S(_15745_), .Y(_157__3_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(data_240__4_), .Y(_15749_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_15749_), .B(_14902__bF_buf12), .S(_15745_), .Y(_157__4_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(data_240__5_), .Y(_15750_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_15750_), .B(_14903__bF_buf12), .S(_15745_), .Y(_157__5_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(data_240__6_), .Y(_15751_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_15751_), .B(_15049__bF_buf0), .S(_15745_), .Y(_157__6_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(data_240__7_), .Y(_15752_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_15752_), .B(_14908__bF_buf12), .S(_15745_), .Y(_157__7_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(data_240__8_), .Y(_15753_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_15753_), .B(_15052__bF_buf13), .S(_15745_), .Y(_157__8_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(data_240__9_), .Y(_15754_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_15754_), .B(_14913__bF_buf14), .S(_15745_), .Y(_157__9_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_15744_), .B(_15739_), .C(data_240__10_), .Y(_15755_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf2), .B(_15745_), .Y(_15756_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_15755_), .B(_15756_), .Y(_157__10_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(data_240__11_), .Y(_15757_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_15757_), .B(_14918__bF_buf12), .S(_15745_), .Y(_157__11_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(data_240__12_), .Y(_15758_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_15758_), .B(_14920__bF_buf12), .S(_15745_), .Y(_157__12_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(data_240__13_), .Y(_15759_) );
MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_15759_), .B(_14924__bF_buf12), .S(_15745_), .Y(_157__13_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(data_240__14_), .Y(_15760_) );
MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_15760_), .B(_15060__bF_buf0), .S(_15745_), .Y(_157__14_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(data_240__15_), .Y(_15761_) );
MUX2X1 MUX2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_15761_), .B(_15062__bF_buf13), .S(_15745_), .Y(_157__15_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(data_239__0_), .Y(_15762_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(_14886__bF_buf0), .Y(_15763_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_15763_), .Y(_15764_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf0), .B(_15764_), .Y(_15765_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(_14947_), .C(_14963__bF_buf2), .Y(_15766_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_15766_), .C(_15005__bF_buf3), .Y(_15767_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_15576_), .B(_15767_), .C(_15765_), .Y(_15768_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_15742_), .B(_15768_), .C(_15120__bF_buf2), .Y(_15769_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_15569_), .B(_15769_), .C(_15564_), .Y(_15770_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_15743_), .C(_15770_), .Y(_15771_) );
MUX2X1 MUX2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_15762_), .B(_14932__bF_buf14), .S(_15771_), .Y(_155__0_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(data_239__1_), .Y(_15772_) );
MUX2X1 MUX2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_15772_), .B(_14894__bF_buf13), .S(_15771_), .Y(_155__1_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(data_239__2_), .Y(_15773_) );
MUX2X1 MUX2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_15773_), .B(_14897__bF_buf13), .S(_15771_), .Y(_155__2_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(data_239__3_), .Y(_15774_) );
MUX2X1 MUX2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_15774_), .B(_14899__bF_buf13), .S(_15771_), .Y(_155__3_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(data_239__4_), .Y(_15775_) );
MUX2X1 MUX2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_15775_), .B(_14902__bF_buf11), .S(_15771_), .Y(_155__4_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(data_239__5_), .Y(_15776_) );
MUX2X1 MUX2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_15776_), .B(_14903__bF_buf11), .S(_15771_), .Y(_155__5_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(data_239__6_), .Y(_15777_) );
MUX2X1 MUX2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_15777_), .B(_15049__bF_buf14), .S(_15771_), .Y(_155__6_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(data_239__7_), .Y(_15778_) );
MUX2X1 MUX2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_15778_), .B(_14908__bF_buf11), .S(_15771_), .Y(_155__7_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(data_239__8_), .Y(_15779_) );
MUX2X1 MUX2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_15779_), .B(_15052__bF_buf12), .S(_15771_), .Y(_155__8_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(data_239__9_), .Y(_15780_) );
MUX2X1 MUX2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_15780_), .B(_14913__bF_buf13), .S(_15771_), .Y(_155__9_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(data_239__10_), .Y(_15781_) );
MUX2X1 MUX2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_15781_), .B(_15055__bF_buf13), .S(_15771_), .Y(_155__10_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(data_239__11_), .Y(_15782_) );
MUX2X1 MUX2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_15782_), .B(_14918__bF_buf11), .S(_15771_), .Y(_155__11_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(data_239__12_), .Y(_15783_) );
MUX2X1 MUX2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_15783_), .B(_14920__bF_buf11), .S(_15771_), .Y(_155__12_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(data_239__13_), .Y(_15784_) );
MUX2X1 MUX2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_15784_), .B(_14924__bF_buf11), .S(_15771_), .Y(_155__13_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(data_239__14_), .Y(_15785_) );
MUX2X1 MUX2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_15785_), .B(_15060__bF_buf14), .S(_15771_), .Y(_155__14_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(data_239__15_), .Y(_15786_) );
MUX2X1 MUX2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_15786_), .B(_15062__bF_buf12), .S(_15771_), .Y(_155__15_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(data_238__0_), .Y(_15787_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_14983_), .Y(_15788_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15005__bF_buf2), .C(_15787_), .Y(_15789_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf1), .B(_15788__bF_buf8), .Y(_15790_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_15790_), .Y(_15791_) );
AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_15791_), .B(_15789_), .Y(_154__0_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(data_238__1_), .Y(_15792_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf2), .B(_15766_), .Y(_15793_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_15575__bF_buf1), .B(_15793__bF_buf5), .Y(_15794_) );
MUX2X1 MUX2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_15792_), .B(_14894__bF_buf12), .S(_15794_), .Y(_154__1_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(data_238__2_), .B(_15790_), .Y(_15795_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf12), .B(_15790_), .C(_15795_), .Y(_154__2_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(data_238__3_), .Y(_15796_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15005__bF_buf0), .C(_15796_), .Y(_15797_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_15790_), .Y(_15798_) );
AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_15798_), .B(_15797_), .Y(_154__3_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(data_238__4_), .Y(_15799_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15005__bF_buf3), .C(_15799_), .Y(_15800_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_15790_), .Y(_15801_) );
AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_15801_), .B(_15800_), .Y(_154__4_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(data_238__5_), .Y(_15802_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15005__bF_buf2), .C(_15802_), .Y(_15803_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf3), .B(_15794_), .C(_15803_), .Y(_15804_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(_15804_), .Y(_154__5_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(data_238__6_), .Y(_15805_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15005__bF_buf1), .C(_15805_), .Y(_15806_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_15790_), .Y(_15807_) );
AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_15807_), .B(_15806_), .Y(_154__6_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(data_238__7_), .Y(_15808_) );
MUX2X1 MUX2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_15808_), .B(_14908__bF_buf10), .S(_15794_), .Y(_154__7_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(data_238__8_), .Y(_15809_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15005__bF_buf0), .C(_15809_), .Y(_15810_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf2), .B(_15794_), .C(_15810_), .Y(_15811_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(_15811_), .Y(_154__8_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(data_238__9_), .Y(_15812_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15005__bF_buf3), .C(_15812_), .Y(_15813_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf3), .B(_15794_), .C(_15813_), .Y(_15814_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_15814_), .Y(_154__9_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(data_238__10_), .Y(_15815_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15005__bF_buf2), .C(_15815_), .Y(_15816_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_15575__bF_buf0), .C(_15793__bF_buf4), .Y(_15817_) );
AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_15816_), .B(_15817_), .Y(_154__10_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(data_238__11_), .Y(_15818_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15005__bF_buf1), .C(_15818_), .Y(_15819_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf3), .B(_15794_), .C(_15819_), .Y(_15820_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(_15820_), .Y(_154__11_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(data_238__12_), .Y(_15821_) );
MUX2X1 MUX2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_15821_), .B(_14920__bF_buf10), .S(_15794_), .Y(_154__12_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(data_238__13_), .B(_15790_), .Y(_15822_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf3), .B(_15794_), .Y(_15823_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_15823_), .B(_15822_), .Y(_154__13_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(data_238__14_), .Y(_15824_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15005__bF_buf0), .C(_15824_), .Y(_15825_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_15575__bF_buf3), .C(_15793__bF_buf3), .Y(_15826_) );
AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_15825_), .B(_15826_), .Y(_154__14_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(data_238__15_), .B(_15790_), .Y(_15827_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf3), .B(_15794_), .Y(_15828_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_15828_), .B(_15827_), .Y(_154__15_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(data_237__0_), .Y(_15829_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf2), .B(_14957_), .C(_15575__bF_buf2), .Y(_15830_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(_15084_), .Y(_15831_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf0), .B(_15831_), .Y(_15832_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_15576_), .B(_15592_), .Y(_15833_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_15830_), .B(_15833_), .C(_15832_), .Y(_15834_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .Y(_15835_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_15835_), .B(_15005__bF_buf3), .C(_15742_), .Y(_15836_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_15836_), .B(_15770_), .Y(_15837_) );
INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(_15837_), .Y(_15838_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15838__bF_buf3), .C(_15829_), .Y(_15839_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(_15830_), .Y(_15840_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_15084_), .B(_15183__bF_buf7), .Y(_15841_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_15576_), .Y(_15842_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_15842_), .B(_15570_), .Y(_15843_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_15840_), .B(_15843_), .C(_15841_), .Y(_15844_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_15837_), .C(_15844_), .Y(_15845_) );
AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_15845_), .B(_15839_), .Y(_153__0_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(data_237__1_), .Y(_15846_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15838__bF_buf2), .C(_15846_), .Y(_15847_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_15837_), .C(_15844_), .Y(_15848_) );
AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_15848_), .B(_15847_), .Y(_153__1_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(data_237__2_), .Y(_15849_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15838__bF_buf1), .C(_15849_), .Y(_15850_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_15838__bF_buf0), .B(_15834__bF_buf1), .Y(_15851_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_15851_), .Y(_15852_) );
AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_15852_), .B(_15850_), .Y(_153__2_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(data_237__3_), .Y(_15853_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf0), .B(_15838__bF_buf3), .C(_15853_), .Y(_15854_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_15837_), .C(_15844_), .Y(_15855_) );
AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_15855_), .B(_15854_), .Y(_153__3_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(data_237__4_), .Y(_15856_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15838__bF_buf2), .C(_15856_), .Y(_15857_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_15837_), .C(_15844_), .Y(_15858_) );
AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_15858_), .B(_15857_), .Y(_153__4_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(data_237__5_), .Y(_15859_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15838__bF_buf1), .C(_15859_), .Y(_15860_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_15837_), .C(_15844_), .Y(_15861_) );
AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_15861_), .B(_15860_), .Y(_153__5_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(data_237__6_), .Y(_15862_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15838__bF_buf0), .C(_15862_), .Y(_15863_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_15851_), .Y(_15864_) );
AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_15864_), .B(_15863_), .Y(_153__6_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(data_237__7_), .Y(_15865_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf1), .B(_15838__bF_buf3), .C(_15865_), .Y(_15866_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_15837_), .C(_15844_), .Y(_15867_) );
AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_15867_), .B(_15866_), .Y(_153__7_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(data_237__8_), .Y(_15868_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf0), .B(_15838__bF_buf2), .C(_15868_), .Y(_15869_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_15851_), .Y(_15870_) );
AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_15870_), .B(_15869_), .Y(_153__8_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(data_237__9_), .Y(_15871_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15838__bF_buf1), .C(_15871_), .Y(_15872_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_15851_), .Y(_15873_) );
AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_15873_), .B(_15872_), .Y(_153__9_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(data_237__10_), .Y(_15874_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15838__bF_buf0), .C(_15874_), .Y(_15875_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_15851_), .Y(_15876_) );
AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_15876_), .B(_15875_), .Y(_153__10_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(data_237__11_), .Y(_15877_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15838__bF_buf3), .C(_15877_), .Y(_15878_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_15837_), .C(_15844_), .Y(_15879_) );
AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_15879_), .B(_15878_), .Y(_153__11_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(data_237__12_), .Y(_15880_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf1), .B(_15838__bF_buf2), .C(_15880_), .Y(_15881_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_15837_), .C(_15844_), .Y(_15882_) );
AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_15882_), .B(_15881_), .Y(_153__12_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(data_237__13_), .Y(_15883_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf0), .B(_15838__bF_buf1), .C(_15883_), .Y(_15884_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_15851_), .Y(_15885_) );
AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_15885_), .B(_15884_), .Y(_153__13_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(data_237__14_), .Y(_15886_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15838__bF_buf0), .C(_15886_), .Y(_15887_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_15851_), .Y(_15888_) );
AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_15888_), .B(_15887_), .Y(_153__14_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(data_237__15_), .Y(_15889_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15838__bF_buf3), .C(_15889_), .Y(_15890_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_15851_), .Y(_15891_) );
AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_15891_), .B(_15890_), .Y(_153__15_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(data_236__0_), .Y(_15892_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_14983_), .B(_15575__bF_buf1), .Y(_15893_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_15763_), .C(_15575__bF_buf0), .Y(_15894_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_15893_), .B(_15742_), .C(_15894_), .Y(_15895_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_15576_), .B(_15895_), .C(_15028_), .Y(_15896_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_15507_), .B(_15511_), .C(_15896_), .Y(_15897_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15005__bF_buf2), .C(_15742_), .Y(_15898_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(_15898_), .Y(_15899_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_15897_), .B(_15074__bF_buf12), .C(_15899_), .Y(_15900_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15900__bF_buf10), .C(_15892_), .Y(_15901_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf9), .B(_15834__bF_buf1), .Y(_15902_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_15902_), .Y(_15903_) );
AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_15903_), .B(_15901_), .Y(_152__0_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(data_236__1_), .Y(_15904_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf0), .B(_15900__bF_buf8), .C(_15904_), .Y(_15905_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_15902_), .Y(_15906_) );
AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_15906_), .B(_15905_), .Y(_152__1_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(data_236__2_), .Y(_15907_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15900__bF_buf7), .C(_15907_), .Y(_15908_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_15902_), .Y(_15909_) );
AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_15909_), .B(_15908_), .Y(_152__2_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(data_236__3_), .Y(_15910_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15900__bF_buf6), .C(_15910_), .Y(_15911_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_15902_), .Y(_15912_) );
AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_15912_), .B(_15911_), .Y(_152__3_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(data_236__4_), .Y(_15913_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15900__bF_buf5), .C(_15913_), .Y(_15914_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_15902_), .Y(_15915_) );
AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_15915_), .B(_15914_), .Y(_152__4_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(data_236__5_), .Y(_15916_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf1), .B(_15900__bF_buf4), .C(_15916_), .Y(_15917_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_15902_), .Y(_15918_) );
AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_15918_), .B(_15917_), .Y(_152__5_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(data_236__6_), .Y(_15919_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf0), .B(_15900__bF_buf3), .C(_15919_), .Y(_15920_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_15902_), .Y(_15921_) );
AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_15921_), .B(_15920_), .Y(_152__6_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(data_236__7_), .Y(_15922_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15900__bF_buf2), .C(_15922_), .Y(_15923_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_15902_), .Y(_15924_) );
AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_15924_), .B(_15923_), .Y(_152__7_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(data_236__8_), .Y(_15925_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15900__bF_buf1), .C(_15925_), .Y(_15926_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_15902_), .Y(_15927_) );
AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_15927_), .B(_15926_), .Y(_152__8_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(data_236__9_), .Y(_15928_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15900__bF_buf0), .C(_15928_), .Y(_15929_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_15902_), .Y(_15930_) );
AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_15930_), .B(_15929_), .Y(_152__9_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(data_236__10_), .Y(_15931_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf1), .B(_15900__bF_buf10), .C(_15931_), .Y(_15932_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_15902_), .Y(_15933_) );
AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_15933_), .B(_15932_), .Y(_152__10_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(data_236__11_), .Y(_15934_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf0), .B(_15900__bF_buf9), .C(_15934_), .Y(_15935_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_15902_), .Y(_15936_) );
AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_15936_), .B(_15935_), .Y(_152__11_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(data_236__12_), .Y(_15937_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf4), .B(_15900__bF_buf8), .C(_15937_), .Y(_15938_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_15902_), .Y(_15939_) );
AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_15939_), .B(_15938_), .Y(_152__12_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(data_236__13_), .Y(_15940_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf3), .B(_15900__bF_buf7), .C(_15940_), .Y(_15941_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_15902_), .Y(_15942_) );
AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_15942_), .B(_15941_), .Y(_152__13_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(data_236__14_), .Y(_15943_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf2), .B(_15900__bF_buf6), .C(_15943_), .Y(_15944_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_15902_), .Y(_15945_) );
AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_15945_), .B(_15944_), .Y(_152__14_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(data_236__15_), .Y(_15946_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_15834__bF_buf1), .B(_15900__bF_buf5), .C(_15946_), .Y(_15947_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf10), .B(_15902_), .Y(_15948_) );
AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_15948_), .B(_15947_), .Y(_152__15_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_15770_), .B(_15183__bF_buf6), .C(_15898_), .Y(_15949_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(_15163_), .Y(_15950_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf3), .B(_14951_), .C(_15950_), .Y(_15951_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .B(_15005__bF_buf1), .C(IDATA_PROG_write_bF_buf0), .Y(_15952_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_15575__bF_buf3), .B(_15951_), .C(_15952_), .Y(_15953_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_15842_), .B(_15120__bF_buf1), .C(_15953_), .Y(_15954_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_15954_), .C(_15074__bF_buf11), .Y(_15955_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf8), .C(data_235__0_), .Y(_15956_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(_15954_), .Y(_15957_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_15957_), .C(_15183__bF_buf5), .Y(_15958_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf4), .B(IDATA_PROG_data_0_bF_buf2), .C(_15958_), .Y(_15959_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_15956_), .B(_15959_), .Y(_151__0_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf7), .C(data_235__1_), .Y(_15960_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf3), .B(IDATA_PROG_data_1_bF_buf3), .C(_15958_), .Y(_15961_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_15960_), .B(_15961_), .Y(_151__1_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(data_235__2_), .Y(_15962_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf2), .C(_15962_), .Y(_15963_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_15955_), .C(_15949__bF_buf6), .Y(_15964_) );
AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_15964_), .B(_15963_), .Y(_151__2_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf5), .C(data_235__3_), .Y(_15965_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf1), .B(IDATA_PROG_data_3_bF_buf3), .C(_15958_), .Y(_15966_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_15965_), .B(_15966_), .Y(_151__3_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf4), .C(data_235__4_), .Y(_15967_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf0), .B(IDATA_PROG_data_4_bF_buf3), .C(_15958_), .Y(_15968_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_15967_), .B(_15968_), .Y(_151__4_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf3), .C(data_235__5_), .Y(_15969_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf10), .B(IDATA_PROG_data_5_bF_buf2), .C(_15958_), .Y(_15970_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_15969_), .B(_15970_), .Y(_151__5_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(data_235__6_), .Y(_15971_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf9), .C(_15971_), .Y(_15972_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_15955_), .C(_15949__bF_buf2), .Y(_15973_) );
AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_15973_), .B(_15972_), .Y(_151__6_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf1), .C(data_235__7_), .Y(_15974_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf8), .B(IDATA_PROG_data_7_bF_buf4), .C(_15958_), .Y(_15975_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_15974_), .B(_15975_), .Y(_151__7_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(data_235__8_), .Y(_15976_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf7), .C(_15976_), .Y(_15977_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_15955_), .C(_15949__bF_buf0), .Y(_15978_) );
AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_15978_), .B(_15977_), .Y(_151__8_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(data_235__9_), .Y(_15979_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf6), .C(_15979_), .Y(_15980_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_15955_), .C(_15949__bF_buf8), .Y(_15981_) );
AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_15981_), .B(_15980_), .Y(_151__9_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(data_235__10_), .Y(_15982_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf5), .C(_15982_), .Y(_15983_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_15955_), .C(_15949__bF_buf7), .Y(_15984_) );
AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_15984_), .B(_15983_), .Y(_151__10_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf6), .C(data_235__11_), .Y(_15985_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf4), .B(IDATA_PROG_data_11_bF_buf2), .C(_15958_), .Y(_15986_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_15985_), .B(_15986_), .Y(_151__11_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_15955_), .B(_15949__bF_buf5), .C(data_235__12_), .Y(_15987_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf3), .B(IDATA_PROG_data_12_bF_buf3), .C(_15958_), .Y(_15988_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_15987_), .B(_15988_), .Y(_151__12_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(data_235__13_), .Y(_15989_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf2), .C(_15989_), .Y(_15990_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_15955_), .C(_15949__bF_buf4), .Y(_15991_) );
AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_15991_), .B(_15990_), .Y(_151__13_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(data_235__14_), .Y(_15992_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf1), .C(_15992_), .Y(_15993_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_15955_), .C(_15949__bF_buf3), .Y(_15994_) );
AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_15994_), .B(_15993_), .Y(_151__14_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(data_235__15_), .Y(_15995_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_15958_), .B(_15900__bF_buf0), .C(_15995_), .Y(_15996_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_15955_), .C(_15949__bF_buf2), .Y(_15997_) );
AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_15997_), .B(_15996_), .Y(_151__15_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(data_234__0_), .Y(_15998_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .B(_14883_), .C(IDATA_PROG_write_bF_buf8), .Y(_15999_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .B(_14882__bF_buf1), .C(_15999_), .Y(_16000_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14952__bF_buf1), .C(_15575__bF_buf2), .Y(_16001_) );
AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_16001_), .B(_15842_), .Y(_16002_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf0), .B(_16000_), .C(_16002_), .Y(_16003_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(_16003_), .Y(_16004_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_16004_), .C(_15183__bF_buf4), .Y(_16005_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf10), .C(_15998_), .Y(_16006_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_16003_), .C(_15074__bF_buf10), .Y(_16007_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_16007_), .C(_15949__bF_buf1), .Y(_16008_) );
AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_16008_), .B(_16006_), .Y(_150__0_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(data_234__1_), .Y(_16009_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf9), .C(_16009_), .Y(_16010_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_16007_), .C(_15949__bF_buf0), .Y(_16011_) );
AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_16011_), .B(_16010_), .Y(_150__1_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(data_234__2_), .Y(_16012_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf8), .C(_16012_), .Y(_16013_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_16007_), .C(_15949__bF_buf8), .Y(_16014_) );
AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_16014_), .B(_16013_), .Y(_150__2_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(data_234__3_), .Y(_16015_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf7), .C(_16015_), .Y(_16016_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_16007_), .C(_15949__bF_buf7), .Y(_16017_) );
AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_16017_), .B(_16016_), .Y(_150__3_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(data_234__4_), .Y(_16018_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf6), .C(_16018_), .Y(_16019_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_16007_), .C(_15949__bF_buf6), .Y(_16020_) );
AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_16020_), .B(_16019_), .Y(_150__4_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(data_234__5_), .Y(_16021_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf5), .C(_16021_), .Y(_16022_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_16007_), .C(_15949__bF_buf5), .Y(_16023_) );
AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_16023_), .B(_16022_), .Y(_150__5_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(data_234__6_), .Y(_16024_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf4), .C(_16024_), .Y(_16025_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_16007_), .C(_15949__bF_buf4), .Y(_16026_) );
AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_16026_), .B(_16025_), .Y(_150__6_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(data_234__7_), .Y(_16027_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf3), .C(_16027_), .Y(_16028_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_16007_), .C(_15949__bF_buf3), .Y(_16029_) );
AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_16029_), .B(_16028_), .Y(_150__7_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(data_234__8_), .Y(_16030_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf2), .C(_16030_), .Y(_16031_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_16007_), .C(_15949__bF_buf2), .Y(_16032_) );
AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_16032_), .B(_16031_), .Y(_150__8_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(data_234__9_), .Y(_16033_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf1), .C(_16033_), .Y(_16034_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_16007_), .C(_15949__bF_buf1), .Y(_16035_) );
AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_16035_), .B(_16034_), .Y(_150__9_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(data_234__10_), .Y(_16036_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf0), .C(_16036_), .Y(_16037_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_16007_), .C(_15949__bF_buf0), .Y(_16038_) );
AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_16038_), .B(_16037_), .Y(_150__10_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(data_234__11_), .Y(_16039_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf10), .C(_16039_), .Y(_16040_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_16007_), .C(_15949__bF_buf8), .Y(_16041_) );
AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_16041_), .B(_16040_), .Y(_150__11_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(data_234__12_), .Y(_16042_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf9), .C(_16042_), .Y(_16043_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_16007_), .C(_15949__bF_buf7), .Y(_16044_) );
AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_16044_), .B(_16043_), .Y(_150__12_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(data_234__13_), .Y(_16045_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf8), .C(_16045_), .Y(_16046_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_16007_), .C(_15949__bF_buf6), .Y(_16047_) );
AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_16047_), .B(_16046_), .Y(_150__13_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(data_234__14_), .Y(_16048_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf7), .C(_16048_), .Y(_16049_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_16007_), .C(_15949__bF_buf5), .Y(_16050_) );
AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_16050_), .B(_16049_), .Y(_150__14_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(data_234__15_), .Y(_16051_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_16005_), .B(_15900__bF_buf6), .C(_16051_), .Y(_16052_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_16007_), .C(_15949__bF_buf4), .Y(_16053_) );
AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_16053_), .B(_16052_), .Y(_150__15_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(data_233__0_), .Y(_16054_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_14989_), .B(IDATA_PROG_addr[0]), .C(_14977__bF_buf3), .Y(_16055_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_15575__bF_buf1), .B(_16055_), .C(_15576_), .Y(_16056_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_16000_), .B(_16056_), .Y(_16057_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_16057_), .Y(_16058_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_16058_), .C(_15183__bF_buf3), .Y(_16059_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf5), .C(_16054_), .Y(_16060_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(_16058_), .Y(_16061_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_16061_), .C(_15074__bF_buf9), .Y(_16062_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_16062_), .C(_15949__bF_buf3), .Y(_16063_) );
AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_16063_), .B(_16060_), .Y(_149__0_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(data_233__1_), .Y(_16064_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf4), .C(_16064_), .Y(_16065_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_16062_), .C(_15949__bF_buf2), .Y(_16066_) );
AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_16066_), .B(_16065_), .Y(_149__1_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(data_233__2_), .Y(_16067_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf3), .C(_16067_), .Y(_16068_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_16062_), .C(_15949__bF_buf1), .Y(_16069_) );
AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_16069_), .B(_16068_), .Y(_149__2_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(data_233__3_), .Y(_16070_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf2), .C(_16070_), .Y(_16071_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_16062_), .C(_15949__bF_buf0), .Y(_16072_) );
AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_16072_), .B(_16071_), .Y(_149__3_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(data_233__4_), .Y(_16073_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf1), .C(_16073_), .Y(_16074_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_16062_), .C(_15949__bF_buf8), .Y(_16075_) );
AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_16075_), .B(_16074_), .Y(_149__4_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(data_233__5_), .Y(_16076_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf0), .C(_16076_), .Y(_16077_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_16062_), .C(_15949__bF_buf7), .Y(_16078_) );
AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_16078_), .B(_16077_), .Y(_149__5_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(data_233__6_), .Y(_16079_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf10), .C(_16079_), .Y(_16080_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_16062_), .C(_15949__bF_buf6), .Y(_16081_) );
AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_16081_), .B(_16080_), .Y(_149__6_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(data_233__7_), .Y(_16082_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf9), .C(_16082_), .Y(_16083_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_16062_), .C(_15949__bF_buf5), .Y(_16084_) );
AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_16084_), .B(_16083_), .Y(_149__7_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(data_233__8_), .Y(_16085_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf8), .C(_16085_), .Y(_16086_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_16062_), .C(_15949__bF_buf4), .Y(_16087_) );
AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_16087_), .B(_16086_), .Y(_149__8_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(data_233__9_), .Y(_16088_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf7), .C(_16088_), .Y(_16089_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_16062_), .C(_15949__bF_buf3), .Y(_16090_) );
AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_16090_), .B(_16089_), .Y(_149__9_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(data_233__10_), .Y(_16091_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf6), .C(_16091_), .Y(_16092_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_16062_), .C(_15949__bF_buf2), .Y(_16093_) );
AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_16093_), .B(_16092_), .Y(_149__10_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(data_233__11_), .Y(_16094_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf5), .C(_16094_), .Y(_16095_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_16062_), .C(_15949__bF_buf1), .Y(_16096_) );
AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_16096_), .B(_16095_), .Y(_149__11_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(data_233__12_), .Y(_16097_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf4), .C(_16097_), .Y(_16098_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_16062_), .C(_15949__bF_buf0), .Y(_16099_) );
AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_16099_), .B(_16098_), .Y(_149__12_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(data_233__13_), .Y(_16100_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf3), .C(_16100_), .Y(_16101_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_16062_), .C(_15949__bF_buf8), .Y(_16102_) );
AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_16102_), .B(_16101_), .Y(_149__13_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(data_233__14_), .Y(_16103_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf2), .C(_16103_), .Y(_16104_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_16062_), .C(_15949__bF_buf7), .Y(_16105_) );
AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_16105_), .B(_16104_), .Y(_149__14_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(data_233__15_), .Y(_16106_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_16059_), .B(_15900__bF_buf1), .C(_16106_), .Y(_16107_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_16062_), .C(_15949__bF_buf6), .Y(_16108_) );
AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_16108_), .B(_16107_), .Y(_149__15_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf3), .B(_14952__bF_buf0), .C(_15575__bF_buf0), .Y(_16109_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_15833_), .B(_16109_), .C(_15832_), .Y(_16110_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf0), .B(_16110_), .Y(_16111_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_16111__bF_buf3), .B(data_232__0_), .Y(_16112_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_16111__bF_buf2), .Y(_16113_) );
AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_16112_), .B(_16113_), .Y(_148__0_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_16111__bF_buf1), .B(data_232__1_), .Y(_16114_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_16111__bF_buf0), .Y(_16115_) );
AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_16114_), .B(_16115_), .Y(_148__1_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(data_232__2_), .Y(_16116_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf10), .C(_16116_), .Y(_16117_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_16111__bF_buf3), .Y(_16118_) );
AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_16118_), .B(_16117_), .Y(_148__2_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_16111__bF_buf2), .B(data_232__3_), .Y(_16119_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_16111__bF_buf1), .Y(_16120_) );
AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_16119_), .B(_16120_), .Y(_148__3_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_16111__bF_buf0), .B(data_232__4_), .Y(_16121_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_16111__bF_buf3), .Y(_16122_) );
AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_16121_), .B(_16122_), .Y(_148__4_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_16111__bF_buf2), .B(data_232__5_), .Y(_16123_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_16111__bF_buf1), .Y(_16124_) );
AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_16123_), .B(_16124_), .Y(_148__5_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(data_232__6_), .Y(_16125_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf9), .C(_16125_), .Y(_16126_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_16111__bF_buf0), .Y(_16127_) );
AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_16127_), .B(_16126_), .Y(_148__6_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(data_232__7_), .Y(_16128_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf8), .C(_16128_), .Y(_16129_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_16111__bF_buf3), .Y(_16130_) );
AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_16130_), .B(_16129_), .Y(_148__7_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(data_232__8_), .Y(_16131_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf7), .C(_16131_), .Y(_16132_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_16111__bF_buf2), .Y(_16133_) );
AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_16133_), .B(_16132_), .Y(_148__8_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(data_232__9_), .Y(_16134_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf6), .C(_16134_), .Y(_16135_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf7), .B(_16111__bF_buf1), .Y(_16136_) );
AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_16136_), .B(_16135_), .Y(_148__9_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(data_232__10_), .Y(_16137_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf5), .C(_16137_), .Y(_16138_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_16111__bF_buf0), .Y(_16139_) );
AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_16139_), .B(_16138_), .Y(_148__10_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_16111__bF_buf3), .B(data_232__11_), .Y(_16140_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_16111__bF_buf2), .Y(_16141_) );
AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_16140_), .B(_16141_), .Y(_148__11_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(data_232__12_), .Y(_16142_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf4), .C(_16142_), .Y(_16143_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_16111__bF_buf1), .Y(_16144_) );
AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_16144_), .B(_16143_), .Y(_148__12_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(data_232__13_), .Y(_16145_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf3), .C(_16145_), .Y(_16146_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_16111__bF_buf0), .Y(_16147_) );
AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_16147_), .B(_16146_), .Y(_148__13_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(data_232__14_), .Y(_16148_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf2), .C(_16148_), .Y(_16149_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_16111__bF_buf3), .Y(_16150_) );
AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_16150_), .B(_16149_), .Y(_148__14_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(data_232__15_), .Y(_16151_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_16110_), .B(_15900__bF_buf1), .C(_16151_), .Y(_16152_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_16111__bF_buf2), .Y(_16153_) );
AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_16153_), .B(_16152_), .Y(_148__15_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(data_231__0_), .Y(_16154_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf2), .B(_15363_), .C(_15575__bF_buf3), .Y(_16155_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14977__bF_buf2), .Y(_16156_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_14976_), .B(_14977__bF_buf1), .Y(_16157_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_16156_), .B(_16157_), .C(_15575__bF_buf2), .Y(_16158_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf0), .B(_15576_), .Y(_16159_) );
AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_16159_), .B(_16158_), .Y(_16160_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf3), .B(_16155_), .C(_16160_), .Y(_16161_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(_16161_), .Y(_16162_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_16162_), .C(_15183__bF_buf2), .Y(_16163_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf0), .C(_16154_), .Y(_16164_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_16161_), .B(_15592_), .C(_15074__bF_buf8), .Y(_16165_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_16165_), .C(_15949__bF_buf5), .Y(_16166_) );
AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_16166_), .B(_16164_), .Y(_147__0_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(data_231__1_), .Y(_16167_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf10), .C(_16167_), .Y(_16168_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_16165_), .C(_15949__bF_buf4), .Y(_16169_) );
AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_16169_), .B(_16168_), .Y(_147__1_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf3), .C(data_231__2_), .Y(_16170_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf9), .B(IDATA_PROG_data_2_bF_buf2), .C(_16163_), .Y(_16171_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_16170_), .B(_16171_), .Y(_147__2_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(data_231__3_), .Y(_16172_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf8), .C(_16172_), .Y(_16173_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_16165_), .C(_15949__bF_buf2), .Y(_16174_) );
AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_16174_), .B(_16173_), .Y(_147__3_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(data_231__4_), .Y(_16175_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf7), .C(_16175_), .Y(_16176_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_16165_), .C(_15949__bF_buf1), .Y(_16177_) );
AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_16177_), .B(_16176_), .Y(_147__4_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(data_231__5_), .Y(_16178_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf6), .C(_16178_), .Y(_16179_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_16165_), .C(_15949__bF_buf0), .Y(_16180_) );
AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_16180_), .B(_16179_), .Y(_147__5_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf8), .C(data_231__6_), .Y(_16181_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf5), .B(IDATA_PROG_data_6_bF_buf2), .C(_16163_), .Y(_16182_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_16181_), .B(_16182_), .Y(_147__6_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(data_231__7_), .Y(_16183_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf4), .C(_16183_), .Y(_16184_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_16165_), .C(_15949__bF_buf7), .Y(_16185_) );
AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(_16185_), .B(_16184_), .Y(_147__7_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf6), .C(data_231__8_), .Y(_16186_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf3), .B(IDATA_PROG_data_8_bF_buf1), .C(_16163_), .Y(_16187_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_16186_), .B(_16187_), .Y(_147__8_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf5), .C(data_231__9_), .Y(_16188_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf2), .B(IDATA_PROG_data_9_bF_buf2), .C(_16163_), .Y(_16189_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_16188_), .B(_16189_), .Y(_147__9_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf4), .C(data_231__10_), .Y(_16190_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf1), .B(IDATA_PROG_data_10_bF_buf1), .C(_16163_), .Y(_16191_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_16190_), .B(_16191_), .Y(_147__10_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(data_231__11_), .Y(_16192_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf0), .C(_16192_), .Y(_16193_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_16165_), .C(_15949__bF_buf3), .Y(_16194_) );
AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_16194_), .B(_16193_), .Y(_147__11_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(data_231__12_), .Y(_16195_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_16163_), .B(_15900__bF_buf10), .C(_16195_), .Y(_16196_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_16165_), .C(_15949__bF_buf2), .Y(_16197_) );
AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_16197_), .B(_16196_), .Y(_147__12_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf1), .C(data_231__13_), .Y(_16198_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf9), .B(IDATA_PROG_data_13_bF_buf2), .C(_16163_), .Y(_16199_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_16198_), .B(_16199_), .Y(_147__13_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf0), .C(data_231__14_), .Y(_16200_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf8), .B(IDATA_PROG_data_14_bF_buf2), .C(_16163_), .Y(_16201_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_16200_), .B(_16201_), .Y(_147__14_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_16165_), .B(_15949__bF_buf8), .C(data_231__15_), .Y(_16202_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf7), .B(IDATA_PROG_data_15_bF_buf2), .C(_16163_), .Y(_16203_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_16202_), .B(_16203_), .Y(_147__15_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_14958_), .Y(_16204_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_16204_), .B(_14965__bF_buf1), .C(_15999_), .Y(_16205_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_15842_), .B(_16205_), .Y(_16206_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf0), .B(_15360_), .C(_15120__bF_buf2), .Y(_16207_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_16206_), .B(_16207_), .Y(_16208_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_16208_), .C(_15074__bF_buf7), .Y(_16209_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_16209_), .B(_15949__bF_buf7), .Y(_16210_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(data_230__0_), .Y(_16211_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_16207_), .B(_16206_), .Y(_16212_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_16212_), .C(_15183__bF_buf1), .Y(_16213_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf6), .C(_16211_), .Y(_16214_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_0_bF_buf1), .C(_16214_), .Y(_16215_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_16215_), .Y(_146__0_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(data_230__1_), .Y(_16216_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf5), .C(_16216_), .Y(_16217_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_1_bF_buf2), .C(_16217_), .Y(_16218_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(_16218_), .Y(_146__1_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(data_230__2_), .Y(_16219_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf4), .C(_16219_), .Y(_16220_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_2_bF_buf1), .C(_16220_), .Y(_16221_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_16221_), .Y(_146__2_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(data_230__3_), .Y(_16222_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf3), .C(_16222_), .Y(_16223_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_3_bF_buf2), .C(_16223_), .Y(_16224_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_16224_), .Y(_146__3_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(data_230__4_), .Y(_16225_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf2), .C(_16225_), .Y(_16226_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_4_bF_buf2), .C(_16226_), .Y(_16227_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_16227_), .Y(_146__4_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(data_230__5_), .Y(_16228_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf1), .C(_16228_), .Y(_16229_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_5_bF_buf1), .C(_16229_), .Y(_16230_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(_16230_), .Y(_146__5_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(data_230__6_), .Y(_16231_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf0), .C(_16231_), .Y(_16232_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_6_bF_buf1), .C(_16232_), .Y(_257_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(_257_), .Y(_146__6_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(data_230__7_), .Y(_258_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf10), .C(_258_), .Y(_259_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_7_bF_buf3), .C(_259_), .Y(_260_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(_260_), .Y(_146__7_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(data_230__8_), .Y(_261_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf9), .C(_261_), .Y(_262_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_8_bF_buf0), .C(_262_), .Y(_263_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(_263_), .Y(_146__8_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(data_230__9_), .Y(_264_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf8), .C(_264_), .Y(_265_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_9_bF_buf1), .C(_265_), .Y(_266_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(_266_), .Y(_146__9_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(data_230__10_), .Y(_267_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf7), .C(_267_), .Y(_268_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_10_bF_buf0), .C(_268_), .Y(_269_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(_269_), .Y(_146__10_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(data_230__11_), .Y(_270_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf6), .C(_270_), .Y(_271_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_11_bF_buf1), .C(_271_), .Y(_272_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(_272_), .Y(_146__11_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(data_230__12_), .Y(_273_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf5), .C(_273_), .Y(_274_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_12_bF_buf2), .C(_274_), .Y(_275_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(_275_), .Y(_146__12_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(data_230__13_), .Y(_276_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf4), .C(_276_), .Y(_277_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_13_bF_buf1), .C(_277_), .Y(_278_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(_278_), .Y(_146__13_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(data_230__14_), .Y(_279_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf3), .C(_279_), .Y(_280_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_14_bF_buf1), .C(_280_), .Y(_281_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(_281_), .Y(_146__14_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(data_230__15_), .Y(_282_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_16213_), .B(_15900__bF_buf2), .C(_282_), .Y(_283_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_16210_), .B(IDATA_PROG_data_15_bF_buf1), .C(_283_), .Y(_284_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(_284_), .Y(_146__15_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(data_229__0_), .Y(_285_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf3), .B(_15453_), .C(_15120__bF_buf1), .Y(_286_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_16206_), .Y(_287_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_287_), .C(_15183__bF_buf0), .Y(_288_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf1), .C(_285_), .Y(_289_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(_287_), .Y(_290_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf6), .B(_15592_), .C(_290_), .Y(_291_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_15949__bF_buf6), .C(_291_), .Y(_292_) );
AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_289_), .Y(_144__0_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(data_229__1_), .Y(_293_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf0), .C(_293_), .Y(_294_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_15949__bF_buf5), .C(_291_), .Y(_295_) );
AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_294_), .Y(_144__1_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(data_229__2_), .Y(_296_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf10), .C(_296_), .Y(_297_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_15949__bF_buf4), .C(_291_), .Y(_298_) );
AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_297_), .Y(_144__2_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(data_229__3_), .Y(_299_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf9), .C(_299_), .Y(_300_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_15949__bF_buf3), .C(_291_), .Y(_301_) );
AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_300_), .Y(_144__3_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(data_229__4_), .Y(_302_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf8), .C(_302_), .Y(_303_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_15949__bF_buf2), .C(_291_), .Y(_304_) );
AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_303_), .Y(_144__4_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(data_229__5_), .Y(_305_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf7), .C(_305_), .Y(_306_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_15949__bF_buf1), .C(_291_), .Y(_307_) );
AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_306_), .Y(_144__5_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(data_229__6_), .Y(_308_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf6), .C(_308_), .Y(_309_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_15949__bF_buf0), .C(_291_), .Y(_310_) );
AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_309_), .Y(_144__6_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(data_229__7_), .Y(_311_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf5), .C(_311_), .Y(_312_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_15949__bF_buf8), .C(_291_), .Y(_313_) );
AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_312_), .Y(_144__7_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(data_229__8_), .Y(_314_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf4), .C(_314_), .Y(_315_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_15949__bF_buf7), .C(_291_), .Y(_316_) );
AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_315_), .Y(_144__8_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(data_229__9_), .Y(_317_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf3), .C(_317_), .Y(_318_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_15949__bF_buf6), .C(_291_), .Y(_319_) );
AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_318_), .Y(_144__9_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(data_229__10_), .Y(_320_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf2), .C(_320_), .Y(_321_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_15949__bF_buf5), .C(_291_), .Y(_322_) );
AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_321_), .Y(_144__10_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(data_229__11_), .Y(_323_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf1), .C(_323_), .Y(_324_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_15949__bF_buf4), .C(_291_), .Y(_325_) );
AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_324_), .Y(_144__11_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(data_229__12_), .Y(_326_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf0), .C(_326_), .Y(_327_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_15949__bF_buf3), .C(_291_), .Y(_328_) );
AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_327_), .Y(_144__12_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(data_229__13_), .Y(_329_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf10), .C(_329_), .Y(_330_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_15949__bF_buf2), .C(_291_), .Y(_331_) );
AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_330_), .Y(_144__13_) );
INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(data_229__14_), .Y(_332_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf9), .C(_332_), .Y(_333_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_15949__bF_buf1), .C(_291_), .Y(_334_) );
AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_333_), .Y(_144__14_) );
INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(data_229__15_), .Y(_335_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_15900__bF_buf8), .C(_335_), .Y(_336_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_15949__bF_buf0), .C(_291_), .Y(_337_) );
AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_336_), .Y(_144__15_) );
INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(data_228__0_), .Y(_338_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_15843_), .B(_15841_), .Y(_339_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14965__bF_buf0), .C(_15575__bF_buf1), .Y(_340_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_341_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_15900__bF_buf7), .Y(_342_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_342__bF_buf4), .Y(_343_) );
MUX2X1 MUX2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_14932__bF_buf5), .S(_343_), .Y(_143__0_) );
INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(data_228__1_), .Y(_344_) );
MUX2X1 MUX2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_14894__bF_buf4), .S(_343_), .Y(_143__1_) );
INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(data_228__2_), .Y(_345_) );
MUX2X1 MUX2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_14897__bF_buf4), .S(_343_), .Y(_143__2_) );
INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(data_228__3_), .Y(_346_) );
MUX2X1 MUX2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_14899__bF_buf4), .S(_343_), .Y(_143__3_) );
INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(data_228__4_), .Y(_347_) );
MUX2X1 MUX2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_14902__bF_buf2), .S(_343_), .Y(_143__4_) );
INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(data_228__5_), .Y(_348_) );
MUX2X1 MUX2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_14903__bF_buf3), .S(_343_), .Y(_143__5_) );
INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(data_228__6_), .Y(_349_) );
MUX2X1 MUX2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_15049__bF_buf5), .S(_343_), .Y(_143__6_) );
INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(data_228__7_), .Y(_350_) );
MUX2X1 MUX2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_14908__bF_buf2), .S(_343_), .Y(_143__7_) );
INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(data_228__8_), .Y(_351_) );
MUX2X1 MUX2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_15052__bF_buf4), .S(_343_), .Y(_143__8_) );
INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(data_228__9_), .Y(_352_) );
MUX2X1 MUX2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_14913__bF_buf5), .S(_343_), .Y(_143__9_) );
INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(data_228__10_), .Y(_353_) );
MUX2X1 MUX2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_15055__bF_buf4), .S(_343_), .Y(_143__10_) );
INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(data_228__11_), .Y(_354_) );
MUX2X1 MUX2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_14918__bF_buf3), .S(_343_), .Y(_143__11_) );
INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(data_228__12_), .Y(_355_) );
MUX2X1 MUX2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_14920__bF_buf2), .S(_343_), .Y(_143__12_) );
INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(data_228__13_), .Y(_356_) );
MUX2X1 MUX2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_14924__bF_buf3), .S(_343_), .Y(_143__13_) );
INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(data_228__14_), .Y(_357_) );
MUX2X1 MUX2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_15060__bF_buf5), .S(_343_), .Y(_143__14_) );
INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(data_228__15_), .Y(_358_) );
MUX2X1 MUX2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_15062__bF_buf4), .S(_343_), .Y(_143__15_) );
INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(data_227__0_), .Y(_359_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_15770_), .B(_15183__bF_buf8), .Y(_360_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_15899_), .B(_340_), .C(_360_), .Y(_361_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_15074__bF_buf5), .Y(_362_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_15575__bF_buf0), .B(_15580_), .Y(_363_) );
INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(_363_), .Y(_364_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf1), .B(_14942__bF_buf1), .C(IDATA_PROG_write_bF_buf6), .Y(_365_) );
INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(_365_), .Y(_366_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_15005__bF_buf2), .C(_366_), .Y(_367_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_364_), .Y(_368_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf0), .B(_368_), .C(_362_), .Y(_369_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf5), .B(_369_), .C(_359_), .Y(_370_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_15001_), .C(_15570_), .Y(_371_) );
INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(_368_), .Y(_372_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_372_), .C(_371_), .Y(_373_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_373_), .C(_342__bF_buf3), .Y(_374_) );
AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_370_), .Y(_142__0_) );
INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(data_227__1_), .Y(_375_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf4), .B(_369_), .C(_375_), .Y(_376_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_373_), .C(_342__bF_buf2), .Y(_377_) );
AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_376_), .Y(_142__1_) );
INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(data_227__2_), .Y(_378_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf3), .B(_369_), .C(_378_), .Y(_379_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_373_), .C(_342__bF_buf1), .Y(_380_) );
AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_379_), .Y(_142__2_) );
INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(data_227__3_), .Y(_381_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf2), .B(_369_), .C(_381_), .Y(_382_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_373_), .C(_342__bF_buf0), .Y(_383_) );
AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_382_), .Y(_142__3_) );
INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(data_227__4_), .Y(_384_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf1), .B(_369_), .C(_384_), .Y(_385_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_373_), .C(_342__bF_buf4), .Y(_386_) );
AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_385_), .Y(_142__4_) );
INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(data_227__5_), .Y(_387_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf0), .B(_369_), .C(_387_), .Y(_388_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_373_), .C(_342__bF_buf3), .Y(_389_) );
AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_388_), .Y(_142__5_) );
INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(data_227__6_), .Y(_390_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf5), .B(_369_), .C(_390_), .Y(_391_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_373_), .C(_342__bF_buf2), .Y(_392_) );
AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_391_), .Y(_142__6_) );
INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(data_227__7_), .Y(_393_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf4), .B(_369_), .C(_393_), .Y(_394_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_373_), .C(_342__bF_buf1), .Y(_395_) );
AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_394_), .Y(_142__7_) );
INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(data_227__8_), .Y(_396_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf3), .B(_369_), .C(_396_), .Y(_397_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_373_), .C(_342__bF_buf0), .Y(_398_) );
AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_397_), .Y(_142__8_) );
INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(data_227__9_), .Y(_399_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf2), .B(_369_), .C(_399_), .Y(_400_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_373_), .C(_342__bF_buf4), .Y(_401_) );
AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_400_), .Y(_142__9_) );
INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(data_227__10_), .Y(_402_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf1), .B(_369_), .C(_402_), .Y(_403_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf3), .B(_373_), .C(_342__bF_buf3), .Y(_404_) );
AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_403_), .Y(_142__10_) );
INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(data_227__11_), .Y(_405_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf0), .B(_369_), .C(_405_), .Y(_406_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_373_), .C(_342__bF_buf2), .Y(_407_) );
AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_406_), .Y(_142__11_) );
INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(data_227__12_), .Y(_408_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf5), .B(_369_), .C(_408_), .Y(_409_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_373_), .C(_342__bF_buf1), .Y(_410_) );
AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_409_), .Y(_142__12_) );
INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(data_227__13_), .Y(_411_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf4), .B(_369_), .C(_411_), .Y(_412_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_373_), .C(_342__bF_buf0), .Y(_413_) );
AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_412_), .Y(_142__13_) );
INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(data_227__14_), .Y(_414_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf3), .B(_369_), .C(_414_), .Y(_415_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_373_), .C(_342__bF_buf4), .Y(_416_) );
AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_415_), .Y(_142__14_) );
INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(data_227__15_), .Y(_417_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf2), .B(_369_), .C(_417_), .Y(_418_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_373_), .C(_342__bF_buf3), .Y(_419_) );
AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_418_), .Y(_142__15_) );
INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(data_226__0_), .Y(_420_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_371_), .Y(_421_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf4), .B(_15575__bF_buf3), .C(_365_), .Y(_422_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_15005__bF_buf1), .C(_422_), .Y(_423_) );
INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(_423_), .Y(_424_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_421_), .Y(_425_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf3), .B(_361__bF_buf1), .C(_420_), .Y(_426_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf0), .B(_425__bF_buf2), .Y(_427_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_427_), .Y(_428_) );
AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_426_), .Y(_141__0_) );
INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(data_226__1_), .Y(_429_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf1), .B(_361__bF_buf5), .C(_429_), .Y(_430_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_427_), .Y(_431_) );
AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_430_), .Y(_141__1_) );
INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(data_226__2_), .Y(_432_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf0), .B(_361__bF_buf4), .C(_432_), .Y(_433_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_427_), .Y(_434_) );
AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_433_), .Y(_141__2_) );
INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(data_226__3_), .Y(_435_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf3), .B(_361__bF_buf3), .C(_435_), .Y(_436_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_427_), .Y(_437_) );
AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_436_), .Y(_141__3_) );
INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(data_226__4_), .Y(_438_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf2), .B(_361__bF_buf2), .C(_438_), .Y(_439_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_427_), .Y(_440_) );
AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_439_), .Y(_141__4_) );
INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(data_226__5_), .Y(_441_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf1), .B(_361__bF_buf1), .C(_441_), .Y(_442_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_427_), .Y(_443_) );
AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_442_), .Y(_141__5_) );
INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(data_226__6_), .Y(_444_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf0), .B(_361__bF_buf0), .C(_444_), .Y(_445_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_427_), .Y(_446_) );
AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_445_), .Y(_141__6_) );
INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(data_226__7_), .Y(_447_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf3), .B(_361__bF_buf5), .C(_447_), .Y(_448_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_427_), .Y(_449_) );
AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_448_), .Y(_141__7_) );
INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(data_226__8_), .Y(_450_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf2), .B(_361__bF_buf4), .C(_450_), .Y(_451_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_427_), .Y(_452_) );
AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_451_), .Y(_141__8_) );
INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(data_226__9_), .Y(_453_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf1), .B(_361__bF_buf3), .C(_453_), .Y(_454_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_427_), .Y(_455_) );
AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_454_), .Y(_141__9_) );
INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(data_226__10_), .Y(_456_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf0), .B(_361__bF_buf2), .C(_456_), .Y(_457_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_427_), .Y(_458_) );
AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_457_), .Y(_141__10_) );
INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(data_226__11_), .Y(_459_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf3), .B(_361__bF_buf1), .C(_459_), .Y(_460_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_427_), .Y(_461_) );
AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_460_), .Y(_141__11_) );
INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(data_226__12_), .Y(_462_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf2), .B(_361__bF_buf0), .C(_462_), .Y(_463_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_427_), .Y(_464_) );
AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_463_), .Y(_141__12_) );
INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(data_226__13_), .Y(_465_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf1), .B(_361__bF_buf5), .C(_465_), .Y(_466_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_427_), .Y(_467_) );
AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_466_), .Y(_141__13_) );
INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(data_226__14_), .Y(_468_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf0), .B(_361__bF_buf4), .C(_468_), .Y(_469_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_427_), .Y(_470_) );
AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_469_), .Y(_141__14_) );
INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(data_226__15_), .Y(_471_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_425__bF_buf3), .B(_361__bF_buf3), .C(_471_), .Y(_472_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf2), .B(_427_), .Y(_473_) );
AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_472_), .Y(_141__15_) );
INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(data_225__0_), .Y(_474_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(_15684_), .Y(_475_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_15005__bF_buf0), .B(_475_), .C(_422_), .Y(_476_) );
INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(_476_), .Y(_477_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf3), .B(_477_), .C(_362_), .Y(_478_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_361__bF_buf2), .Y(_479_) );
MUX2X1 MUX2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_474_), .S(_479_), .Y(_140__0_) );
INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(data_225__1_), .Y(_480_) );
MUX2X1 MUX2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_480_), .S(_479_), .Y(_140__1_) );
INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(data_225__2_), .Y(_481_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf1), .B(_478_), .C(_481_), .Y(_482_) );
NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_476_), .C(_371_), .Y(_483_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_483_), .C(_342__bF_buf2), .Y(_484_) );
AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_482_), .Y(_140__2_) );
INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(data_225__3_), .Y(_485_) );
MUX2X1 MUX2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_485_), .S(_479_), .Y(_140__3_) );
INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(data_225__4_), .Y(_486_) );
MUX2X1 MUX2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_486_), .S(_479_), .Y(_140__4_) );
INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(data_225__5_), .Y(_487_) );
MUX2X1 MUX2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_487_), .S(_479_), .Y(_140__5_) );
INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(data_225__6_), .Y(_488_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf0), .B(_478_), .C(_488_), .Y(_489_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_483_), .C(_342__bF_buf1), .Y(_490_) );
AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_489_), .Y(_140__6_) );
INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(data_225__7_), .Y(_491_) );
MUX2X1 MUX2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_491_), .S(_479_), .Y(_140__7_) );
INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(data_225__8_), .Y(_492_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf5), .B(_478_), .C(_492_), .Y(_493_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_483_), .C(_342__bF_buf0), .Y(_494_) );
AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_493_), .Y(_140__8_) );
INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(data_225__9_), .Y(_495_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf4), .B(_478_), .C(_495_), .Y(_496_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_483_), .C(_342__bF_buf4), .Y(_497_) );
AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_496_), .Y(_140__9_) );
INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(data_225__10_), .Y(_498_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf3), .B(_478_), .C(_498_), .Y(_499_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_483_), .C(_342__bF_buf3), .Y(_500_) );
AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_499_), .Y(_140__10_) );
INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(data_225__11_), .Y(_501_) );
MUX2X1 MUX2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_501_), .S(_479_), .Y(_140__11_) );
INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(data_225__12_), .Y(_502_) );
MUX2X1 MUX2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_502_), .S(_479_), .Y(_140__12_) );
INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(data_225__13_), .Y(_503_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf2), .B(_478_), .C(_503_), .Y(_504_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_483_), .C(_342__bF_buf2), .Y(_505_) );
AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_504_), .Y(_140__13_) );
INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(data_225__14_), .Y(_506_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf1), .B(_478_), .C(_506_), .Y(_507_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_483_), .C(_342__bF_buf1), .Y(_508_) );
AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_507_), .Y(_140__14_) );
INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(data_225__15_), .Y(_509_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf0), .B(_478_), .C(_509_), .Y(_510_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_483_), .C(_342__bF_buf0), .Y(_511_) );
AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_510_), .Y(_140__15_) );
INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(data_224__0_), .Y(_512_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf3), .B(_14975_), .C(_15575__bF_buf2), .Y(_513_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf0), .B(_15006__bF_buf0), .C(_513_), .Y(_514_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_15028_), .Y(_515_) );
INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(_515_), .Y(_516_) );
NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_15592_), .B(_516_), .C(_15074__bF_buf4), .Y(_517_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_517_), .C(_15949__bF_buf8), .Y(_518_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf3), .B(_14882__bF_buf15_bF_buf2), .C(_512_), .Y(_519_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14_bF_buf2), .B(_518__bF_buf2), .Y(_520_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_520_), .Y(_521_) );
AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_519_), .Y(_139__0_) );
INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(data_224__1_), .Y(_522_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf1), .B(_14882__bF_buf13_bF_buf2), .C(_522_), .Y(_523_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_520_), .Y(_524_) );
AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_523_), .Y(_139__1_) );
INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(data_224__2_), .Y(_525_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf0), .B(_14882__bF_buf12), .C(_525_), .Y(_526_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_520_), .Y(_527_) );
AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_526_), .Y(_139__2_) );
INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(data_224__3_), .Y(_528_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf3), .B(_14882__bF_buf11), .C(_528_), .Y(_529_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_520_), .Y(_530_) );
AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_529_), .Y(_139__3_) );
INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(data_224__4_), .Y(_531_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf2), .B(_14882__bF_buf10), .C(_531_), .Y(_532_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_520_), .Y(_533_) );
AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_532_), .Y(_139__4_) );
INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(data_224__5_), .Y(_534_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf1), .B(_14882__bF_buf9), .C(_534_), .Y(_535_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_520_), .Y(_536_) );
AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_535_), .Y(_139__5_) );
INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(data_224__6_), .Y(_537_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf0), .B(_14882__bF_buf8), .C(_537_), .Y(_538_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_520_), .Y(_539_) );
AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_538_), .Y(_139__6_) );
INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(data_224__7_), .Y(_540_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf3), .B(_14882__bF_buf7), .C(_540_), .Y(_541_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_15570_), .B(_515_), .C(_15183__bF_buf7), .Y(_542_) );
NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_15900__bF_buf6), .B(_341_), .C(_542_), .Y(_543_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf5), .B(_14908__bF_buf12), .C(_543_), .Y(_544_) );
AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_541_), .Y(_139__7_) );
INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(data_224__8_), .Y(_545_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf2), .B(_14882__bF_buf6), .C(_545_), .Y(_546_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_520_), .Y(_547_) );
AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_546_), .Y(_139__8_) );
INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(data_224__9_), .Y(_548_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf1), .B(_14882__bF_buf5), .C(_548_), .Y(_549_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_520_), .Y(_550_) );
AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_549_), .Y(_139__9_) );
INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(data_224__10_), .Y(_551_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf0), .B(_14882__bF_buf4), .C(_551_), .Y(_552_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_520_), .Y(_553_) );
AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_552_), .Y(_139__10_) );
INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(data_224__11_), .Y(_554_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf3), .B(_14882__bF_buf3), .C(_554_), .Y(_555_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_520_), .Y(_556_) );
AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_555_), .Y(_139__11_) );
INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(data_224__12_), .Y(_557_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf2), .B(_14882__bF_buf2), .C(_557_), .Y(_558_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_14920__bF_buf12), .C(_543_), .Y(_559_) );
AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_558_), .Y(_139__12_) );
INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(data_224__13_), .Y(_560_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf1), .B(_14882__bF_buf1), .C(_560_), .Y(_561_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_520_), .Y(_562_) );
AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_561_), .Y(_139__13_) );
INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(data_224__14_), .Y(_563_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf0), .B(_14882__bF_buf0), .C(_563_), .Y(_564_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_520_), .Y(_565_) );
AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_564_), .Y(_139__14_) );
INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(data_224__15_), .Y(_566_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_518__bF_buf3), .B(_14882__bF_buf15_bF_buf1), .C(_566_), .Y(_567_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_520_), .Y(_568_) );
AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_567_), .Y(_139__15_) );
INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(data_223__0_), .Y(_569_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf3), .B(_14942__bF_buf3), .C(_15766_), .Y(_570_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(_570_), .Y(_571_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_15006__bF_buf4), .C(_513_), .Y(_572_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_515_), .Y(_573_) );
INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(_573_), .Y(_574_) );
NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_574_), .C(_371_), .Y(_575_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf3), .B(_575_), .Y(_576_) );
MUX2X1 MUX2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_14932__bF_buf0), .S(_576_), .Y(_138__0_) );
INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(data_223__1_), .Y(_577_) );
MUX2X1 MUX2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_14894__bF_buf14), .S(_576_), .Y(_138__1_) );
INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(data_223__2_), .Y(_578_) );
MUX2X1 MUX2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_14897__bF_buf14), .S(_576_), .Y(_138__2_) );
INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(data_223__3_), .Y(_579_) );
MUX2X1 MUX2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_14899__bF_buf14), .S(_576_), .Y(_138__3_) );
INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(data_223__4_), .Y(_580_) );
MUX2X1 MUX2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_14902__bF_buf11), .S(_576_), .Y(_138__4_) );
INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(data_223__5_), .Y(_581_) );
MUX2X1 MUX2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_14903__bF_buf12), .S(_576_), .Y(_138__5_) );
INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(data_223__6_), .Y(_582_) );
MUX2X1 MUX2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_15049__bF_buf0), .S(_576_), .Y(_138__6_) );
INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(data_223__7_), .Y(_583_) );
MUX2X1 MUX2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_14908__bF_buf11), .S(_576_), .Y(_138__7_) );
INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(data_223__8_), .Y(_584_) );
MUX2X1 MUX2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_15052__bF_buf13), .S(_576_), .Y(_138__8_) );
INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(data_223__9_), .Y(_585_) );
MUX2X1 MUX2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_14913__bF_buf0), .S(_576_), .Y(_138__9_) );
INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(data_223__10_), .Y(_586_) );
MUX2X1 MUX2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_15055__bF_buf13), .S(_576_), .Y(_138__10_) );
INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(data_223__11_), .Y(_587_) );
MUX2X1 MUX2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_14918__bF_buf12), .S(_576_), .Y(_138__11_) );
INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(data_223__12_), .Y(_588_) );
MUX2X1 MUX2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_14920__bF_buf11), .S(_576_), .Y(_138__12_) );
INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(data_223__13_), .Y(_589_) );
MUX2X1 MUX2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_14924__bF_buf12), .S(_576_), .Y(_138__13_) );
INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(data_223__14_), .Y(_590_) );
MUX2X1 MUX2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_15060__bF_buf0), .S(_576_), .Y(_138__14_) );
INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(data_223__15_), .Y(_591_) );
MUX2X1 MUX2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_15062__bF_buf13), .S(_576_), .Y(_138__15_) );
INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf3), .Y(_592_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_15793__bF_buf2), .Y(_593_) );
INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(data_222__0_), .Y(_594_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15006__bF_buf2), .C(_594_), .Y(_595_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf0), .B(_593_), .C(_595_), .Y(_596_) );
INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(_596_), .Y(_137__0_) );
INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(data_222__1_), .Y(_597_) );
MUX2X1 MUX2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_14894__bF_buf13), .S(_593_), .Y(_137__1_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf1), .B(_15788__bF_buf7), .Y(_598_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(data_222__2_), .B(_598_), .Y(_599_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf13), .B(_598_), .C(_599_), .Y(_137__2_) );
INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(data_222__3_), .Y(_600_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15006__bF_buf0), .C(_600_), .Y(_601_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_598_), .Y(_602_) );
AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_601_), .Y(_137__3_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(data_222__4_), .B(_598_), .Y(_603_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_598_), .C(_603_), .Y(_137__4_) );
INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(data_222__5_), .Y(_604_) );
MUX2X1 MUX2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_14903__bF_buf11), .S(_593_), .Y(_137__5_) );
INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(data_222__6_), .Y(_605_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15006__bF_buf4), .C(_605_), .Y(_606_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_592_), .C(_15793__bF_buf1), .Y(_607_) );
AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_607_), .Y(_137__6_) );
INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(data_222__7_), .Y(_608_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15006__bF_buf3), .C(_608_), .Y(_609_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_592_), .C(_15793__bF_buf0), .Y(_610_) );
AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_610_), .Y(_137__7_) );
INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(data_222__8_), .Y(_611_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15006__bF_buf2), .C(_611_), .Y(_612_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf4), .B(_593_), .C(_612_), .Y(_613_) );
INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(_613_), .Y(_137__8_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(data_222__9_), .B(_598_), .Y(_614_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf14), .B(_598_), .C(_614_), .Y(_137__9_) );
INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(data_222__10_), .Y(_615_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15006__bF_buf1), .C(_615_), .Y(_616_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf4), .B(_593_), .C(_616_), .Y(_617_) );
INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(_617_), .Y(_137__10_) );
INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(data_222__11_), .Y(_618_) );
MUX2X1 MUX2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_14918__bF_buf11), .S(_593_), .Y(_137__11_) );
INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(data_222__12_), .Y(_619_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15006__bF_buf0), .C(_619_), .Y(_620_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf1), .B(_593_), .C(_620_), .Y(_621_) );
INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(_621_), .Y(_137__12_) );
INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(data_222__13_), .Y(_622_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15006__bF_buf4), .C(_622_), .Y(_623_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf0), .B(_593_), .C(_623_), .Y(_624_) );
INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(_624_), .Y(_137__13_) );
INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(data_222__14_), .Y(_625_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15006__bF_buf3), .C(_625_), .Y(_626_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf0), .B(_593_), .C(_626_), .Y(_627_) );
INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(_627_), .Y(_137__14_) );
INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(data_222__15_), .Y(_628_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15006__bF_buf2), .C(_628_), .Y(_629_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_592_), .C(_15793__bF_buf5), .Y(_630_) );
AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_630_), .Y(_137__15_) );
INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(data_221__0_), .Y(_631_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf2), .B(_573_), .C(_362_), .Y(_632_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf5), .B(_542_), .C(_632_), .Y(_633_) );
NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_15841_), .B(_341_), .C(_15900__bF_buf5), .Y(_634_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf1), .B(_15034_), .C(_15570_), .Y(_635_) );
INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(_635_), .Y(_636_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_15835_), .B(_15006__bF_buf0), .C(_513_), .Y(_637_) );
INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(_637_), .Y(_638_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_638_), .C(_634_), .Y(_639_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_631_), .Y(_640_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_543_), .Y(_641_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_15832_), .B(_340_), .C(_15949__bF_buf7), .Y(_642_) );
NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_637_), .C(_642_), .Y(_643_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_641_), .C(_643_), .Y(_644_) );
AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_640_), .Y(_136__0_) );
INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(data_221__1_), .Y(_645_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_645_), .Y(_646_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_641_), .C(_643_), .Y(_647_) );
AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_646_), .Y(_136__1_) );
INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(data_221__2_), .Y(_648_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_643_), .Y(_649_) );
MUX2X1 MUX2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_14897__bF_buf12), .S(_649_), .Y(_136__2_) );
INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(data_221__3_), .Y(_650_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_650_), .Y(_651_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_641_), .C(_643_), .Y(_652_) );
AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_651_), .Y(_136__3_) );
INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(data_221__4_), .Y(_653_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_653_), .Y(_654_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_641_), .C(_643_), .Y(_655_) );
AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_654_), .Y(_136__4_) );
INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(data_221__5_), .Y(_656_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_656_), .Y(_657_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_641_), .C(_643_), .Y(_658_) );
AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_657_), .Y(_136__5_) );
INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(data_221__6_), .Y(_659_) );
MUX2X1 MUX2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_15049__bF_buf13), .S(_649_), .Y(_136__6_) );
INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(data_221__7_), .Y(_660_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_660_), .Y(_661_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_641_), .C(_643_), .Y(_662_) );
AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_661_), .Y(_136__7_) );
INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(data_221__8_), .Y(_663_) );
MUX2X1 MUX2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_15052__bF_buf12), .S(_649_), .Y(_136__8_) );
INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(data_221__9_), .Y(_664_) );
MUX2X1 MUX2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_14913__bF_buf13), .S(_649_), .Y(_136__9_) );
INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(data_221__10_), .Y(_665_) );
MUX2X1 MUX2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_15055__bF_buf12), .S(_649_), .Y(_136__10_) );
INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(data_221__11_), .Y(_666_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_666_), .Y(_667_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_641_), .C(_643_), .Y(_668_) );
AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_667_), .Y(_136__11_) );
INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(data_221__12_), .Y(_669_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_633_), .C(_669_), .Y(_670_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_641_), .C(_643_), .Y(_671_) );
AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_670_), .Y(_136__12_) );
INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(data_221__13_), .Y(_672_) );
MUX2X1 MUX2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_14924__bF_buf11), .S(_649_), .Y(_136__13_) );
INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(data_221__14_), .Y(_673_) );
MUX2X1 MUX2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_15060__bF_buf14), .S(_649_), .Y(_136__14_) );
INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(data_221__15_), .Y(_674_) );
MUX2X1 MUX2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_15062__bF_buf11), .S(_649_), .Y(_136__15_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_634_), .Y(_675_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15006__bF_buf4), .C(_513_), .Y(_676_) );
INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(_676_), .Y(_677_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_677_), .C(_518__bF_buf2), .Y(_678_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf7), .B(_675_), .Y(_679_) );
INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(data_220__0_), .Y(_680_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_675_), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_0_bF_buf4), .C(_681_), .Y(_682_) );
INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(_682_), .Y(_135__0_) );
INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(data_220__1_), .Y(_683_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf5), .B(_675_), .C(_683_), .Y(_684_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_1_bF_buf1), .C(_684_), .Y(_685_) );
INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(_685_), .Y(_135__1_) );
INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(data_220__2_), .Y(_686_) );
MUX2X1 MUX2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_14897__bF_buf11), .S(_679_), .Y(_135__2_) );
INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(data_220__3_), .Y(_687_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf4), .B(_675_), .C(_687_), .Y(_688_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_3_bF_buf1), .C(_688_), .Y(_689_) );
INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(_689_), .Y(_135__3_) );
INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(data_220__4_), .Y(_690_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf3), .B(_675_), .C(_690_), .Y(_691_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_4_bF_buf1), .C(_691_), .Y(_692_) );
INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(_692_), .Y(_135__4_) );
INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(data_220__5_), .Y(_693_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_675_), .C(_693_), .Y(_694_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_5_bF_buf0), .C(_694_), .Y(_695_) );
INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(_695_), .Y(_135__5_) );
INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(data_220__6_), .Y(_696_) );
MUX2X1 MUX2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_15049__bF_buf12), .S(_679_), .Y(_135__6_) );
INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(data_220__7_), .Y(_697_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf1), .B(_675_), .C(_697_), .Y(_698_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_7_bF_buf2), .C(_698_), .Y(_699_) );
INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(_699_), .Y(_135__7_) );
INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(data_220__8_), .Y(_700_) );
MUX2X1 MUX2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_15052__bF_buf11), .S(_679_), .Y(_135__8_) );
INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(data_220__9_), .Y(_701_) );
MUX2X1 MUX2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_14913__bF_buf12), .S(_679_), .Y(_135__9_) );
INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(data_220__10_), .Y(_702_) );
MUX2X1 MUX2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_15055__bF_buf11), .S(_679_), .Y(_135__10_) );
INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(data_220__11_), .Y(_703_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf0), .B(_675_), .C(_703_), .Y(_704_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_11_bF_buf0), .C(_704_), .Y(_705_) );
INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_135__11_) );
INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(data_220__12_), .Y(_706_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf7), .B(_675_), .C(_706_), .Y(_707_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(IDATA_PROG_data_12_bF_buf0), .C(_707_), .Y(_708_) );
INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(_708_), .Y(_135__12_) );
INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(data_220__13_), .Y(_709_) );
MUX2X1 MUX2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_14924__bF_buf10), .S(_679_), .Y(_135__13_) );
INVX1 INVX1_596 ( .gnd(gnd), .vdd(vdd), .A(data_220__14_), .Y(_710_) );
MUX2X1 MUX2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_15060__bF_buf13), .S(_679_), .Y(_135__14_) );
INVX1 INVX1_597 ( .gnd(gnd), .vdd(vdd), .A(data_220__15_), .Y(_711_) );
MUX2X1 MUX2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_15062__bF_buf10), .S(_679_), .Y(_135__15_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .B(_15006__bF_buf3), .C(IDATA_PROG_write_bF_buf2), .Y(_712_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_15951_), .C(_712_), .Y(_713_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_713_), .C(_342__bF_buf4), .Y(_714_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_714_), .Y(_715_) );
INVX1 INVX1_598 ( .gnd(gnd), .vdd(vdd), .A(data_219__0_), .Y(_716_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf5), .B(_714_), .C(_716_), .Y(_717_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_0_bF_buf3), .C(_717_), .Y(_718_) );
INVX1 INVX1_599 ( .gnd(gnd), .vdd(vdd), .A(_718_), .Y(_133__0_) );
INVX1 INVX1_600 ( .gnd(gnd), .vdd(vdd), .A(data_219__1_), .Y(_719_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf4), .B(_714_), .C(_719_), .Y(_720_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_1_bF_buf0), .C(_720_), .Y(_721_) );
INVX1 INVX1_601 ( .gnd(gnd), .vdd(vdd), .A(_721_), .Y(_133__1_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_678__bF_buf3), .Y(_722_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(data_219__2_), .B(_722_), .Y(_723_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_722_), .C(_723_), .Y(_133__2_) );
INVX1 INVX1_602 ( .gnd(gnd), .vdd(vdd), .A(data_219__3_), .Y(_724_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_714_), .C(_724_), .Y(_725_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_3_bF_buf0), .C(_725_), .Y(_726_) );
INVX1 INVX1_603 ( .gnd(gnd), .vdd(vdd), .A(_726_), .Y(_133__3_) );
INVX1 INVX1_604 ( .gnd(gnd), .vdd(vdd), .A(data_219__4_), .Y(_727_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf1), .B(_714_), .C(_727_), .Y(_728_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_4_bF_buf0), .C(_728_), .Y(_729_) );
INVX1 INVX1_605 ( .gnd(gnd), .vdd(vdd), .A(_729_), .Y(_133__4_) );
INVX1 INVX1_606 ( .gnd(gnd), .vdd(vdd), .A(data_219__5_), .Y(_730_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf0), .B(_714_), .C(_730_), .Y(_731_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_5_bF_buf4), .C(_731_), .Y(_732_) );
INVX1 INVX1_607 ( .gnd(gnd), .vdd(vdd), .A(_732_), .Y(_133__5_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(data_219__6_), .B(_722_), .Y(_733_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_722_), .C(_733_), .Y(_133__6_) );
INVX1 INVX1_608 ( .gnd(gnd), .vdd(vdd), .A(data_219__7_), .Y(_734_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf7), .B(_714_), .C(_734_), .Y(_735_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_7_bF_buf1), .C(_735_), .Y(_736_) );
INVX1 INVX1_609 ( .gnd(gnd), .vdd(vdd), .A(_736_), .Y(_133__7_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(data_219__8_), .B(_722_), .Y(_737_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_722_), .C(_737_), .Y(_133__8_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(data_219__9_), .B(_722_), .Y(_738_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_722_), .C(_738_), .Y(_133__9_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(data_219__10_), .B(_722_), .Y(_739_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_722_), .C(_739_), .Y(_133__10_) );
INVX1 INVX1_610 ( .gnd(gnd), .vdd(vdd), .A(data_219__11_), .Y(_740_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_714_), .C(_740_), .Y(_741_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_11_bF_buf4), .C(_741_), .Y(_742_) );
INVX1 INVX1_611 ( .gnd(gnd), .vdd(vdd), .A(_742_), .Y(_133__11_) );
INVX1 INVX1_612 ( .gnd(gnd), .vdd(vdd), .A(data_219__12_), .Y(_743_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf5), .B(_714_), .C(_743_), .Y(_744_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(IDATA_PROG_data_12_bF_buf4), .C(_744_), .Y(_745_) );
INVX1 INVX1_613 ( .gnd(gnd), .vdd(vdd), .A(_745_), .Y(_133__12_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(data_219__13_), .B(_722_), .Y(_746_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_722_), .C(_746_), .Y(_133__13_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(data_219__14_), .B(_722_), .Y(_747_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_722_), .C(_747_), .Y(_133__14_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(data_219__15_), .B(_722_), .Y(_748_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_722_), .C(_748_), .Y(_133__15_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_14964_), .Y(_749_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_749_), .Y(_750_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14_bF_buf1), .B(_592_), .Y(_751_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf2), .B(_15160_), .C(_750_), .D(_751_), .Y(_752_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf4), .B(_592_), .C(_752_), .Y(_753_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_753_), .C(_342__bF_buf3), .Y(_754_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf4), .B(_754_), .Y(_755_) );
INVX1 INVX1_614 ( .gnd(gnd), .vdd(vdd), .A(data_218__0_), .Y(_756_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf3), .B(_754_), .C(_756_), .Y(_757_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_0_bF_buf2), .C(_757_), .Y(_758_) );
INVX1 INVX1_615 ( .gnd(gnd), .vdd(vdd), .A(_758_), .Y(_132__0_) );
INVX1 INVX1_616 ( .gnd(gnd), .vdd(vdd), .A(data_218__1_), .Y(_759_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_754_), .C(_759_), .Y(_760_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_1_bF_buf4), .C(_760_), .Y(_761_) );
INVX1 INVX1_617 ( .gnd(gnd), .vdd(vdd), .A(_761_), .Y(_132__1_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_678__bF_buf1), .Y(_762_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(data_218__2_), .B(_762_), .Y(_763_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_762_), .C(_763_), .Y(_132__2_) );
INVX1 INVX1_618 ( .gnd(gnd), .vdd(vdd), .A(data_218__3_), .Y(_764_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf0), .B(_754_), .C(_764_), .Y(_765_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_3_bF_buf4), .C(_765_), .Y(_766_) );
INVX1 INVX1_619 ( .gnd(gnd), .vdd(vdd), .A(_766_), .Y(_132__3_) );
INVX1 INVX1_620 ( .gnd(gnd), .vdd(vdd), .A(data_218__4_), .Y(_767_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf7), .B(_754_), .C(_767_), .Y(_768_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_4_bF_buf4), .C(_768_), .Y(_769_) );
INVX1 INVX1_621 ( .gnd(gnd), .vdd(vdd), .A(_769_), .Y(_132__4_) );
INVX1 INVX1_622 ( .gnd(gnd), .vdd(vdd), .A(data_218__5_), .Y(_770_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_754_), .C(_770_), .Y(_771_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_5_bF_buf3), .C(_771_), .Y(_772_) );
INVX1 INVX1_623 ( .gnd(gnd), .vdd(vdd), .A(_772_), .Y(_132__5_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(data_218__6_), .B(_762_), .Y(_773_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_762_), .C(_773_), .Y(_132__6_) );
INVX1 INVX1_624 ( .gnd(gnd), .vdd(vdd), .A(data_218__7_), .Y(_774_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf5), .B(_754_), .C(_774_), .Y(_775_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_7_bF_buf0), .C(_775_), .Y(_776_) );
INVX1 INVX1_625 ( .gnd(gnd), .vdd(vdd), .A(_776_), .Y(_132__7_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(data_218__8_), .B(_762_), .Y(_777_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_762_), .C(_777_), .Y(_132__8_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(data_218__9_), .B(_762_), .Y(_778_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_762_), .C(_778_), .Y(_132__9_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(data_218__10_), .B(_762_), .Y(_779_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_762_), .C(_779_), .Y(_132__10_) );
INVX1 INVX1_626 ( .gnd(gnd), .vdd(vdd), .A(data_218__11_), .Y(_780_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf4), .B(_754_), .C(_780_), .Y(_781_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_11_bF_buf3), .C(_781_), .Y(_782_) );
INVX1 INVX1_627 ( .gnd(gnd), .vdd(vdd), .A(_782_), .Y(_132__11_) );
INVX1 INVX1_628 ( .gnd(gnd), .vdd(vdd), .A(data_218__12_), .Y(_783_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf3), .B(_754_), .C(_783_), .Y(_784_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(IDATA_PROG_data_12_bF_buf3), .C(_784_), .Y(_785_) );
INVX1 INVX1_629 ( .gnd(gnd), .vdd(vdd), .A(_785_), .Y(_132__12_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(data_218__13_), .B(_762_), .Y(_786_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_762_), .C(_786_), .Y(_132__13_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(data_218__14_), .B(_762_), .Y(_787_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_762_), .C(_787_), .Y(_132__14_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(data_218__15_), .B(_762_), .Y(_788_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_762_), .C(_788_), .Y(_132__15_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_16055_), .B(_749_), .Y(_789_) );
INVX1 INVX1_630 ( .gnd(gnd), .vdd(vdd), .A(_789_), .Y(_790_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf13_bF_buf1), .B(_592_), .C(_790_), .Y(_791_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_791_), .C(_342__bF_buf2), .Y(_792_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_792_), .Y(_793_) );
INVX1 INVX1_631 ( .gnd(gnd), .vdd(vdd), .A(data_217__0_), .Y(_794_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf1), .B(_792_), .C(_794_), .Y(_795_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_0_bF_buf1), .C(_795_), .Y(_796_) );
INVX1 INVX1_632 ( .gnd(gnd), .vdd(vdd), .A(_796_), .Y(_131__0_) );
INVX1 INVX1_633 ( .gnd(gnd), .vdd(vdd), .A(data_217__1_), .Y(_797_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf0), .B(_792_), .C(_797_), .Y(_798_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_1_bF_buf3), .C(_798_), .Y(_799_) );
INVX1 INVX1_634 ( .gnd(gnd), .vdd(vdd), .A(_799_), .Y(_131__1_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_678__bF_buf7), .Y(_800_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(data_217__2_), .B(_800_), .Y(_801_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_800_), .C(_801_), .Y(_131__2_) );
INVX1 INVX1_635 ( .gnd(gnd), .vdd(vdd), .A(data_217__3_), .Y(_802_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_792_), .C(_802_), .Y(_803_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_3_bF_buf3), .C(_803_), .Y(_804_) );
INVX1 INVX1_636 ( .gnd(gnd), .vdd(vdd), .A(_804_), .Y(_131__3_) );
INVX1 INVX1_637 ( .gnd(gnd), .vdd(vdd), .A(data_217__4_), .Y(_805_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf5), .B(_792_), .C(_805_), .Y(_806_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_4_bF_buf3), .C(_806_), .Y(_807_) );
INVX1 INVX1_638 ( .gnd(gnd), .vdd(vdd), .A(_807_), .Y(_131__4_) );
INVX1 INVX1_639 ( .gnd(gnd), .vdd(vdd), .A(data_217__5_), .Y(_808_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf4), .B(_792_), .C(_808_), .Y(_809_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_5_bF_buf2), .C(_809_), .Y(_810_) );
INVX1 INVX1_640 ( .gnd(gnd), .vdd(vdd), .A(_810_), .Y(_131__5_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(data_217__6_), .B(_800_), .Y(_811_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_800_), .C(_811_), .Y(_131__6_) );
INVX1 INVX1_641 ( .gnd(gnd), .vdd(vdd), .A(data_217__7_), .Y(_812_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf3), .B(_792_), .C(_812_), .Y(_813_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_7_bF_buf5), .C(_813_), .Y(_814_) );
INVX1 INVX1_642 ( .gnd(gnd), .vdd(vdd), .A(_814_), .Y(_131__7_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(data_217__8_), .B(_800_), .Y(_815_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_800_), .C(_815_), .Y(_131__8_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(data_217__9_), .B(_800_), .Y(_816_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_800_), .C(_816_), .Y(_131__9_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(data_217__10_), .B(_800_), .Y(_817_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_800_), .C(_817_), .Y(_131__10_) );
INVX1 INVX1_643 ( .gnd(gnd), .vdd(vdd), .A(data_217__11_), .Y(_818_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_792_), .C(_818_), .Y(_819_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_11_bF_buf2), .C(_819_), .Y(_820_) );
INVX1 INVX1_644 ( .gnd(gnd), .vdd(vdd), .A(_820_), .Y(_131__11_) );
INVX1 INVX1_645 ( .gnd(gnd), .vdd(vdd), .A(data_217__12_), .Y(_821_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf1), .B(_792_), .C(_821_), .Y(_822_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(IDATA_PROG_data_12_bF_buf2), .C(_822_), .Y(_823_) );
INVX1 INVX1_646 ( .gnd(gnd), .vdd(vdd), .A(_823_), .Y(_131__12_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(data_217__13_), .B(_800_), .Y(_824_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_800_), .C(_824_), .Y(_131__13_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(data_217__14_), .B(_800_), .Y(_825_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_800_), .C(_825_), .Y(_131__14_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(data_217__15_), .B(_800_), .Y(_826_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_800_), .C(_826_), .Y(_131__15_) );
INVX1 INVX1_647 ( .gnd(gnd), .vdd(vdd), .A(data_216__0_), .Y(_827_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf3), .B(_592_), .C(_15592_), .Y(_828_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_14977__bF_buf0), .B(_15006__bF_buf1), .C(_828_), .Y(_829_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_829_), .Y(_830_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf0), .B(_830_), .Y(_831_) );
MUX2X1 MUX2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_827_), .S(_831_), .Y(_130__0_) );
INVX1 INVX1_648 ( .gnd(gnd), .vdd(vdd), .A(data_216__1_), .Y(_832_) );
MUX2X1 MUX2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_832_), .S(_831_), .Y(_130__1_) );
INVX1 INVX1_649 ( .gnd(gnd), .vdd(vdd), .A(data_216__2_), .Y(_833_) );
MUX2X1 MUX2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_833_), .S(_831_), .Y(_130__2_) );
INVX1 INVX1_650 ( .gnd(gnd), .vdd(vdd), .A(data_216__3_), .Y(_834_) );
MUX2X1 MUX2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_834_), .S(_831_), .Y(_130__3_) );
INVX1 INVX1_651 ( .gnd(gnd), .vdd(vdd), .A(data_216__4_), .Y(_835_) );
MUX2X1 MUX2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_835_), .S(_831_), .Y(_130__4_) );
INVX1 INVX1_652 ( .gnd(gnd), .vdd(vdd), .A(data_216__5_), .Y(_836_) );
MUX2X1 MUX2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_836_), .S(_831_), .Y(_130__5_) );
INVX1 INVX1_653 ( .gnd(gnd), .vdd(vdd), .A(data_216__6_), .Y(_837_) );
MUX2X1 MUX2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_837_), .S(_831_), .Y(_130__6_) );
INVX1 INVX1_654 ( .gnd(gnd), .vdd(vdd), .A(data_216__7_), .Y(_838_) );
MUX2X1 MUX2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_838_), .S(_831_), .Y(_130__7_) );
INVX1 INVX1_655 ( .gnd(gnd), .vdd(vdd), .A(data_216__8_), .Y(_839_) );
MUX2X1 MUX2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_839_), .S(_831_), .Y(_130__8_) );
INVX1 INVX1_656 ( .gnd(gnd), .vdd(vdd), .A(data_216__9_), .Y(_840_) );
MUX2X1 MUX2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_840_), .S(_831_), .Y(_130__9_) );
INVX1 INVX1_657 ( .gnd(gnd), .vdd(vdd), .A(data_216__10_), .Y(_841_) );
MUX2X1 MUX2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_841_), .S(_831_), .Y(_130__10_) );
INVX1 INVX1_658 ( .gnd(gnd), .vdd(vdd), .A(data_216__11_), .Y(_842_) );
MUX2X1 MUX2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_842_), .S(_831_), .Y(_130__11_) );
INVX1 INVX1_659 ( .gnd(gnd), .vdd(vdd), .A(data_216__12_), .Y(_843_) );
MUX2X1 MUX2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_843_), .S(_831_), .Y(_130__12_) );
INVX1 INVX1_660 ( .gnd(gnd), .vdd(vdd), .A(data_216__13_), .Y(_844_) );
MUX2X1 MUX2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_844_), .S(_831_), .Y(_130__13_) );
INVX1 INVX1_661 ( .gnd(gnd), .vdd(vdd), .A(data_216__14_), .Y(_845_) );
MUX2X1 MUX2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_845_), .S(_831_), .Y(_130__14_) );
INVX1 INVX1_662 ( .gnd(gnd), .vdd(vdd), .A(data_216__15_), .Y(_846_) );
MUX2X1 MUX2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_846_), .S(_831_), .Y(_130__15_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_14977__bF_buf3), .B(IDATA_PROG_addr[1]), .C(IDATA_PROG_write_bF_buf0), .Y(_847_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_15364_), .Y(_848_) );
INVX1 INVX1_663 ( .gnd(gnd), .vdd(vdd), .A(_848_), .Y(_849_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf12), .B(_592_), .C(_849_), .Y(_850_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_850_), .C(_342__bF_buf1), .Y(_851_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf7), .B(_851_), .Y(_852_) );
INVX1 INVX1_664 ( .gnd(gnd), .vdd(vdd), .A(data_215__0_), .Y(_853_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_851_), .C(_853_), .Y(_854_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_0_bF_buf0), .C(_854_), .Y(_855_) );
INVX1 INVX1_665 ( .gnd(gnd), .vdd(vdd), .A(_855_), .Y(_129__0_) );
INVX1 INVX1_666 ( .gnd(gnd), .vdd(vdd), .A(data_215__1_), .Y(_856_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf5), .B(_851_), .C(_856_), .Y(_857_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_1_bF_buf2), .C(_857_), .Y(_858_) );
INVX1 INVX1_667 ( .gnd(gnd), .vdd(vdd), .A(_858_), .Y(_129__1_) );
INVX1 INVX1_668 ( .gnd(gnd), .vdd(vdd), .A(data_215__2_), .Y(_859_) );
MUX2X1 MUX2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_14897__bF_buf6), .S(_852_), .Y(_129__2_) );
INVX1 INVX1_669 ( .gnd(gnd), .vdd(vdd), .A(data_215__3_), .Y(_860_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf4), .B(_851_), .C(_860_), .Y(_861_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_3_bF_buf2), .C(_861_), .Y(_862_) );
INVX1 INVX1_670 ( .gnd(gnd), .vdd(vdd), .A(_862_), .Y(_129__3_) );
INVX1 INVX1_671 ( .gnd(gnd), .vdd(vdd), .A(data_215__4_), .Y(_863_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf3), .B(_851_), .C(_863_), .Y(_864_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_4_bF_buf2), .C(_864_), .Y(_865_) );
INVX1 INVX1_672 ( .gnd(gnd), .vdd(vdd), .A(_865_), .Y(_129__4_) );
INVX1 INVX1_673 ( .gnd(gnd), .vdd(vdd), .A(data_215__5_), .Y(_866_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_851_), .C(_866_), .Y(_867_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_5_bF_buf1), .C(_867_), .Y(_868_) );
INVX1 INVX1_674 ( .gnd(gnd), .vdd(vdd), .A(_868_), .Y(_129__5_) );
INVX1 INVX1_675 ( .gnd(gnd), .vdd(vdd), .A(data_215__6_), .Y(_869_) );
MUX2X1 MUX2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_15049__bF_buf7), .S(_852_), .Y(_129__6_) );
INVX1 INVX1_676 ( .gnd(gnd), .vdd(vdd), .A(data_215__7_), .Y(_870_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf1), .B(_851_), .C(_870_), .Y(_871_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_7_bF_buf4), .C(_871_), .Y(_872_) );
INVX1 INVX1_677 ( .gnd(gnd), .vdd(vdd), .A(_872_), .Y(_129__7_) );
INVX1 INVX1_678 ( .gnd(gnd), .vdd(vdd), .A(data_215__8_), .Y(_873_) );
MUX2X1 MUX2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_15052__bF_buf6), .S(_852_), .Y(_129__8_) );
INVX1 INVX1_679 ( .gnd(gnd), .vdd(vdd), .A(data_215__9_), .Y(_874_) );
MUX2X1 MUX2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_14913__bF_buf7), .S(_852_), .Y(_129__9_) );
INVX1 INVX1_680 ( .gnd(gnd), .vdd(vdd), .A(data_215__10_), .Y(_875_) );
MUX2X1 MUX2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_15055__bF_buf6), .S(_852_), .Y(_129__10_) );
INVX1 INVX1_681 ( .gnd(gnd), .vdd(vdd), .A(data_215__11_), .Y(_876_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf0), .B(_851_), .C(_876_), .Y(_877_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_11_bF_buf1), .C(_877_), .Y(_878_) );
INVX1 INVX1_682 ( .gnd(gnd), .vdd(vdd), .A(_878_), .Y(_129__11_) );
INVX1 INVX1_683 ( .gnd(gnd), .vdd(vdd), .A(data_215__12_), .Y(_879_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf7), .B(_851_), .C(_879_), .Y(_880_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(IDATA_PROG_data_12_bF_buf1), .C(_880_), .Y(_881_) );
INVX1 INVX1_684 ( .gnd(gnd), .vdd(vdd), .A(_881_), .Y(_129__12_) );
INVX1 INVX1_685 ( .gnd(gnd), .vdd(vdd), .A(data_215__13_), .Y(_882_) );
MUX2X1 MUX2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_882_), .B(_14924__bF_buf5), .S(_852_), .Y(_129__13_) );
INVX1 INVX1_686 ( .gnd(gnd), .vdd(vdd), .A(data_215__14_), .Y(_883_) );
MUX2X1 MUX2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_15060__bF_buf8), .S(_852_), .Y(_129__14_) );
INVX1 INVX1_687 ( .gnd(gnd), .vdd(vdd), .A(data_215__15_), .Y(_884_) );
MUX2X1 MUX2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_15062__bF_buf5), .S(_852_), .Y(_129__15_) );
INVX1 INVX1_688 ( .gnd(gnd), .vdd(vdd), .A(data_214__0_), .Y(_885_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_361__bF_buf4), .Y(_886_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_16204_), .Y(_887_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(_15360_), .Y(_888_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf2), .B(_888_), .C(_592_), .Y(_889_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_751_), .C(_889_), .Y(_890_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_890_), .B(_371_), .Y(_891_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_886_), .Y(_892_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf6), .B(_892_), .Y(_893_) );
MUX2X1 MUX2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_885_), .S(_893__bF_buf3), .Y(_128__0_) );
INVX1 INVX1_689 ( .gnd(gnd), .vdd(vdd), .A(data_214__1_), .Y(_894_) );
MUX2X1 MUX2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_894_), .S(_893__bF_buf2), .Y(_128__1_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(data_214__2_), .B(_893__bF_buf1), .Y(_895_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_893__bF_buf0), .C(_895_), .Y(_128__2_) );
INVX1 INVX1_690 ( .gnd(gnd), .vdd(vdd), .A(data_214__3_), .Y(_896_) );
MUX2X1 MUX2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_896_), .S(_893__bF_buf3), .Y(_128__3_) );
INVX1 INVX1_691 ( .gnd(gnd), .vdd(vdd), .A(data_214__4_), .Y(_897_) );
MUX2X1 MUX2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_897_), .S(_893__bF_buf2), .Y(_128__4_) );
INVX1 INVX1_692 ( .gnd(gnd), .vdd(vdd), .A(data_214__5_), .Y(_898_) );
MUX2X1 MUX2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_898_), .S(_893__bF_buf1), .Y(_128__5_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(data_214__6_), .B(_893__bF_buf0), .Y(_899_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_893__bF_buf3), .C(_899_), .Y(_128__6_) );
INVX1 INVX1_693 ( .gnd(gnd), .vdd(vdd), .A(data_214__7_), .Y(_900_) );
MUX2X1 MUX2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_900_), .S(_893__bF_buf2), .Y(_128__7_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(data_214__8_), .B(_893__bF_buf1), .Y(_901_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_893__bF_buf0), .C(_901_), .Y(_128__8_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(data_214__9_), .B(_893__bF_buf3), .Y(_902_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_893__bF_buf2), .C(_902_), .Y(_128__9_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(data_214__10_), .B(_893__bF_buf1), .Y(_903_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_893__bF_buf0), .C(_903_), .Y(_128__10_) );
INVX1 INVX1_694 ( .gnd(gnd), .vdd(vdd), .A(data_214__11_), .Y(_904_) );
MUX2X1 MUX2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_904_), .S(_893__bF_buf3), .Y(_128__11_) );
INVX1 INVX1_695 ( .gnd(gnd), .vdd(vdd), .A(data_214__12_), .Y(_905_) );
MUX2X1 MUX2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_905_), .S(_893__bF_buf2), .Y(_128__12_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(data_214__13_), .B(_893__bF_buf1), .Y(_906_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_893__bF_buf0), .C(_906_), .Y(_128__13_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(data_214__14_), .B(_893__bF_buf3), .Y(_907_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_893__bF_buf2), .C(_907_), .Y(_128__14_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(data_214__15_), .B(_893__bF_buf1), .Y(_908_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_893__bF_buf0), .C(_908_), .Y(_128__15_) );
INVX1 INVX1_696 ( .gnd(gnd), .vdd(vdd), .A(data_213__0_), .Y(_909_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_14958_), .B(_15006__bF_buf0), .C(IDATA_PROG_write_bF_buf8), .Y(_910_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[0]), .B(_14977__bF_buf2), .C(_15509_), .Y(_911_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_911_), .C(_910_), .Y(_912_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_912_), .C(_886_), .Y(_913_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_913__bF_buf3), .B(_678__bF_buf5), .Y(_914_) );
NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf4), .B(_678__bF_buf4), .C(_913__bF_buf2), .Y(_915_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_914_), .C(_915_), .Y(_127__0_) );
INVX1 INVX1_697 ( .gnd(gnd), .vdd(vdd), .A(data_213__1_), .Y(_916_) );
NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf1), .B(_678__bF_buf3), .C(_913__bF_buf1), .Y(_917_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_914_), .C(_917_), .Y(_127__1_) );
INVX1 INVX1_698 ( .gnd(gnd), .vdd(vdd), .A(data_213__2_), .Y(_918_) );
NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf0), .B(_678__bF_buf2), .C(_913__bF_buf0), .Y(_919_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_914_), .C(_919_), .Y(_127__2_) );
INVX1 INVX1_699 ( .gnd(gnd), .vdd(vdd), .A(data_213__3_), .Y(_920_) );
NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf1), .B(_678__bF_buf1), .C(_913__bF_buf3), .Y(_921_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(_914_), .C(_921_), .Y(_127__3_) );
INVX1 INVX1_700 ( .gnd(gnd), .vdd(vdd), .A(data_213__4_), .Y(_922_) );
NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf1), .B(_678__bF_buf0), .C(_913__bF_buf2), .Y(_923_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_914_), .C(_923_), .Y(_127__4_) );
INVX1 INVX1_701 ( .gnd(gnd), .vdd(vdd), .A(data_213__5_), .Y(_924_) );
NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf0), .B(_678__bF_buf7), .C(_913__bF_buf1), .Y(_925_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_914_), .C(_925_), .Y(_127__5_) );
INVX1 INVX1_702 ( .gnd(gnd), .vdd(vdd), .A(data_213__6_), .Y(_926_) );
NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf0), .B(_678__bF_buf6), .C(_913__bF_buf0), .Y(_927_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_914_), .C(_927_), .Y(_127__6_) );
INVX1 INVX1_703 ( .gnd(gnd), .vdd(vdd), .A(data_213__7_), .Y(_928_) );
NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf3), .B(_678__bF_buf5), .C(_913__bF_buf3), .Y(_929_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_914_), .C(_929_), .Y(_127__7_) );
INVX1 INVX1_704 ( .gnd(gnd), .vdd(vdd), .A(data_213__8_), .Y(_930_) );
NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf3), .B(_678__bF_buf4), .C(_913__bF_buf2), .Y(_931_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_914_), .C(_931_), .Y(_127__8_) );
INVX1 INVX1_705 ( .gnd(gnd), .vdd(vdd), .A(data_213__9_), .Y(_932_) );
NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf0), .B(_678__bF_buf3), .C(_913__bF_buf1), .Y(_933_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_914_), .C(_933_), .Y(_127__9_) );
INVX1 INVX1_706 ( .gnd(gnd), .vdd(vdd), .A(data_213__10_), .Y(_934_) );
NOR3X1 NOR3X1_50 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf3), .B(_678__bF_buf2), .C(_913__bF_buf0), .Y(_935_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_914_), .C(_935_), .Y(_127__10_) );
INVX1 INVX1_707 ( .gnd(gnd), .vdd(vdd), .A(data_213__11_), .Y(_936_) );
NOR3X1 NOR3X1_51 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf0), .B(_678__bF_buf1), .C(_913__bF_buf3), .Y(_937_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_914_), .C(_937_), .Y(_127__11_) );
INVX1 INVX1_708 ( .gnd(gnd), .vdd(vdd), .A(data_213__12_), .Y(_938_) );
NOR3X1 NOR3X1_52 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf0), .B(_678__bF_buf0), .C(_913__bF_buf2), .Y(_939_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_914_), .C(_939_), .Y(_127__12_) );
INVX1 INVX1_709 ( .gnd(gnd), .vdd(vdd), .A(data_213__13_), .Y(_940_) );
NOR3X1 NOR3X1_53 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf4), .B(_678__bF_buf7), .C(_913__bF_buf1), .Y(_941_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_914_), .C(_941_), .Y(_127__13_) );
INVX1 INVX1_710 ( .gnd(gnd), .vdd(vdd), .A(data_213__14_), .Y(_942_) );
NOR3X1 NOR3X1_54 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf4), .B(_678__bF_buf6), .C(_913__bF_buf0), .Y(_943_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_914_), .C(_943_), .Y(_127__14_) );
INVX1 INVX1_711 ( .gnd(gnd), .vdd(vdd), .A(data_213__15_), .Y(_944_) );
NOR3X1 NOR3X1_55 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf0), .B(_678__bF_buf5), .C(_913__bF_buf3), .Y(_945_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_914_), .C(_945_), .Y(_127__15_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_15508_), .B(_15006__bF_buf4), .C(_828_), .Y(_946_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_361__bF_buf3), .B(_946_), .Y(_947_) );
NOR3X1 NOR3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_15841_), .C(_678__bF_buf4), .Y(_948_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(data_212__0_), .B(_948__bF_buf4), .Y(_949_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_948__bF_buf3), .C(_949_), .Y(_126__0_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(data_212__1_), .B(_948__bF_buf2), .Y(_950_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_948__bF_buf1), .C(_950_), .Y(_126__1_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(data_212__2_), .B(_948__bF_buf0), .Y(_951_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_948__bF_buf4), .C(_951_), .Y(_126__2_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(data_212__3_), .B(_948__bF_buf3), .Y(_952_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_948__bF_buf2), .C(_952_), .Y(_126__3_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(data_212__4_), .B(_948__bF_buf1), .Y(_953_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_948__bF_buf0), .C(_953_), .Y(_126__4_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(data_212__5_), .B(_948__bF_buf4), .Y(_954_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_948__bF_buf3), .C(_954_), .Y(_126__5_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(data_212__6_), .B(_948__bF_buf2), .Y(_955_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_948__bF_buf1), .C(_955_), .Y(_126__6_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(data_212__7_), .B(_948__bF_buf0), .Y(_956_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_948__bF_buf4), .C(_956_), .Y(_126__7_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(data_212__8_), .B(_948__bF_buf3), .Y(_957_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_948__bF_buf2), .C(_957_), .Y(_126__8_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(data_212__9_), .B(_948__bF_buf1), .Y(_958_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_948__bF_buf0), .C(_958_), .Y(_126__9_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(data_212__10_), .B(_948__bF_buf4), .Y(_959_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_948__bF_buf3), .C(_959_), .Y(_126__10_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(data_212__11_), .B(_948__bF_buf2), .Y(_960_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_948__bF_buf1), .C(_960_), .Y(_126__11_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(data_212__12_), .B(_948__bF_buf0), .Y(_961_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_948__bF_buf4), .C(_961_), .Y(_126__12_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(data_212__13_), .B(_948__bF_buf3), .Y(_962_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_948__bF_buf2), .C(_962_), .Y(_126__13_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(data_212__14_), .B(_948__bF_buf1), .Y(_963_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_948__bF_buf0), .C(_963_), .Y(_126__14_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(data_212__15_), .B(_948__bF_buf4), .Y(_964_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_948__bF_buf3), .C(_964_), .Y(_126__15_) );
INVX1 INVX1_712 ( .gnd(gnd), .vdd(vdd), .A(data_211__0_), .Y(_965_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf3), .B(_15034_), .C(IDATA_PROG_write_bF_buf7), .Y(_966_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf3), .B(_15025__bF_buf2), .C(_15006__bF_buf3), .D(_15571_), .Y(_967_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_967_), .Y(_968_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_15006__bF_buf2), .B(_15581_), .C(_968_), .Y(_969_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_15025__bF_buf1), .C(_15026_), .Y(_970_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_15023_), .Y(_971_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_15183__bF_buf6), .Y(_972_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_969_), .Y(_973_) );
NOR3X1 NOR3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_973_), .C(_678__bF_buf3), .Y(_974_) );
MUX2X1 MUX2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_965_), .S(_974__bF_buf3), .Y(_125__0_) );
INVX1 INVX1_713 ( .gnd(gnd), .vdd(vdd), .A(data_211__1_), .Y(_975_) );
MUX2X1 MUX2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_975_), .S(_974__bF_buf2), .Y(_125__1_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(data_211__2_), .B(_974__bF_buf1), .Y(_976_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_974__bF_buf0), .C(_976_), .Y(_125__2_) );
INVX1 INVX1_714 ( .gnd(gnd), .vdd(vdd), .A(data_211__3_), .Y(_977_) );
MUX2X1 MUX2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_977_), .S(_974__bF_buf3), .Y(_125__3_) );
INVX1 INVX1_715 ( .gnd(gnd), .vdd(vdd), .A(data_211__4_), .Y(_978_) );
MUX2X1 MUX2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_978_), .S(_974__bF_buf2), .Y(_125__4_) );
INVX1 INVX1_716 ( .gnd(gnd), .vdd(vdd), .A(data_211__5_), .Y(_979_) );
MUX2X1 MUX2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_979_), .S(_974__bF_buf1), .Y(_125__5_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(data_211__6_), .B(_974__bF_buf0), .Y(_980_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_974__bF_buf3), .C(_980_), .Y(_125__6_) );
INVX1 INVX1_717 ( .gnd(gnd), .vdd(vdd), .A(data_211__7_), .Y(_981_) );
MUX2X1 MUX2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_981_), .S(_974__bF_buf2), .Y(_125__7_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(data_211__8_), .B(_974__bF_buf1), .Y(_982_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_974__bF_buf0), .C(_982_), .Y(_125__8_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(data_211__9_), .B(_974__bF_buf3), .Y(_983_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_974__bF_buf2), .C(_983_), .Y(_125__9_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(data_211__10_), .B(_974__bF_buf1), .Y(_984_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf3), .B(_974__bF_buf0), .C(_984_), .Y(_125__10_) );
INVX1 INVX1_718 ( .gnd(gnd), .vdd(vdd), .A(data_211__11_), .Y(_985_) );
MUX2X1 MUX2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_985_), .S(_974__bF_buf3), .Y(_125__11_) );
INVX1 INVX1_719 ( .gnd(gnd), .vdd(vdd), .A(data_211__12_), .Y(_986_) );
MUX2X1 MUX2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_986_), .S(_974__bF_buf2), .Y(_125__12_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(data_211__13_), .B(_974__bF_buf1), .Y(_987_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_974__bF_buf0), .C(_987_), .Y(_125__13_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(data_211__14_), .B(_974__bF_buf3), .Y(_988_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf5), .B(_974__bF_buf2), .C(_988_), .Y(_125__14_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(data_211__15_), .B(_974__bF_buf1), .Y(_989_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf2), .B(_974__bF_buf0), .C(_989_), .Y(_125__15_) );
INVX1 INVX1_720 ( .gnd(gnd), .vdd(vdd), .A(data_210__0_), .Y(_990_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_967_), .Y(_991_) );
INVX1 INVX1_721 ( .gnd(gnd), .vdd(vdd), .A(_966_), .Y(_992_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_15006__bF_buf1), .C(_992_), .Y(_993_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_993_), .Y(_994_) );
NOR3X1 NOR3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_678__bF_buf2), .B(_947_), .C(_994_), .Y(_995_) );
MUX2X1 MUX2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_990_), .S(_995__bF_buf3), .Y(_124__0_) );
INVX1 INVX1_722 ( .gnd(gnd), .vdd(vdd), .A(data_210__1_), .Y(_996_) );
MUX2X1 MUX2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_996_), .S(_995__bF_buf2), .Y(_124__1_) );
INVX1 INVX1_723 ( .gnd(gnd), .vdd(vdd), .A(data_210__2_), .Y(_997_) );
NOR3X1 NOR3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_676_), .C(_543_), .Y(_998_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_361__bF_buf2), .Y(_999_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_998_), .Y(_1000_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_994_), .C(_997_), .Y(_1001_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_995__bF_buf1), .Y(_1002_) );
AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1002_), .Y(_124__2_) );
INVX1 INVX1_724 ( .gnd(gnd), .vdd(vdd), .A(data_210__3_), .Y(_1003_) );
MUX2X1 MUX2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_1003_), .S(_995__bF_buf0), .Y(_124__3_) );
INVX1 INVX1_725 ( .gnd(gnd), .vdd(vdd), .A(data_210__4_), .Y(_1004_) );
MUX2X1 MUX2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_1004_), .S(_995__bF_buf3), .Y(_124__4_) );
INVX1 INVX1_726 ( .gnd(gnd), .vdd(vdd), .A(data_210__5_), .Y(_1005_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_994_), .C(_1005_), .Y(_1006_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_995__bF_buf2), .Y(_1007_) );
AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_1007_), .Y(_124__5_) );
INVX1 INVX1_727 ( .gnd(gnd), .vdd(vdd), .A(data_210__6_), .Y(_1008_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_994_), .C(_1008_), .Y(_1009_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_995__bF_buf1), .Y(_1010_) );
AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .B(_1010_), .Y(_124__6_) );
INVX1 INVX1_728 ( .gnd(gnd), .vdd(vdd), .A(data_210__7_), .Y(_1011_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_994_), .C(_1011_), .Y(_1012_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_995__bF_buf0), .Y(_1013_) );
AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_1012_), .B(_1013_), .Y(_124__7_) );
INVX1 INVX1_729 ( .gnd(gnd), .vdd(vdd), .A(data_210__8_), .Y(_1014_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_994_), .C(_1014_), .Y(_1015_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_995__bF_buf3), .Y(_1016_) );
AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .B(_1016_), .Y(_124__8_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_995__bF_buf2), .Y(_1017_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(data_210__9_), .B(_995__bF_buf1), .C(_1017_), .Y(_1018_) );
INVX1 INVX1_730 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .Y(_124__9_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_995__bF_buf0), .Y(_1019_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(data_210__10_), .B(_995__bF_buf3), .C(_1019_), .Y(_1020_) );
INVX1 INVX1_731 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .Y(_124__10_) );
INVX1 INVX1_732 ( .gnd(gnd), .vdd(vdd), .A(data_210__11_), .Y(_1021_) );
MUX2X1 MUX2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_1021_), .S(_995__bF_buf2), .Y(_124__11_) );
INVX1 INVX1_733 ( .gnd(gnd), .vdd(vdd), .A(data_210__12_), .Y(_1022_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_994_), .C(_1022_), .Y(_1023_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_995__bF_buf1), .Y(_1024_) );
AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1024_), .Y(_124__12_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_995__bF_buf0), .Y(_1025_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(data_210__13_), .B(_995__bF_buf3), .C(_1025_), .Y(_1026_) );
INVX1 INVX1_734 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .Y(_124__13_) );
INVX1 INVX1_735 ( .gnd(gnd), .vdd(vdd), .A(data_210__14_), .Y(_1027_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_994_), .C(_1027_), .Y(_1028_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_995__bF_buf2), .Y(_1029_) );
AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1029_), .Y(_124__14_) );
INVX1 INVX1_736 ( .gnd(gnd), .vdd(vdd), .A(data_210__15_), .Y(_1030_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_994_), .C(_1030_), .Y(_1031_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_995__bF_buf1), .Y(_1032_) );
AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .B(_1032_), .Y(_124__15_) );
INVX1 INVX1_737 ( .gnd(gnd), .vdd(vdd), .A(data_209__0_), .Y(_1033_) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(_972_), .Y(_1034_) );
INVX1 INVX1_738 ( .gnd(gnd), .vdd(vdd), .A(_993_), .Y(_1035_) );
INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf0), .Y(_1036_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf1), .B(_1036__bF_buf3), .C(_15684_), .D(_592_), .Y(_1037_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1037_), .C(_1034_), .Y(_1038_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1038_), .C(_1033_), .Y(_1039_) );
NOR3X1 NOR3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_1038_), .C(_678__bF_buf1), .Y(_1040_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_1040__bF_buf3), .Y(_1041_) );
AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1041_), .Y(_122__0_) );
INVX1 INVX1_739 ( .gnd(gnd), .vdd(vdd), .A(data_209__1_), .Y(_1042_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1038_), .C(_1042_), .Y(_1043_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_1040__bF_buf2), .Y(_1044_) );
AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .B(_1044_), .Y(_122__1_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(data_209__2_), .B(_1040__bF_buf1), .Y(_1045_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_1040__bF_buf0), .C(_1045_), .Y(_122__2_) );
INVX1 INVX1_740 ( .gnd(gnd), .vdd(vdd), .A(data_209__3_), .Y(_1046_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1038_), .C(_1046_), .Y(_1047_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_1040__bF_buf3), .Y(_1048_) );
AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .B(_1048_), .Y(_122__3_) );
INVX1 INVX1_741 ( .gnd(gnd), .vdd(vdd), .A(data_209__4_), .Y(_1049_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1038_), .C(_1049_), .Y(_1050_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_1040__bF_buf2), .Y(_1051_) );
AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1051_), .Y(_122__4_) );
INVX1 INVX1_742 ( .gnd(gnd), .vdd(vdd), .A(data_209__5_), .Y(_1052_) );
MUX2X1 MUX2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_1052_), .S(_1040__bF_buf1), .Y(_122__5_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(data_209__6_), .B(_1040__bF_buf0), .Y(_1053_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_1040__bF_buf3), .C(_1053_), .Y(_122__6_) );
INVX1 INVX1_743 ( .gnd(gnd), .vdd(vdd), .A(data_209__7_), .Y(_1054_) );
MUX2X1 MUX2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_1054_), .S(_1040__bF_buf2), .Y(_122__7_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(data_209__8_), .B(_1040__bF_buf1), .Y(_1055_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_1040__bF_buf0), .C(_1055_), .Y(_122__8_) );
INVX1 INVX1_744 ( .gnd(gnd), .vdd(vdd), .A(data_209__9_), .Y(_1056_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1038_), .C(_1056_), .Y(_1057_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_1040__bF_buf3), .Y(_1058_) );
AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1058_), .Y(_122__9_) );
INVX1 INVX1_745 ( .gnd(gnd), .vdd(vdd), .A(data_209__10_), .Y(_1059_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1038_), .C(_1059_), .Y(_1060_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_1040__bF_buf2), .Y(_1061_) );
AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_1061_), .Y(_122__10_) );
INVX1 INVX1_746 ( .gnd(gnd), .vdd(vdd), .A(data_209__11_), .Y(_1062_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1038_), .C(_1062_), .Y(_1063_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_1040__bF_buf1), .Y(_1064_) );
AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1064_), .Y(_122__11_) );
INVX1 INVX1_747 ( .gnd(gnd), .vdd(vdd), .A(data_209__12_), .Y(_1065_) );
MUX2X1 MUX2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_1065_), .S(_1040__bF_buf0), .Y(_122__12_) );
INVX1 INVX1_748 ( .gnd(gnd), .vdd(vdd), .A(data_209__13_), .Y(_1066_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1038_), .C(_1066_), .Y(_1067_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_1040__bF_buf3), .Y(_1068_) );
AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .B(_1068_), .Y(_122__13_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(data_209__14_), .B(_1040__bF_buf2), .Y(_1069_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_1040__bF_buf1), .C(_1069_), .Y(_122__14_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(data_209__15_), .B(_1040__bF_buf0), .Y(_1070_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_1040__bF_buf3), .C(_1070_), .Y(_122__15_) );
INVX1 INVX1_749 ( .gnd(gnd), .vdd(vdd), .A(data_208__0_), .Y(_1071_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_14883_), .B(_15064_), .C(_15026_), .Y(_1072_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf2), .B(_14975_), .C(_592_), .Y(_1073_) );
INVX1 INVX1_750 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .Y(_1074_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1074_), .Y(_1075_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_15023_), .B(_15074__bF_buf3), .Y(_1076_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1076_), .Y(_1077_) );
INVX1 INVX1_751 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .Y(_1078_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_999_), .B(_1078_), .C(_998_), .Y(_1079_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf3), .B(_14882__bF_buf11), .C(_1071_), .Y(_1080_) );
NOR3X1 NOR3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_1077_), .C(_678__bF_buf0), .Y(_1081_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(IDATA_PROG_write_bF_buf6), .C(_1081_), .Y(_1082_) );
AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1082_), .Y(_121__0_) );
INVX1 INVX1_752 ( .gnd(gnd), .vdd(vdd), .A(data_208__1_), .Y(_1083_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf2), .B(_14882__bF_buf10), .C(_1083_), .Y(_1084_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf5), .B(_14894__bF_buf5), .C(_1081_), .Y(_1085_) );
AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1085_), .Y(_121__1_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_1081_), .Y(_1086_) );
INVX1 INVX1_753 ( .gnd(gnd), .vdd(vdd), .A(data_208__2_), .Y(_1087_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf1), .B(_14882__bF_buf9), .C(_1087_), .Y(_1088_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf3), .B(_1086_), .C(_1088_), .Y(_1089_) );
INVX1 INVX1_754 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .Y(_121__2_) );
INVX1 INVX1_755 ( .gnd(gnd), .vdd(vdd), .A(data_208__3_), .Y(_1090_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf0), .B(_14882__bF_buf8), .C(_1090_), .Y(_1091_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf3), .B(_14899__bF_buf5), .C(_1081_), .Y(_1092_) );
AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .B(_1092_), .Y(_121__3_) );
INVX1 INVX1_756 ( .gnd(gnd), .vdd(vdd), .A(data_208__4_), .Y(_1093_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf3), .B(_14882__bF_buf7), .C(_1093_), .Y(_1094_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_14902__bF_buf2), .C(_1081_), .Y(_1095_) );
AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1095_), .Y(_121__4_) );
INVX1 INVX1_757 ( .gnd(gnd), .vdd(vdd), .A(data_208__5_), .Y(_1096_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf2), .B(_14882__bF_buf6), .C(_1096_), .Y(_1097_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_14903__bF_buf3), .C(_1081_), .Y(_1098_) );
AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .B(_1098_), .Y(_121__5_) );
INVX1 INVX1_758 ( .gnd(gnd), .vdd(vdd), .A(data_208__6_), .Y(_1099_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf1), .B(_14882__bF_buf5), .C(_1099_), .Y(_1100_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf4), .B(_1086_), .C(_1100_), .Y(_1101_) );
INVX1 INVX1_759 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_121__6_) );
INVX1 INVX1_760 ( .gnd(gnd), .vdd(vdd), .A(data_208__7_), .Y(_1102_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf0), .B(_14882__bF_buf4), .C(_1102_), .Y(_1103_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf0), .B(_14908__bF_buf2), .C(_1081_), .Y(_1104_) );
AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1104_), .Y(_121__7_) );
INVX1 INVX1_761 ( .gnd(gnd), .vdd(vdd), .A(data_208__8_), .Y(_1105_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf3), .B(_14882__bF_buf3), .C(_1105_), .Y(_1106_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf2), .B(_1086_), .C(_1106_), .Y(_1107_) );
INVX1 INVX1_762 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .Y(_121__8_) );
INVX1 INVX1_763 ( .gnd(gnd), .vdd(vdd), .A(data_208__9_), .Y(_1108_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf2), .B(_14882__bF_buf2), .C(_1108_), .Y(_1109_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf4), .B(_1086_), .C(_1109_), .Y(_1110_) );
INVX1 INVX1_764 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .Y(_121__9_) );
INVX1 INVX1_765 ( .gnd(gnd), .vdd(vdd), .A(data_208__10_), .Y(_1111_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf1), .B(_14882__bF_buf1), .C(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf2), .B(_1086_), .C(_1112_), .Y(_1113_) );
INVX1 INVX1_766 ( .gnd(gnd), .vdd(vdd), .A(_1113_), .Y(_121__10_) );
INVX1 INVX1_767 ( .gnd(gnd), .vdd(vdd), .A(data_208__11_), .Y(_1114_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf0), .B(_14882__bF_buf0), .C(_1114_), .Y(_1115_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .B(_14918__bF_buf3), .C(_1081_), .Y(_1116_) );
AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1116_), .Y(_121__11_) );
INVX1 INVX1_768 ( .gnd(gnd), .vdd(vdd), .A(data_208__12_), .Y(_1117_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf3), .B(_14882__bF_buf15_bF_buf0), .C(_1117_), .Y(_1118_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_14920__bF_buf3), .C(_1081_), .Y(_1119_) );
AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1119_), .Y(_121__12_) );
INVX1 INVX1_769 ( .gnd(gnd), .vdd(vdd), .A(data_208__13_), .Y(_1120_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf2), .B(_14882__bF_buf14_bF_buf0), .C(_1120_), .Y(_1121_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf3), .B(_1086_), .C(_1121_), .Y(_1122_) );
INVX1 INVX1_770 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .Y(_121__13_) );
INVX1 INVX1_771 ( .gnd(gnd), .vdd(vdd), .A(data_208__14_), .Y(_1123_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf1), .B(_14882__bF_buf13_bF_buf0), .C(_1123_), .Y(_1124_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf3), .B(_1086_), .C(_1124_), .Y(_1125_) );
INVX1 INVX1_772 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .Y(_121__14_) );
INVX1 INVX1_773 ( .gnd(gnd), .vdd(vdd), .A(data_208__15_), .Y(_1126_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_1079__bF_buf0), .B(_14882__bF_buf12), .C(_1126_), .Y(_1127_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf5), .B(_1086_), .C(_1127_), .Y(_1128_) );
INVX1 INVX1_774 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .Y(_121__15_) );
INVX1 INVX1_775 ( .gnd(gnd), .vdd(vdd), .A(data_207__0_), .Y(_1129_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_15025__bF_buf4), .C(_1073_), .Y(_1130_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_972_), .Y(_1131_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1131_), .Y(_1132_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .Y(_1133_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_1133_), .Y(_1134_) );
MUX2X1 MUX2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_14932__bF_buf6), .S(_1134_), .Y(_120__0_) );
INVX1 INVX1_776 ( .gnd(gnd), .vdd(vdd), .A(data_207__1_), .Y(_1135_) );
MUX2X1 MUX2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_14894__bF_buf4), .S(_1134_), .Y(_120__1_) );
INVX1 INVX1_777 ( .gnd(gnd), .vdd(vdd), .A(data_207__2_), .Y(_1136_) );
MUX2X1 MUX2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_14897__bF_buf0), .S(_1134_), .Y(_120__2_) );
INVX1 INVX1_778 ( .gnd(gnd), .vdd(vdd), .A(data_207__3_), .Y(_1137_) );
MUX2X1 MUX2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_14899__bF_buf4), .S(_1134_), .Y(_120__3_) );
INVX1 INVX1_779 ( .gnd(gnd), .vdd(vdd), .A(data_207__4_), .Y(_1138_) );
MUX2X1 MUX2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_14902__bF_buf1), .S(_1134_), .Y(_120__4_) );
INVX1 INVX1_780 ( .gnd(gnd), .vdd(vdd), .A(data_207__5_), .Y(_1139_) );
MUX2X1 MUX2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_14903__bF_buf2), .S(_1134_), .Y(_120__5_) );
INVX1 INVX1_781 ( .gnd(gnd), .vdd(vdd), .A(data_207__6_), .Y(_1140_) );
MUX2X1 MUX2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_15049__bF_buf1), .S(_1134_), .Y(_120__6_) );
INVX1 INVX1_782 ( .gnd(gnd), .vdd(vdd), .A(data_207__7_), .Y(_1141_) );
MUX2X1 MUX2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_14908__bF_buf1), .S(_1134_), .Y(_120__7_) );
INVX1 INVX1_783 ( .gnd(gnd), .vdd(vdd), .A(data_207__8_), .Y(_1142_) );
MUX2X1 MUX2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_15052__bF_buf0), .S(_1134_), .Y(_120__8_) );
INVX1 INVX1_784 ( .gnd(gnd), .vdd(vdd), .A(data_207__9_), .Y(_1143_) );
MUX2X1 MUX2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_14913__bF_buf1), .S(_1134_), .Y(_120__9_) );
INVX1 INVX1_785 ( .gnd(gnd), .vdd(vdd), .A(data_207__10_), .Y(_1144_) );
MUX2X1 MUX2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_15055__bF_buf0), .S(_1134_), .Y(_120__10_) );
INVX1 INVX1_786 ( .gnd(gnd), .vdd(vdd), .A(data_207__11_), .Y(_1145_) );
MUX2X1 MUX2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(_14918__bF_buf2), .S(_1134_), .Y(_120__11_) );
INVX1 INVX1_787 ( .gnd(gnd), .vdd(vdd), .A(data_207__12_), .Y(_1146_) );
MUX2X1 MUX2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .B(_14920__bF_buf2), .S(_1134_), .Y(_120__12_) );
INVX1 INVX1_788 ( .gnd(gnd), .vdd(vdd), .A(data_207__13_), .Y(_1147_) );
MUX2X1 MUX2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_14924__bF_buf13), .S(_1134_), .Y(_120__13_) );
INVX1 INVX1_789 ( .gnd(gnd), .vdd(vdd), .A(data_207__14_), .Y(_1148_) );
MUX2X1 MUX2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_15060__bF_buf2), .S(_1134_), .Y(_120__14_) );
INVX1 INVX1_790 ( .gnd(gnd), .vdd(vdd), .A(data_207__15_), .Y(_1149_) );
MUX2X1 MUX2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_15062__bF_buf13), .S(_1134_), .Y(_120__15_) );
INVX1 INVX1_791 ( .gnd(gnd), .vdd(vdd), .A(data_206__0_), .Y(_1150_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15025__bF_buf3), .C(_1150_), .Y(_1151_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf2), .B(_15788__bF_buf6), .Y(_1152_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_1152_), .Y(_1153_) );
AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1151_), .Y(_119__0_) );
INVX1 INVX1_792 ( .gnd(gnd), .vdd(vdd), .A(data_206__1_), .Y(_1154_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15025__bF_buf1), .C(_1154_), .Y(_1155_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_1152_), .Y(_1156_) );
AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .B(_1155_), .Y(_119__1_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(data_206__2_), .B(_1152_), .Y(_1157_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_1152_), .C(_1157_), .Y(_119__2_) );
INVX1 INVX1_793 ( .gnd(gnd), .vdd(vdd), .A(data_206__3_), .Y(_1158_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15025__bF_buf0), .C(_1158_), .Y(_1159_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_1036__bF_buf2), .C(_15793__bF_buf4), .Y(_1160_) );
AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1160_), .Y(_119__3_) );
INVX1 INVX1_794 ( .gnd(gnd), .vdd(vdd), .A(data_206__4_), .Y(_1161_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1036__bF_buf1), .B(_15793__bF_buf3), .Y(_1162_) );
MUX2X1 MUX2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(_14902__bF_buf0), .S(_1162_), .Y(_119__4_) );
INVX1 INVX1_795 ( .gnd(gnd), .vdd(vdd), .A(data_206__5_), .Y(_1163_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15025__bF_buf4), .C(_1163_), .Y(_1164_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_1152_), .Y(_1165_) );
AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1164_), .Y(_119__5_) );
INVX1 INVX1_796 ( .gnd(gnd), .vdd(vdd), .A(data_206__6_), .Y(_1166_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15025__bF_buf3), .C(_1166_), .Y(_1167_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf0), .B(_1036__bF_buf0), .C(_15793__bF_buf2), .Y(_1168_) );
AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_1168_), .Y(_119__6_) );
INVX1 INVX1_797 ( .gnd(gnd), .vdd(vdd), .A(data_206__7_), .Y(_1169_) );
MUX2X1 MUX2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_14908__bF_buf0), .S(_1162_), .Y(_119__7_) );
INVX1 INVX1_798 ( .gnd(gnd), .vdd(vdd), .A(data_206__8_), .Y(_1170_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15025__bF_buf2), .C(_1170_), .Y(_1171_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_1036__bF_buf3), .C(_15793__bF_buf1), .Y(_1172_) );
AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1172_), .Y(_119__8_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(data_206__9_), .B(_1152_), .Y(_1173_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_1152_), .C(_1173_), .Y(_119__9_) );
INVX1 INVX1_799 ( .gnd(gnd), .vdd(vdd), .A(data_206__10_), .Y(_1174_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15025__bF_buf1), .C(_1174_), .Y(_1175_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_1152_), .Y(_1176_) );
AND2X2 AND2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1175_), .Y(_119__10_) );
INVX1 INVX1_800 ( .gnd(gnd), .vdd(vdd), .A(data_206__11_), .Y(_1177_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15025__bF_buf0), .C(_1177_), .Y(_1178_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_1152_), .Y(_1179_) );
AND2X2 AND2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_1178_), .Y(_119__11_) );
INVX1 INVX1_801 ( .gnd(gnd), .vdd(vdd), .A(data_206__12_), .Y(_1180_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15025__bF_buf4), .C(_1180_), .Y(_1181_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_1152_), .Y(_1182_) );
AND2X2 AND2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1181_), .Y(_119__12_) );
INVX1 INVX1_802 ( .gnd(gnd), .vdd(vdd), .A(data_206__13_), .Y(_1183_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15025__bF_buf3), .C(_1183_), .Y(_1184_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_1036__bF_buf2), .C(_15793__bF_buf0), .Y(_1185_) );
AND2X2 AND2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1185_), .Y(_119__13_) );
INVX1 INVX1_803 ( .gnd(gnd), .vdd(vdd), .A(data_206__14_), .Y(_1186_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15025__bF_buf2), .C(_1186_), .Y(_1187_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_1036__bF_buf1), .C(_15793__bF_buf5), .Y(_1188_) );
AND2X2 AND2X2_378 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1188_), .Y(_119__14_) );
INVX1 INVX1_804 ( .gnd(gnd), .vdd(vdd), .A(data_206__15_), .Y(_1189_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15025__bF_buf1), .C(_1189_), .Y(_1190_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_1036__bF_buf0), .C(_15793__bF_buf4), .Y(_1191_) );
AND2X2 AND2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_1191_), .Y(_119__15_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1081_), .Y(_1192_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1036__bF_buf3), .B(_15078_), .C(_966_), .Y(_1193_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1193_), .C(_1034_), .Y(_1194_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1194_), .B(_1000__bF_buf3), .Y(_1195_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__0_), .Y(_1196_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1077_), .C(_1132_), .Y(_1197_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1194_), .Y(_1198_) );
NOR3X1 NOR3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_0_bF_buf3), .C(_1198_), .Y(_1199_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_1199_), .Y(_118__0_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__1_), .Y(_1200_) );
NOR3X1 NOR3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_1_bF_buf0), .C(_1198_), .Y(_1201_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_1201_), .Y(_118__1_) );
INVX1 INVX1_805 ( .gnd(gnd), .vdd(vdd), .A(data_205__2_), .Y(_1202_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .Y(_1203_) );
MUX2X1 MUX2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(_14897__bF_buf13), .S(_1203_), .Y(_118__2_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__3_), .Y(_1204_) );
NOR3X1 NOR3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_3_bF_buf0), .C(_1198_), .Y(_1205_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1205_), .Y(_118__3_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__4_), .Y(_1206_) );
NOR3X1 NOR3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_4_bF_buf0), .C(_1198_), .Y(_1207_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_1207_), .Y(_118__4_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__5_), .Y(_1208_) );
NOR3X1 NOR3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_5_bF_buf4), .C(_1198_), .Y(_1209_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_1209_), .Y(_118__5_) );
INVX1 INVX1_806 ( .gnd(gnd), .vdd(vdd), .A(data_205__6_), .Y(_1210_) );
MUX2X1 MUX2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(_15049__bF_buf14), .S(_1203_), .Y(_118__6_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__7_), .Y(_1211_) );
NOR3X1 NOR3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_7_bF_buf2), .C(_1198_), .Y(_1212_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1212_), .Y(_118__7_) );
INVX1 INVX1_807 ( .gnd(gnd), .vdd(vdd), .A(data_205__8_), .Y(_1213_) );
MUX2X1 MUX2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .B(_15052__bF_buf12), .S(_1203_), .Y(_118__8_) );
INVX1 INVX1_808 ( .gnd(gnd), .vdd(vdd), .A(data_205__9_), .Y(_1214_) );
MUX2X1 MUX2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_14913__bF_buf14), .S(_1203_), .Y(_118__9_) );
INVX1 INVX1_809 ( .gnd(gnd), .vdd(vdd), .A(data_205__10_), .Y(_1215_) );
MUX2X1 MUX2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_15055__bF_buf12), .S(_1203_), .Y(_118__10_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__11_), .Y(_1216_) );
NOR3X1 NOR3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_11_bF_buf4), .C(_1198_), .Y(_1217_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1216_), .B(_1217_), .Y(_118__11_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1192_), .C(data_205__12_), .Y(_1218_) );
NOR3X1 NOR3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(IDATA_PROG_data_12_bF_buf4), .C(_1198_), .Y(_1219_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1218_), .B(_1219_), .Y(_118__12_) );
INVX1 INVX1_810 ( .gnd(gnd), .vdd(vdd), .A(data_205__13_), .Y(_1220_) );
MUX2X1 MUX2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_14924__bF_buf11), .S(_1203_), .Y(_118__13_) );
INVX1 INVX1_811 ( .gnd(gnd), .vdd(vdd), .A(data_205__14_), .Y(_1221_) );
MUX2X1 MUX2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_15060__bF_buf0), .S(_1203_), .Y(_118__14_) );
INVX1 INVX1_812 ( .gnd(gnd), .vdd(vdd), .A(data_205__15_), .Y(_1222_) );
MUX2X1 MUX2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_15062__bF_buf11), .S(_1203_), .Y(_118__15_) );
INVX1 INVX1_813 ( .gnd(gnd), .vdd(vdd), .A(data_204__0_), .Y(_1223_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15025__bF_buf0), .C(_1073_), .Y(_1224_) );
NOR3X1 NOR3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1224_), .C(_1081_), .Y(_1225_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_15025__bF_buf4), .C(_1225__bF_buf6), .Y(_1226_) );
INVX1 INVX1_814 ( .gnd(gnd), .vdd(vdd), .A(_970_), .Y(_1227_) );
NOR3X1 NOR3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_15074__bF_buf2), .C(_678__bF_buf7), .Y(_1228_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1227_), .B(_15082_), .C(_1228_), .Y(_1229_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf4), .C(_1223_), .Y(_1230_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_15035_), .B(_1036__bF_buf2), .C(_1229__bF_buf3), .Y(_1231_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_1225__bF_buf5), .C(_1231_), .Y(_1232_) );
AND2X2 AND2X2_380 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1232_), .Y(_117__0_) );
INVX1 INVX1_815 ( .gnd(gnd), .vdd(vdd), .A(data_204__1_), .Y(_1233_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1225__bF_buf4), .B(_1231_), .Y(_1234_) );
MUX2X1 MUX2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_14894__bF_buf2), .S(_1234_), .Y(_117__1_) );
INVX1 INVX1_816 ( .gnd(gnd), .vdd(vdd), .A(data_204__2_), .Y(_1235_) );
MUX2X1 MUX2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1235_), .B(_14897__bF_buf12), .S(_1234_), .Y(_117__2_) );
INVX1 INVX1_817 ( .gnd(gnd), .vdd(vdd), .A(data_204__3_), .Y(_1236_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf2), .C(_1236_), .Y(_1237_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_1225__bF_buf3), .C(_1231_), .Y(_1238_) );
AND2X2 AND2X2_381 ( .gnd(gnd), .vdd(vdd), .A(_1237_), .B(_1238_), .Y(_117__3_) );
INVX1 INVX1_818 ( .gnd(gnd), .vdd(vdd), .A(data_204__4_), .Y(_1239_) );
MUX2X1 MUX2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_14902__bF_buf13), .S(_1234_), .Y(_117__4_) );
INVX1 INVX1_819 ( .gnd(gnd), .vdd(vdd), .A(data_204__5_), .Y(_1240_) );
MUX2X1 MUX2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_14903__bF_buf0), .S(_1234_), .Y(_117__5_) );
INVX1 INVX1_820 ( .gnd(gnd), .vdd(vdd), .A(data_204__6_), .Y(_1241_) );
MUX2X1 MUX2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_15049__bF_buf13), .S(_1234_), .Y(_117__6_) );
INVX1 INVX1_821 ( .gnd(gnd), .vdd(vdd), .A(data_204__7_), .Y(_1242_) );
MUX2X1 MUX2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .B(_14908__bF_buf13), .S(_1234_), .Y(_117__7_) );
INVX1 INVX1_822 ( .gnd(gnd), .vdd(vdd), .A(data_204__8_), .Y(_1243_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf1), .C(_1243_), .Y(_1244_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1229__bF_buf0), .B(_1226_), .Y(_1245_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_1245_), .Y(_1246_) );
AND2X2 AND2X2_382 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1244_), .Y(_117__8_) );
INVX1 INVX1_823 ( .gnd(gnd), .vdd(vdd), .A(data_204__9_), .Y(_1247_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf4), .C(_1247_), .Y(_1248_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_1245_), .Y(_1249_) );
AND2X2 AND2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .B(_1248_), .Y(_117__9_) );
INVX1 INVX1_824 ( .gnd(gnd), .vdd(vdd), .A(data_204__10_), .Y(_1250_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf3), .C(_1250_), .Y(_1251_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_1245_), .Y(_1252_) );
AND2X2 AND2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_1252_), .B(_1251_), .Y(_117__10_) );
INVX1 INVX1_825 ( .gnd(gnd), .vdd(vdd), .A(data_204__11_), .Y(_1253_) );
MUX2X1 MUX2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1253_), .B(_14918__bF_buf0), .S(_1234_), .Y(_117__11_) );
INVX1 INVX1_826 ( .gnd(gnd), .vdd(vdd), .A(data_204__12_), .Y(_1254_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf2), .C(_1254_), .Y(_1255_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_1225__bF_buf2), .C(_1231_), .Y(_1256_) );
AND2X2 AND2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(_1256_), .Y(_117__12_) );
INVX1 INVX1_827 ( .gnd(gnd), .vdd(vdd), .A(data_204__13_), .Y(_1257_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf1), .C(_1257_), .Y(_1258_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_1245_), .Y(_1259_) );
AND2X2 AND2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_1259_), .B(_1258_), .Y(_117__13_) );
INVX1 INVX1_828 ( .gnd(gnd), .vdd(vdd), .A(data_204__14_), .Y(_1260_) );
MUX2X1 MUX2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_15060__bF_buf14), .S(_1234_), .Y(_117__14_) );
INVX1 INVX1_829 ( .gnd(gnd), .vdd(vdd), .A(data_204__15_), .Y(_1261_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1229__bF_buf0), .C(_1261_), .Y(_1262_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf10), .B(_1245_), .Y(_1263_) );
AND2X2 AND2X2_387 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_1262_), .Y(_117__15_) );
INVX1 INVX1_830 ( .gnd(gnd), .vdd(vdd), .A(data_203__0_), .Y(_1264_) );
INVX1 INVX1_831 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .Y(_1265_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_1265_), .C(_1079__bF_buf3), .Y(_1266_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .B(_15025__bF_buf3), .C(IDATA_PROG_write_bF_buf5), .Y(_1267_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1036__bF_buf1), .B(_15951_), .C(_1267_), .Y(_1268_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1034_), .Y(_1269_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1269_), .Y(_1270_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1270_), .C(_1264_), .Y(_1271_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1269_), .B(_1000__bF_buf4), .Y(_1272_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_1272_), .C(_1225__bF_buf1), .Y(_1273_) );
AND2X2 AND2X2_388 ( .gnd(gnd), .vdd(vdd), .A(_1271_), .B(_1273_), .Y(_116__0_) );
INVX1 INVX1_832 ( .gnd(gnd), .vdd(vdd), .A(data_203__1_), .Y(_1274_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1270_), .C(_1274_), .Y(_1275_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_1272_), .C(_1225__bF_buf0), .Y(_1276_) );
AND2X2 AND2X2_389 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1276_), .Y(_116__1_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_1266__bF_buf3), .Y(_1277_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(data_203__2_), .B(_1277_), .Y(_1278_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_1277_), .C(_1278_), .Y(_116__2_) );
INVX1 INVX1_833 ( .gnd(gnd), .vdd(vdd), .A(data_203__3_), .Y(_1279_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1270_), .C(_1279_), .Y(_1280_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_1272_), .C(_1225__bF_buf6), .Y(_1281_) );
AND2X2 AND2X2_390 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1281_), .Y(_116__3_) );
INVX1 INVX1_834 ( .gnd(gnd), .vdd(vdd), .A(data_203__4_), .Y(_1282_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1270_), .C(_1282_), .Y(_1283_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_1272_), .C(_1225__bF_buf5), .Y(_1284_) );
AND2X2 AND2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1284_), .Y(_116__4_) );
INVX1 INVX1_835 ( .gnd(gnd), .vdd(vdd), .A(data_203__5_), .Y(_1285_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1270_), .C(_1285_), .Y(_1286_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_1272_), .C(_1225__bF_buf4), .Y(_1287_) );
AND2X2 AND2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1287_), .Y(_116__5_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(data_203__6_), .B(_1277_), .Y(_1288_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_1277_), .C(_1288_), .Y(_116__6_) );
INVX1 INVX1_836 ( .gnd(gnd), .vdd(vdd), .A(data_203__7_), .Y(_1289_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1270_), .C(_1289_), .Y(_1290_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_1272_), .C(_1225__bF_buf3), .Y(_1291_) );
AND2X2 AND2X2_393 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1291_), .Y(_116__7_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(data_203__8_), .B(_1277_), .Y(_1292_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_1277_), .C(_1292_), .Y(_116__8_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(data_203__9_), .B(_1277_), .Y(_1293_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_1277_), .C(_1293_), .Y(_116__9_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(data_203__10_), .B(_1277_), .Y(_1294_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_1277_), .C(_1294_), .Y(_116__10_) );
INVX1 INVX1_837 ( .gnd(gnd), .vdd(vdd), .A(data_203__11_), .Y(_1295_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1270_), .C(_1295_), .Y(_1296_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_1272_), .C(_1225__bF_buf2), .Y(_1297_) );
AND2X2 AND2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_1297_), .Y(_116__11_) );
INVX1 INVX1_838 ( .gnd(gnd), .vdd(vdd), .A(data_203__12_), .Y(_1298_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1270_), .C(_1298_), .Y(_1299_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_1272_), .C(_1225__bF_buf1), .Y(_1300_) );
AND2X2 AND2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1300_), .Y(_116__12_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(data_203__13_), .B(_1277_), .Y(_1301_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_1277_), .C(_1301_), .Y(_116__13_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(data_203__14_), .B(_1277_), .Y(_1302_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_1277_), .C(_1302_), .Y(_116__14_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(data_203__15_), .B(_1277_), .Y(_1303_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_1277_), .C(_1303_), .Y(_116__15_) );
INVX1 INVX1_839 ( .gnd(gnd), .vdd(vdd), .A(data_202__0_), .Y(_1304_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_15064_), .B(_14883_), .C(IDATA_PROG_write_bF_buf4), .Y(_1305_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .Y(_1306_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14952__bF_buf3), .C(_1036__bF_buf0), .Y(_1307_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_1306_), .C(_1307_), .Y(_1308_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_1308_), .Y(_1309_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1309_), .Y(_1310_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1310_), .C(_1304_), .Y(_1311_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1000__bF_buf2), .Y(_1312_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_1312_), .C(_1225__bF_buf0), .Y(_1313_) );
AND2X2 AND2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1313_), .Y(_115__0_) );
INVX1 INVX1_840 ( .gnd(gnd), .vdd(vdd), .A(data_202__1_), .Y(_1314_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1225__bF_buf6), .Y(_1315_) );
MUX2X1 MUX2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_14894__bF_buf0), .S(_1315_), .Y(_115__1_) );
INVX1 INVX1_841 ( .gnd(gnd), .vdd(vdd), .A(data_202__2_), .Y(_1316_) );
MUX2X1 MUX2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_14897__bF_buf10), .S(_1315_), .Y(_115__2_) );
INVX1 INVX1_842 ( .gnd(gnd), .vdd(vdd), .A(data_202__3_), .Y(_1317_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1310_), .C(_1317_), .Y(_1318_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_1312_), .C(_1225__bF_buf5), .Y(_1319_) );
AND2X2 AND2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1319_), .Y(_115__3_) );
INVX1 INVX1_843 ( .gnd(gnd), .vdd(vdd), .A(data_202__4_), .Y(_1320_) );
MUX2X1 MUX2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_14902__bF_buf11), .S(_1315_), .Y(_115__4_) );
INVX1 INVX1_844 ( .gnd(gnd), .vdd(vdd), .A(data_202__5_), .Y(_1321_) );
MUX2X1 MUX2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_14903__bF_buf12), .S(_1315_), .Y(_115__5_) );
INVX1 INVX1_845 ( .gnd(gnd), .vdd(vdd), .A(data_202__6_), .Y(_1322_) );
MUX2X1 MUX2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(_15049__bF_buf11), .S(_1315_), .Y(_115__6_) );
INVX1 INVX1_846 ( .gnd(gnd), .vdd(vdd), .A(data_202__7_), .Y(_1323_) );
MUX2X1 MUX2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_14908__bF_buf11), .S(_1315_), .Y(_115__7_) );
INVX1 INVX1_847 ( .gnd(gnd), .vdd(vdd), .A(data_202__8_), .Y(_1324_) );
MUX2X1 MUX2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(_15052__bF_buf9), .S(_1315_), .Y(_115__8_) );
INVX1 INVX1_848 ( .gnd(gnd), .vdd(vdd), .A(data_202__9_), .Y(_1325_) );
MUX2X1 MUX2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_14913__bF_buf11), .S(_1315_), .Y(_115__9_) );
INVX1 INVX1_849 ( .gnd(gnd), .vdd(vdd), .A(data_202__10_), .Y(_1326_) );
MUX2X1 MUX2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(_15055__bF_buf9), .S(_1315_), .Y(_115__10_) );
INVX1 INVX1_850 ( .gnd(gnd), .vdd(vdd), .A(data_202__11_), .Y(_1327_) );
MUX2X1 MUX2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1327_), .B(_14918__bF_buf12), .S(_1315_), .Y(_115__11_) );
INVX1 INVX1_851 ( .gnd(gnd), .vdd(vdd), .A(data_202__12_), .Y(_1328_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1310_), .C(_1328_), .Y(_1329_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_1312_), .C(_1225__bF_buf4), .Y(_1330_) );
AND2X2 AND2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1330_), .Y(_115__12_) );
INVX1 INVX1_852 ( .gnd(gnd), .vdd(vdd), .A(data_202__13_), .Y(_1331_) );
MUX2X1 MUX2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .B(_14924__bF_buf8), .S(_1315_), .Y(_115__13_) );
INVX1 INVX1_853 ( .gnd(gnd), .vdd(vdd), .A(data_202__14_), .Y(_1332_) );
MUX2X1 MUX2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_15060__bF_buf12), .S(_1315_), .Y(_115__14_) );
INVX1 INVX1_854 ( .gnd(gnd), .vdd(vdd), .A(data_202__15_), .Y(_1333_) );
MUX2X1 MUX2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_15062__bF_buf8), .S(_1315_), .Y(_115__15_) );
INVX1 INVX1_855 ( .gnd(gnd), .vdd(vdd), .A(data_201__0_), .Y(_1334_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_678__bF_buf6), .Y(_1335_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1335_), .Y(_1336_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_789_), .Y(_1337_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1337_), .B(_1336_), .Y(_1338_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1225__bF_buf3), .B(_1338_), .Y(_1339_) );
MUX2X1 MUX2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .B(_14932__bF_buf1), .S(_1339_), .Y(_114__0_) );
INVX1 INVX1_856 ( .gnd(gnd), .vdd(vdd), .A(data_201__1_), .Y(_1340_) );
MUX2X1 MUX2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_14894__bF_buf14), .S(_1339_), .Y(_114__1_) );
INVX1 INVX1_857 ( .gnd(gnd), .vdd(vdd), .A(data_201__2_), .Y(_1341_) );
MUX2X1 MUX2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_14897__bF_buf9), .S(_1339_), .Y(_114__2_) );
INVX1 INVX1_858 ( .gnd(gnd), .vdd(vdd), .A(data_201__3_), .Y(_1342_) );
MUX2X1 MUX2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_14899__bF_buf14), .S(_1339_), .Y(_114__3_) );
INVX1 INVX1_859 ( .gnd(gnd), .vdd(vdd), .A(data_201__4_), .Y(_1343_) );
MUX2X1 MUX2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_14902__bF_buf10), .S(_1339_), .Y(_114__4_) );
INVX1 INVX1_860 ( .gnd(gnd), .vdd(vdd), .A(data_201__5_), .Y(_1344_) );
MUX2X1 MUX2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_14903__bF_buf11), .S(_1339_), .Y(_114__5_) );
INVX1 INVX1_861 ( .gnd(gnd), .vdd(vdd), .A(data_201__6_), .Y(_1345_) );
MUX2X1 MUX2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_15049__bF_buf10), .S(_1339_), .Y(_114__6_) );
INVX1 INVX1_862 ( .gnd(gnd), .vdd(vdd), .A(data_201__7_), .Y(_1346_) );
MUX2X1 MUX2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_14908__bF_buf10), .S(_1339_), .Y(_114__7_) );
INVX1 INVX1_863 ( .gnd(gnd), .vdd(vdd), .A(data_201__8_), .Y(_1347_) );
MUX2X1 MUX2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_15052__bF_buf8), .S(_1339_), .Y(_114__8_) );
INVX1 INVX1_864 ( .gnd(gnd), .vdd(vdd), .A(data_201__9_), .Y(_1348_) );
MUX2X1 MUX2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_14913__bF_buf10), .S(_1339_), .Y(_114__9_) );
INVX1 INVX1_865 ( .gnd(gnd), .vdd(vdd), .A(data_201__10_), .Y(_1349_) );
MUX2X1 MUX2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1349_), .B(_15055__bF_buf8), .S(_1339_), .Y(_114__10_) );
INVX1 INVX1_866 ( .gnd(gnd), .vdd(vdd), .A(data_201__11_), .Y(_1350_) );
MUX2X1 MUX2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_14918__bF_buf11), .S(_1339_), .Y(_114__11_) );
INVX1 INVX1_867 ( .gnd(gnd), .vdd(vdd), .A(data_201__12_), .Y(_1351_) );
MUX2X1 MUX2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1351_), .B(_14920__bF_buf11), .S(_1339_), .Y(_114__12_) );
INVX1 INVX1_868 ( .gnd(gnd), .vdd(vdd), .A(data_201__13_), .Y(_1352_) );
MUX2X1 MUX2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_14924__bF_buf7), .S(_1339_), .Y(_114__13_) );
INVX1 INVX1_869 ( .gnd(gnd), .vdd(vdd), .A(data_201__14_), .Y(_1353_) );
MUX2X1 MUX2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1353_), .B(_15060__bF_buf11), .S(_1339_), .Y(_114__14_) );
INVX1 INVX1_870 ( .gnd(gnd), .vdd(vdd), .A(data_201__15_), .Y(_1354_) );
MUX2X1 MUX2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(_15062__bF_buf7), .S(_1339_), .Y(_114__15_) );
INVX1 INVX1_871 ( .gnd(gnd), .vdd(vdd), .A(data_200__0_), .Y(_1355_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf1), .B(_14952__bF_buf2), .C(_1036__bF_buf3), .Y(_1356_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1225__bF_buf2), .Y(_1357_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf4), .C(_1355_), .Y(_1358_) );
INVX1 INVX1_872 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .Y(_1359_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1359_), .B(_1229__bF_buf3), .Y(_1360_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_1225__bF_buf1), .C(_1360_), .Y(_1361_) );
AND2X2 AND2X2_399 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1361_), .Y(_113__0_) );
INVX1 INVX1_873 ( .gnd(gnd), .vdd(vdd), .A(data_200__1_), .Y(_1362_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf2), .C(_1362_), .Y(_1363_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_1225__bF_buf0), .C(_1360_), .Y(_1364_) );
AND2X2 AND2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1364_), .Y(_113__1_) );
INVX1 INVX1_874 ( .gnd(gnd), .vdd(vdd), .A(data_200__2_), .Y(_1365_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1229__bF_buf1), .B(_1357_), .Y(_1366_) );
MUX2X1 MUX2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_1365_), .S(_1366_), .Y(_113__2_) );
INVX1 INVX1_875 ( .gnd(gnd), .vdd(vdd), .A(data_200__3_), .Y(_1367_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf0), .C(_1367_), .Y(_1368_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_1225__bF_buf6), .C(_1360_), .Y(_1369_) );
AND2X2 AND2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(_1369_), .Y(_113__3_) );
INVX1 INVX1_876 ( .gnd(gnd), .vdd(vdd), .A(data_200__4_), .Y(_1370_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf4), .C(_1370_), .Y(_1371_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_1225__bF_buf5), .C(_1360_), .Y(_1372_) );
AND2X2 AND2X2_402 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .B(_1372_), .Y(_113__4_) );
INVX1 INVX1_877 ( .gnd(gnd), .vdd(vdd), .A(data_200__5_), .Y(_1373_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf3), .C(_1373_), .Y(_1374_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_1225__bF_buf4), .C(_1360_), .Y(_1375_) );
AND2X2 AND2X2_403 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .B(_1375_), .Y(_113__5_) );
INVX1 INVX1_878 ( .gnd(gnd), .vdd(vdd), .A(data_200__6_), .Y(_1376_) );
MUX2X1 MUX2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_1376_), .S(_1366_), .Y(_113__6_) );
INVX1 INVX1_879 ( .gnd(gnd), .vdd(vdd), .A(data_200__7_), .Y(_1377_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf2), .C(_1377_), .Y(_1378_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_1225__bF_buf3), .C(_1360_), .Y(_1379_) );
AND2X2 AND2X2_404 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .B(_1379_), .Y(_113__7_) );
INVX1 INVX1_880 ( .gnd(gnd), .vdd(vdd), .A(data_200__8_), .Y(_1380_) );
MUX2X1 MUX2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_1380_), .S(_1366_), .Y(_113__8_) );
INVX1 INVX1_881 ( .gnd(gnd), .vdd(vdd), .A(data_200__9_), .Y(_1381_) );
MUX2X1 MUX2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_1381_), .S(_1366_), .Y(_113__9_) );
INVX1 INVX1_882 ( .gnd(gnd), .vdd(vdd), .A(data_200__10_), .Y(_1382_) );
MUX2X1 MUX2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_1382_), .S(_1366_), .Y(_113__10_) );
INVX1 INVX1_883 ( .gnd(gnd), .vdd(vdd), .A(data_200__11_), .Y(_1383_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf1), .C(_1383_), .Y(_1384_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_1225__bF_buf2), .C(_1360_), .Y(_1385_) );
AND2X2 AND2X2_405 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1385_), .Y(_113__11_) );
INVX1 INVX1_884 ( .gnd(gnd), .vdd(vdd), .A(data_200__12_), .Y(_1386_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1229__bF_buf0), .C(_1386_), .Y(_1387_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_1225__bF_buf1), .C(_1360_), .Y(_1388_) );
AND2X2 AND2X2_406 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_1388_), .Y(_113__12_) );
INVX1 INVX1_885 ( .gnd(gnd), .vdd(vdd), .A(data_200__13_), .Y(_1389_) );
MUX2X1 MUX2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_1389_), .S(_1366_), .Y(_113__13_) );
INVX1 INVX1_886 ( .gnd(gnd), .vdd(vdd), .A(data_200__14_), .Y(_1390_) );
MUX2X1 MUX2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_1390_), .S(_1366_), .Y(_113__14_) );
INVX1 INVX1_887 ( .gnd(gnd), .vdd(vdd), .A(data_200__15_), .Y(_1391_) );
MUX2X1 MUX2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_1391_), .S(_1366_), .Y(_113__15_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_1306_), .C(_1034_), .Y(_1392_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1392_), .Y(_1393_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1266__bF_buf5), .Y(_1394_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(data_199__0_), .B(_1394_), .Y(_1395_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_1394_), .C(_1395_), .Y(_110__0_) );
INVX1 INVX1_888 ( .gnd(gnd), .vdd(vdd), .A(data_199__1_), .Y(_1396_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1393_), .C(_1396_), .Y(_1397_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .B(_1000__bF_buf0), .Y(_1398_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_1398_), .C(_1225__bF_buf0), .Y(_1399_) );
AND2X2 AND2X2_407 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1399_), .Y(_110__1_) );
INVX1 INVX1_889 ( .gnd(gnd), .vdd(vdd), .A(data_199__2_), .Y(_1400_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_1225__bF_buf6), .Y(_1401_) );
MUX2X1 MUX2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_14897__bF_buf7), .S(_1401_), .Y(_110__2_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(data_199__3_), .B(_1394_), .Y(_1402_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_1394_), .C(_1402_), .Y(_110__3_) );
INVX1 INVX1_890 ( .gnd(gnd), .vdd(vdd), .A(data_199__4_), .Y(_1403_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1393_), .C(_1403_), .Y(_1404_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_1398_), .C(_1225__bF_buf5), .Y(_1405_) );
AND2X2 AND2X2_408 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1405_), .Y(_110__4_) );
INVX1 INVX1_891 ( .gnd(gnd), .vdd(vdd), .A(data_199__5_), .Y(_1406_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1393_), .C(_1406_), .Y(_1407_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_1398_), .C(_1225__bF_buf4), .Y(_1408_) );
AND2X2 AND2X2_409 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1408_), .Y(_110__5_) );
INVX1 INVX1_892 ( .gnd(gnd), .vdd(vdd), .A(data_199__6_), .Y(_1409_) );
MUX2X1 MUX2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_15049__bF_buf8), .S(_1401_), .Y(_110__6_) );
INVX1 INVX1_893 ( .gnd(gnd), .vdd(vdd), .A(data_199__7_), .Y(_1410_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1393_), .C(_1410_), .Y(_1411_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_1398_), .C(_1225__bF_buf3), .Y(_1412_) );
AND2X2 AND2X2_410 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_1412_), .Y(_110__7_) );
INVX1 INVX1_894 ( .gnd(gnd), .vdd(vdd), .A(data_199__8_), .Y(_1413_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1393_), .C(_1413_), .Y(_1414_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_1394_), .Y(_1415_) );
AND2X2 AND2X2_411 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_1414_), .Y(_110__8_) );
INVX1 INVX1_895 ( .gnd(gnd), .vdd(vdd), .A(data_199__9_), .Y(_1416_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1393_), .C(_1416_), .Y(_1417_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_1394_), .Y(_1418_) );
AND2X2 AND2X2_412 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1417_), .Y(_110__9_) );
INVX1 INVX1_896 ( .gnd(gnd), .vdd(vdd), .A(data_199__10_), .Y(_1419_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1393_), .C(_1419_), .Y(_1420_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_1394_), .Y(_1421_) );
AND2X2 AND2X2_413 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1420_), .Y(_110__10_) );
INVX1 INVX1_897 ( .gnd(gnd), .vdd(vdd), .A(data_199__11_), .Y(_1422_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1393_), .C(_1422_), .Y(_1423_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_1398_), .C(_1225__bF_buf2), .Y(_1424_) );
AND2X2 AND2X2_414 ( .gnd(gnd), .vdd(vdd), .A(_1423_), .B(_1424_), .Y(_110__11_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(data_199__12_), .B(_1394_), .Y(_1425_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_1394_), .C(_1425_), .Y(_110__12_) );
INVX1 INVX1_898 ( .gnd(gnd), .vdd(vdd), .A(data_199__13_), .Y(_1426_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1393_), .C(_1426_), .Y(_1427_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_1394_), .Y(_1428_) );
AND2X2 AND2X2_415 ( .gnd(gnd), .vdd(vdd), .A(_1428_), .B(_1427_), .Y(_110__13_) );
INVX1 INVX1_899 ( .gnd(gnd), .vdd(vdd), .A(data_199__14_), .Y(_1429_) );
MUX2X1 MUX2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1429_), .B(_15060__bF_buf9), .S(_1401_), .Y(_110__14_) );
INVX1 INVX1_900 ( .gnd(gnd), .vdd(vdd), .A(data_199__15_), .Y(_1430_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1393_), .C(_1430_), .Y(_1431_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_1394_), .Y(_1432_) );
AND2X2 AND2X2_416 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(_1431_), .Y(_110__15_) );
INVX1 INVX1_901 ( .gnd(gnd), .vdd(vdd), .A(data_198__0_), .Y(_1433_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_16204_), .B(_14965__bF_buf0), .C(_1305_), .Y(_1434_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_15360_), .B(_15025__bF_buf2), .C(_1434_), .Y(_1435_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_1435_), .Y(_1436_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1436_), .Y(_1437_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1437_), .C(_1433_), .Y(_1438_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1000__bF_buf3), .Y(_1439_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_1439_), .C(_1225__bF_buf1), .Y(_1440_) );
AND2X2 AND2X2_417 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1440_), .Y(_109__0_) );
INVX1 INVX1_902 ( .gnd(gnd), .vdd(vdd), .A(data_198__1_), .Y(_1441_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1437_), .C(_1441_), .Y(_1442_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_1439_), .C(_1225__bF_buf0), .Y(_1443_) );
AND2X2 AND2X2_418 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1443_), .Y(_109__1_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1437_), .B(_1266__bF_buf4), .Y(_1444_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(data_198__2_), .B(_1444_), .Y(_1445_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_1444_), .C(_1445_), .Y(_109__2_) );
INVX1 INVX1_903 ( .gnd(gnd), .vdd(vdd), .A(data_198__3_), .Y(_1446_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1437_), .C(_1446_), .Y(_1447_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_1439_), .C(_1225__bF_buf6), .Y(_1448_) );
AND2X2 AND2X2_419 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1448_), .Y(_109__3_) );
INVX1 INVX1_904 ( .gnd(gnd), .vdd(vdd), .A(data_198__4_), .Y(_1449_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1437_), .C(_1449_), .Y(_1450_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_1439_), .C(_1225__bF_buf5), .Y(_1451_) );
AND2X2 AND2X2_420 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1451_), .Y(_109__4_) );
INVX1 INVX1_905 ( .gnd(gnd), .vdd(vdd), .A(data_198__5_), .Y(_1452_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1437_), .C(_1452_), .Y(_1453_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_1439_), .C(_1225__bF_buf4), .Y(_1454_) );
AND2X2 AND2X2_421 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1454_), .Y(_109__5_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(data_198__6_), .B(_1444_), .Y(_1455_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_1444_), .C(_1455_), .Y(_109__6_) );
INVX1 INVX1_906 ( .gnd(gnd), .vdd(vdd), .A(data_198__7_), .Y(_1456_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1437_), .C(_1456_), .Y(_1457_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_1439_), .C(_1225__bF_buf3), .Y(_1458_) );
AND2X2 AND2X2_422 ( .gnd(gnd), .vdd(vdd), .A(_1457_), .B(_1458_), .Y(_109__7_) );
INVX1 INVX1_907 ( .gnd(gnd), .vdd(vdd), .A(data_198__8_), .Y(_1459_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1437_), .C(_1459_), .Y(_1460_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_1444_), .Y(_1461_) );
AND2X2 AND2X2_423 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_1460_), .Y(_109__8_) );
INVX1 INVX1_908 ( .gnd(gnd), .vdd(vdd), .A(data_198__9_), .Y(_1462_) );
OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1437_), .C(_1462_), .Y(_1463_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf7), .B(_1444_), .Y(_1464_) );
AND2X2 AND2X2_424 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1463_), .Y(_109__9_) );
INVX1 INVX1_909 ( .gnd(gnd), .vdd(vdd), .A(data_198__10_), .Y(_1465_) );
OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1437_), .C(_1465_), .Y(_1466_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_1444_), .Y(_1467_) );
AND2X2 AND2X2_425 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_1466_), .Y(_109__10_) );
INVX1 INVX1_910 ( .gnd(gnd), .vdd(vdd), .A(data_198__11_), .Y(_1468_) );
OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1437_), .C(_1468_), .Y(_1469_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_1439_), .C(_1225__bF_buf2), .Y(_1470_) );
AND2X2 AND2X2_426 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1470_), .Y(_109__11_) );
INVX1 INVX1_911 ( .gnd(gnd), .vdd(vdd), .A(data_198__12_), .Y(_1471_) );
OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1437_), .C(_1471_), .Y(_1472_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_1439_), .C(_1225__bF_buf1), .Y(_1473_) );
AND2X2 AND2X2_427 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .B(_1473_), .Y(_109__12_) );
INVX1 INVX1_912 ( .gnd(gnd), .vdd(vdd), .A(data_198__13_), .Y(_1474_) );
OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1437_), .C(_1474_), .Y(_1475_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_1444_), .Y(_1476_) );
AND2X2 AND2X2_428 ( .gnd(gnd), .vdd(vdd), .A(_1476_), .B(_1475_), .Y(_109__13_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(data_198__14_), .B(_1444_), .Y(_1477_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_1444_), .C(_1477_), .Y(_109__14_) );
INVX1 INVX1_913 ( .gnd(gnd), .vdd(vdd), .A(data_198__15_), .Y(_1478_) );
OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1437_), .C(_1478_), .Y(_1479_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_1444_), .Y(_1480_) );
AND2X2 AND2X2_429 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1479_), .Y(_109__15_) );
INVX1 INVX1_914 ( .gnd(gnd), .vdd(vdd), .A(data_197__0_), .Y(_1481_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_15509_), .B(_887_), .Y(_1482_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf1), .B(_15453_), .Y(_1483_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .B(_1482_), .C(_1483_), .Y(_1484_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1484_), .C(_1335_), .Y(_1485_) );
OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1485_), .C(_1481_), .Y(_1486_) );
INVX1 INVX1_915 ( .gnd(gnd), .vdd(vdd), .A(_1482_), .Y(_1487_) );
OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(_1306_), .C(_1034_), .Y(_1488_) );
NOR3X1 NOR3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1488_), .C(_1000__bF_buf2), .Y(_1489_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_1489_), .C(_1225__bF_buf0), .Y(_1490_) );
AND2X2 AND2X2_430 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .B(_1490_), .Y(_108__0_) );
INVX1 INVX1_916 ( .gnd(gnd), .vdd(vdd), .A(data_197__1_), .Y(_1491_) );
OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1485_), .C(_1491_), .Y(_1492_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_1489_), .C(_1225__bF_buf6), .Y(_1493_) );
AND2X2 AND2X2_431 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1493_), .Y(_108__1_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_1266__bF_buf2), .Y(_1494_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(data_197__2_), .B(_1494_), .Y(_1495_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_1494_), .C(_1495_), .Y(_108__2_) );
INVX1 INVX1_917 ( .gnd(gnd), .vdd(vdd), .A(data_197__3_), .Y(_1496_) );
OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf1), .B(_1485_), .C(_1496_), .Y(_1497_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_1489_), .C(_1225__bF_buf5), .Y(_1498_) );
AND2X2 AND2X2_432 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .B(_1498_), .Y(_108__3_) );
INVX1 INVX1_918 ( .gnd(gnd), .vdd(vdd), .A(data_197__4_), .Y(_1499_) );
OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf0), .B(_1485_), .C(_1499_), .Y(_1500_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_1489_), .C(_1225__bF_buf4), .Y(_1501_) );
AND2X2 AND2X2_433 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1501_), .Y(_108__4_) );
INVX1 INVX1_919 ( .gnd(gnd), .vdd(vdd), .A(data_197__5_), .Y(_1502_) );
OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf5), .B(_1485_), .C(_1502_), .Y(_1503_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_1489_), .C(_1225__bF_buf3), .Y(_1504_) );
AND2X2 AND2X2_434 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .B(_1504_), .Y(_108__5_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(data_197__6_), .B(_1494_), .Y(_1505_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_1494_), .C(_1505_), .Y(_108__6_) );
INVX1 INVX1_920 ( .gnd(gnd), .vdd(vdd), .A(data_197__7_), .Y(_1506_) );
OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf4), .B(_1485_), .C(_1506_), .Y(_1507_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_1489_), .C(_1225__bF_buf2), .Y(_1508_) );
AND2X2 AND2X2_435 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .B(_1508_), .Y(_108__7_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(data_197__8_), .B(_1494_), .Y(_1509_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_1494_), .C(_1509_), .Y(_108__8_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(data_197__9_), .B(_1494_), .Y(_1510_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_1494_), .C(_1510_), .Y(_108__9_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(data_197__10_), .B(_1494_), .Y(_1511_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_1494_), .C(_1511_), .Y(_108__10_) );
INVX1 INVX1_921 ( .gnd(gnd), .vdd(vdd), .A(data_197__11_), .Y(_1512_) );
OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf3), .B(_1485_), .C(_1512_), .Y(_1513_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_1489_), .C(_1225__bF_buf1), .Y(_1514_) );
AND2X2 AND2X2_436 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(_1514_), .Y(_108__11_) );
INVX1 INVX1_922 ( .gnd(gnd), .vdd(vdd), .A(data_197__12_), .Y(_1515_) );
OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_1266__bF_buf2), .B(_1485_), .C(_1515_), .Y(_1516_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_1489_), .C(_1225__bF_buf0), .Y(_1517_) );
AND2X2 AND2X2_437 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1517_), .Y(_108__12_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(data_197__13_), .B(_1494_), .Y(_1518_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_1494_), .C(_1518_), .Y(_108__13_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(data_197__14_), .B(_1494_), .Y(_1519_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_1494_), .C(_1519_), .Y(_108__14_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(data_197__15_), .B(_1494_), .Y(_1520_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_1494_), .C(_1520_), .Y(_108__15_) );
INVX1 INVX1_923 ( .gnd(gnd), .vdd(vdd), .A(data_196__0_), .Y(_1521_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(_1229__bF_buf4), .Y(_1522_) );
OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14965__bF_buf3), .C(_1036__bF_buf2), .Y(_1523_) );
INVX1 INVX1_924 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .Y(_1524_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1266__bF_buf1), .Y(_1525_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1525__bF_buf4), .Y(_1526_) );
MUX2X1 MUX2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_14932__bF_buf11), .S(_1526_), .Y(_107__0_) );
INVX1 INVX1_925 ( .gnd(gnd), .vdd(vdd), .A(data_196__1_), .Y(_1527_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1225__bF_buf6), .Y(_1528_) );
OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf5), .B(_1229__bF_buf3), .C(_1527_), .Y(_1529_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_1522_), .C(_1525__bF_buf3), .Y(_1530_) );
AND2X2 AND2X2_438 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1529_), .Y(_107__1_) );
INVX1 INVX1_926 ( .gnd(gnd), .vdd(vdd), .A(data_196__2_), .Y(_1531_) );
OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1229__bF_buf2), .C(_1531_), .Y(_1532_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1229__bF_buf1), .B(_1528__bF_buf3), .Y(_1533_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_1533_), .Y(_1534_) );
AND2X2 AND2X2_439 ( .gnd(gnd), .vdd(vdd), .A(_1534_), .B(_1532_), .Y(_107__2_) );
INVX1 INVX1_927 ( .gnd(gnd), .vdd(vdd), .A(data_196__3_), .Y(_1535_) );
MUX2X1 MUX2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_14899__bF_buf9), .S(_1526_), .Y(_107__3_) );
INVX1 INVX1_928 ( .gnd(gnd), .vdd(vdd), .A(data_196__4_), .Y(_1536_) );
OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf2), .B(_1229__bF_buf0), .C(_1536_), .Y(_1537_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_1522_), .C(_1525__bF_buf2), .Y(_1538_) );
AND2X2 AND2X2_440 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1537_), .Y(_107__4_) );
INVX1 INVX1_929 ( .gnd(gnd), .vdd(vdd), .A(data_196__5_), .Y(_1539_) );
OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf1), .B(_1229__bF_buf4), .C(_1539_), .Y(_1540_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_1522_), .C(_1525__bF_buf1), .Y(_1541_) );
AND2X2 AND2X2_441 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1540_), .Y(_107__5_) );
INVX1 INVX1_930 ( .gnd(gnd), .vdd(vdd), .A(data_196__6_), .Y(_1542_) );
OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf0), .B(_1229__bF_buf3), .C(_1542_), .Y(_1543_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_1533_), .Y(_1544_) );
AND2X2 AND2X2_442 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1543_), .Y(_107__6_) );
INVX1 INVX1_931 ( .gnd(gnd), .vdd(vdd), .A(data_196__7_), .Y(_1545_) );
OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf5), .B(_1229__bF_buf2), .C(_1545_), .Y(_1546_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_1522_), .C(_1525__bF_buf0), .Y(_1547_) );
AND2X2 AND2X2_443 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1546_), .Y(_107__7_) );
INVX1 INVX1_932 ( .gnd(gnd), .vdd(vdd), .A(data_196__8_), .Y(_1548_) );
MUX2X1 MUX2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_15052__bF_buf3), .S(_1526_), .Y(_107__8_) );
INVX1 INVX1_933 ( .gnd(gnd), .vdd(vdd), .A(data_196__9_), .Y(_1549_) );
MUX2X1 MUX2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_14913__bF_buf5), .S(_1526_), .Y(_107__9_) );
INVX1 INVX1_934 ( .gnd(gnd), .vdd(vdd), .A(data_196__10_), .Y(_1550_) );
MUX2X1 MUX2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_15055__bF_buf3), .S(_1526_), .Y(_107__10_) );
INVX1 INVX1_935 ( .gnd(gnd), .vdd(vdd), .A(data_196__11_), .Y(_1551_) );
OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1229__bF_buf1), .C(_1551_), .Y(_1552_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_1522_), .C(_1525__bF_buf4), .Y(_1553_) );
AND2X2 AND2X2_444 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1552_), .Y(_107__11_) );
INVX1 INVX1_936 ( .gnd(gnd), .vdd(vdd), .A(data_196__12_), .Y(_1554_) );
MUX2X1 MUX2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_14920__bF_buf6), .S(_1526_), .Y(_107__12_) );
INVX1 INVX1_937 ( .gnd(gnd), .vdd(vdd), .A(data_196__13_), .Y(_1555_) );
MUX2X1 MUX2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_14924__bF_buf2), .S(_1526_), .Y(_107__13_) );
INVX1 INVX1_938 ( .gnd(gnd), .vdd(vdd), .A(data_196__14_), .Y(_1556_) );
OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf3), .B(_1229__bF_buf0), .C(_1556_), .Y(_1557_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_1533_), .Y(_1558_) );
AND2X2 AND2X2_445 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1557_), .Y(_107__14_) );
INVX1 INVX1_939 ( .gnd(gnd), .vdd(vdd), .A(data_196__15_), .Y(_1559_) );
MUX2X1 MUX2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_15062__bF_buf2), .S(_1526_), .Y(_107__15_) );
INVX1 INVX1_940 ( .gnd(gnd), .vdd(vdd), .A(data_195__0_), .Y(_1560_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_14884_), .B(_14938_), .Y(_1561_) );
INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .Y(_1562_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_15035_), .C(_14882__bF_buf11), .Y(_1563_) );
OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_15025__bF_buf0), .C(_1563_), .Y(_1564_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1036__bF_buf1), .B(_15580_), .C(_1564_), .Y(_1565_) );
OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf2), .B(_1562__bF_buf3), .C(_1565_), .Y(_1566_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1335_), .Y(_1567_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .B(_1566_), .Y(_1568_) );
OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf2), .B(_1568_), .C(_1560_), .Y(_1569_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(_1567_), .Y(_1570_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_1570_), .C(_1525__bF_buf3), .Y(_1571_) );
AND2X2 AND2X2_446 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1569_), .Y(_106__0_) );
INVX1 INVX1_941 ( .gnd(gnd), .vdd(vdd), .A(data_195__1_), .Y(_1572_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1525__bF_buf2), .Y(_1573_) );
MUX2X1 MUX2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_14894__bF_buf8), .S(_1573_), .Y(_106__1_) );
INVX1 INVX1_942 ( .gnd(gnd), .vdd(vdd), .A(data_195__2_), .Y(_1574_) );
MUX2X1 MUX2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1574_), .B(_14897__bF_buf3), .S(_1573_), .Y(_106__2_) );
INVX1 INVX1_943 ( .gnd(gnd), .vdd(vdd), .A(data_195__3_), .Y(_1575_) );
OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf1), .B(_1568_), .C(_1575_), .Y(_1576_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_1570_), .C(_1525__bF_buf1), .Y(_1577_) );
AND2X2 AND2X2_447 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1576_), .Y(_106__3_) );
INVX1 INVX1_944 ( .gnd(gnd), .vdd(vdd), .A(data_195__4_), .Y(_1578_) );
MUX2X1 MUX2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1578_), .B(_14902__bF_buf4), .S(_1573_), .Y(_106__4_) );
INVX1 INVX1_945 ( .gnd(gnd), .vdd(vdd), .A(data_195__5_), .Y(_1579_) );
MUX2X1 MUX2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_14903__bF_buf5), .S(_1573_), .Y(_106__5_) );
INVX1 INVX1_946 ( .gnd(gnd), .vdd(vdd), .A(data_195__6_), .Y(_1580_) );
MUX2X1 MUX2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_15049__bF_buf4), .S(_1573_), .Y(_106__6_) );
INVX1 INVX1_947 ( .gnd(gnd), .vdd(vdd), .A(data_195__7_), .Y(_1581_) );
MUX2X1 MUX2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(_14908__bF_buf4), .S(_1573_), .Y(_106__7_) );
INVX1 INVX1_948 ( .gnd(gnd), .vdd(vdd), .A(data_195__8_), .Y(_1582_) );
OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf0), .B(_1568_), .C(_1582_), .Y(_1583_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1568_), .B(_1528__bF_buf5), .Y(_1584_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_1584_), .Y(_1585_) );
AND2X2 AND2X2_448 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1583_), .Y(_106__8_) );
INVX1 INVX1_949 ( .gnd(gnd), .vdd(vdd), .A(data_195__9_), .Y(_1586_) );
OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1568_), .C(_1586_), .Y(_1587_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_1584_), .Y(_1588_) );
AND2X2 AND2X2_449 ( .gnd(gnd), .vdd(vdd), .A(_1588_), .B(_1587_), .Y(_106__9_) );
INVX1 INVX1_950 ( .gnd(gnd), .vdd(vdd), .A(data_195__10_), .Y(_1589_) );
OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf3), .B(_1568_), .C(_1589_), .Y(_1590_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_1584_), .Y(_1591_) );
AND2X2 AND2X2_450 ( .gnd(gnd), .vdd(vdd), .A(_1591_), .B(_1590_), .Y(_106__10_) );
INVX1 INVX1_951 ( .gnd(gnd), .vdd(vdd), .A(data_195__11_), .Y(_1592_) );
MUX2X1 MUX2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1592_), .B(_14918__bF_buf5), .S(_1573_), .Y(_106__11_) );
INVX1 INVX1_952 ( .gnd(gnd), .vdd(vdd), .A(data_195__12_), .Y(_1593_) );
OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf2), .B(_1568_), .C(_1593_), .Y(_1594_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_1570_), .C(_1525__bF_buf0), .Y(_1595_) );
AND2X2 AND2X2_451 ( .gnd(gnd), .vdd(vdd), .A(_1595_), .B(_1594_), .Y(_106__12_) );
INVX1 INVX1_953 ( .gnd(gnd), .vdd(vdd), .A(data_195__13_), .Y(_1596_) );
OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf1), .B(_1568_), .C(_1596_), .Y(_1597_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_1584_), .Y(_1598_) );
AND2X2 AND2X2_452 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .B(_1597_), .Y(_106__13_) );
INVX1 INVX1_954 ( .gnd(gnd), .vdd(vdd), .A(data_195__14_), .Y(_1599_) );
MUX2X1 MUX2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_15060__bF_buf5), .S(_1573_), .Y(_106__14_) );
INVX1 INVX1_955 ( .gnd(gnd), .vdd(vdd), .A(data_195__15_), .Y(_1600_) );
OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf0), .B(_1568_), .C(_1600_), .Y(_1601_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_1584_), .Y(_1602_) );
AND2X2 AND2X2_453 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1601_), .Y(_106__15_) );
INVX1 INVX1_956 ( .gnd(gnd), .vdd(vdd), .A(data_194__0_), .Y(_1603_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .Y(_1604_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf4), .B(_15571_), .Y(_1605_) );
INVX1 INVX1_957 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1606_) );
OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_1562__bF_buf2), .B(_14942__bF_buf2), .C(IDATA_PROG_write_bF_buf3), .Y(_1607_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf1), .B(_1036__bF_buf0), .C(_1607_), .Y(_1608_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .B(_1608_), .C(_1335_), .Y(_1609_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .B(_1609_), .Y(_1610_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1610_), .B(_1525__bF_buf4), .Y(_1611_) );
MUX2X1 MUX2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1603_), .B(_14932__bF_buf9), .S(_1611_), .Y(_105__0_) );
INVX1 INVX1_958 ( .gnd(gnd), .vdd(vdd), .A(data_194__1_), .Y(_1612_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_1604_), .Y(_1613_) );
OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf5), .B(_1613_), .C(_1612_), .Y(_1614_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_1610_), .C(_1525__bF_buf3), .Y(_1615_) );
AND2X2 AND2X2_454 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1614_), .Y(_105__1_) );
INVX1 INVX1_959 ( .gnd(gnd), .vdd(vdd), .A(data_194__2_), .Y(_1616_) );
OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1613_), .C(_1616_), .Y(_1617_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1613_), .B(_1528__bF_buf3), .Y(_1618_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_1618_), .Y(_1619_) );
AND2X2 AND2X2_455 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(_1617_), .Y(_105__2_) );
INVX1 INVX1_960 ( .gnd(gnd), .vdd(vdd), .A(data_194__3_), .Y(_1620_) );
MUX2X1 MUX2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_14899__bF_buf7), .S(_1611_), .Y(_105__3_) );
INVX1 INVX1_961 ( .gnd(gnd), .vdd(vdd), .A(data_194__4_), .Y(_1621_) );
OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf2), .B(_1613_), .C(_1621_), .Y(_1622_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_1610_), .C(_1525__bF_buf2), .Y(_1623_) );
AND2X2 AND2X2_456 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1622_), .Y(_105__4_) );
INVX1 INVX1_962 ( .gnd(gnd), .vdd(vdd), .A(data_194__5_), .Y(_1624_) );
OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf1), .B(_1613_), .C(_1624_), .Y(_1625_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_1610_), .C(_1525__bF_buf1), .Y(_1626_) );
AND2X2 AND2X2_457 ( .gnd(gnd), .vdd(vdd), .A(_1626_), .B(_1625_), .Y(_105__5_) );
INVX1 INVX1_963 ( .gnd(gnd), .vdd(vdd), .A(data_194__6_), .Y(_1627_) );
OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf0), .B(_1613_), .C(_1627_), .Y(_1628_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_1618_), .Y(_1629_) );
AND2X2 AND2X2_458 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1628_), .Y(_105__6_) );
INVX1 INVX1_964 ( .gnd(gnd), .vdd(vdd), .A(data_194__7_), .Y(_1630_) );
OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf5), .B(_1613_), .C(_1630_), .Y(_1631_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_1610_), .C(_1525__bF_buf0), .Y(_1632_) );
AND2X2 AND2X2_459 ( .gnd(gnd), .vdd(vdd), .A(_1632_), .B(_1631_), .Y(_105__7_) );
INVX1 INVX1_965 ( .gnd(gnd), .vdd(vdd), .A(data_194__8_), .Y(_1633_) );
MUX2X1 MUX2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(_15052__bF_buf1), .S(_1611_), .Y(_105__8_) );
INVX1 INVX1_966 ( .gnd(gnd), .vdd(vdd), .A(data_194__9_), .Y(_1634_) );
MUX2X1 MUX2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_14913__bF_buf3), .S(_1611_), .Y(_105__9_) );
INVX1 INVX1_967 ( .gnd(gnd), .vdd(vdd), .A(data_194__10_), .Y(_1635_) );
MUX2X1 MUX2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_15055__bF_buf1), .S(_1611_), .Y(_105__10_) );
INVX1 INVX1_968 ( .gnd(gnd), .vdd(vdd), .A(data_194__11_), .Y(_1636_) );
OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1613_), .C(_1636_), .Y(_1637_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_1610_), .C(_1525__bF_buf4), .Y(_1638_) );
AND2X2 AND2X2_460 ( .gnd(gnd), .vdd(vdd), .A(_1638_), .B(_1637_), .Y(_105__11_) );
INVX1 INVX1_969 ( .gnd(gnd), .vdd(vdd), .A(data_194__12_), .Y(_1639_) );
MUX2X1 MUX2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_14920__bF_buf4), .S(_1611_), .Y(_105__12_) );
INVX1 INVX1_970 ( .gnd(gnd), .vdd(vdd), .A(data_194__13_), .Y(_1640_) );
MUX2X1 MUX2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1640_), .B(_14924__bF_buf0), .S(_1611_), .Y(_105__13_) );
INVX1 INVX1_971 ( .gnd(gnd), .vdd(vdd), .A(data_194__14_), .Y(_1641_) );
OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf3), .B(_1613_), .C(_1641_), .Y(_1642_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_1618_), .Y(_1643_) );
AND2X2 AND2X2_461 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1642_), .Y(_105__14_) );
INVX1 INVX1_972 ( .gnd(gnd), .vdd(vdd), .A(data_194__15_), .Y(_1644_) );
MUX2X1 MUX2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_15062__bF_buf0), .S(_1611_), .Y(_105__15_) );
INVX1 INVX1_973 ( .gnd(gnd), .vdd(vdd), .A(data_193__0_), .Y(_1645_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_15025__bF_buf3), .B(_475_), .Y(_1646_) );
INVX1 INVX1_974 ( .gnd(gnd), .vdd(vdd), .A(_1646_), .Y(_1647_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1647_), .C(_1335_), .Y(_1648_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1604_), .Y(_1649_) );
OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf2), .B(_1649_), .C(_1645_), .Y(_1650_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .B(_1648_), .Y(_1651_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_1651_), .C(_1525__bF_buf3), .Y(_1652_) );
AND2X2 AND2X2_462 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1650_), .Y(_104__0_) );
INVX1 INVX1_975 ( .gnd(gnd), .vdd(vdd), .A(data_193__1_), .Y(_1653_) );
OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf1), .B(_1649_), .C(_1653_), .Y(_1654_) );
NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_1651_), .C(_1525__bF_buf2), .Y(_1655_) );
AND2X2 AND2X2_463 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1654_), .Y(_104__1_) );
INVX1 INVX1_976 ( .gnd(gnd), .vdd(vdd), .A(data_193__2_), .Y(_1656_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .B(_1525__bF_buf1), .Y(_1657_) );
MUX2X1 MUX2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_14897__bF_buf1), .S(_1657_), .Y(_104__2_) );
INVX1 INVX1_977 ( .gnd(gnd), .vdd(vdd), .A(data_193__3_), .Y(_1658_) );
OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf0), .B(_1649_), .C(_1658_), .Y(_1659_) );
NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_1651_), .C(_1525__bF_buf0), .Y(_1660_) );
AND2X2 AND2X2_464 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1659_), .Y(_104__3_) );
INVX1 INVX1_978 ( .gnd(gnd), .vdd(vdd), .A(data_193__4_), .Y(_1661_) );
OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf5), .B(_1649_), .C(_1661_), .Y(_1662_) );
NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_1651_), .C(_1525__bF_buf4), .Y(_1663_) );
AND2X2 AND2X2_465 ( .gnd(gnd), .vdd(vdd), .A(_1663_), .B(_1662_), .Y(_104__4_) );
INVX1 INVX1_979 ( .gnd(gnd), .vdd(vdd), .A(data_193__5_), .Y(_1664_) );
OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1649_), .C(_1664_), .Y(_1665_) );
NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_1651_), .C(_1525__bF_buf3), .Y(_1666_) );
AND2X2 AND2X2_466 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1665_), .Y(_104__5_) );
INVX1 INVX1_980 ( .gnd(gnd), .vdd(vdd), .A(data_193__6_), .Y(_1667_) );
MUX2X1 MUX2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_15049__bF_buf2), .S(_1657_), .Y(_104__6_) );
INVX1 INVX1_981 ( .gnd(gnd), .vdd(vdd), .A(data_193__7_), .Y(_1668_) );
OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf3), .B(_1649_), .C(_1668_), .Y(_1669_) );
NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_1651_), .C(_1525__bF_buf2), .Y(_1670_) );
AND2X2 AND2X2_467 ( .gnd(gnd), .vdd(vdd), .A(_1670_), .B(_1669_), .Y(_104__7_) );
INVX1 INVX1_982 ( .gnd(gnd), .vdd(vdd), .A(data_193__8_), .Y(_1671_) );
MUX2X1 MUX2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1671_), .B(_15052__bF_buf0), .S(_1657_), .Y(_104__8_) );
INVX1 INVX1_983 ( .gnd(gnd), .vdd(vdd), .A(data_193__9_), .Y(_1672_) );
MUX2X1 MUX2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1672_), .B(_14913__bF_buf2), .S(_1657_), .Y(_104__9_) );
INVX1 INVX1_984 ( .gnd(gnd), .vdd(vdd), .A(data_193__10_), .Y(_1673_) );
MUX2X1 MUX2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1673_), .B(_15055__bF_buf0), .S(_1657_), .Y(_104__10_) );
INVX1 INVX1_985 ( .gnd(gnd), .vdd(vdd), .A(data_193__11_), .Y(_1674_) );
OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf2), .B(_1649_), .C(_1674_), .Y(_1675_) );
NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_1651_), .C(_1525__bF_buf1), .Y(_1676_) );
AND2X2 AND2X2_468 ( .gnd(gnd), .vdd(vdd), .A(_1676_), .B(_1675_), .Y(_104__11_) );
INVX1 INVX1_986 ( .gnd(gnd), .vdd(vdd), .A(data_193__12_), .Y(_1677_) );
OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf1), .B(_1649_), .C(_1677_), .Y(_1678_) );
NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_1651_), .C(_1525__bF_buf0), .Y(_1679_) );
AND2X2 AND2X2_469 ( .gnd(gnd), .vdd(vdd), .A(_1679_), .B(_1678_), .Y(_104__12_) );
INVX1 INVX1_987 ( .gnd(gnd), .vdd(vdd), .A(data_193__13_), .Y(_1680_) );
MUX2X1 MUX2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1680_), .B(_14924__bF_buf13), .S(_1657_), .Y(_104__13_) );
INVX1 INVX1_988 ( .gnd(gnd), .vdd(vdd), .A(data_193__14_), .Y(_1681_) );
MUX2X1 MUX2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .B(_15060__bF_buf3), .S(_1657_), .Y(_104__14_) );
INVX1 INVX1_989 ( .gnd(gnd), .vdd(vdd), .A(data_193__15_), .Y(_1682_) );
MUX2X1 MUX2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .B(_15062__bF_buf13), .S(_1657_), .Y(_104__15_) );
INVX1 INVX1_990 ( .gnd(gnd), .vdd(vdd), .A(data_192__0_), .Y(_1683_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_15183__bF_buf5), .B(_1335_), .Y(_1684_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_14975_), .B(_14978__bF_buf0), .Y(_1685_) );
OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14945_), .C(_15021_), .Y(_1686_) );
INVX1 INVX1_991 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .Y(_1687_) );
OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_14884_), .B(_14938_), .C(_1687_), .Y(_1688_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_1688_), .Y(_1689_) );
OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_15025__bF_buf2), .C(_1689_), .Y(_1690_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1690_), .B(_1684_), .Y(_1691_) );
NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1225__bF_buf5), .B(_1523_), .C(_1691_), .Y(_1692_) );
OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf10), .C(_1683_), .Y(_1693_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf9), .B(_1692_), .Y(_1694_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_1694__bF_buf3), .Y(_1695_) );
AND2X2 AND2X2_470 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_1693_), .Y(_103__0_) );
INVX1 INVX1_992 ( .gnd(gnd), .vdd(vdd), .A(data_192__1_), .Y(_1696_) );
OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf8), .C(_1696_), .Y(_1697_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_1694__bF_buf2), .Y(_1698_) );
AND2X2 AND2X2_471 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_1697_), .Y(_103__1_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(data_192__2_), .B(_1694__bF_buf1), .Y(_1699_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_1694__bF_buf0), .C(_1699_), .Y(_103__2_) );
INVX1 INVX1_993 ( .gnd(gnd), .vdd(vdd), .A(data_192__3_), .Y(_1700_) );
OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf7), .C(_1700_), .Y(_1701_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_1694__bF_buf3), .Y(_1702_) );
AND2X2 AND2X2_472 ( .gnd(gnd), .vdd(vdd), .A(_1702_), .B(_1701_), .Y(_103__3_) );
INVX1 INVX1_994 ( .gnd(gnd), .vdd(vdd), .A(data_192__4_), .Y(_1703_) );
OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf6), .C(_1703_), .Y(_1704_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_1694__bF_buf2), .Y(_1705_) );
AND2X2 AND2X2_473 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .B(_1704_), .Y(_103__4_) );
INVX1 INVX1_995 ( .gnd(gnd), .vdd(vdd), .A(data_192__5_), .Y(_1706_) );
OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf5), .C(_1706_), .Y(_1707_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_1694__bF_buf1), .Y(_1708_) );
AND2X2 AND2X2_474 ( .gnd(gnd), .vdd(vdd), .A(_1708_), .B(_1707_), .Y(_103__5_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(data_192__6_), .B(_1694__bF_buf0), .Y(_1709_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_1694__bF_buf3), .C(_1709_), .Y(_103__6_) );
INVX1 INVX1_996 ( .gnd(gnd), .vdd(vdd), .A(data_192__7_), .Y(_1710_) );
OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf4), .C(_1710_), .Y(_1711_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_1694__bF_buf2), .Y(_1712_) );
AND2X2 AND2X2_475 ( .gnd(gnd), .vdd(vdd), .A(_1712_), .B(_1711_), .Y(_103__7_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(data_192__8_), .B(_1694__bF_buf1), .Y(_1713_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_1694__bF_buf0), .C(_1713_), .Y(_103__8_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(data_192__9_), .B(_1694__bF_buf3), .Y(_1714_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_1694__bF_buf2), .C(_1714_), .Y(_103__9_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(data_192__10_), .B(_1694__bF_buf1), .Y(_1715_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_1694__bF_buf0), .C(_1715_), .Y(_103__10_) );
INVX1 INVX1_997 ( .gnd(gnd), .vdd(vdd), .A(data_192__11_), .Y(_1716_) );
OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf3), .C(_1716_), .Y(_1717_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_1694__bF_buf3), .Y(_1718_) );
AND2X2 AND2X2_476 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .B(_1717_), .Y(_103__11_) );
INVX1 INVX1_998 ( .gnd(gnd), .vdd(vdd), .A(data_192__12_), .Y(_1719_) );
OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_14882__bF_buf2), .C(_1719_), .Y(_1720_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_1694__bF_buf2), .Y(_1721_) );
AND2X2 AND2X2_477 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(_1720_), .Y(_103__12_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(data_192__13_), .B(_1694__bF_buf1), .Y(_1722_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_1694__bF_buf0), .C(_1722_), .Y(_103__13_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(data_192__14_), .B(_1694__bF_buf3), .Y(_1723_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_1694__bF_buf2), .C(_1723_), .Y(_103__14_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(data_192__15_), .B(_1694__bF_buf1), .Y(_1724_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_1694__bF_buf0), .C(_1724_), .Y(_103__15_) );
INVX1 INVX1_999 ( .gnd(gnd), .vdd(vdd), .A(data_191__0_), .Y(_1725_) );
OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf4), .B(_14975_), .C(_1036__bF_buf3), .Y(_1726_) );
OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_1562__bF_buf1), .C(_1726_), .Y(_1727_) );
INVX1 INVX1_1000 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .Y(_1728_) );
NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1728_), .C(_1335_), .Y(_1729_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1228_), .C(_1729_), .Y(_1730_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_1730_), .Y(_1731_) );
MUX2X1 MUX2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(_14932__bF_buf6), .S(_1731_), .Y(_102__0_) );
INVX1 INVX1_1001 ( .gnd(gnd), .vdd(vdd), .A(data_191__1_), .Y(_1732_) );
MUX2X1 MUX2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1732_), .B(_14894__bF_buf4), .S(_1731_), .Y(_102__1_) );
MUX2X1 MUX2X1_284 ( .gnd(gnd), .vdd(vdd), .A(data_191__2_), .B(IDATA_PROG_data_2_bF_buf2), .S(_1731_), .Y(_1733_) );
INVX1 INVX1_1002 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .Y(_102__2_) );
INVX1 INVX1_1003 ( .gnd(gnd), .vdd(vdd), .A(data_191__3_), .Y(_1734_) );
MUX2X1 MUX2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .B(_14899__bF_buf4), .S(_1731_), .Y(_102__3_) );
INVX1 INVX1_1004 ( .gnd(gnd), .vdd(vdd), .A(data_191__4_), .Y(_1735_) );
MUX2X1 MUX2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(_14902__bF_buf0), .S(_1731_), .Y(_102__4_) );
INVX1 INVX1_1005 ( .gnd(gnd), .vdd(vdd), .A(data_191__5_), .Y(_1736_) );
MUX2X1 MUX2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_14903__bF_buf1), .S(_1731_), .Y(_102__5_) );
MUX2X1 MUX2X1_288 ( .gnd(gnd), .vdd(vdd), .A(data_191__6_), .B(IDATA_PROG_data_6_bF_buf3), .S(_1731_), .Y(_1737_) );
INVX1 INVX1_1006 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .Y(_102__6_) );
INVX1 INVX1_1007 ( .gnd(gnd), .vdd(vdd), .A(data_191__7_), .Y(_1738_) );
MUX2X1 MUX2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1738_), .B(_14908__bF_buf0), .S(_1731_), .Y(_102__7_) );
MUX2X1 MUX2X1_290 ( .gnd(gnd), .vdd(vdd), .A(data_191__8_), .B(IDATA_PROG_data_8_bF_buf1), .S(_1731_), .Y(_1739_) );
INVX1 INVX1_1008 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .Y(_102__8_) );
MUX2X1 MUX2X1_291 ( .gnd(gnd), .vdd(vdd), .A(data_191__9_), .B(IDATA_PROG_data_9_bF_buf3), .S(_1731_), .Y(_1740_) );
INVX1 INVX1_1009 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .Y(_102__9_) );
MUX2X1 MUX2X1_292 ( .gnd(gnd), .vdd(vdd), .A(data_191__10_), .B(IDATA_PROG_data_10_bF_buf1), .S(_1731_), .Y(_1741_) );
INVX1 INVX1_1010 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .Y(_102__10_) );
INVX1 INVX1_1011 ( .gnd(gnd), .vdd(vdd), .A(data_191__11_), .Y(_1742_) );
MUX2X1 MUX2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1742_), .B(_14918__bF_buf1), .S(_1731_), .Y(_102__11_) );
INVX1 INVX1_1012 ( .gnd(gnd), .vdd(vdd), .A(data_191__12_), .Y(_1743_) );
MUX2X1 MUX2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(_14920__bF_buf1), .S(_1731_), .Y(_102__12_) );
MUX2X1 MUX2X1_295 ( .gnd(gnd), .vdd(vdd), .A(data_191__13_), .B(IDATA_PROG_data_13_bF_buf2), .S(_1731_), .Y(_1744_) );
INVX1 INVX1_1013 ( .gnd(gnd), .vdd(vdd), .A(_1744_), .Y(_102__13_) );
MUX2X1 MUX2X1_296 ( .gnd(gnd), .vdd(vdd), .A(data_191__14_), .B(IDATA_PROG_data_14_bF_buf2), .S(_1731_), .Y(_1745_) );
INVX1 INVX1_1014 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .Y(_102__14_) );
MUX2X1 MUX2X1_297 ( .gnd(gnd), .vdd(vdd), .A(data_191__15_), .B(IDATA_PROG_data_15_bF_buf4), .S(_1731_), .Y(_1746_) );
INVX1 INVX1_1015 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .Y(_102__15_) );
INVX1 INVX1_1016 ( .gnd(gnd), .vdd(vdd), .A(data_190__0_), .Y(_1747_) );
OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_1562__bF_buf0), .C(_1747_), .Y(_1748_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1562__bF_buf3), .B(_15788__bF_buf3), .Y(_1749_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_1749_), .Y(_1750_) );
AND2X2 AND2X2_478 ( .gnd(gnd), .vdd(vdd), .A(_1750_), .B(_1748_), .Y(_101__0_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_15793__bF_buf3), .Y(_1751_) );
INVX1 INVX1_1017 ( .gnd(gnd), .vdd(vdd), .A(data_190__1_), .Y(_1752_) );
OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_1562__bF_buf2), .C(_1752_), .Y(_1753_) );
OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf4), .B(_1751_), .C(_1753_), .Y(_1754_) );
INVX1 INVX1_1018 ( .gnd(gnd), .vdd(vdd), .A(_1754_), .Y(_101__1_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(data_190__2_), .B(_1749_), .Y(_1755_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_1749_), .C(_1755_), .Y(_101__2_) );
INVX1 INVX1_1019 ( .gnd(gnd), .vdd(vdd), .A(data_190__3_), .Y(_1756_) );
MUX2X1 MUX2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .B(_14899__bF_buf3), .S(_1751_), .Y(_101__3_) );
INVX1 INVX1_1020 ( .gnd(gnd), .vdd(vdd), .A(data_190__4_), .Y(_1757_) );
MUX2X1 MUX2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(_14902__bF_buf13), .S(_1751_), .Y(_101__4_) );
INVX1 INVX1_1021 ( .gnd(gnd), .vdd(vdd), .A(data_190__5_), .Y(_1758_) );
OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_1562__bF_buf1), .C(_1758_), .Y(_1759_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_1749_), .Y(_1760_) );
AND2X2 AND2X2_479 ( .gnd(gnd), .vdd(vdd), .A(_1760_), .B(_1759_), .Y(_101__5_) );
INVX1 INVX1_1022 ( .gnd(gnd), .vdd(vdd), .A(data_190__6_), .Y(_1761_) );
OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_1562__bF_buf0), .C(_1761_), .Y(_1762_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf0), .B(_1749_), .Y(_1763_) );
AND2X2 AND2X2_480 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(_1762_), .Y(_101__6_) );
INVX1 INVX1_1023 ( .gnd(gnd), .vdd(vdd), .A(data_190__7_), .Y(_1764_) );
MUX2X1 MUX2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1764_), .B(_14908__bF_buf13), .S(_1751_), .Y(_101__7_) );
INVX1 INVX1_1024 ( .gnd(gnd), .vdd(vdd), .A(data_190__8_), .Y(_1765_) );
OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_1562__bF_buf3), .C(_1765_), .Y(_1766_) );
OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf0), .B(_1751_), .C(_1766_), .Y(_1767_) );
INVX1 INVX1_1025 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .Y(_101__8_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(data_190__9_), .B(_1749_), .Y(_1768_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_1749_), .C(_1768_), .Y(_101__9_) );
INVX1 INVX1_1026 ( .gnd(gnd), .vdd(vdd), .A(data_190__10_), .Y(_1769_) );
OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_1562__bF_buf2), .C(_1769_), .Y(_1770_) );
OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf0), .B(_1751_), .C(_1770_), .Y(_1771_) );
INVX1 INVX1_1027 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .Y(_101__10_) );
INVX1 INVX1_1028 ( .gnd(gnd), .vdd(vdd), .A(data_190__11_), .Y(_1772_) );
OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_1562__bF_buf1), .C(_1772_), .Y(_1773_) );
OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf3), .B(_1751_), .C(_1773_), .Y(_1774_) );
INVX1 INVX1_1029 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .Y(_101__11_) );
INVX1 INVX1_1030 ( .gnd(gnd), .vdd(vdd), .A(data_190__12_), .Y(_1775_) );
MUX2X1 MUX2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1775_), .B(_14920__bF_buf0), .S(_1751_), .Y(_101__12_) );
INVX1 INVX1_1031 ( .gnd(gnd), .vdd(vdd), .A(data_190__13_), .Y(_1776_) );
OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_1562__bF_buf0), .C(_1776_), .Y(_1777_) );
OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf1), .B(_1751_), .C(_1777_), .Y(_1778_) );
INVX1 INVX1_1032 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .Y(_101__13_) );
INVX1 INVX1_1033 ( .gnd(gnd), .vdd(vdd), .A(data_190__14_), .Y(_1779_) );
OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_1562__bF_buf3), .C(_1779_), .Y(_1780_) );
NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_1561_), .C(_15793__bF_buf2), .Y(_1781_) );
AND2X2 AND2X2_481 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1781_), .Y(_101__14_) );
INVX1 INVX1_1034 ( .gnd(gnd), .vdd(vdd), .A(data_190__15_), .Y(_1782_) );
OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_1562__bF_buf2), .C(_1782_), .Y(_1783_) );
NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_1561_), .C(_15793__bF_buf1), .Y(_1784_) );
AND2X2 AND2X2_482 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1784_), .Y(_101__15_) );
INVX1 INVX1_1035 ( .gnd(gnd), .vdd(vdd), .A(data_189__0_), .Y(_1785_) );
INVX1 INVX1_1036 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .Y(_1786_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .B(_1000__bF_buf1), .Y(_1787_) );
OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_15025__bF_buf1), .C(_1563_), .Y(_1788_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_15078_), .C(_1788_), .Y(_1789_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_1787_), .Y(_1790_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1790_), .B(_1528__bF_buf0), .Y(_1791_) );
NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_1786_), .C(_1791_), .Y(_1792_) );
MUX2X1 MUX2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1785_), .B(_14932__bF_buf4), .S(_1792_), .Y(_99__0_) );
INVX1 INVX1_1037 ( .gnd(gnd), .vdd(vdd), .A(data_189__1_), .Y(_1793_) );
MUX2X1 MUX2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1793_), .B(_14894__bF_buf3), .S(_1792_), .Y(_99__1_) );
INVX1 INVX1_1038 ( .gnd(gnd), .vdd(vdd), .A(data_189__2_), .Y(_1794_) );
MUX2X1 MUX2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_14897__bF_buf13), .S(_1792_), .Y(_99__2_) );
INVX1 INVX1_1039 ( .gnd(gnd), .vdd(vdd), .A(data_189__3_), .Y(_1795_) );
MUX2X1 MUX2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1795_), .B(_14899__bF_buf2), .S(_1792_), .Y(_99__3_) );
INVX1 INVX1_1040 ( .gnd(gnd), .vdd(vdd), .A(data_189__4_), .Y(_1796_) );
MUX2X1 MUX2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1796_), .B(_14902__bF_buf12), .S(_1792_), .Y(_99__4_) );
INVX1 INVX1_1041 ( .gnd(gnd), .vdd(vdd), .A(data_189__5_), .Y(_1797_) );
MUX2X1 MUX2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1797_), .B(_14903__bF_buf13), .S(_1792_), .Y(_99__5_) );
INVX1 INVX1_1042 ( .gnd(gnd), .vdd(vdd), .A(data_189__6_), .Y(_1798_) );
MUX2X1 MUX2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_15049__bF_buf14), .S(_1792_), .Y(_99__6_) );
INVX1 INVX1_1043 ( .gnd(gnd), .vdd(vdd), .A(data_189__7_), .Y(_1799_) );
MUX2X1 MUX2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1799_), .B(_14908__bF_buf12), .S(_1792_), .Y(_99__7_) );
INVX1 INVX1_1044 ( .gnd(gnd), .vdd(vdd), .A(data_189__8_), .Y(_1800_) );
MUX2X1 MUX2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1800_), .B(_15052__bF_buf12), .S(_1792_), .Y(_99__8_) );
INVX1 INVX1_1045 ( .gnd(gnd), .vdd(vdd), .A(data_189__9_), .Y(_1801_) );
MUX2X1 MUX2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1801_), .B(_14913__bF_buf14), .S(_1792_), .Y(_99__9_) );
INVX1 INVX1_1046 ( .gnd(gnd), .vdd(vdd), .A(data_189__10_), .Y(_1802_) );
MUX2X1 MUX2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_15055__bF_buf12), .S(_1792_), .Y(_99__10_) );
INVX1 INVX1_1047 ( .gnd(gnd), .vdd(vdd), .A(data_189__11_), .Y(_1803_) );
MUX2X1 MUX2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_14918__bF_buf0), .S(_1792_), .Y(_99__11_) );
INVX1 INVX1_1048 ( .gnd(gnd), .vdd(vdd), .A(data_189__12_), .Y(_1804_) );
MUX2X1 MUX2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .B(_14920__bF_buf13), .S(_1792_), .Y(_99__12_) );
INVX1 INVX1_1049 ( .gnd(gnd), .vdd(vdd), .A(data_189__13_), .Y(_1805_) );
MUX2X1 MUX2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(_14924__bF_buf11), .S(_1792_), .Y(_99__13_) );
INVX1 INVX1_1050 ( .gnd(gnd), .vdd(vdd), .A(data_189__14_), .Y(_1806_) );
MUX2X1 MUX2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1806_), .B(_15060__bF_buf0), .S(_1792_), .Y(_99__14_) );
INVX1 INVX1_1051 ( .gnd(gnd), .vdd(vdd), .A(data_189__15_), .Y(_1807_) );
MUX2X1 MUX2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1807_), .B(_15062__bF_buf10), .S(_1792_), .Y(_99__15_) );
OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_1562__bF_buf1), .C(_1726_), .Y(_1808_) );
INVX1 INVX1_1052 ( .gnd(gnd), .vdd(vdd), .A(_1808_), .Y(_1809_) );
NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1786_), .B(_1809_), .C(_1692_), .Y(_1810_) );
OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf1), .B(_14957_), .C(_1561_), .Y(_1811_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_15082_), .B(_1228_), .Y(_1812_) );
INVX1 INVX1_1053 ( .gnd(gnd), .vdd(vdd), .A(_1812__bF_buf3), .Y(_1813_) );
NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1811_), .B(_1813_), .C(_1525__bF_buf4), .Y(_1814_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .B(_1810__bF_buf7), .Y(_1815_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(data_188__0_), .B(_1815__bF_buf3), .Y(_1816_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_1815__bF_buf2), .C(_1816_), .Y(_98__0_) );
INVX1 INVX1_1054 ( .gnd(gnd), .vdd(vdd), .A(data_188__1_), .Y(_1817_) );
MUX2X1 MUX2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_1817_), .S(_1815__bF_buf1), .Y(_98__1_) );
INVX1 INVX1_1055 ( .gnd(gnd), .vdd(vdd), .A(data_188__2_), .Y(_1818_) );
MUX2X1 MUX2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf12), .B(_1818_), .S(_1815__bF_buf0), .Y(_98__2_) );
INVX1 INVX1_1056 ( .gnd(gnd), .vdd(vdd), .A(data_188__3_), .Y(_1819_) );
MUX2X1 MUX2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_1819_), .S(_1815__bF_buf3), .Y(_98__3_) );
INVX1 INVX1_1057 ( .gnd(gnd), .vdd(vdd), .A(data_188__4_), .Y(_1820_) );
MUX2X1 MUX2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_1820_), .S(_1815__bF_buf2), .Y(_98__4_) );
INVX1 INVX1_1058 ( .gnd(gnd), .vdd(vdd), .A(data_188__5_), .Y(_1821_) );
MUX2X1 MUX2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_1821_), .S(_1815__bF_buf1), .Y(_98__5_) );
INVX1 INVX1_1059 ( .gnd(gnd), .vdd(vdd), .A(data_188__6_), .Y(_1822_) );
MUX2X1 MUX2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_1822_), .S(_1815__bF_buf0), .Y(_98__6_) );
INVX1 INVX1_1060 ( .gnd(gnd), .vdd(vdd), .A(data_188__7_), .Y(_1823_) );
MUX2X1 MUX2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_1823_), .S(_1815__bF_buf3), .Y(_98__7_) );
INVX1 INVX1_1061 ( .gnd(gnd), .vdd(vdd), .A(data_188__8_), .Y(_1824_) );
MUX2X1 MUX2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_1824_), .S(_1815__bF_buf2), .Y(_98__8_) );
INVX1 INVX1_1062 ( .gnd(gnd), .vdd(vdd), .A(data_188__9_), .Y(_1825_) );
MUX2X1 MUX2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_1825_), .S(_1815__bF_buf1), .Y(_98__9_) );
INVX1 INVX1_1063 ( .gnd(gnd), .vdd(vdd), .A(data_188__10_), .Y(_1826_) );
MUX2X1 MUX2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_1826_), .S(_1815__bF_buf0), .Y(_98__10_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(data_188__11_), .B(_1815__bF_buf3), .Y(_1827_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_1815__bF_buf2), .C(_1827_), .Y(_98__11_) );
INVX1 INVX1_1064 ( .gnd(gnd), .vdd(vdd), .A(data_188__12_), .Y(_1828_) );
MUX2X1 MUX2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_1828_), .S(_1815__bF_buf1), .Y(_98__12_) );
INVX1 INVX1_1065 ( .gnd(gnd), .vdd(vdd), .A(data_188__13_), .Y(_1829_) );
MUX2X1 MUX2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_1829_), .S(_1815__bF_buf0), .Y(_98__13_) );
INVX1 INVX1_1066 ( .gnd(gnd), .vdd(vdd), .A(data_188__14_), .Y(_1830_) );
MUX2X1 MUX2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf14), .B(_1830_), .S(_1815__bF_buf3), .Y(_98__14_) );
INVX1 INVX1_1067 ( .gnd(gnd), .vdd(vdd), .A(data_188__15_), .Y(_1831_) );
MUX2X1 MUX2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_1831_), .S(_1815__bF_buf2), .Y(_98__15_) );
NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1726_), .C(_1228_), .Y(_1832_) );
NOR3X1 NOR3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1832_), .C(_1266__bF_buf0), .Y(_1833_) );
NOR3X1 NOR3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1808_), .C(_1833_), .Y(_1834_) );
OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_1562__bF_buf0), .B(_15160_), .C(IDATA_PROG_write_bF_buf1), .Y(_1835_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_15951_), .C(_1835_), .Y(_1836_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1836_), .B(_1787_), .Y(_1837_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_1528__bF_buf5), .Y(_1838_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__0_), .Y(_1839_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_1528__bF_buf4), .B(_1837_), .Y(_1840_) );
NOR3X1 NOR3X1_75 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf2), .B(_1840_), .C(_1810__bF_buf6), .Y(_1841_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1841_), .Y(_97__0_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__1_), .Y(_1842_) );
NOR3X1 NOR3X1_76 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf3), .B(_1840_), .C(_1810__bF_buf5), .Y(_1843_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_1843_), .Y(_97__1_) );
INVX1 INVX1_1068 ( .gnd(gnd), .vdd(vdd), .A(data_187__2_), .Y(_1844_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1840_), .B(_1810__bF_buf4), .Y(_1845_) );
MUX2X1 MUX2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_1844_), .S(_1845_), .Y(_97__2_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__3_), .Y(_1846_) );
NOR3X1 NOR3X1_77 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf4), .B(_1840_), .C(_1810__bF_buf3), .Y(_1847_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1846_), .B(_1847_), .Y(_97__3_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__4_), .Y(_1848_) );
NOR3X1 NOR3X1_78 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf4), .B(_1840_), .C(_1810__bF_buf2), .Y(_1849_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1849_), .Y(_97__4_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__5_), .Y(_1850_) );
NOR3X1 NOR3X1_79 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf3), .B(_1840_), .C(_1810__bF_buf1), .Y(_1851_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1851_), .Y(_97__5_) );
INVX1 INVX1_1069 ( .gnd(gnd), .vdd(vdd), .A(data_187__6_), .Y(_1852_) );
MUX2X1 MUX2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_1852_), .S(_1845_), .Y(_97__6_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__7_), .Y(_1853_) );
NOR3X1 NOR3X1_80 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf1), .B(_1840_), .C(_1810__bF_buf0), .Y(_1854_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_1854_), .Y(_97__7_) );
INVX1 INVX1_1070 ( .gnd(gnd), .vdd(vdd), .A(data_187__8_), .Y(_1855_) );
MUX2X1 MUX2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_1855_), .S(_1845_), .Y(_97__8_) );
INVX1 INVX1_1071 ( .gnd(gnd), .vdd(vdd), .A(data_187__9_), .Y(_1856_) );
MUX2X1 MUX2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_1856_), .S(_1845_), .Y(_97__9_) );
INVX1 INVX1_1072 ( .gnd(gnd), .vdd(vdd), .A(data_187__10_), .Y(_1857_) );
MUX2X1 MUX2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_1857_), .S(_1845_), .Y(_97__10_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__11_), .Y(_1858_) );
NOR3X1 NOR3X1_81 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf2), .B(_1840_), .C(_1810__bF_buf7), .Y(_1859_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1858_), .B(_1859_), .Y(_97__11_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1838_), .B(_1834_), .C(data_187__12_), .Y(_1860_) );
NOR3X1 NOR3X1_82 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf3), .B(_1840_), .C(_1810__bF_buf6), .Y(_1861_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_1861_), .Y(_97__12_) );
INVX1 INVX1_1073 ( .gnd(gnd), .vdd(vdd), .A(data_187__13_), .Y(_1862_) );
MUX2X1 MUX2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_1862_), .S(_1845_), .Y(_97__13_) );
INVX1 INVX1_1074 ( .gnd(gnd), .vdd(vdd), .A(data_187__14_), .Y(_1863_) );
MUX2X1 MUX2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_1863_), .S(_1845_), .Y(_97__14_) );
INVX1 INVX1_1075 ( .gnd(gnd), .vdd(vdd), .A(data_187__15_), .Y(_1864_) );
MUX2X1 MUX2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_1864_), .S(_1845_), .Y(_97__15_) );
INVX1 INVX1_1076 ( .gnd(gnd), .vdd(vdd), .A(data_186__0_), .Y(_1865_) );
OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14884_), .C(IDATA_PROG_write_bF_buf0), .Y(_1866_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .Y(_1867_) );
OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14952__bF_buf0), .C(_1561_), .Y(_1868_) );
OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_1867_), .C(_1868_), .Y(_1869_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1869_), .B(_1604_), .Y(_1870_) );
NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_1870_), .C(_1525__bF_buf3), .Y(_1871_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1871_), .B(_1810__bF_buf5), .Y(_1872_) );
MUX2X1 MUX2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_1865_), .S(_1872_), .Y(_96__0_) );
INVX1 INVX1_1077 ( .gnd(gnd), .vdd(vdd), .A(data_186__1_), .Y(_1873_) );
MUX2X1 MUX2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_1873_), .S(_1872_), .Y(_96__1_) );
INVX1 INVX1_1078 ( .gnd(gnd), .vdd(vdd), .A(data_186__2_), .Y(_1874_) );
MUX2X1 MUX2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_1874_), .S(_1872_), .Y(_96__2_) );
INVX1 INVX1_1079 ( .gnd(gnd), .vdd(vdd), .A(data_186__3_), .Y(_1875_) );
MUX2X1 MUX2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_1875_), .S(_1872_), .Y(_96__3_) );
INVX1 INVX1_1080 ( .gnd(gnd), .vdd(vdd), .A(data_186__4_), .Y(_1876_) );
MUX2X1 MUX2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_1876_), .S(_1872_), .Y(_96__4_) );
INVX1 INVX1_1081 ( .gnd(gnd), .vdd(vdd), .A(data_186__5_), .Y(_1877_) );
MUX2X1 MUX2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_1877_), .S(_1872_), .Y(_96__5_) );
INVX1 INVX1_1082 ( .gnd(gnd), .vdd(vdd), .A(data_186__6_), .Y(_1878_) );
MUX2X1 MUX2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_1878_), .S(_1872_), .Y(_96__6_) );
INVX1 INVX1_1083 ( .gnd(gnd), .vdd(vdd), .A(data_186__7_), .Y(_1879_) );
MUX2X1 MUX2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_1879_), .S(_1872_), .Y(_96__7_) );
INVX1 INVX1_1084 ( .gnd(gnd), .vdd(vdd), .A(data_186__8_), .Y(_1880_) );
MUX2X1 MUX2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_1880_), .S(_1872_), .Y(_96__8_) );
INVX1 INVX1_1085 ( .gnd(gnd), .vdd(vdd), .A(data_186__9_), .Y(_1881_) );
MUX2X1 MUX2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_1881_), .S(_1872_), .Y(_96__9_) );
INVX1 INVX1_1086 ( .gnd(gnd), .vdd(vdd), .A(data_186__10_), .Y(_1882_) );
MUX2X1 MUX2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_1882_), .S(_1872_), .Y(_96__10_) );
INVX1 INVX1_1087 ( .gnd(gnd), .vdd(vdd), .A(data_186__11_), .Y(_1883_) );
MUX2X1 MUX2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_1883_), .S(_1872_), .Y(_96__11_) );
INVX1 INVX1_1088 ( .gnd(gnd), .vdd(vdd), .A(data_186__12_), .Y(_1884_) );
MUX2X1 MUX2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_1884_), .S(_1872_), .Y(_96__12_) );
INVX1 INVX1_1089 ( .gnd(gnd), .vdd(vdd), .A(data_186__13_), .Y(_1885_) );
MUX2X1 MUX2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_1885_), .S(_1872_), .Y(_96__13_) );
INVX1 INVX1_1090 ( .gnd(gnd), .vdd(vdd), .A(data_186__14_), .Y(_1886_) );
MUX2X1 MUX2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_1886_), .S(_1872_), .Y(_96__14_) );
INVX1 INVX1_1091 ( .gnd(gnd), .vdd(vdd), .A(data_186__15_), .Y(_1887_) );
MUX2X1 MUX2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_1887_), .S(_1872_), .Y(_96__15_) );
INVX1 INVX1_1092 ( .gnd(gnd), .vdd(vdd), .A(data_185__0_), .Y(_1888_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .B(_1528__bF_buf3), .Y(_1889_) );
OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_1867_), .C(_1889_), .Y(_1890_) );
OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf3), .B(_1810__bF_buf4), .C(_1888_), .Y(_1891_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1810__bF_buf3), .B(_1890__bF_buf2), .Y(_1892_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_1892_), .Y(_1893_) );
AND2X2 AND2X2_483 ( .gnd(gnd), .vdd(vdd), .A(_1893_), .B(_1891_), .Y(_95__0_) );
INVX1 INVX1_1093 ( .gnd(gnd), .vdd(vdd), .A(data_185__1_), .Y(_1894_) );
OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf1), .B(_1810__bF_buf2), .C(_1894_), .Y(_1895_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_1892_), .Y(_1896_) );
AND2X2 AND2X2_484 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(_1895_), .Y(_95__1_) );
INVX1 INVX1_1094 ( .gnd(gnd), .vdd(vdd), .A(data_185__2_), .Y(_1897_) );
OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf0), .B(_1810__bF_buf1), .C(_1897_), .Y(_1898_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_1892_), .Y(_1899_) );
AND2X2 AND2X2_485 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .B(_1898_), .Y(_95__2_) );
INVX1 INVX1_1095 ( .gnd(gnd), .vdd(vdd), .A(data_185__3_), .Y(_1900_) );
OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf3), .B(_1810__bF_buf0), .C(_1900_), .Y(_1901_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_1892_), .Y(_1902_) );
AND2X2 AND2X2_486 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .B(_1901_), .Y(_95__3_) );
INVX1 INVX1_1096 ( .gnd(gnd), .vdd(vdd), .A(data_185__4_), .Y(_1903_) );
OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf2), .B(_1810__bF_buf7), .C(_1903_), .Y(_1904_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_1892_), .Y(_1905_) );
AND2X2 AND2X2_487 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_1904_), .Y(_95__4_) );
INVX1 INVX1_1097 ( .gnd(gnd), .vdd(vdd), .A(data_185__5_), .Y(_1906_) );
OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf1), .B(_1810__bF_buf6), .C(_1906_), .Y(_1907_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_1892_), .Y(_1908_) );
AND2X2 AND2X2_488 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_1907_), .Y(_95__5_) );
INVX1 INVX1_1098 ( .gnd(gnd), .vdd(vdd), .A(data_185__6_), .Y(_1909_) );
OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf0), .B(_1810__bF_buf5), .C(_1909_), .Y(_1910_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_1892_), .Y(_1911_) );
AND2X2 AND2X2_489 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .B(_1910_), .Y(_95__6_) );
INVX1 INVX1_1099 ( .gnd(gnd), .vdd(vdd), .A(data_185__7_), .Y(_1912_) );
OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf3), .B(_1810__bF_buf4), .C(_1912_), .Y(_1913_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_1892_), .Y(_1914_) );
AND2X2 AND2X2_490 ( .gnd(gnd), .vdd(vdd), .A(_1914_), .B(_1913_), .Y(_95__7_) );
INVX1 INVX1_1100 ( .gnd(gnd), .vdd(vdd), .A(data_185__8_), .Y(_1915_) );
OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf2), .B(_1810__bF_buf3), .C(_1915_), .Y(_1916_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_1892_), .Y(_1917_) );
AND2X2 AND2X2_491 ( .gnd(gnd), .vdd(vdd), .A(_1917_), .B(_1916_), .Y(_95__8_) );
INVX1 INVX1_1101 ( .gnd(gnd), .vdd(vdd), .A(data_185__9_), .Y(_1918_) );
OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf1), .B(_1810__bF_buf2), .C(_1918_), .Y(_1919_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_1892_), .Y(_1920_) );
AND2X2 AND2X2_492 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_1919_), .Y(_95__9_) );
INVX1 INVX1_1102 ( .gnd(gnd), .vdd(vdd), .A(data_185__10_), .Y(_1921_) );
OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf0), .B(_1810__bF_buf1), .C(_1921_), .Y(_1922_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_1892_), .Y(_1923_) );
AND2X2 AND2X2_493 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_1922_), .Y(_95__10_) );
INVX1 INVX1_1103 ( .gnd(gnd), .vdd(vdd), .A(data_185__11_), .Y(_1924_) );
OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf3), .B(_1810__bF_buf0), .C(_1924_), .Y(_1925_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_1892_), .Y(_1926_) );
AND2X2 AND2X2_494 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_1925_), .Y(_95__11_) );
INVX1 INVX1_1104 ( .gnd(gnd), .vdd(vdd), .A(data_185__12_), .Y(_1927_) );
OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf2), .B(_1810__bF_buf7), .C(_1927_), .Y(_1928_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_1892_), .Y(_1929_) );
AND2X2 AND2X2_495 ( .gnd(gnd), .vdd(vdd), .A(_1929_), .B(_1928_), .Y(_95__12_) );
INVX1 INVX1_1105 ( .gnd(gnd), .vdd(vdd), .A(data_185__13_), .Y(_1930_) );
OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf1), .B(_1810__bF_buf6), .C(_1930_), .Y(_1931_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_1892_), .Y(_1932_) );
AND2X2 AND2X2_496 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1931_), .Y(_95__13_) );
INVX1 INVX1_1106 ( .gnd(gnd), .vdd(vdd), .A(data_185__14_), .Y(_1933_) );
OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf0), .B(_1810__bF_buf5), .C(_1933_), .Y(_1934_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_1892_), .Y(_1935_) );
AND2X2 AND2X2_497 ( .gnd(gnd), .vdd(vdd), .A(_1935_), .B(_1934_), .Y(_95__14_) );
INVX1 INVX1_1107 ( .gnd(gnd), .vdd(vdd), .A(data_185__15_), .Y(_1936_) );
OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_1890__bF_buf3), .B(_1810__bF_buf4), .C(_1936_), .Y(_1937_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_1892_), .Y(_1938_) );
AND2X2 AND2X2_498 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1937_), .Y(_95__15_) );
INVX1 INVX1_1108 ( .gnd(gnd), .vdd(vdd), .A(data_184__0_), .Y(_1939_) );
OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf2), .B(_14952__bF_buf4), .C(_1561_), .Y(_1940_) );
NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1813_), .B(_1940_), .C(_1525__bF_buf2), .Y(_1941_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_1810__bF_buf3), .Y(_1942_) );
MUX2X1 MUX2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_1939_), .S(_1942__bF_buf3), .Y(_94__0_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(data_184__1_), .B(_1942__bF_buf2), .Y(_1943_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_1942__bF_buf1), .C(_1943_), .Y(_94__1_) );
INVX1 INVX1_1109 ( .gnd(gnd), .vdd(vdd), .A(data_184__2_), .Y(_1944_) );
MUX2X1 MUX2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_1944_), .S(_1942__bF_buf0), .Y(_94__2_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(data_184__3_), .B(_1942__bF_buf3), .Y(_1945_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_1942__bF_buf2), .C(_1945_), .Y(_94__3_) );
NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(data_184__4_), .B(_1942__bF_buf1), .Y(_1946_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_1942__bF_buf0), .C(_1946_), .Y(_94__4_) );
NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(data_184__5_), .B(_1942__bF_buf3), .Y(_1947_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_1942__bF_buf2), .C(_1947_), .Y(_94__5_) );
INVX1 INVX1_1110 ( .gnd(gnd), .vdd(vdd), .A(data_184__6_), .Y(_1948_) );
MUX2X1 MUX2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_1948_), .S(_1942__bF_buf1), .Y(_94__6_) );
NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(data_184__7_), .B(_1942__bF_buf0), .Y(_1949_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_1942__bF_buf3), .C(_1949_), .Y(_94__7_) );
INVX1 INVX1_1111 ( .gnd(gnd), .vdd(vdd), .A(data_184__8_), .Y(_1950_) );
MUX2X1 MUX2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_1950_), .S(_1942__bF_buf2), .Y(_94__8_) );
INVX1 INVX1_1112 ( .gnd(gnd), .vdd(vdd), .A(data_184__9_), .Y(_1951_) );
MUX2X1 MUX2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_1951_), .S(_1942__bF_buf1), .Y(_94__9_) );
INVX1 INVX1_1113 ( .gnd(gnd), .vdd(vdd), .A(data_184__10_), .Y(_1952_) );
MUX2X1 MUX2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_1952_), .S(_1942__bF_buf0), .Y(_94__10_) );
INVX1 INVX1_1114 ( .gnd(gnd), .vdd(vdd), .A(data_184__11_), .Y(_1953_) );
MUX2X1 MUX2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_1953_), .S(_1942__bF_buf3), .Y(_94__11_) );
NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(data_184__12_), .B(_1942__bF_buf2), .Y(_1954_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_1942__bF_buf1), .C(_1954_), .Y(_94__12_) );
INVX1 INVX1_1115 ( .gnd(gnd), .vdd(vdd), .A(data_184__13_), .Y(_1955_) );
MUX2X1 MUX2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_1955_), .S(_1942__bF_buf0), .Y(_94__13_) );
INVX1 INVX1_1116 ( .gnd(gnd), .vdd(vdd), .A(data_184__14_), .Y(_1956_) );
MUX2X1 MUX2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_1956_), .S(_1942__bF_buf3), .Y(_94__14_) );
INVX1 INVX1_1117 ( .gnd(gnd), .vdd(vdd), .A(data_184__15_), .Y(_1957_) );
MUX2X1 MUX2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_1957_), .S(_1942__bF_buf2), .Y(_94__15_) );
INVX1 INVX1_1118 ( .gnd(gnd), .vdd(vdd), .A(data_183__0_), .Y(_1958_) );
OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_1867_), .C(_1889_), .Y(_1959_) );
NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1810__bF_buf2), .B(_1959_), .Y(_1960_) );
MUX2X1 MUX2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_1958_), .S(_1960_), .Y(_93__0_) );
INVX1 INVX1_1119 ( .gnd(gnd), .vdd(vdd), .A(data_183__1_), .Y(_1961_) );
MUX2X1 MUX2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_1961_), .S(_1960_), .Y(_93__1_) );
INVX1 INVX1_1120 ( .gnd(gnd), .vdd(vdd), .A(data_183__2_), .Y(_1962_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .B(_1810__bF_buf1), .Y(_1963_) );
NOR3X1 NOR3X1_83 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf1), .B(_1810__bF_buf0), .C(_1959_), .Y(_1964_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(_1963_), .C(_1964_), .Y(_93__2_) );
INVX1 INVX1_1121 ( .gnd(gnd), .vdd(vdd), .A(data_183__3_), .Y(_1965_) );
MUX2X1 MUX2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_1965_), .S(_1960_), .Y(_93__3_) );
INVX1 INVX1_1122 ( .gnd(gnd), .vdd(vdd), .A(data_183__4_), .Y(_1966_) );
MUX2X1 MUX2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_1966_), .S(_1960_), .Y(_93__4_) );
INVX1 INVX1_1123 ( .gnd(gnd), .vdd(vdd), .A(data_183__5_), .Y(_1967_) );
MUX2X1 MUX2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_1967_), .S(_1960_), .Y(_93__5_) );
INVX1 INVX1_1124 ( .gnd(gnd), .vdd(vdd), .A(data_183__6_), .Y(_1968_) );
NOR3X1 NOR3X1_84 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf2), .B(_1810__bF_buf7), .C(_1959_), .Y(_1969_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1968_), .B(_1963_), .C(_1969_), .Y(_93__6_) );
INVX1 INVX1_1125 ( .gnd(gnd), .vdd(vdd), .A(data_183__7_), .Y(_1970_) );
MUX2X1 MUX2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_1970_), .S(_1960_), .Y(_93__7_) );
INVX1 INVX1_1126 ( .gnd(gnd), .vdd(vdd), .A(data_183__8_), .Y(_1971_) );
OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .B(_1810__bF_buf6), .C(_1971_), .Y(_1972_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_1960_), .Y(_1973_) );
AND2X2 AND2X2_499 ( .gnd(gnd), .vdd(vdd), .A(_1973_), .B(_1972_), .Y(_93__8_) );
INVX1 INVX1_1127 ( .gnd(gnd), .vdd(vdd), .A(data_183__9_), .Y(_1974_) );
NOR3X1 NOR3X1_85 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf2), .B(_1810__bF_buf5), .C(_1959_), .Y(_1975_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1974_), .B(_1963_), .C(_1975_), .Y(_93__9_) );
INVX1 INVX1_1128 ( .gnd(gnd), .vdd(vdd), .A(data_183__10_), .Y(_1976_) );
NOR3X1 NOR3X1_86 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf4), .B(_1810__bF_buf4), .C(_1959_), .Y(_1977_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_1963_), .C(_1977_), .Y(_93__10_) );
INVX1 INVX1_1129 ( .gnd(gnd), .vdd(vdd), .A(data_183__11_), .Y(_1978_) );
OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .B(_1810__bF_buf3), .C(_1978_), .Y(_1979_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_1960_), .Y(_1980_) );
AND2X2 AND2X2_500 ( .gnd(gnd), .vdd(vdd), .A(_1980_), .B(_1979_), .Y(_93__11_) );
INVX1 INVX1_1130 ( .gnd(gnd), .vdd(vdd), .A(data_183__12_), .Y(_1981_) );
MUX2X1 MUX2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_1981_), .S(_1960_), .Y(_93__12_) );
INVX1 INVX1_1131 ( .gnd(gnd), .vdd(vdd), .A(data_183__13_), .Y(_1982_) );
NOR3X1 NOR3X1_87 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf0), .B(_1810__bF_buf2), .C(_1959_), .Y(_1983_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1982_), .B(_1963_), .C(_1983_), .Y(_93__13_) );
INVX1 INVX1_1132 ( .gnd(gnd), .vdd(vdd), .A(data_183__14_), .Y(_1984_) );
NOR3X1 NOR3X1_88 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf1), .B(_1810__bF_buf1), .C(_1959_), .Y(_1985_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1984_), .B(_1963_), .C(_1985_), .Y(_93__14_) );
INVX1 INVX1_1133 ( .gnd(gnd), .vdd(vdd), .A(data_183__15_), .Y(_1986_) );
NOR3X1 NOR3X1_89 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf3), .B(_1810__bF_buf0), .C(_1959_), .Y(_1987_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_1963_), .C(_1987_), .Y(_93__15_) );
INVX1 INVX1_1134 ( .gnd(gnd), .vdd(vdd), .A(data_182__0_), .Y(_1988_) );
OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(_14977__bF_buf1), .C(_15509_), .Y(_1989_) );
OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_1989_), .B(_16204_), .C(_1866_), .Y(_1990_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1889_), .Y(_1991_) );
NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1810__bF_buf7), .B(_1991_), .Y(_1992_) );
MUX2X1 MUX2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_1988_), .S(_1992_), .Y(_92__0_) );
INVX1 INVX1_1135 ( .gnd(gnd), .vdd(vdd), .A(data_182__1_), .Y(_1993_) );
OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf6), .C(_1993_), .Y(_1994_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_1992_), .Y(_1995_) );
AND2X2 AND2X2_501 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .B(_1994_), .Y(_92__1_) );
INVX1 INVX1_1136 ( .gnd(gnd), .vdd(vdd), .A(data_182__2_), .Y(_1996_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf5), .Y(_1997_) );
NOR3X1 NOR3X1_90 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf0), .B(_1810__bF_buf4), .C(_1991_), .Y(_1998_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_1997_), .C(_1998_), .Y(_92__2_) );
INVX1 INVX1_1137 ( .gnd(gnd), .vdd(vdd), .A(data_182__3_), .Y(_1999_) );
MUX2X1 MUX2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_1999_), .S(_1992_), .Y(_92__3_) );
INVX1 INVX1_1138 ( .gnd(gnd), .vdd(vdd), .A(data_182__4_), .Y(_2000_) );
OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf3), .C(_2000_), .Y(_2001_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_1992_), .Y(_2002_) );
AND2X2 AND2X2_502 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2001_), .Y(_92__4_) );
INVX1 INVX1_1139 ( .gnd(gnd), .vdd(vdd), .A(data_182__5_), .Y(_2003_) );
OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf2), .C(_2003_), .Y(_2004_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_1992_), .Y(_2005_) );
AND2X2 AND2X2_503 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .B(_2004_), .Y(_92__5_) );
INVX1 INVX1_1140 ( .gnd(gnd), .vdd(vdd), .A(data_182__6_), .Y(_2006_) );
NOR3X1 NOR3X1_91 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf1), .B(_1810__bF_buf1), .C(_1991_), .Y(_2007_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_1997_), .C(_2007_), .Y(_92__6_) );
INVX1 INVX1_1141 ( .gnd(gnd), .vdd(vdd), .A(data_182__7_), .Y(_2008_) );
OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf0), .C(_2008_), .Y(_2009_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_1992_), .Y(_2010_) );
AND2X2 AND2X2_504 ( .gnd(gnd), .vdd(vdd), .A(_2010_), .B(_2009_), .Y(_92__7_) );
INVX1 INVX1_1142 ( .gnd(gnd), .vdd(vdd), .A(data_182__8_), .Y(_2011_) );
NOR3X1 NOR3X1_92 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf4), .B(_1810__bF_buf7), .C(_1991_), .Y(_2012_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_2011_), .B(_1997_), .C(_2012_), .Y(_92__8_) );
INVX1 INVX1_1143 ( .gnd(gnd), .vdd(vdd), .A(data_182__9_), .Y(_2013_) );
OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf6), .C(_2013_), .Y(_2014_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_1992_), .Y(_2015_) );
AND2X2 AND2X2_505 ( .gnd(gnd), .vdd(vdd), .A(_2015_), .B(_2014_), .Y(_92__9_) );
INVX1 INVX1_1144 ( .gnd(gnd), .vdd(vdd), .A(data_182__10_), .Y(_2016_) );
OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf5), .C(_2016_), .Y(_2017_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_1992_), .Y(_2018_) );
AND2X2 AND2X2_506 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .B(_2017_), .Y(_92__10_) );
INVX1 INVX1_1145 ( .gnd(gnd), .vdd(vdd), .A(data_182__11_), .Y(_2019_) );
MUX2X1 MUX2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_2019_), .S(_1992_), .Y(_92__11_) );
INVX1 INVX1_1146 ( .gnd(gnd), .vdd(vdd), .A(data_182__12_), .Y(_2020_) );
MUX2X1 MUX2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_2020_), .S(_1992_), .Y(_92__12_) );
INVX1 INVX1_1147 ( .gnd(gnd), .vdd(vdd), .A(data_182__13_), .Y(_2021_) );
OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf4), .C(_2021_), .Y(_2022_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_1992_), .Y(_2023_) );
AND2X2 AND2X2_507 ( .gnd(gnd), .vdd(vdd), .A(_2023_), .B(_2022_), .Y(_92__13_) );
INVX1 INVX1_1148 ( .gnd(gnd), .vdd(vdd), .A(data_182__14_), .Y(_2024_) );
NOR3X1 NOR3X1_93 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf0), .B(_1810__bF_buf3), .C(_1991_), .Y(_2025_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_1997_), .C(_2025_), .Y(_92__14_) );
INVX1 INVX1_1149 ( .gnd(gnd), .vdd(vdd), .A(data_182__15_), .Y(_2026_) );
OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_1991_), .B(_1810__bF_buf2), .C(_2026_), .Y(_2027_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_1992_), .Y(_2028_) );
AND2X2 AND2X2_508 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_2027_), .Y(_92__15_) );
INVX1 INVX1_1150 ( .gnd(gnd), .vdd(vdd), .A(data_181__0_), .Y(_2029_) );
NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_16204_), .B(_911_), .Y(_2030_) );
OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_2030_), .C(_1889_), .Y(_2031_) );
OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_1810__bF_buf1), .C(_2029_), .Y(_2032_) );
NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1810__bF_buf0), .B(_2031_), .Y(_2033_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_2033_), .Y(_2034_) );
AND2X2 AND2X2_509 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .B(_2032_), .Y(_91__0_) );
INVX1 INVX1_1151 ( .gnd(gnd), .vdd(vdd), .A(data_181__1_), .Y(_2035_) );
MUX2X1 MUX2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_2035_), .S(_2033_), .Y(_91__1_) );
INVX1 INVX1_1152 ( .gnd(gnd), .vdd(vdd), .A(data_181__2_), .Y(_2036_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_1810__bF_buf7), .Y(_2037_) );
NOR3X1 NOR3X1_94 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf3), .B(_1810__bF_buf6), .C(_2031_), .Y(_2038_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_2037_), .C(_2038_), .Y(_91__2_) );
INVX1 INVX1_1153 ( .gnd(gnd), .vdd(vdd), .A(data_181__3_), .Y(_2039_) );
MUX2X1 MUX2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_2039_), .S(_2033_), .Y(_91__3_) );
INVX1 INVX1_1154 ( .gnd(gnd), .vdd(vdd), .A(data_181__4_), .Y(_2040_) );
MUX2X1 MUX2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_2040_), .S(_2033_), .Y(_91__4_) );
INVX1 INVX1_1155 ( .gnd(gnd), .vdd(vdd), .A(data_181__5_), .Y(_2041_) );
MUX2X1 MUX2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_2041_), .S(_2033_), .Y(_91__5_) );
INVX1 INVX1_1156 ( .gnd(gnd), .vdd(vdd), .A(data_181__6_), .Y(_2042_) );
OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_1810__bF_buf5), .C(_2042_), .Y(_2043_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_2033_), .Y(_2044_) );
AND2X2 AND2X2_510 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(_2043_), .Y(_91__6_) );
INVX1 INVX1_1157 ( .gnd(gnd), .vdd(vdd), .A(data_181__7_), .Y(_2045_) );
MUX2X1 MUX2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_2045_), .S(_2033_), .Y(_91__7_) );
INVX1 INVX1_1158 ( .gnd(gnd), .vdd(vdd), .A(data_181__8_), .Y(_2046_) );
NOR3X1 NOR3X1_95 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf3), .B(_1810__bF_buf4), .C(_2031_), .Y(_2047_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(_2037_), .C(_2047_), .Y(_91__8_) );
INVX1 INVX1_1159 ( .gnd(gnd), .vdd(vdd), .A(data_181__9_), .Y(_2048_) );
NOR3X1 NOR3X1_96 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf1), .B(_1810__bF_buf3), .C(_2031_), .Y(_2049_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(_2037_), .C(_2049_), .Y(_91__9_) );
INVX1 INVX1_1160 ( .gnd(gnd), .vdd(vdd), .A(data_181__10_), .Y(_2050_) );
NOR3X1 NOR3X1_97 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf3), .B(_1810__bF_buf2), .C(_2031_), .Y(_2051_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(_2037_), .C(_2051_), .Y(_91__10_) );
INVX1 INVX1_1161 ( .gnd(gnd), .vdd(vdd), .A(data_181__11_), .Y(_2052_) );
MUX2X1 MUX2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_2052_), .S(_2033_), .Y(_91__11_) );
INVX1 INVX1_1162 ( .gnd(gnd), .vdd(vdd), .A(data_181__12_), .Y(_2053_) );
MUX2X1 MUX2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_2053_), .S(_2033_), .Y(_91__12_) );
INVX1 INVX1_1163 ( .gnd(gnd), .vdd(vdd), .A(data_181__13_), .Y(_2054_) );
NOR3X1 NOR3X1_98 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf4), .B(_1810__bF_buf1), .C(_2031_), .Y(_2055_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2037_), .C(_2055_), .Y(_91__13_) );
INVX1 INVX1_1164 ( .gnd(gnd), .vdd(vdd), .A(data_181__14_), .Y(_2056_) );
NOR3X1 NOR3X1_99 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf4), .B(_1810__bF_buf0), .C(_2031_), .Y(_2057_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .B(_2037_), .C(_2057_), .Y(_91__14_) );
INVX1 INVX1_1165 ( .gnd(gnd), .vdd(vdd), .A(data_181__15_), .Y(_2058_) );
NOR3X1 NOR3X1_100 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf2), .B(_1810__bF_buf7), .C(_2031_), .Y(_2059_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(_2037_), .C(_2059_), .Y(_91__15_) );
INVX1 INVX1_1166 ( .gnd(gnd), .vdd(vdd), .A(data_180__0_), .Y(_2060_) );
OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14965__bF_buf1), .C(_1561_), .Y(_2061_) );
AND2X2 AND2X2_511 ( .gnd(gnd), .vdd(vdd), .A(_1525__bF_buf1), .B(_2061_), .Y(_2062_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_1834_), .Y(_2063_) );
OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf3), .B(_1812__bF_buf2), .C(_2060_), .Y(_2064_) );
NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1812__bF_buf1), .B(_2063__bF_buf2), .Y(_2065_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_2065__bF_buf3), .Y(_2066_) );
AND2X2 AND2X2_512 ( .gnd(gnd), .vdd(vdd), .A(_2066_), .B(_2064_), .Y(_90__0_) );
INVX1 INVX1_1167 ( .gnd(gnd), .vdd(vdd), .A(data_180__1_), .Y(_2067_) );
OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf1), .B(_1812__bF_buf0), .C(_2067_), .Y(_2068_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_2065__bF_buf2), .Y(_2069_) );
AND2X2 AND2X2_513 ( .gnd(gnd), .vdd(vdd), .A(_2069_), .B(_2068_), .Y(_90__1_) );
INVX1 INVX1_1168 ( .gnd(gnd), .vdd(vdd), .A(data_180__2_), .Y(_2070_) );
OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf0), .B(_1812__bF_buf3), .C(_2070_), .Y(_2071_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_2065__bF_buf1), .Y(_2072_) );
AND2X2 AND2X2_514 ( .gnd(gnd), .vdd(vdd), .A(_2072_), .B(_2071_), .Y(_90__2_) );
INVX1 INVX1_1169 ( .gnd(gnd), .vdd(vdd), .A(data_180__3_), .Y(_2073_) );
OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf3), .B(_1812__bF_buf2), .C(_2073_), .Y(_2074_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_2065__bF_buf0), .Y(_2075_) );
AND2X2 AND2X2_515 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .B(_2074_), .Y(_90__3_) );
INVX1 INVX1_1170 ( .gnd(gnd), .vdd(vdd), .A(data_180__4_), .Y(_2076_) );
OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf2), .B(_1812__bF_buf1), .C(_2076_), .Y(_2077_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_2065__bF_buf3), .Y(_2078_) );
AND2X2 AND2X2_516 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2077_), .Y(_90__4_) );
INVX1 INVX1_1171 ( .gnd(gnd), .vdd(vdd), .A(data_180__5_), .Y(_2079_) );
OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf1), .B(_1812__bF_buf0), .C(_2079_), .Y(_2080_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_2065__bF_buf2), .Y(_2081_) );
AND2X2 AND2X2_517 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .B(_2080_), .Y(_90__5_) );
INVX1 INVX1_1172 ( .gnd(gnd), .vdd(vdd), .A(data_180__6_), .Y(_2082_) );
OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf0), .B(_1812__bF_buf3), .C(_2082_), .Y(_2083_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_2065__bF_buf1), .Y(_2084_) );
AND2X2 AND2X2_518 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2083_), .Y(_90__6_) );
INVX1 INVX1_1173 ( .gnd(gnd), .vdd(vdd), .A(data_180__7_), .Y(_2085_) );
OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf3), .B(_1812__bF_buf2), .C(_2085_), .Y(_2086_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_2065__bF_buf0), .Y(_2087_) );
AND2X2 AND2X2_519 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(_2086_), .Y(_90__7_) );
INVX1 INVX1_1174 ( .gnd(gnd), .vdd(vdd), .A(data_180__8_), .Y(_2088_) );
OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf2), .B(_1812__bF_buf1), .C(_2088_), .Y(_2089_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_2065__bF_buf3), .Y(_2090_) );
AND2X2 AND2X2_520 ( .gnd(gnd), .vdd(vdd), .A(_2090_), .B(_2089_), .Y(_90__8_) );
INVX1 INVX1_1175 ( .gnd(gnd), .vdd(vdd), .A(data_180__9_), .Y(_2091_) );
OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf1), .B(_1812__bF_buf0), .C(_2091_), .Y(_2092_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf7), .B(_2065__bF_buf2), .Y(_2093_) );
AND2X2 AND2X2_521 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_2092_), .Y(_90__9_) );
INVX1 INVX1_1176 ( .gnd(gnd), .vdd(vdd), .A(data_180__10_), .Y(_2094_) );
OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf0), .B(_1812__bF_buf3), .C(_2094_), .Y(_2095_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_2065__bF_buf1), .Y(_2096_) );
AND2X2 AND2X2_522 ( .gnd(gnd), .vdd(vdd), .A(_2096_), .B(_2095_), .Y(_90__10_) );
INVX1 INVX1_1177 ( .gnd(gnd), .vdd(vdd), .A(data_180__11_), .Y(_2097_) );
OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf3), .B(_1812__bF_buf2), .C(_2097_), .Y(_2098_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_2065__bF_buf0), .Y(_2099_) );
AND2X2 AND2X2_523 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_2098_), .Y(_90__11_) );
INVX1 INVX1_1178 ( .gnd(gnd), .vdd(vdd), .A(data_180__12_), .Y(_2100_) );
OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf2), .B(_1812__bF_buf1), .C(_2100_), .Y(_2101_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_2065__bF_buf3), .Y(_2102_) );
AND2X2 AND2X2_524 ( .gnd(gnd), .vdd(vdd), .A(_2102_), .B(_2101_), .Y(_90__12_) );
INVX1 INVX1_1179 ( .gnd(gnd), .vdd(vdd), .A(data_180__13_), .Y(_2103_) );
OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf1), .B(_1812__bF_buf0), .C(_2103_), .Y(_2104_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_2065__bF_buf2), .Y(_2105_) );
AND2X2 AND2X2_525 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2104_), .Y(_90__13_) );
INVX1 INVX1_1180 ( .gnd(gnd), .vdd(vdd), .A(data_180__14_), .Y(_2106_) );
OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_2063__bF_buf0), .B(_1812__bF_buf3), .C(_2106_), .Y(_2107_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_2065__bF_buf1), .Y(_2108_) );
AND2X2 AND2X2_526 ( .gnd(gnd), .vdd(vdd), .A(_2108_), .B(_2107_), .Y(_90__14_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_2065__bF_buf0), .B(data_180__15_), .Y(_2109_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_2065__bF_buf3), .Y(_2110_) );
AND2X2 AND2X2_527 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2110_), .Y(_90__15_) );
INVX1 INVX1_1181 ( .gnd(gnd), .vdd(vdd), .A(data_179__0_), .Y(_2111_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2061_), .B(_1525__bF_buf0), .Y(_2112_) );
NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2112_), .B(_1810__bF_buf6), .Y(_2113_) );
OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf2), .B(_15034_), .C(IDATA_PROG_write_bF_buf8), .Y(_2114_) );
INVX1 INVX1_1182 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .Y(_2115_) );
OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_1562__bF_buf3), .C(_2115_), .Y(_2116_) );
OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(_14942__bF_buf1), .C(_1686_), .Y(_2117_) );
OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf1), .B(_15019__bF_buf1), .C(_2117_), .Y(_2118_) );
NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2118_), .Y(_2119_) );
OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_1562__bF_buf2), .B(_15581_), .C(_2119_), .Y(_2120_) );
NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_1684_), .Y(_2121_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(_2113_), .Y(_2122_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2122_), .Y(_2123_) );
AND2X2 AND2X2_528 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2121_), .Y(_2124_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_2124_), .Y(_2125_) );
AND2X2 AND2X2_529 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(_2123_), .Y(_88__0_) );
INVX1 INVX1_1183 ( .gnd(gnd), .vdd(vdd), .A(data_179__1_), .Y(_2126_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .B(_2122_), .Y(_2127_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_2124_), .Y(_2128_) );
AND2X2 AND2X2_530 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2127_), .Y(_88__1_) );
INVX1 INVX1_1184 ( .gnd(gnd), .vdd(vdd), .A(data_179__2_), .Y(_2129_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(_2122_), .Y(_2130_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_2124_), .Y(_2131_) );
AND2X2 AND2X2_531 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(_2130_), .Y(_88__2_) );
INVX1 INVX1_1185 ( .gnd(gnd), .vdd(vdd), .A(data_179__3_), .Y(_2132_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_2122_), .Y(_2133_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_2124_), .Y(_2134_) );
AND2X2 AND2X2_532 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(_2133_), .Y(_88__3_) );
INVX1 INVX1_1186 ( .gnd(gnd), .vdd(vdd), .A(data_179__4_), .Y(_2135_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2122_), .Y(_2136_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_2124_), .Y(_2137_) );
AND2X2 AND2X2_533 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(_2136_), .Y(_88__4_) );
INVX1 INVX1_1187 ( .gnd(gnd), .vdd(vdd), .A(data_179__5_), .Y(_2138_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2138_), .B(_2122_), .Y(_2139_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_2124_), .Y(_2140_) );
AND2X2 AND2X2_534 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .B(_2139_), .Y(_88__5_) );
INVX1 INVX1_1188 ( .gnd(gnd), .vdd(vdd), .A(data_179__6_), .Y(_2141_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(_2122_), .Y(_2142_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_2124_), .Y(_2143_) );
AND2X2 AND2X2_535 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2142_), .Y(_88__6_) );
INVX1 INVX1_1189 ( .gnd(gnd), .vdd(vdd), .A(data_179__7_), .Y(_2144_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2144_), .B(_2122_), .Y(_2145_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_2124_), .Y(_2146_) );
AND2X2 AND2X2_536 ( .gnd(gnd), .vdd(vdd), .A(_2146_), .B(_2145_), .Y(_88__7_) );
INVX1 INVX1_1190 ( .gnd(gnd), .vdd(vdd), .A(data_179__8_), .Y(_2147_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(_2122_), .Y(_2148_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_2124_), .Y(_2149_) );
AND2X2 AND2X2_537 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_2148_), .Y(_88__8_) );
INVX1 INVX1_1191 ( .gnd(gnd), .vdd(vdd), .A(data_179__9_), .Y(_2150_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2122_), .Y(_2151_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_2124_), .Y(_2152_) );
AND2X2 AND2X2_538 ( .gnd(gnd), .vdd(vdd), .A(_2152_), .B(_2151_), .Y(_88__9_) );
INVX1 INVX1_1192 ( .gnd(gnd), .vdd(vdd), .A(data_179__10_), .Y(_2153_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(_2122_), .Y(_2154_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_2124_), .Y(_2155_) );
AND2X2 AND2X2_539 ( .gnd(gnd), .vdd(vdd), .A(_2155_), .B(_2154_), .Y(_88__10_) );
INVX1 INVX1_1193 ( .gnd(gnd), .vdd(vdd), .A(data_179__11_), .Y(_2156_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2122_), .Y(_2157_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_2124_), .Y(_2158_) );
AND2X2 AND2X2_540 ( .gnd(gnd), .vdd(vdd), .A(_2158_), .B(_2157_), .Y(_88__11_) );
INVX1 INVX1_1194 ( .gnd(gnd), .vdd(vdd), .A(data_179__12_), .Y(_2159_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(_2122_), .Y(_2160_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_2124_), .Y(_2161_) );
AND2X2 AND2X2_541 ( .gnd(gnd), .vdd(vdd), .A(_2161_), .B(_2160_), .Y(_88__12_) );
INVX1 INVX1_1195 ( .gnd(gnd), .vdd(vdd), .A(data_179__13_), .Y(_2162_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2162_), .B(_2122_), .Y(_2163_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_2124_), .Y(_2164_) );
AND2X2 AND2X2_542 ( .gnd(gnd), .vdd(vdd), .A(_2164_), .B(_2163_), .Y(_88__13_) );
INVX1 INVX1_1196 ( .gnd(gnd), .vdd(vdd), .A(data_179__14_), .Y(_2165_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .B(_2122_), .Y(_2166_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_2124_), .Y(_2167_) );
AND2X2 AND2X2_543 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2166_), .Y(_88__14_) );
INVX1 INVX1_1197 ( .gnd(gnd), .vdd(vdd), .A(data_179__15_), .Y(_2168_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2168_), .B(_2122_), .Y(_2169_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf2), .B(_2124_), .Y(_2170_) );
AND2X2 AND2X2_544 ( .gnd(gnd), .vdd(vdd), .A(_2170_), .B(_2169_), .Y(_88__15_) );
INVX1 INVX1_1198 ( .gnd(gnd), .vdd(vdd), .A(data_178__0_), .Y(_2171_) );
OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_1562__bF_buf1), .C(_2119_), .Y(_2172_) );
NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_2172_), .B(_1684_), .Y(_2173_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_2173_), .B(_2113_), .Y(_2174_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2174_), .Y(_2175_) );
AND2X2 AND2X2_545 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2173_), .Y(_2176_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_2176_), .Y(_2177_) );
AND2X2 AND2X2_546 ( .gnd(gnd), .vdd(vdd), .A(_2177_), .B(_2175_), .Y(_87__0_) );
INVX1 INVX1_1199 ( .gnd(gnd), .vdd(vdd), .A(data_178__1_), .Y(_2178_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2178_), .B(_2174_), .Y(_2179_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_2176_), .Y(_2180_) );
AND2X2 AND2X2_547 ( .gnd(gnd), .vdd(vdd), .A(_2180_), .B(_2179_), .Y(_87__1_) );
INVX1 INVX1_1200 ( .gnd(gnd), .vdd(vdd), .A(data_178__2_), .Y(_2181_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2181_), .B(_2174_), .Y(_2182_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_2176_), .Y(_2183_) );
AND2X2 AND2X2_548 ( .gnd(gnd), .vdd(vdd), .A(_2183_), .B(_2182_), .Y(_87__2_) );
INVX1 INVX1_1201 ( .gnd(gnd), .vdd(vdd), .A(data_178__3_), .Y(_2184_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2184_), .B(_2174_), .Y(_2185_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_2176_), .Y(_2186_) );
AND2X2 AND2X2_549 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2185_), .Y(_87__3_) );
INVX1 INVX1_1202 ( .gnd(gnd), .vdd(vdd), .A(data_178__4_), .Y(_2187_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2187_), .B(_2174_), .Y(_2188_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_2176_), .Y(_2189_) );
AND2X2 AND2X2_550 ( .gnd(gnd), .vdd(vdd), .A(_2189_), .B(_2188_), .Y(_87__4_) );
INVX1 INVX1_1203 ( .gnd(gnd), .vdd(vdd), .A(data_178__5_), .Y(_2190_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .B(_2174_), .Y(_2191_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_2176_), .Y(_2192_) );
AND2X2 AND2X2_551 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .B(_2191_), .Y(_87__5_) );
INVX1 INVX1_1204 ( .gnd(gnd), .vdd(vdd), .A(data_178__6_), .Y(_2193_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2174_), .Y(_2194_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_2176_), .Y(_2195_) );
AND2X2 AND2X2_552 ( .gnd(gnd), .vdd(vdd), .A(_2195_), .B(_2194_), .Y(_87__6_) );
INVX1 INVX1_1205 ( .gnd(gnd), .vdd(vdd), .A(data_178__7_), .Y(_2196_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2196_), .B(_2174_), .Y(_2197_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_2176_), .Y(_2198_) );
AND2X2 AND2X2_553 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .B(_2197_), .Y(_87__7_) );
INVX1 INVX1_1206 ( .gnd(gnd), .vdd(vdd), .A(data_178__8_), .Y(_2199_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2199_), .B(_2174_), .Y(_2200_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_2176_), .Y(_2201_) );
AND2X2 AND2X2_554 ( .gnd(gnd), .vdd(vdd), .A(_2201_), .B(_2200_), .Y(_87__8_) );
INVX1 INVX1_1207 ( .gnd(gnd), .vdd(vdd), .A(data_178__9_), .Y(_2202_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2202_), .B(_2174_), .Y(_2203_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_2176_), .Y(_2204_) );
AND2X2 AND2X2_555 ( .gnd(gnd), .vdd(vdd), .A(_2204_), .B(_2203_), .Y(_87__9_) );
INVX1 INVX1_1208 ( .gnd(gnd), .vdd(vdd), .A(data_178__10_), .Y(_2205_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2205_), .B(_2174_), .Y(_2206_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf3), .B(_2176_), .Y(_2207_) );
AND2X2 AND2X2_556 ( .gnd(gnd), .vdd(vdd), .A(_2207_), .B(_2206_), .Y(_87__10_) );
INVX1 INVX1_1209 ( .gnd(gnd), .vdd(vdd), .A(data_178__11_), .Y(_2208_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2174_), .Y(_2209_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_2176_), .Y(_2210_) );
AND2X2 AND2X2_557 ( .gnd(gnd), .vdd(vdd), .A(_2210_), .B(_2209_), .Y(_87__11_) );
INVX1 INVX1_1210 ( .gnd(gnd), .vdd(vdd), .A(data_178__12_), .Y(_2211_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2211_), .B(_2174_), .Y(_2212_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_2176_), .Y(_2213_) );
AND2X2 AND2X2_558 ( .gnd(gnd), .vdd(vdd), .A(_2213_), .B(_2212_), .Y(_87__12_) );
INVX1 INVX1_1211 ( .gnd(gnd), .vdd(vdd), .A(data_178__13_), .Y(_2214_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2174_), .Y(_2215_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_2176_), .Y(_2216_) );
AND2X2 AND2X2_559 ( .gnd(gnd), .vdd(vdd), .A(_2216_), .B(_2215_), .Y(_87__13_) );
INVX1 INVX1_1212 ( .gnd(gnd), .vdd(vdd), .A(data_178__14_), .Y(_2217_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2217_), .B(_2174_), .Y(_2218_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_2176_), .Y(_2219_) );
AND2X2 AND2X2_560 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .B(_2218_), .Y(_87__14_) );
INVX1 INVX1_1213 ( .gnd(gnd), .vdd(vdd), .A(data_178__15_), .Y(_2220_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_2220_), .B(_2174_), .Y(_2221_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_2176_), .Y(_2222_) );
AND2X2 AND2X2_561 ( .gnd(gnd), .vdd(vdd), .A(_2222_), .B(_2221_), .Y(_87__15_) );
INVX1 INVX1_1214 ( .gnd(gnd), .vdd(vdd), .A(data_177__0_), .Y(_2223_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_15684_), .C(_2114_), .Y(_2224_) );
OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_1562__bF_buf0), .C(_2224_), .Y(_2225_) );
NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2225_), .Y(_2226_) );
AND2X2 AND2X2_562 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2226_), .Y(_2227_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2227_), .B(_2113_), .Y(_2228_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2223_), .B(_2228_), .Y(_2229_) );
AND2X2 AND2X2_563 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2227_), .Y(_2230_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_2230_), .Y(_2231_) );
AND2X2 AND2X2_564 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .B(_2229_), .Y(_86__0_) );
INVX1 INVX1_1215 ( .gnd(gnd), .vdd(vdd), .A(data_177__1_), .Y(_2232_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2228_), .Y(_2233_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_2230_), .Y(_2234_) );
AND2X2 AND2X2_565 ( .gnd(gnd), .vdd(vdd), .A(_2234_), .B(_2233_), .Y(_86__1_) );
INVX1 INVX1_1216 ( .gnd(gnd), .vdd(vdd), .A(data_177__2_), .Y(_2235_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(_2228_), .Y(_2236_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_2230_), .Y(_2237_) );
AND2X2 AND2X2_566 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_2236_), .Y(_86__2_) );
INVX1 INVX1_1217 ( .gnd(gnd), .vdd(vdd), .A(data_177__3_), .Y(_2238_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_2238_), .B(_2228_), .Y(_2239_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_2230_), .Y(_2240_) );
AND2X2 AND2X2_567 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .B(_2239_), .Y(_86__3_) );
INVX1 INVX1_1218 ( .gnd(gnd), .vdd(vdd), .A(data_177__4_), .Y(_2241_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2241_), .B(_2228_), .Y(_2242_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_2230_), .Y(_2243_) );
AND2X2 AND2X2_568 ( .gnd(gnd), .vdd(vdd), .A(_2243_), .B(_2242_), .Y(_86__4_) );
INVX1 INVX1_1219 ( .gnd(gnd), .vdd(vdd), .A(data_177__5_), .Y(_2244_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .B(_2228_), .Y(_2245_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_2230_), .Y(_2246_) );
AND2X2 AND2X2_569 ( .gnd(gnd), .vdd(vdd), .A(_2246_), .B(_2245_), .Y(_86__5_) );
INVX1 INVX1_1220 ( .gnd(gnd), .vdd(vdd), .A(data_177__6_), .Y(_2247_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2247_), .B(_2228_), .Y(_2248_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_2230_), .Y(_2249_) );
AND2X2 AND2X2_570 ( .gnd(gnd), .vdd(vdd), .A(_2249_), .B(_2248_), .Y(_86__6_) );
INVX1 INVX1_1221 ( .gnd(gnd), .vdd(vdd), .A(data_177__7_), .Y(_2250_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2250_), .B(_2228_), .Y(_2251_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_2230_), .Y(_2252_) );
AND2X2 AND2X2_571 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .B(_2251_), .Y(_86__7_) );
INVX1 INVX1_1222 ( .gnd(gnd), .vdd(vdd), .A(data_177__8_), .Y(_2253_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2253_), .B(_2228_), .Y(_2254_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_2230_), .Y(_2255_) );
AND2X2 AND2X2_572 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .B(_2254_), .Y(_86__8_) );
INVX1 INVX1_1223 ( .gnd(gnd), .vdd(vdd), .A(data_177__9_), .Y(_2256_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2256_), .B(_2228_), .Y(_2257_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_2230_), .Y(_2258_) );
AND2X2 AND2X2_573 ( .gnd(gnd), .vdd(vdd), .A(_2258_), .B(_2257_), .Y(_86__9_) );
INVX1 INVX1_1224 ( .gnd(gnd), .vdd(vdd), .A(data_177__10_), .Y(_2259_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_2259_), .B(_2228_), .Y(_2260_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_2230_), .Y(_2261_) );
AND2X2 AND2X2_574 ( .gnd(gnd), .vdd(vdd), .A(_2261_), .B(_2260_), .Y(_86__10_) );
INVX1 INVX1_1225 ( .gnd(gnd), .vdd(vdd), .A(data_177__11_), .Y(_2262_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_2262_), .B(_2228_), .Y(_2263_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_2230_), .Y(_2264_) );
AND2X2 AND2X2_575 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .B(_2263_), .Y(_86__11_) );
INVX1 INVX1_1226 ( .gnd(gnd), .vdd(vdd), .A(data_177__12_), .Y(_2265_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .B(_2228_), .Y(_2266_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_2230_), .Y(_2267_) );
AND2X2 AND2X2_576 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2266_), .Y(_86__12_) );
INVX1 INVX1_1227 ( .gnd(gnd), .vdd(vdd), .A(data_177__13_), .Y(_2268_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2268_), .B(_2228_), .Y(_2269_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_2230_), .Y(_2270_) );
AND2X2 AND2X2_577 ( .gnd(gnd), .vdd(vdd), .A(_2270_), .B(_2269_), .Y(_86__13_) );
INVX1 INVX1_1228 ( .gnd(gnd), .vdd(vdd), .A(data_177__14_), .Y(_2271_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2271_), .B(_2228_), .Y(_2272_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_2230_), .Y(_2273_) );
AND2X2 AND2X2_578 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_2272_), .Y(_86__14_) );
INVX1 INVX1_1229 ( .gnd(gnd), .vdd(vdd), .A(data_177__15_), .Y(_2274_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2274_), .B(_2228_), .Y(_2275_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_2230_), .Y(_2276_) );
AND2X2 AND2X2_579 ( .gnd(gnd), .vdd(vdd), .A(_2276_), .B(_2275_), .Y(_86__15_) );
OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_1562__bF_buf3), .C(_1687_), .Y(_2277_) );
NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_2277_), .B(_1684_), .Y(_2278_) );
NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_2278_), .C(_1834_), .Y(_2279_) );
NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf1), .B(_2279_), .Y(_2280_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_2280__bF_buf4), .Y(_2281_) );
OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(data_176__0_), .B(_2280__bF_buf3), .C(_2281_), .Y(_2282_) );
INVX1 INVX1_1230 ( .gnd(gnd), .vdd(vdd), .A(_2282_), .Y(_85__0_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_2280__bF_buf2), .Y(_2283_) );
OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(data_176__1_), .B(_2280__bF_buf1), .C(_2283_), .Y(_2284_) );
INVX1 INVX1_1231 ( .gnd(gnd), .vdd(vdd), .A(_2284_), .Y(_85__1_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_2280__bF_buf0), .Y(_2285_) );
OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(data_176__2_), .B(_2280__bF_buf4), .C(_2285_), .Y(_2286_) );
INVX1 INVX1_1232 ( .gnd(gnd), .vdd(vdd), .A(_2286_), .Y(_85__2_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_2280__bF_buf3), .Y(_2287_) );
OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(data_176__3_), .B(_2280__bF_buf2), .C(_2287_), .Y(_2288_) );
INVX1 INVX1_1233 ( .gnd(gnd), .vdd(vdd), .A(_2288_), .Y(_85__3_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_2280__bF_buf1), .Y(_2289_) );
OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(data_176__4_), .B(_2280__bF_buf0), .C(_2289_), .Y(_2290_) );
INVX1 INVX1_1234 ( .gnd(gnd), .vdd(vdd), .A(_2290_), .Y(_85__4_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_2280__bF_buf4), .Y(_2291_) );
OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(data_176__5_), .B(_2280__bF_buf3), .C(_2291_), .Y(_2292_) );
INVX1 INVX1_1235 ( .gnd(gnd), .vdd(vdd), .A(_2292_), .Y(_85__5_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_2280__bF_buf2), .Y(_2293_) );
OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(data_176__6_), .B(_2280__bF_buf1), .C(_2293_), .Y(_2294_) );
INVX1 INVX1_1236 ( .gnd(gnd), .vdd(vdd), .A(_2294_), .Y(_85__6_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_2280__bF_buf0), .Y(_2295_) );
OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(data_176__7_), .B(_2280__bF_buf4), .C(_2295_), .Y(_2296_) );
INVX1 INVX1_1237 ( .gnd(gnd), .vdd(vdd), .A(_2296_), .Y(_85__7_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_2280__bF_buf3), .Y(_2297_) );
OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(data_176__8_), .B(_2280__bF_buf2), .C(_2297_), .Y(_2298_) );
INVX1 INVX1_1238 ( .gnd(gnd), .vdd(vdd), .A(_2298_), .Y(_85__8_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_2280__bF_buf1), .Y(_2299_) );
OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(data_176__9_), .B(_2280__bF_buf0), .C(_2299_), .Y(_2300_) );
INVX1 INVX1_1239 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .Y(_85__9_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_2280__bF_buf4), .Y(_2301_) );
OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(data_176__10_), .B(_2280__bF_buf3), .C(_2301_), .Y(_2302_) );
INVX1 INVX1_1240 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .Y(_85__10_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_2280__bF_buf2), .Y(_2303_) );
OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(data_176__11_), .B(_2280__bF_buf1), .C(_2303_), .Y(_2304_) );
INVX1 INVX1_1241 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .Y(_85__11_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_2280__bF_buf0), .Y(_2305_) );
OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(data_176__12_), .B(_2280__bF_buf4), .C(_2305_), .Y(_2306_) );
INVX1 INVX1_1242 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .Y(_85__12_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_2280__bF_buf3), .Y(_2307_) );
OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(data_176__13_), .B(_2280__bF_buf2), .C(_2307_), .Y(_2308_) );
INVX1 INVX1_1243 ( .gnd(gnd), .vdd(vdd), .A(_2308_), .Y(_85__13_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf5), .B(_2280__bF_buf1), .Y(_2309_) );
OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(data_176__14_), .B(_2280__bF_buf0), .C(_2309_), .Y(_2310_) );
INVX1 INVX1_1244 ( .gnd(gnd), .vdd(vdd), .A(_2310_), .Y(_85__14_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_2280__bF_buf4), .Y(_2311_) );
OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(data_176__15_), .B(_2280__bF_buf3), .C(_2311_), .Y(_2312_) );
INVX1 INVX1_1245 ( .gnd(gnd), .vdd(vdd), .A(_2312_), .Y(_85__15_) );
OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_14950_), .B(_14954_), .C(_14963__bF_buf0), .Y(_2313_) );
OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14940_), .C(_14974_), .Y(_2314_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_2313_), .C(_2314_), .Y(_2315_) );
INVX4 INVX4_9 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf0), .Y(_2316_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_14983_), .B(_2316_), .Y(_2317_) );
NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .B(_2315_), .C(_2317_), .Y(_2318_) );
NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf0), .B(_2318_), .Y(_2319_) );
NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(data_175__0_), .B(_2319__bF_buf4), .Y(_2320_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_2319__bF_buf3), .C(_2320_), .Y(_84__0_) );
NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(data_175__1_), .B(_2319__bF_buf2), .Y(_2321_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_2319__bF_buf1), .C(_2321_), .Y(_84__1_) );
NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(data_175__2_), .B(_2319__bF_buf0), .Y(_2322_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_2319__bF_buf4), .C(_2322_), .Y(_84__2_) );
NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(data_175__3_), .B(_2319__bF_buf3), .Y(_2323_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_2319__bF_buf2), .C(_2323_), .Y(_84__3_) );
NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(data_175__4_), .B(_2319__bF_buf1), .Y(_2324_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_2319__bF_buf0), .C(_2324_), .Y(_84__4_) );
NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(data_175__5_), .B(_2319__bF_buf4), .Y(_2325_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_2319__bF_buf3), .C(_2325_), .Y(_84__5_) );
NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(data_175__6_), .B(_2319__bF_buf2), .Y(_2326_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_2319__bF_buf1), .C(_2326_), .Y(_84__6_) );
NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(data_175__7_), .B(_2319__bF_buf0), .Y(_2327_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_2319__bF_buf4), .C(_2327_), .Y(_84__7_) );
NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(data_175__8_), .B(_2319__bF_buf3), .Y(_2328_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_2319__bF_buf2), .C(_2328_), .Y(_84__8_) );
NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(data_175__9_), .B(_2319__bF_buf1), .Y(_2329_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_2319__bF_buf0), .C(_2329_), .Y(_84__9_) );
NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(data_175__10_), .B(_2319__bF_buf4), .Y(_2330_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_2319__bF_buf3), .C(_2330_), .Y(_84__10_) );
NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(data_175__11_), .B(_2319__bF_buf2), .Y(_2331_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_2319__bF_buf1), .C(_2331_), .Y(_84__11_) );
NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(data_175__12_), .B(_2319__bF_buf0), .Y(_2332_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_2319__bF_buf4), .C(_2332_), .Y(_84__12_) );
NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(data_175__13_), .B(_2319__bF_buf3), .Y(_2333_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_2319__bF_buf2), .C(_2333_), .Y(_84__13_) );
NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(data_175__14_), .B(_2319__bF_buf1), .Y(_2334_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_2319__bF_buf0), .C(_2334_), .Y(_84__14_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_2319__bF_buf4), .Y(_2335_) );
OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(data_175__15_), .B(_2319__bF_buf3), .C(_2335_), .Y(_2336_) );
INVX1 INVX1_1246 ( .gnd(gnd), .vdd(vdd), .A(_2336_), .Y(_84__15_) );
INVX1 INVX1_1247 ( .gnd(gnd), .vdd(vdd), .A(data_174__0_), .Y(_2337_) );
OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15019__bF_buf3), .C(_2337_), .Y(_2338_) );
NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf2), .B(_15788__bF_buf2), .Y(_2339_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_2339__bF_buf3), .Y(_2340_) );
AND2X2 AND2X2_580 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2338_), .Y(_83__0_) );
INVX1 INVX1_1248 ( .gnd(gnd), .vdd(vdd), .A(data_174__1_), .Y(_2341_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_15793__bF_buf0), .B(_2316_), .Y(_2342_) );
MUX2X1 MUX2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_14894__bF_buf4), .S(_2342_), .Y(_83__1_) );
NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(data_174__2_), .B(_2339__bF_buf2), .Y(_2343_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_2339__bF_buf1), .C(_2343_), .Y(_83__2_) );
INVX1 INVX1_1249 ( .gnd(gnd), .vdd(vdd), .A(data_174__3_), .Y(_2344_) );
OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15019__bF_buf1), .C(_2344_), .Y(_2345_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_2339__bF_buf0), .Y(_2346_) );
AND2X2 AND2X2_581 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2345_), .Y(_83__3_) );
INVX1 INVX1_1250 ( .gnd(gnd), .vdd(vdd), .A(data_174__4_), .Y(_2347_) );
OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15019__bF_buf0), .C(_2347_), .Y(_2348_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_2339__bF_buf3), .Y(_2349_) );
AND2X2 AND2X2_582 ( .gnd(gnd), .vdd(vdd), .A(_2349_), .B(_2348_), .Y(_83__4_) );
INVX1 INVX1_1251 ( .gnd(gnd), .vdd(vdd), .A(data_174__5_), .Y(_2350_) );
OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15019__bF_buf3), .C(_2350_), .Y(_2351_) );
NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_2339__bF_buf2), .Y(_2352_) );
AND2X2 AND2X2_583 ( .gnd(gnd), .vdd(vdd), .A(_2352_), .B(_2351_), .Y(_83__5_) );
INVX1 INVX1_1252 ( .gnd(gnd), .vdd(vdd), .A(data_174__6_), .Y(_2353_) );
OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15019__bF_buf2), .C(_2353_), .Y(_2354_) );
NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_2339__bF_buf1), .Y(_2355_) );
AND2X2 AND2X2_584 ( .gnd(gnd), .vdd(vdd), .A(_2355_), .B(_2354_), .Y(_83__6_) );
INVX1 INVX1_1253 ( .gnd(gnd), .vdd(vdd), .A(data_174__7_), .Y(_2356_) );
OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15019__bF_buf1), .C(_2356_), .Y(_2357_) );
NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_2339__bF_buf0), .Y(_2358_) );
AND2X2 AND2X2_585 ( .gnd(gnd), .vdd(vdd), .A(_2358_), .B(_2357_), .Y(_83__7_) );
INVX1 INVX1_1254 ( .gnd(gnd), .vdd(vdd), .A(data_174__8_), .Y(_2359_) );
OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15019__bF_buf0), .C(_2359_), .Y(_2360_) );
NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_2339__bF_buf3), .Y(_2361_) );
AND2X2 AND2X2_586 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .B(_2360_), .Y(_83__8_) );
NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(data_174__9_), .B(_2339__bF_buf2), .Y(_2362_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_2339__bF_buf1), .C(_2362_), .Y(_83__9_) );
NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(data_174__10_), .B(_2339__bF_buf0), .Y(_2363_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_2339__bF_buf3), .C(_2363_), .Y(_83__10_) );
NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(data_174__11_), .B(_2339__bF_buf2), .Y(_2364_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_2339__bF_buf1), .C(_2364_), .Y(_83__11_) );
INVX1 INVX1_1255 ( .gnd(gnd), .vdd(vdd), .A(data_174__12_), .Y(_2365_) );
OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15019__bF_buf3), .C(_2365_), .Y(_2366_) );
NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_2339__bF_buf0), .Y(_2367_) );
AND2X2 AND2X2_587 ( .gnd(gnd), .vdd(vdd), .A(_2367_), .B(_2366_), .Y(_83__12_) );
INVX1 INVX1_1256 ( .gnd(gnd), .vdd(vdd), .A(data_174__13_), .Y(_2368_) );
OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15019__bF_buf2), .C(_2368_), .Y(_2369_) );
NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_15793__bF_buf5), .C(_2316_), .Y(_2370_) );
AND2X2 AND2X2_588 ( .gnd(gnd), .vdd(vdd), .A(_2369_), .B(_2370_), .Y(_83__13_) );
NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(data_174__14_), .B(_2339__bF_buf3), .Y(_2371_) );
NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf3), .B(_2342_), .Y(_2372_) );
NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2371_), .Y(_83__14_) );
NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(data_174__15_), .B(_2339__bF_buf2), .Y(_2373_) );
NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf1), .B(_2342_), .Y(_2374_) );
NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2374_), .B(_2373_), .Y(_83__15_) );
INVX1 INVX1_1257 ( .gnd(gnd), .vdd(vdd), .A(data_173__0_), .Y(_2375_) );
NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .B(_2316_), .Y(_2376_) );
INVX1 INVX1_1258 ( .gnd(gnd), .vdd(vdd), .A(_2278_), .Y(_2377_) );
NOR3X1 NOR3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_2112_), .B(_2377_), .C(_1810__bF_buf5), .Y(_2378_) );
INVX1 INVX1_1259 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .Y(_2379_) );
NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2378_), .Y(_2380_) );
NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .B(_15739_), .Y(_2381_) );
NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2381_), .B(_1000__bF_buf0), .Y(_2382_) );
INVX1 INVX1_1260 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .Y(_2383_) );
OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf3), .B(_14975_), .C(_1561_), .Y(_2384_) );
OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_15019__bF_buf1), .C(_2384_), .Y(_2385_) );
NOR3X1 NOR3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_2383_), .B(_2385_), .C(_2063__bF_buf3), .Y(_2386_) );
NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2376_), .B(_2386_), .C(_2380_), .Y(_2387_) );
MUX2X1 MUX2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2375_), .B(_14932__bF_buf4), .S(_2387__bF_buf3), .Y(_82__0_) );
INVX1 INVX1_1261 ( .gnd(gnd), .vdd(vdd), .A(data_173__1_), .Y(_2388_) );
MUX2X1 MUX2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2388_), .B(_14894__bF_buf3), .S(_2387__bF_buf2), .Y(_82__1_) );
INVX1 INVX1_1262 ( .gnd(gnd), .vdd(vdd), .A(data_173__2_), .Y(_2389_) );
MUX2X1 MUX2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_14897__bF_buf0), .S(_2387__bF_buf1), .Y(_82__2_) );
INVX1 INVX1_1263 ( .gnd(gnd), .vdd(vdd), .A(data_173__3_), .Y(_2390_) );
NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2390_), .B(_2387__bF_buf0), .Y(_2391_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_2387__bF_buf3), .Y(_2392_) );
NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_2392_), .Y(_2393_) );
AND2X2 AND2X2_589 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .B(_2391_), .Y(_82__3_) );
INVX1 INVX1_1264 ( .gnd(gnd), .vdd(vdd), .A(data_173__4_), .Y(_2394_) );
MUX2X1 MUX2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2394_), .B(_14902__bF_buf11), .S(_2387__bF_buf2), .Y(_82__4_) );
INVX1 INVX1_1265 ( .gnd(gnd), .vdd(vdd), .A(data_173__5_), .Y(_2395_) );
MUX2X1 MUX2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2395_), .B(_14903__bF_buf12), .S(_2387__bF_buf1), .Y(_82__5_) );
INVX1 INVX1_1266 ( .gnd(gnd), .vdd(vdd), .A(data_173__6_), .Y(_2396_) );
MUX2X1 MUX2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2396_), .B(_15049__bF_buf0), .S(_2387__bF_buf0), .Y(_82__6_) );
INVX1 INVX1_1267 ( .gnd(gnd), .vdd(vdd), .A(data_173__7_), .Y(_2397_) );
NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2387__bF_buf3), .Y(_2398_) );
NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_2392_), .Y(_2399_) );
AND2X2 AND2X2_590 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .B(_2398_), .Y(_82__7_) );
INVX1 INVX1_1268 ( .gnd(gnd), .vdd(vdd), .A(data_173__8_), .Y(_2400_) );
NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .B(_2387__bF_buf2), .Y(_2401_) );
NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_2392_), .Y(_2402_) );
AND2X2 AND2X2_591 ( .gnd(gnd), .vdd(vdd), .A(_2402_), .B(_2401_), .Y(_82__8_) );
INVX1 INVX1_1269 ( .gnd(gnd), .vdd(vdd), .A(data_173__9_), .Y(_2403_) );
NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2403_), .B(_2387__bF_buf1), .Y(_2404_) );
NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_2392_), .Y(_2405_) );
AND2X2 AND2X2_592 ( .gnd(gnd), .vdd(vdd), .A(_2405_), .B(_2404_), .Y(_82__9_) );
INVX1 INVX1_1270 ( .gnd(gnd), .vdd(vdd), .A(data_173__10_), .Y(_2406_) );
MUX2X1 MUX2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2406_), .B(_15055__bF_buf12), .S(_2387__bF_buf0), .Y(_82__10_) );
INVX1 INVX1_1271 ( .gnd(gnd), .vdd(vdd), .A(data_173__11_), .Y(_2407_) );
MUX2X1 MUX2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2407_), .B(_14918__bF_buf13), .S(_2387__bF_buf3), .Y(_82__11_) );
INVX1 INVX1_1272 ( .gnd(gnd), .vdd(vdd), .A(data_173__12_), .Y(_2408_) );
MUX2X1 MUX2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .B(_14920__bF_buf12), .S(_2387__bF_buf2), .Y(_82__12_) );
INVX1 INVX1_1273 ( .gnd(gnd), .vdd(vdd), .A(data_173__13_), .Y(_2409_) );
NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(_2387__bF_buf1), .Y(_2410_) );
NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_2392_), .Y(_2411_) );
AND2X2 AND2X2_593 ( .gnd(gnd), .vdd(vdd), .A(_2411_), .B(_2410_), .Y(_82__13_) );
INVX1 INVX1_1274 ( .gnd(gnd), .vdd(vdd), .A(data_173__14_), .Y(_2412_) );
MUX2X1 MUX2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2412_), .B(_15060__bF_buf3), .S(_2387__bF_buf0), .Y(_82__14_) );
INVX1 INVX1_1275 ( .gnd(gnd), .vdd(vdd), .A(data_173__15_), .Y(_2413_) );
NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(_2387__bF_buf3), .Y(_2414_) );
NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_2392_), .Y(_2415_) );
AND2X2 AND2X2_594 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .B(_2414_), .Y(_82__15_) );
INVX1 INVX1_1276 ( .gnd(gnd), .vdd(vdd), .A(data_172__0_), .Y(_2416_) );
OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_14981_), .B(_14983_), .C(_2316_), .Y(_2417_) );
NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2417_), .B(_2386_), .C(_2380_), .Y(_2418_) );
NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2416_), .B(_2418__bF_buf3), .Y(_2419_) );
INVX4 INVX4_10 ( .gnd(gnd), .vdd(vdd), .A(_2418__bF_buf2), .Y(_2420_) );
NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_2420_), .Y(_2421_) );
AND2X2 AND2X2_595 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(_2419_), .Y(_81__0_) );
INVX1 INVX1_1277 ( .gnd(gnd), .vdd(vdd), .A(data_172__1_), .Y(_2422_) );
NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2422_), .B(_2418__bF_buf1), .Y(_2423_) );
NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_2420_), .Y(_2424_) );
AND2X2 AND2X2_596 ( .gnd(gnd), .vdd(vdd), .A(_2424_), .B(_2423_), .Y(_81__1_) );
INVX1 INVX1_1278 ( .gnd(gnd), .vdd(vdd), .A(data_172__2_), .Y(_2425_) );
NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2425_), .B(_2418__bF_buf0), .Y(_2426_) );
NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_2420_), .Y(_2427_) );
AND2X2 AND2X2_597 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(_2426_), .Y(_81__2_) );
INVX1 INVX1_1279 ( .gnd(gnd), .vdd(vdd), .A(data_172__3_), .Y(_2428_) );
MUX2X1 MUX2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2428_), .B(_14899__bF_buf1), .S(_2418__bF_buf3), .Y(_81__3_) );
INVX1 INVX1_1280 ( .gnd(gnd), .vdd(vdd), .A(data_172__4_), .Y(_2429_) );
NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2418__bF_buf2), .Y(_2430_) );
NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_2420_), .Y(_2431_) );
AND2X2 AND2X2_598 ( .gnd(gnd), .vdd(vdd), .A(_2431_), .B(_2430_), .Y(_81__4_) );
INVX1 INVX1_1281 ( .gnd(gnd), .vdd(vdd), .A(data_172__5_), .Y(_2432_) );
NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2432_), .B(_2418__bF_buf1), .Y(_2433_) );
NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_2420_), .Y(_2434_) );
AND2X2 AND2X2_599 ( .gnd(gnd), .vdd(vdd), .A(_2434_), .B(_2433_), .Y(_81__5_) );
INVX1 INVX1_1282 ( .gnd(gnd), .vdd(vdd), .A(data_172__6_), .Y(_2435_) );
NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2435_), .B(_2418__bF_buf0), .Y(_2436_) );
NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_2420_), .Y(_2437_) );
AND2X2 AND2X2_600 ( .gnd(gnd), .vdd(vdd), .A(_2437_), .B(_2436_), .Y(_81__6_) );
INVX1 INVX1_1283 ( .gnd(gnd), .vdd(vdd), .A(data_172__7_), .Y(_2438_) );
MUX2X1 MUX2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2438_), .B(_14908__bF_buf10), .S(_2418__bF_buf3), .Y(_81__7_) );
INVX1 INVX1_1284 ( .gnd(gnd), .vdd(vdd), .A(data_172__8_), .Y(_2439_) );
MUX2X1 MUX2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2439_), .B(_15052__bF_buf11), .S(_2418__bF_buf2), .Y(_81__8_) );
INVX1 INVX1_1285 ( .gnd(gnd), .vdd(vdd), .A(data_172__9_), .Y(_2440_) );
MUX2X1 MUX2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2440_), .B(_14913__bF_buf14), .S(_2418__bF_buf1), .Y(_81__9_) );
INVX1 INVX1_1286 ( .gnd(gnd), .vdd(vdd), .A(data_172__10_), .Y(_2441_) );
NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2441_), .B(_2418__bF_buf0), .Y(_2442_) );
NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_2420_), .Y(_2443_) );
AND2X2 AND2X2_601 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2442_), .Y(_81__10_) );
INVX1 INVX1_1287 ( .gnd(gnd), .vdd(vdd), .A(data_172__11_), .Y(_2444_) );
NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(_2418__bF_buf3), .Y(_2445_) );
NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_2420_), .Y(_2446_) );
AND2X2 AND2X2_602 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2445_), .Y(_81__11_) );
INVX1 INVX1_1288 ( .gnd(gnd), .vdd(vdd), .A(data_172__12_), .Y(_2447_) );
NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2447_), .B(_2418__bF_buf2), .Y(_2448_) );
NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_2420_), .Y(_2449_) );
AND2X2 AND2X2_603 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2448_), .Y(_81__12_) );
INVX1 INVX1_1289 ( .gnd(gnd), .vdd(vdd), .A(data_172__13_), .Y(_2450_) );
MUX2X1 MUX2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(_14924__bF_buf10), .S(_2418__bF_buf1), .Y(_81__13_) );
INVX1 INVX1_1290 ( .gnd(gnd), .vdd(vdd), .A(data_172__14_), .Y(_2451_) );
NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2418__bF_buf0), .Y(_2452_) );
NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_2420_), .Y(_2453_) );
AND2X2 AND2X2_604 ( .gnd(gnd), .vdd(vdd), .A(_2453_), .B(_2452_), .Y(_81__14_) );
INVX1 INVX1_1291 ( .gnd(gnd), .vdd(vdd), .A(data_172__15_), .Y(_2454_) );
MUX2X1 MUX2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2454_), .B(_15062__bF_buf10), .S(_2418__bF_buf3), .Y(_81__15_) );
INVX1 INVX1_1292 ( .gnd(gnd), .vdd(vdd), .A(data_171__0_), .Y(_2455_) );
OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_15019__bF_buf0), .C(_2384_), .Y(_2456_) );
NOR3X1 NOR3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2456_), .C(_2378_), .Y(_2457_) );
INVX1 INVX1_1293 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .Y(_2458_) );
INVX1 INVX1_1294 ( .gnd(gnd), .vdd(vdd), .A(_15951_), .Y(_2459_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_2316_), .B(_15161_), .C(_14882__bF_buf15_bF_buf3), .Y(_2460_) );
OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_15019__bF_buf3), .C(_2460_), .Y(_2461_) );
NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2458_), .B(_2461_), .Y(_2462_) );
AND2X2 AND2X2_605 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2462_), .Y(_2463_) );
NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2463_), .B(_2113_), .Y(_2464_) );
INVX1 INVX1_1295 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .Y(_2465_) );
NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_2465_), .Y(_2466_) );
MUX2X1 MUX2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_14932__bF_buf2), .S(_2466_), .Y(_80__0_) );
INVX1 INVX1_1296 ( .gnd(gnd), .vdd(vdd), .A(data_171__1_), .Y(_2467_) );
MUX2X1 MUX2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(_14894__bF_buf1), .S(_2466_), .Y(_80__1_) );
INVX1 INVX1_1297 ( .gnd(gnd), .vdd(vdd), .A(data_171__2_), .Y(_2468_) );
MUX2X1 MUX2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2468_), .B(_14897__bF_buf13), .S(_2466_), .Y(_80__2_) );
INVX1 INVX1_1298 ( .gnd(gnd), .vdd(vdd), .A(_2456_), .Y(_2469_) );
NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2318_), .B(_2469_), .C(_2279_), .Y(_2470_) );
NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2470_), .Y(_2471_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_2465_), .C(data_171__3_), .Y(_2472_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_2471__bF_buf3), .C(_2472_), .Y(_80__3_) );
NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(data_171__4_), .B(_2471__bF_buf2), .Y(_2473_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_2471__bF_buf1), .C(_2473_), .Y(_80__4_) );
INVX1 INVX1_1299 ( .gnd(gnd), .vdd(vdd), .A(data_171__5_), .Y(_2474_) );
MUX2X1 MUX2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_2474_), .S(_2471__bF_buf0), .Y(_80__5_) );
NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(data_171__6_), .B(_2471__bF_buf3), .Y(_2475_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_2471__bF_buf2), .C(_2475_), .Y(_80__6_) );
NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(data_171__7_), .B(_2471__bF_buf1), .Y(_2476_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_2471__bF_buf0), .C(_2476_), .Y(_80__7_) );
INVX1 INVX1_1300 ( .gnd(gnd), .vdd(vdd), .A(data_171__8_), .Y(_2477_) );
MUX2X1 MUX2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_2477_), .S(_2471__bF_buf3), .Y(_80__8_) );
NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(data_171__9_), .B(_2471__bF_buf2), .Y(_2478_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_2471__bF_buf1), .C(_2478_), .Y(_80__9_) );
NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(data_171__10_), .B(_2471__bF_buf0), .Y(_2479_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_2471__bF_buf3), .C(_2479_), .Y(_80__10_) );
NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(data_171__11_), .B(_2471__bF_buf2), .Y(_2480_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_2471__bF_buf1), .C(_2480_), .Y(_80__11_) );
INVX1 INVX1_1301 ( .gnd(gnd), .vdd(vdd), .A(data_171__12_), .Y(_2481_) );
MUX2X1 MUX2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_2481_), .S(_2471__bF_buf0), .Y(_80__12_) );
NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(data_171__13_), .B(_2471__bF_buf3), .Y(_2482_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_2471__bF_buf2), .C(_2482_), .Y(_80__13_) );
NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(data_171__14_), .B(_2471__bF_buf1), .Y(_2483_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_2471__bF_buf0), .C(_2483_), .Y(_80__14_) );
NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(data_171__15_), .B(_2471__bF_buf3), .Y(_2484_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_2471__bF_buf2), .C(_2484_), .Y(_80__15_) );
INVX1 INVX1_1302 ( .gnd(gnd), .vdd(vdd), .A(data_170__0_), .Y(_2485_) );
NOR3X1 NOR3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_2458_), .B(_2112_), .C(_1810__bF_buf4), .Y(_2486_) );
OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14945_), .C(IDATA_PROG_write_bF_buf7), .Y(_2487_) );
INVX1 INVX1_1303 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .Y(_2488_) );
OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14952__bF_buf3), .C(_2316_), .Y(_2489_) );
OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_2488_), .C(_2489_), .Y(_2490_) );
NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2490_), .B(_1684_), .Y(_2491_) );
AND2X2 AND2X2_606 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(_2491_), .Y(_2492_) );
NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2492_), .B(_2457_), .Y(_2493_) );
MUX2X1 MUX2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2485_), .B(_14932__bF_buf1), .S(_2493_), .Y(_79__0_) );
INVX1 INVX1_1304 ( .gnd(gnd), .vdd(vdd), .A(data_170__1_), .Y(_2494_) );
MUX2X1 MUX2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2494_), .B(_14894__bF_buf0), .S(_2493_), .Y(_79__1_) );
INVX1 INVX1_1305 ( .gnd(gnd), .vdd(vdd), .A(data_170__2_), .Y(_2495_) );
MUX2X1 MUX2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .B(_14897__bF_buf12), .S(_2493_), .Y(_79__2_) );
NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .B(_2486_), .Y(_2496_) );
NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .B(_2470_), .Y(_2497_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2492_), .B(_2457_), .C(data_170__3_), .Y(_2498_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_2497__bF_buf3), .C(_2498_), .Y(_79__3_) );
NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(data_170__4_), .B(_2497__bF_buf2), .Y(_2499_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_2497__bF_buf1), .C(_2499_), .Y(_79__4_) );
NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(data_170__5_), .B(_2497__bF_buf0), .Y(_2500_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_2497__bF_buf3), .C(_2500_), .Y(_79__5_) );
NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(data_170__6_), .B(_2497__bF_buf2), .Y(_2501_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_2497__bF_buf1), .C(_2501_), .Y(_79__6_) );
NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(data_170__7_), .B(_2497__bF_buf0), .Y(_2502_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_2497__bF_buf3), .C(_2502_), .Y(_79__7_) );
INVX1 INVX1_1306 ( .gnd(gnd), .vdd(vdd), .A(data_170__8_), .Y(_2503_) );
MUX2X1 MUX2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_2503_), .S(_2497__bF_buf2), .Y(_79__8_) );
INVX1 INVX1_1307 ( .gnd(gnd), .vdd(vdd), .A(data_170__9_), .Y(_2504_) );
MUX2X1 MUX2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_2504_), .S(_2497__bF_buf1), .Y(_79__9_) );
NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(data_170__10_), .B(_2497__bF_buf0), .Y(_2505_) );
AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_2497__bF_buf3), .C(_2505_), .Y(_79__10_) );
NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(data_170__11_), .B(_2497__bF_buf2), .Y(_2506_) );
AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_2497__bF_buf1), .C(_2506_), .Y(_79__11_) );
NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(data_170__12_), .B(_2497__bF_buf0), .Y(_2507_) );
AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_2497__bF_buf3), .C(_2507_), .Y(_79__12_) );
NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(data_170__13_), .B(_2497__bF_buf2), .Y(_2508_) );
AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_2497__bF_buf1), .C(_2508_), .Y(_79__13_) );
NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(data_170__14_), .B(_2497__bF_buf0), .Y(_2509_) );
AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_2497__bF_buf3), .C(_2509_), .Y(_79__14_) );
NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(data_170__15_), .B(_2497__bF_buf2), .Y(_2510_) );
AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_2497__bF_buf1), .C(_2510_), .Y(_79__15_) );
OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_16055_), .C(_2487_), .Y(_2511_) );
NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2511_), .C(_2486_), .Y(_2512_) );
NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2512_), .Y(_2513_) );
NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(data_169__0_), .B(_2513__bF_buf3), .Y(_2514_) );
AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_2513__bF_buf2), .C(_2514_), .Y(_77__0_) );
INVX1 INVX1_1308 ( .gnd(gnd), .vdd(vdd), .A(data_169__1_), .Y(_2515_) );
MUX2X1 MUX2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_2515_), .S(_2513__bF_buf1), .Y(_77__1_) );
INVX1 INVX1_1309 ( .gnd(gnd), .vdd(vdd), .A(data_169__2_), .Y(_2516_) );
MUX2X1 MUX2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_2516_), .S(_2513__bF_buf0), .Y(_77__2_) );
INVX1 INVX1_1310 ( .gnd(gnd), .vdd(vdd), .A(data_169__3_), .Y(_2517_) );
MUX2X1 MUX2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_2517_), .S(_2513__bF_buf3), .Y(_77__3_) );
INVX1 INVX1_1311 ( .gnd(gnd), .vdd(vdd), .A(data_169__4_), .Y(_2518_) );
MUX2X1 MUX2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_2518_), .S(_2513__bF_buf2), .Y(_77__4_) );
NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(data_169__5_), .B(_2513__bF_buf1), .Y(_2519_) );
AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_2513__bF_buf0), .C(_2519_), .Y(_77__5_) );
INVX1 INVX1_1312 ( .gnd(gnd), .vdd(vdd), .A(data_169__6_), .Y(_2520_) );
MUX2X1 MUX2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_2520_), .S(_2513__bF_buf3), .Y(_77__6_) );
NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(data_169__7_), .B(_2513__bF_buf2), .Y(_2521_) );
AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_2513__bF_buf1), .C(_2521_), .Y(_77__7_) );
NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(data_169__8_), .B(_2513__bF_buf0), .Y(_2522_) );
AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_2513__bF_buf3), .C(_2522_), .Y(_77__8_) );
NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(data_169__9_), .B(_2513__bF_buf2), .Y(_2523_) );
AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_2513__bF_buf1), .C(_2523_), .Y(_77__9_) );
INVX1 INVX1_1313 ( .gnd(gnd), .vdd(vdd), .A(data_169__10_), .Y(_2524_) );
MUX2X1 MUX2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_2524_), .S(_2513__bF_buf0), .Y(_77__10_) );
INVX1 INVX1_1314 ( .gnd(gnd), .vdd(vdd), .A(data_169__11_), .Y(_2525_) );
MUX2X1 MUX2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_2525_), .S(_2513__bF_buf3), .Y(_77__11_) );
NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(data_169__12_), .B(_2513__bF_buf2), .Y(_2526_) );
AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_2513__bF_buf1), .C(_2526_), .Y(_77__12_) );
NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(data_169__13_), .B(_2513__bF_buf0), .Y(_2527_) );
AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_2513__bF_buf3), .C(_2527_), .Y(_77__13_) );
INVX1 INVX1_1315 ( .gnd(gnd), .vdd(vdd), .A(data_169__14_), .Y(_2528_) );
MUX2X1 MUX2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf14), .B(_2528_), .S(_2513__bF_buf2), .Y(_77__14_) );
NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(data_169__15_), .B(_2513__bF_buf1), .Y(_2529_) );
AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_2513__bF_buf0), .C(_2529_), .Y(_77__15_) );
OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf0), .B(_14952__bF_buf2), .C(_2316_), .Y(_2530_) );
NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .B(_2530_), .C(_2113_), .Y(_2531_) );
NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .B(_2470_), .Y(_2532_) );
NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(data_168__0_), .B(_2532__bF_buf3), .Y(_2533_) );
AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_2532__bF_buf2), .C(_2533_), .Y(_76__0_) );
INVX1 INVX1_1316 ( .gnd(gnd), .vdd(vdd), .A(data_168__1_), .Y(_2534_) );
MUX2X1 MUX2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_2534_), .S(_2532__bF_buf1), .Y(_76__1_) );
NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(data_168__2_), .B(_2532__bF_buf0), .Y(_2535_) );
AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_2532__bF_buf3), .C(_2535_), .Y(_76__2_) );
NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(data_168__3_), .B(_2532__bF_buf2), .Y(_2536_) );
AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_2532__bF_buf1), .C(_2536_), .Y(_76__3_) );
INVX1 INVX1_1317 ( .gnd(gnd), .vdd(vdd), .A(data_168__4_), .Y(_2537_) );
MUX2X1 MUX2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_2537_), .S(_2532__bF_buf0), .Y(_76__4_) );
NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(data_168__5_), .B(_2532__bF_buf3), .Y(_2538_) );
AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_2532__bF_buf2), .C(_2538_), .Y(_76__5_) );
INVX1 INVX1_1318 ( .gnd(gnd), .vdd(vdd), .A(data_168__6_), .Y(_2539_) );
MUX2X1 MUX2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_2539_), .S(_2532__bF_buf1), .Y(_76__6_) );
INVX1 INVX1_1319 ( .gnd(gnd), .vdd(vdd), .A(data_168__7_), .Y(_2540_) );
MUX2X1 MUX2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_2540_), .S(_2532__bF_buf0), .Y(_76__7_) );
NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(data_168__8_), .B(_2532__bF_buf3), .Y(_2541_) );
AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_2532__bF_buf2), .C(_2541_), .Y(_76__8_) );
NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(data_168__9_), .B(_2532__bF_buf1), .Y(_2542_) );
AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_2532__bF_buf0), .C(_2542_), .Y(_76__9_) );
INVX1 INVX1_1320 ( .gnd(gnd), .vdd(vdd), .A(data_168__10_), .Y(_2543_) );
MUX2X1 MUX2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_2543_), .S(_2532__bF_buf3), .Y(_76__10_) );
INVX1 INVX1_1321 ( .gnd(gnd), .vdd(vdd), .A(data_168__11_), .Y(_2544_) );
MUX2X1 MUX2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_2544_), .S(_2532__bF_buf2), .Y(_76__11_) );
NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(data_168__12_), .B(_2532__bF_buf1), .Y(_2545_) );
AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_2532__bF_buf0), .C(_2545_), .Y(_76__12_) );
INVX1 INVX1_1322 ( .gnd(gnd), .vdd(vdd), .A(data_168__13_), .Y(_2546_) );
MUX2X1 MUX2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_2546_), .S(_2532__bF_buf3), .Y(_76__13_) );
INVX1 INVX1_1323 ( .gnd(gnd), .vdd(vdd), .A(data_168__14_), .Y(_2547_) );
MUX2X1 MUX2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_2547_), .S(_2532__bF_buf2), .Y(_76__14_) );
INVX1 INVX1_1324 ( .gnd(gnd), .vdd(vdd), .A(data_168__15_), .Y(_2548_) );
MUX2X1 MUX2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_2548_), .S(_2532__bF_buf1), .Y(_76__15_) );
INVX1 INVX1_1325 ( .gnd(gnd), .vdd(vdd), .A(data_167__0_), .Y(_2549_) );
OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_15364_), .B(_847_), .C(_2487_), .Y(_2550_) );
NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2550_), .C(_2486_), .Y(_2551_) );
NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2551_), .Y(_2552_) );
MUX2X1 MUX2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_2549_), .S(_2552__bF_buf3), .Y(_75__0_) );
INVX1 INVX1_1326 ( .gnd(gnd), .vdd(vdd), .A(data_167__1_), .Y(_2553_) );
MUX2X1 MUX2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_2553_), .S(_2552__bF_buf2), .Y(_75__1_) );
NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(data_167__2_), .B(_2552__bF_buf1), .Y(_2554_) );
AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_2552__bF_buf0), .C(_2554_), .Y(_75__2_) );
INVX1 INVX1_1327 ( .gnd(gnd), .vdd(vdd), .A(data_167__3_), .Y(_2555_) );
MUX2X1 MUX2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_2555_), .S(_2552__bF_buf3), .Y(_75__3_) );
INVX1 INVX1_1328 ( .gnd(gnd), .vdd(vdd), .A(data_167__4_), .Y(_2556_) );
MUX2X1 MUX2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_2556_), .S(_2552__bF_buf2), .Y(_75__4_) );
INVX1 INVX1_1329 ( .gnd(gnd), .vdd(vdd), .A(data_167__5_), .Y(_2557_) );
MUX2X1 MUX2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_2557_), .S(_2552__bF_buf1), .Y(_75__5_) );
INVX1 INVX1_1330 ( .gnd(gnd), .vdd(vdd), .A(data_167__6_), .Y(_2558_) );
MUX2X1 MUX2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_2558_), .S(_2552__bF_buf0), .Y(_75__6_) );
NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(data_167__7_), .B(_2552__bF_buf3), .Y(_2559_) );
AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_2552__bF_buf2), .C(_2559_), .Y(_75__7_) );
INVX1 INVX1_1331 ( .gnd(gnd), .vdd(vdd), .A(data_167__8_), .Y(_2560_) );
MUX2X1 MUX2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_2560_), .S(_2552__bF_buf1), .Y(_75__8_) );
NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(data_167__9_), .B(_2552__bF_buf0), .Y(_2561_) );
AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_2552__bF_buf3), .C(_2561_), .Y(_75__9_) );
INVX1 INVX1_1332 ( .gnd(gnd), .vdd(vdd), .A(data_167__10_), .Y(_2562_) );
MUX2X1 MUX2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_2562_), .S(_2552__bF_buf2), .Y(_75__10_) );
INVX1 INVX1_1333 ( .gnd(gnd), .vdd(vdd), .A(data_167__11_), .Y(_2563_) );
MUX2X1 MUX2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_2563_), .S(_2552__bF_buf1), .Y(_75__11_) );
INVX1 INVX1_1334 ( .gnd(gnd), .vdd(vdd), .A(data_167__12_), .Y(_2564_) );
MUX2X1 MUX2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_2564_), .S(_2552__bF_buf0), .Y(_75__12_) );
INVX1 INVX1_1335 ( .gnd(gnd), .vdd(vdd), .A(data_167__13_), .Y(_2565_) );
MUX2X1 MUX2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_2565_), .S(_2552__bF_buf3), .Y(_75__13_) );
INVX1 INVX1_1336 ( .gnd(gnd), .vdd(vdd), .A(data_167__14_), .Y(_2566_) );
MUX2X1 MUX2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_2566_), .S(_2552__bF_buf2), .Y(_75__14_) );
NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(data_167__15_), .B(_2552__bF_buf1), .Y(_2567_) );
AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_2552__bF_buf0), .C(_2567_), .Y(_75__15_) );
INVX1 INVX1_1337 ( .gnd(gnd), .vdd(vdd), .A(data_166__0_), .Y(_2568_) );
OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_2314_), .C(_1686_), .Y(_2569_) );
OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(_2488_), .C(_2569_), .Y(_2570_) );
NOR3X1 NOR3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1684_), .B(_2570_), .C(_2063__bF_buf2), .Y(_2571_) );
NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2457_), .Y(_2572_) );
MUX2X1 MUX2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2568_), .B(_14932__bF_buf12), .S(_2572_), .Y(_74__0_) );
AND2X2 AND2X2_607 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_2571_), .Y(_2573_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf3), .B(data_166__1_), .Y(_2574_) );
NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_2573__bF_buf2), .Y(_2575_) );
AND2X2 AND2X2_608 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .B(_2575_), .Y(_74__1_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf1), .B(data_166__2_), .Y(_2576_) );
NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_2573__bF_buf0), .Y(_2577_) );
AND2X2 AND2X2_609 ( .gnd(gnd), .vdd(vdd), .A(_2576_), .B(_2577_), .Y(_74__2_) );
AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2457_), .C(data_166__3_), .Y(_2578_) );
AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_2573__bF_buf3), .C(_2578_), .Y(_74__3_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf2), .B(data_166__4_), .Y(_2579_) );
NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_2573__bF_buf1), .Y(_2580_) );
AND2X2 AND2X2_610 ( .gnd(gnd), .vdd(vdd), .A(_2579_), .B(_2580_), .Y(_74__4_) );
INVX1 INVX1_1338 ( .gnd(gnd), .vdd(vdd), .A(data_166__5_), .Y(_2581_) );
MUX2X1 MUX2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .B(_14903__bF_buf5), .S(_2572_), .Y(_74__5_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf0), .B(data_166__6_), .Y(_2582_) );
NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_2573__bF_buf3), .Y(_2583_) );
AND2X2 AND2X2_611 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .B(_2583_), .Y(_74__6_) );
INVX1 INVX1_1339 ( .gnd(gnd), .vdd(vdd), .A(data_166__7_), .Y(_2584_) );
MUX2X1 MUX2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .B(_14908__bF_buf4), .S(_2572_), .Y(_74__7_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf2), .B(data_166__8_), .Y(_2585_) );
NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_2573__bF_buf1), .Y(_2586_) );
AND2X2 AND2X2_612 ( .gnd(gnd), .vdd(vdd), .A(_2585_), .B(_2586_), .Y(_74__8_) );
INVX1 INVX1_1340 ( .gnd(gnd), .vdd(vdd), .A(data_166__9_), .Y(_2587_) );
MUX2X1 MUX2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_14913__bF_buf8), .S(_2572_), .Y(_74__9_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf0), .B(data_166__10_), .Y(_2588_) );
NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_2573__bF_buf3), .Y(_2589_) );
AND2X2 AND2X2_613 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2589_), .Y(_74__10_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf2), .B(data_166__11_), .Y(_2590_) );
NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_2573__bF_buf1), .Y(_2591_) );
AND2X2 AND2X2_614 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(_2591_), .Y(_74__11_) );
INVX1 INVX1_1341 ( .gnd(gnd), .vdd(vdd), .A(data_166__12_), .Y(_2592_) );
MUX2X1 MUX2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2592_), .B(_14920__bF_buf5), .S(_2572_), .Y(_74__12_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf0), .B(data_166__13_), .Y(_2593_) );
NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_2573__bF_buf3), .Y(_2594_) );
AND2X2 AND2X2_615 ( .gnd(gnd), .vdd(vdd), .A(_2593_), .B(_2594_), .Y(_74__13_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_2573__bF_buf2), .B(data_166__14_), .Y(_2595_) );
NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_2573__bF_buf1), .Y(_2596_) );
AND2X2 AND2X2_616 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(_2596_), .Y(_74__14_) );
INVX1 INVX1_1342 ( .gnd(gnd), .vdd(vdd), .A(data_166__15_), .Y(_2597_) );
MUX2X1 MUX2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_15062__bF_buf4), .S(_2572_), .Y(_74__15_) );
NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf2), .B(_15453_), .Y(_2598_) );
AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .B(_1482_), .C(_2598_), .Y(_2599_) );
NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2599_), .C(_2486_), .Y(_2600_) );
NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2600_), .Y(_2601_) );
NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(data_165__0_), .B(_2601__bF_buf4), .Y(_2602_) );
AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_2601__bF_buf3), .C(_2602_), .Y(_73__0_) );
NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(data_165__1_), .B(_2601__bF_buf2), .Y(_2603_) );
AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_2601__bF_buf1), .C(_2603_), .Y(_73__1_) );
NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(data_165__2_), .B(_2601__bF_buf0), .Y(_2604_) );
AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_2601__bF_buf4), .C(_2604_), .Y(_73__2_) );
INVX1 INVX1_1343 ( .gnd(gnd), .vdd(vdd), .A(data_165__3_), .Y(_2605_) );
MUX2X1 MUX2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_2605_), .S(_2601__bF_buf3), .Y(_73__3_) );
NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(data_165__4_), .B(_2601__bF_buf2), .Y(_2606_) );
AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_2601__bF_buf1), .C(_2606_), .Y(_73__4_) );
NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(data_165__5_), .B(_2601__bF_buf0), .Y(_2607_) );
AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_2601__bF_buf4), .C(_2607_), .Y(_73__5_) );
NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(data_165__6_), .B(_2601__bF_buf3), .Y(_2608_) );
AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_2601__bF_buf2), .C(_2608_), .Y(_73__6_) );
INVX1 INVX1_1344 ( .gnd(gnd), .vdd(vdd), .A(data_165__7_), .Y(_2609_) );
MUX2X1 MUX2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_2609_), .S(_2601__bF_buf1), .Y(_73__7_) );
NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(data_165__8_), .B(_2601__bF_buf0), .Y(_2610_) );
AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_2601__bF_buf4), .C(_2610_), .Y(_73__8_) );
INVX1 INVX1_1345 ( .gnd(gnd), .vdd(vdd), .A(data_165__9_), .Y(_2611_) );
MUX2X1 MUX2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf7), .B(_2611_), .S(_2601__bF_buf3), .Y(_73__9_) );
NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(data_165__10_), .B(_2601__bF_buf2), .Y(_2612_) );
AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_2601__bF_buf1), .C(_2612_), .Y(_73__10_) );
NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(data_165__11_), .B(_2601__bF_buf0), .Y(_2613_) );
AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_2601__bF_buf4), .C(_2613_), .Y(_73__11_) );
NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(data_165__12_), .B(_2601__bF_buf3), .Y(_2614_) );
AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_2601__bF_buf2), .C(_2614_), .Y(_73__12_) );
NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(data_165__13_), .B(_2601__bF_buf1), .Y(_2615_) );
AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_2601__bF_buf0), .C(_2615_), .Y(_73__13_) );
NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(data_165__14_), .B(_2601__bF_buf4), .Y(_2616_) );
AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_2601__bF_buf3), .C(_2616_), .Y(_73__14_) );
INVX1 INVX1_1346 ( .gnd(gnd), .vdd(vdd), .A(data_165__15_), .Y(_2617_) );
MUX2X1 MUX2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_2617_), .S(_2601__bF_buf2), .Y(_73__15_) );
INVX1 INVX1_1347 ( .gnd(gnd), .vdd(vdd), .A(data_164__0_), .Y(_2618_) );
NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .B(_2113_), .Y(_2619_) );
OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14965__bF_buf3), .C(_2316_), .Y(_2620_) );
NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .B(_2620_), .C(_2380_), .Y(_2621_) );
OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf7), .B(_2619__bF_buf3), .C(_2618_), .Y(_2622_) );
NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_2619__bF_buf2), .B(_2621__bF_buf6), .Y(_2623_) );
NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_2623_), .Y(_2624_) );
AND2X2 AND2X2_617 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .B(_2622_), .Y(_72__0_) );
INVX1 INVX1_1348 ( .gnd(gnd), .vdd(vdd), .A(data_164__1_), .Y(_2625_) );
OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf5), .B(_2619__bF_buf1), .C(_2625_), .Y(_2626_) );
NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_2623_), .Y(_2627_) );
AND2X2 AND2X2_618 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .B(_2626_), .Y(_72__1_) );
INVX1 INVX1_1349 ( .gnd(gnd), .vdd(vdd), .A(data_164__2_), .Y(_2628_) );
OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf4), .B(_2619__bF_buf0), .C(_2628_), .Y(_2629_) );
NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_2623_), .Y(_2630_) );
AND2X2 AND2X2_619 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2629_), .Y(_72__2_) );
INVX1 INVX1_1350 ( .gnd(gnd), .vdd(vdd), .A(data_164__3_), .Y(_2631_) );
OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf3), .B(_2619__bF_buf3), .C(_2631_), .Y(_2632_) );
NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_2623_), .Y(_2633_) );
AND2X2 AND2X2_620 ( .gnd(gnd), .vdd(vdd), .A(_2633_), .B(_2632_), .Y(_72__3_) );
INVX1 INVX1_1351 ( .gnd(gnd), .vdd(vdd), .A(data_164__4_), .Y(_2634_) );
OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf2), .B(_2619__bF_buf2), .C(_2634_), .Y(_2635_) );
NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_2623_), .Y(_2636_) );
AND2X2 AND2X2_621 ( .gnd(gnd), .vdd(vdd), .A(_2636_), .B(_2635_), .Y(_72__4_) );
INVX1 INVX1_1352 ( .gnd(gnd), .vdd(vdd), .A(data_164__5_), .Y(_2637_) );
OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf1), .B(_2619__bF_buf1), .C(_2637_), .Y(_2638_) );
NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_2623_), .Y(_2639_) );
AND2X2 AND2X2_622 ( .gnd(gnd), .vdd(vdd), .A(_2639_), .B(_2638_), .Y(_72__5_) );
INVX1 INVX1_1353 ( .gnd(gnd), .vdd(vdd), .A(data_164__6_), .Y(_2640_) );
OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf0), .B(_2619__bF_buf0), .C(_2640_), .Y(_2641_) );
NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_2623_), .Y(_2642_) );
AND2X2 AND2X2_623 ( .gnd(gnd), .vdd(vdd), .A(_2642_), .B(_2641_), .Y(_72__6_) );
INVX1 INVX1_1354 ( .gnd(gnd), .vdd(vdd), .A(data_164__7_), .Y(_2643_) );
OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf7), .B(_2619__bF_buf3), .C(_2643_), .Y(_2644_) );
NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_2623_), .Y(_2645_) );
AND2X2 AND2X2_624 ( .gnd(gnd), .vdd(vdd), .A(_2645_), .B(_2644_), .Y(_72__7_) );
INVX1 INVX1_1355 ( .gnd(gnd), .vdd(vdd), .A(data_164__8_), .Y(_2646_) );
OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf6), .B(_2619__bF_buf2), .C(_2646_), .Y(_2647_) );
NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_2623_), .Y(_2648_) );
AND2X2 AND2X2_625 ( .gnd(gnd), .vdd(vdd), .A(_2648_), .B(_2647_), .Y(_72__8_) );
INVX1 INVX1_1356 ( .gnd(gnd), .vdd(vdd), .A(data_164__9_), .Y(_2649_) );
OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf5), .B(_2619__bF_buf1), .C(_2649_), .Y(_2650_) );
NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_2623_), .Y(_2651_) );
AND2X2 AND2X2_626 ( .gnd(gnd), .vdd(vdd), .A(_2651_), .B(_2650_), .Y(_72__9_) );
INVX1 INVX1_1357 ( .gnd(gnd), .vdd(vdd), .A(data_164__10_), .Y(_2652_) );
OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf4), .B(_2619__bF_buf0), .C(_2652_), .Y(_2653_) );
NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf3), .B(_2623_), .Y(_2654_) );
AND2X2 AND2X2_627 ( .gnd(gnd), .vdd(vdd), .A(_2654_), .B(_2653_), .Y(_72__10_) );
INVX1 INVX1_1358 ( .gnd(gnd), .vdd(vdd), .A(data_164__11_), .Y(_2655_) );
OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf3), .B(_2619__bF_buf3), .C(_2655_), .Y(_2656_) );
NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_2623_), .Y(_2657_) );
AND2X2 AND2X2_628 ( .gnd(gnd), .vdd(vdd), .A(_2657_), .B(_2656_), .Y(_72__11_) );
INVX1 INVX1_1359 ( .gnd(gnd), .vdd(vdd), .A(data_164__12_), .Y(_2658_) );
OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf2), .B(_2619__bF_buf2), .C(_2658_), .Y(_2659_) );
NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_2623_), .Y(_2660_) );
AND2X2 AND2X2_629 ( .gnd(gnd), .vdd(vdd), .A(_2660_), .B(_2659_), .Y(_72__12_) );
INVX1 INVX1_1360 ( .gnd(gnd), .vdd(vdd), .A(data_164__13_), .Y(_2661_) );
OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf1), .B(_2619__bF_buf1), .C(_2661_), .Y(_2662_) );
NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_2623_), .Y(_2663_) );
AND2X2 AND2X2_630 ( .gnd(gnd), .vdd(vdd), .A(_2663_), .B(_2662_), .Y(_72__13_) );
INVX1 INVX1_1361 ( .gnd(gnd), .vdd(vdd), .A(data_164__14_), .Y(_2664_) );
OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf0), .B(_2619__bF_buf0), .C(_2664_), .Y(_2665_) );
NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_2623_), .Y(_2666_) );
AND2X2 AND2X2_631 ( .gnd(gnd), .vdd(vdd), .A(_2666_), .B(_2665_), .Y(_72__14_) );
INVX1 INVX1_1362 ( .gnd(gnd), .vdd(vdd), .A(data_164__15_), .Y(_2667_) );
OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf7), .B(_2619__bF_buf3), .C(_2667_), .Y(_2668_) );
NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf2), .B(_2623_), .Y(_2669_) );
AND2X2 AND2X2_632 ( .gnd(gnd), .vdd(vdd), .A(_2669_), .B(_2668_), .Y(_72__15_) );
INVX1 INVX1_1363 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2670_) );
NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_2670_), .B(_2470_), .Y(_2671_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .Y(_2672_) );
OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_2672_), .B(_15763_), .C(_14941_), .Y(_2673_) );
OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_15571_), .B(_15019__bF_buf1), .C(_2673_), .Y(_2674_) );
INVX1 INVX1_1364 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .Y(_2675_) );
OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf0), .B(_15581_), .C(_2675_), .Y(_2676_) );
OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf2), .B(_15034_), .C(IDATA_PROG_write_bF_buf6), .Y(_2677_) );
NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2677_), .B(_1684_), .Y(_2678_) );
NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2113_), .Y(_2679_) );
NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2679_), .Y(_2680_) );
NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2680_), .B(_2671_), .Y(_2681_) );
INVX1 INVX1_1365 ( .gnd(gnd), .vdd(vdd), .A(data_163__0_), .Y(_2682_) );
INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(_2680_), .Y(_2683_) );
OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf6), .C(_2682_), .Y(_2684_) );
OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf1), .B(_2681_), .C(_2684_), .Y(_2685_) );
INVX1 INVX1_1366 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .Y(_71__0_) );
INVX1 INVX1_1367 ( .gnd(gnd), .vdd(vdd), .A(data_163__1_), .Y(_2686_) );
OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf5), .C(_2686_), .Y(_2687_) );
OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf2), .B(_2681_), .C(_2687_), .Y(_2688_) );
INVX1 INVX1_1368 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .Y(_71__1_) );
INVX1 INVX1_1369 ( .gnd(gnd), .vdd(vdd), .A(data_163__2_), .Y(_2689_) );
OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf4), .C(_2689_), .Y(_2690_) );
OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf2), .B(_2681_), .C(_2690_), .Y(_2691_) );
INVX1 INVX1_1370 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .Y(_71__2_) );
INVX1 INVX1_1371 ( .gnd(gnd), .vdd(vdd), .A(data_163__3_), .Y(_2692_) );
OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf3), .C(_2692_), .Y(_2693_) );
NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_2680_), .C(_2671_), .Y(_2694_) );
AND2X2 AND2X2_633 ( .gnd(gnd), .vdd(vdd), .A(_2693_), .B(_2694_), .Y(_71__3_) );
INVX1 INVX1_1372 ( .gnd(gnd), .vdd(vdd), .A(data_163__4_), .Y(_2695_) );
OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf2), .C(_2695_), .Y(_2696_) );
OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf3), .B(_2681_), .C(_2696_), .Y(_2697_) );
INVX1 INVX1_1373 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .Y(_71__4_) );
INVX1 INVX1_1374 ( .gnd(gnd), .vdd(vdd), .A(data_163__5_), .Y(_2698_) );
OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf1), .C(_2698_), .Y(_2699_) );
OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf2), .B(_2681_), .C(_2699_), .Y(_2700_) );
INVX1 INVX1_1375 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .Y(_71__5_) );
INVX1 INVX1_1376 ( .gnd(gnd), .vdd(vdd), .A(data_163__6_), .Y(_2701_) );
OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf0), .C(_2701_), .Y(_2702_) );
OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf0), .B(_2681_), .C(_2702_), .Y(_2703_) );
INVX1 INVX1_1377 ( .gnd(gnd), .vdd(vdd), .A(_2703_), .Y(_71__6_) );
INVX1 INVX1_1378 ( .gnd(gnd), .vdd(vdd), .A(data_163__7_), .Y(_2704_) );
OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf7), .C(_2704_), .Y(_2705_) );
OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf0), .B(_2681_), .C(_2705_), .Y(_2706_) );
INVX1 INVX1_1379 ( .gnd(gnd), .vdd(vdd), .A(_2706_), .Y(_71__7_) );
INVX1 INVX1_1380 ( .gnd(gnd), .vdd(vdd), .A(data_163__8_), .Y(_2707_) );
OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf6), .C(_2707_), .Y(_2708_) );
OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf2), .B(_2681_), .C(_2708_), .Y(_2709_) );
INVX1 INVX1_1381 ( .gnd(gnd), .vdd(vdd), .A(_2709_), .Y(_71__8_) );
INVX1 INVX1_1382 ( .gnd(gnd), .vdd(vdd), .A(data_163__9_), .Y(_2710_) );
OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf5), .C(_2710_), .Y(_2711_) );
OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf0), .B(_2681_), .C(_2711_), .Y(_2712_) );
INVX1 INVX1_1383 ( .gnd(gnd), .vdd(vdd), .A(_2712_), .Y(_71__9_) );
INVX1 INVX1_1384 ( .gnd(gnd), .vdd(vdd), .A(data_163__10_), .Y(_2713_) );
OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf4), .C(_2713_), .Y(_2714_) );
OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf2), .B(_2681_), .C(_2714_), .Y(_2715_) );
INVX1 INVX1_1385 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .Y(_71__10_) );
INVX1 INVX1_1386 ( .gnd(gnd), .vdd(vdd), .A(data_163__11_), .Y(_2716_) );
OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf3), .C(_2716_), .Y(_2717_) );
OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf1), .B(_2681_), .C(_2717_), .Y(_2718_) );
INVX1 INVX1_1387 ( .gnd(gnd), .vdd(vdd), .A(_2718_), .Y(_71__11_) );
INVX1 INVX1_1388 ( .gnd(gnd), .vdd(vdd), .A(data_163__12_), .Y(_2719_) );
OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf2), .C(_2719_), .Y(_2720_) );
OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf2), .B(_2681_), .C(_2720_), .Y(_2721_) );
INVX1 INVX1_1389 ( .gnd(gnd), .vdd(vdd), .A(_2721_), .Y(_71__12_) );
INVX1 INVX1_1390 ( .gnd(gnd), .vdd(vdd), .A(data_163__13_), .Y(_2722_) );
OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf1), .C(_2722_), .Y(_2723_) );
OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf3), .B(_2681_), .C(_2723_), .Y(_2724_) );
INVX1 INVX1_1391 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .Y(_71__13_) );
INVX1 INVX1_1392 ( .gnd(gnd), .vdd(vdd), .A(data_163__14_), .Y(_2725_) );
OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf0), .C(_2725_), .Y(_2726_) );
OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf2), .B(_2681_), .C(_2726_), .Y(_2727_) );
INVX1 INVX1_1393 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .Y(_71__14_) );
INVX1 INVX1_1394 ( .gnd(gnd), .vdd(vdd), .A(data_163__15_), .Y(_2728_) );
OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2621__bF_buf7), .C(_2728_), .Y(_2729_) );
OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf0), .B(_2681_), .C(_2729_), .Y(_2730_) );
INVX1 INVX1_1395 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .Y(_71__15_) );
NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2113_), .Y(_2731_) );
INVX1 INVX1_1396 ( .gnd(gnd), .vdd(vdd), .A(_2677_), .Y(_2732_) );
OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_15019__bF_buf3), .C(_2732_), .Y(_2733_) );
INVX1 INVX1_1397 ( .gnd(gnd), .vdd(vdd), .A(_2733_), .Y(_2734_) );
NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_2675_), .Y(_2735_) );
NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_2735_), .B(_2731_), .Y(_2736_) );
NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(_2671_), .Y(_2737_) );
INVX1 INVX1_1398 ( .gnd(gnd), .vdd(vdd), .A(data_162__0_), .Y(_2738_) );
INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .Y(_2739_) );
OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf6), .C(_2738_), .Y(_2740_) );
OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf0), .B(_2737_), .C(_2740_), .Y(_2741_) );
INVX1 INVX1_1399 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .Y(_70__0_) );
INVX1 INVX1_1400 ( .gnd(gnd), .vdd(vdd), .A(data_162__1_), .Y(_2742_) );
OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf5), .C(_2742_), .Y(_2743_) );
OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf1), .B(_2737_), .C(_2743_), .Y(_2744_) );
INVX1 INVX1_1401 ( .gnd(gnd), .vdd(vdd), .A(_2744_), .Y(_70__1_) );
INVX1 INVX1_1402 ( .gnd(gnd), .vdd(vdd), .A(data_162__2_), .Y(_2745_) );
OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf4), .C(_2745_), .Y(_2746_) );
OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf1), .B(_2737_), .C(_2746_), .Y(_2747_) );
INVX1 INVX1_1403 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .Y(_70__2_) );
INVX1 INVX1_1404 ( .gnd(gnd), .vdd(vdd), .A(data_162__3_), .Y(_2748_) );
OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf3), .C(_2748_), .Y(_2749_) );
NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_2736_), .C(_2671_), .Y(_2750_) );
AND2X2 AND2X2_634 ( .gnd(gnd), .vdd(vdd), .A(_2749_), .B(_2750_), .Y(_70__3_) );
INVX1 INVX1_1405 ( .gnd(gnd), .vdd(vdd), .A(data_162__4_), .Y(_2751_) );
OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf2), .C(_2751_), .Y(_2752_) );
OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf2), .B(_2737_), .C(_2752_), .Y(_2753_) );
INVX1 INVX1_1406 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .Y(_70__4_) );
INVX1 INVX1_1407 ( .gnd(gnd), .vdd(vdd), .A(data_162__5_), .Y(_2754_) );
OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf1), .C(_2754_), .Y(_2755_) );
OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf1), .B(_2737_), .C(_2755_), .Y(_2756_) );
INVX1 INVX1_1408 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .Y(_70__5_) );
INVX1 INVX1_1409 ( .gnd(gnd), .vdd(vdd), .A(data_162__6_), .Y(_2757_) );
OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf0), .C(_2757_), .Y(_2758_) );
OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf4), .B(_2737_), .C(_2758_), .Y(_2759_) );
INVX1 INVX1_1410 ( .gnd(gnd), .vdd(vdd), .A(_2759_), .Y(_70__6_) );
INVX1 INVX1_1411 ( .gnd(gnd), .vdd(vdd), .A(data_162__7_), .Y(_2760_) );
OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf7), .C(_2760_), .Y(_2761_) );
OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf5), .B(_2737_), .C(_2761_), .Y(_2762_) );
INVX1 INVX1_1412 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .Y(_70__7_) );
INVX1 INVX1_1413 ( .gnd(gnd), .vdd(vdd), .A(data_162__8_), .Y(_2763_) );
OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf6), .C(_2763_), .Y(_2764_) );
OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf1), .B(_2737_), .C(_2764_), .Y(_2765_) );
INVX1 INVX1_1414 ( .gnd(gnd), .vdd(vdd), .A(_2765_), .Y(_70__8_) );
INVX1 INVX1_1415 ( .gnd(gnd), .vdd(vdd), .A(data_162__9_), .Y(_2766_) );
OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf5), .C(_2766_), .Y(_2767_) );
OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf4), .B(_2737_), .C(_2767_), .Y(_2768_) );
INVX1 INVX1_1416 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .Y(_70__9_) );
INVX1 INVX1_1417 ( .gnd(gnd), .vdd(vdd), .A(data_162__10_), .Y(_2769_) );
OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf4), .C(_2769_), .Y(_2770_) );
OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf1), .B(_2737_), .C(_2770_), .Y(_2771_) );
INVX1 INVX1_1418 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .Y(_70__10_) );
INVX1 INVX1_1419 ( .gnd(gnd), .vdd(vdd), .A(data_162__11_), .Y(_2772_) );
OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf3), .C(_2772_), .Y(_2773_) );
OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf0), .B(_2737_), .C(_2773_), .Y(_2774_) );
INVX1 INVX1_1420 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .Y(_70__11_) );
INVX1 INVX1_1421 ( .gnd(gnd), .vdd(vdd), .A(data_162__12_), .Y(_2775_) );
OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf2), .C(_2775_), .Y(_2776_) );
OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf1), .B(_2737_), .C(_2776_), .Y(_2777_) );
INVX1 INVX1_1422 ( .gnd(gnd), .vdd(vdd), .A(_2777_), .Y(_70__12_) );
INVX1 INVX1_1423 ( .gnd(gnd), .vdd(vdd), .A(data_162__13_), .Y(_2778_) );
OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf1), .C(_2778_), .Y(_2779_) );
OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf2), .B(_2737_), .C(_2779_), .Y(_2780_) );
INVX1 INVX1_1424 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .Y(_70__13_) );
INVX1 INVX1_1425 ( .gnd(gnd), .vdd(vdd), .A(data_162__14_), .Y(_2781_) );
OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf0), .C(_2781_), .Y(_2782_) );
OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf1), .B(_2737_), .C(_2782_), .Y(_2783_) );
INVX1 INVX1_1426 ( .gnd(gnd), .vdd(vdd), .A(_2783_), .Y(_70__14_) );
INVX1 INVX1_1427 ( .gnd(gnd), .vdd(vdd), .A(data_162__15_), .Y(_2784_) );
OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2621__bF_buf7), .C(_2784_), .Y(_2785_) );
OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf5), .B(_2737_), .C(_2785_), .Y(_2786_) );
INVX1 INVX1_1428 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .Y(_70__15_) );
INVX1 INVX1_1429 ( .gnd(gnd), .vdd(vdd), .A(data_161__0_), .Y(_2787_) );
INVX1 INVX1_1430 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2788_) );
OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_15019__bF_buf2), .B(_475_), .C(_2673_), .Y(_2789_) );
NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_2733_), .B(_2789_), .Y(_2790_) );
NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_2788_), .Y(_2791_) );
OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf3), .B(_2621__bF_buf6), .C(_2787_), .Y(_2792_) );
NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf5), .B(_2791__bF_buf2), .Y(_2793_) );
NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_2793_), .Y(_2794_) );
AND2X2 AND2X2_635 ( .gnd(gnd), .vdd(vdd), .A(_2794_), .B(_2792_), .Y(_69__0_) );
INVX1 INVX1_1431 ( .gnd(gnd), .vdd(vdd), .A(data_161__1_), .Y(_2795_) );
OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf1), .B(_2621__bF_buf4), .C(_2795_), .Y(_2796_) );
NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_2793_), .Y(_2797_) );
AND2X2 AND2X2_636 ( .gnd(gnd), .vdd(vdd), .A(_2797_), .B(_2796_), .Y(_69__1_) );
INVX1 INVX1_1432 ( .gnd(gnd), .vdd(vdd), .A(data_161__2_), .Y(_2798_) );
OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf0), .B(_2621__bF_buf3), .C(_2798_), .Y(_2799_) );
NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_2793_), .Y(_2800_) );
AND2X2 AND2X2_637 ( .gnd(gnd), .vdd(vdd), .A(_2800_), .B(_2799_), .Y(_69__2_) );
INVX1 INVX1_1433 ( .gnd(gnd), .vdd(vdd), .A(data_161__3_), .Y(_2801_) );
OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf3), .B(_2621__bF_buf2), .C(_2801_), .Y(_2802_) );
AND2X2 AND2X2_638 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_2790_), .Y(_2803_) );
NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_2671_), .C(_2803_), .Y(_2804_) );
AND2X2 AND2X2_639 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .B(_2802_), .Y(_69__3_) );
INVX1 INVX1_1434 ( .gnd(gnd), .vdd(vdd), .A(data_161__4_), .Y(_2805_) );
OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf2), .B(_2621__bF_buf1), .C(_2805_), .Y(_2806_) );
NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_2793_), .Y(_2807_) );
AND2X2 AND2X2_640 ( .gnd(gnd), .vdd(vdd), .A(_2807_), .B(_2806_), .Y(_69__4_) );
INVX1 INVX1_1435 ( .gnd(gnd), .vdd(vdd), .A(data_161__5_), .Y(_2808_) );
OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf1), .B(_2621__bF_buf0), .C(_2808_), .Y(_2809_) );
NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_2793_), .Y(_2810_) );
AND2X2 AND2X2_641 ( .gnd(gnd), .vdd(vdd), .A(_2810_), .B(_2809_), .Y(_69__5_) );
INVX1 INVX1_1436 ( .gnd(gnd), .vdd(vdd), .A(data_161__6_), .Y(_2811_) );
OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf0), .B(_2621__bF_buf7), .C(_2811_), .Y(_2812_) );
NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_2793_), .Y(_2813_) );
AND2X2 AND2X2_642 ( .gnd(gnd), .vdd(vdd), .A(_2813_), .B(_2812_), .Y(_69__6_) );
INVX1 INVX1_1437 ( .gnd(gnd), .vdd(vdd), .A(data_161__7_), .Y(_2814_) );
OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf3), .B(_2621__bF_buf6), .C(_2814_), .Y(_2815_) );
NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_2793_), .Y(_2816_) );
AND2X2 AND2X2_643 ( .gnd(gnd), .vdd(vdd), .A(_2816_), .B(_2815_), .Y(_69__7_) );
INVX1 INVX1_1438 ( .gnd(gnd), .vdd(vdd), .A(data_161__8_), .Y(_2817_) );
OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf2), .B(_2621__bF_buf5), .C(_2817_), .Y(_2818_) );
NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_2793_), .Y(_2819_) );
AND2X2 AND2X2_644 ( .gnd(gnd), .vdd(vdd), .A(_2819_), .B(_2818_), .Y(_69__8_) );
INVX1 INVX1_1439 ( .gnd(gnd), .vdd(vdd), .A(data_161__9_), .Y(_2820_) );
OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf1), .B(_2621__bF_buf4), .C(_2820_), .Y(_2821_) );
NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_2793_), .Y(_2822_) );
AND2X2 AND2X2_645 ( .gnd(gnd), .vdd(vdd), .A(_2822_), .B(_2821_), .Y(_69__9_) );
INVX1 INVX1_1440 ( .gnd(gnd), .vdd(vdd), .A(data_161__10_), .Y(_2823_) );
OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf0), .B(_2621__bF_buf3), .C(_2823_), .Y(_2824_) );
NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_2793_), .Y(_2825_) );
AND2X2 AND2X2_646 ( .gnd(gnd), .vdd(vdd), .A(_2825_), .B(_2824_), .Y(_69__10_) );
INVX1 INVX1_1441 ( .gnd(gnd), .vdd(vdd), .A(data_161__11_), .Y(_2826_) );
OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf3), .B(_2621__bF_buf2), .C(_2826_), .Y(_2827_) );
NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_2793_), .Y(_2828_) );
AND2X2 AND2X2_647 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .B(_2827_), .Y(_69__11_) );
INVX1 INVX1_1442 ( .gnd(gnd), .vdd(vdd), .A(data_161__12_), .Y(_2829_) );
OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf2), .B(_2621__bF_buf1), .C(_2829_), .Y(_2830_) );
NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_2793_), .Y(_2831_) );
AND2X2 AND2X2_648 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_2830_), .Y(_69__12_) );
INVX1 INVX1_1443 ( .gnd(gnd), .vdd(vdd), .A(data_161__13_), .Y(_2832_) );
OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf1), .B(_2621__bF_buf0), .C(_2832_), .Y(_2833_) );
NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_2793_), .Y(_2834_) );
AND2X2 AND2X2_649 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2833_), .Y(_69__13_) );
INVX1 INVX1_1444 ( .gnd(gnd), .vdd(vdd), .A(data_161__14_), .Y(_2835_) );
OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf0), .B(_2621__bF_buf7), .C(_2835_), .Y(_2836_) );
NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_2793_), .Y(_2837_) );
AND2X2 AND2X2_650 ( .gnd(gnd), .vdd(vdd), .A(_2837_), .B(_2836_), .Y(_69__14_) );
INVX1 INVX1_1445 ( .gnd(gnd), .vdd(vdd), .A(data_161__15_), .Y(_2838_) );
OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_2791__bF_buf3), .B(_2621__bF_buf6), .C(_2838_), .Y(_2839_) );
NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_2793_), .Y(_2840_) );
AND2X2 AND2X2_651 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(_2839_), .Y(_69__15_) );
INVX1 INVX1_1446 ( .gnd(gnd), .vdd(vdd), .A(data_160__0_), .Y(_2841_) );
OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_15019__bF_buf1), .C(_15021_), .Y(_2842_) );
INVX1 INVX1_1447 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .Y(_2843_) );
NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_2843_), .C(_2113_), .Y(_2844_) );
NOR3X1 NOR3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_2670_), .B(_2844_), .C(_2470_), .Y(_2845_) );
NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf5), .B(_2845_), .Y(_2846_) );
MUX2X1 MUX2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2841_), .B(_14932__bF_buf8), .S(_2846_), .Y(_68__0_) );
INVX1 INVX1_1448 ( .gnd(gnd), .vdd(vdd), .A(data_160__1_), .Y(_2847_) );
MUX2X1 MUX2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_14894__bF_buf7), .S(_2846_), .Y(_68__1_) );
INVX1 INVX1_1449 ( .gnd(gnd), .vdd(vdd), .A(data_160__2_), .Y(_2848_) );
MUX2X1 MUX2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2848_), .B(_14897__bF_buf4), .S(_2846_), .Y(_68__2_) );
INVX1 INVX1_1450 ( .gnd(gnd), .vdd(vdd), .A(data_160__3_), .Y(_2849_) );
INVX1 INVX1_1451 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .Y(_2850_) );
NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_2620_), .C(_2850_), .Y(_2851_) );
OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_2851_), .B(_14882__bF_buf14_bF_buf3), .C(_2849_), .Y(_2852_) );
NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_14899__bF_buf4), .C(_2845_), .Y(_2853_) );
AND2X2 AND2X2_652 ( .gnd(gnd), .vdd(vdd), .A(_2852_), .B(_2853_), .Y(_68__3_) );
INVX1 INVX1_1452 ( .gnd(gnd), .vdd(vdd), .A(data_160__4_), .Y(_2854_) );
MUX2X1 MUX2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2854_), .B(_14902__bF_buf0), .S(_2846_), .Y(_68__4_) );
INVX1 INVX1_1453 ( .gnd(gnd), .vdd(vdd), .A(data_160__5_), .Y(_2855_) );
MUX2X1 MUX2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_14903__bF_buf1), .S(_2846_), .Y(_68__5_) );
INVX1 INVX1_1454 ( .gnd(gnd), .vdd(vdd), .A(data_160__6_), .Y(_2856_) );
MUX2X1 MUX2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2856_), .B(_15049__bF_buf4), .S(_2846_), .Y(_68__6_) );
INVX1 INVX1_1455 ( .gnd(gnd), .vdd(vdd), .A(data_160__7_), .Y(_2857_) );
MUX2X1 MUX2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_14908__bF_buf0), .S(_2846_), .Y(_68__7_) );
INVX1 INVX1_1456 ( .gnd(gnd), .vdd(vdd), .A(data_160__8_), .Y(_2858_) );
MUX2X1 MUX2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2858_), .B(_15052__bF_buf1), .S(_2846_), .Y(_68__8_) );
INVX1 INVX1_1457 ( .gnd(gnd), .vdd(vdd), .A(data_160__9_), .Y(_2859_) );
MUX2X1 MUX2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .B(_14913__bF_buf4), .S(_2846_), .Y(_68__9_) );
INVX1 INVX1_1458 ( .gnd(gnd), .vdd(vdd), .A(data_160__10_), .Y(_2860_) );
MUX2X1 MUX2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2860_), .B(_15055__bF_buf1), .S(_2846_), .Y(_68__10_) );
INVX1 INVX1_1459 ( .gnd(gnd), .vdd(vdd), .A(data_160__11_), .Y(_2861_) );
MUX2X1 MUX2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2861_), .B(_14918__bF_buf2), .S(_2846_), .Y(_68__11_) );
INVX1 INVX1_1460 ( .gnd(gnd), .vdd(vdd), .A(data_160__12_), .Y(_2862_) );
MUX2X1 MUX2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .B(_14920__bF_buf1), .S(_2846_), .Y(_68__12_) );
INVX1 INVX1_1461 ( .gnd(gnd), .vdd(vdd), .A(data_160__13_), .Y(_2863_) );
MUX2X1 MUX2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_2863_), .B(_14924__bF_buf0), .S(_2846_), .Y(_68__13_) );
INVX1 INVX1_1462 ( .gnd(gnd), .vdd(vdd), .A(data_160__14_), .Y(_2864_) );
MUX2X1 MUX2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .B(_15060__bF_buf7), .S(_2846_), .Y(_68__14_) );
INVX1 INVX1_1463 ( .gnd(gnd), .vdd(vdd), .A(data_160__15_), .Y(_2865_) );
MUX2X1 MUX2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2865_), .B(_15062__bF_buf0), .S(_2846_), .Y(_68__15_) );
OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf2), .B(_14975_), .C(_2316_), .Y(_2866_) );
OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_15066__bF_buf1), .C(_2866_), .Y(_2867_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .B(_2867_), .Y(_2868_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf5), .B(_2868_), .Y(_2869_) );
OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .B(_2842_), .C(IDATA_PROG_write_bF_buf3), .Y(_2870_) );
NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .B(_2869_), .Y(_2871_) );
NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(data_159__0_), .B(_2871__bF_buf4), .Y(_2872_) );
AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_2871__bF_buf3), .C(_2872_), .Y(_66__0_) );
NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(data_159__1_), .B(_2871__bF_buf2), .Y(_2873_) );
AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_2871__bF_buf1), .C(_2873_), .Y(_66__1_) );
NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(data_159__2_), .B(_2871__bF_buf0), .Y(_2874_) );
AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_2871__bF_buf4), .C(_2874_), .Y(_66__2_) );
NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(data_159__3_), .B(_2871__bF_buf3), .Y(_2875_) );
AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_2871__bF_buf2), .C(_2875_), .Y(_66__3_) );
NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(data_159__4_), .B(_2871__bF_buf1), .Y(_2876_) );
AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_2871__bF_buf0), .C(_2876_), .Y(_66__4_) );
NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(data_159__5_), .B(_2871__bF_buf4), .Y(_2877_) );
AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_2871__bF_buf3), .C(_2877_), .Y(_66__5_) );
NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(data_159__6_), .B(_2871__bF_buf2), .Y(_2878_) );
AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_2871__bF_buf1), .C(_2878_), .Y(_66__6_) );
NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(data_159__7_), .B(_2871__bF_buf0), .Y(_2879_) );
AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_2871__bF_buf4), .C(_2879_), .Y(_66__7_) );
NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(data_159__8_), .B(_2871__bF_buf3), .Y(_2880_) );
AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_2871__bF_buf2), .C(_2880_), .Y(_66__8_) );
NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(data_159__9_), .B(_2871__bF_buf1), .Y(_2881_) );
AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_2871__bF_buf0), .C(_2881_), .Y(_66__9_) );
NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(data_159__10_), .B(_2871__bF_buf4), .Y(_2882_) );
AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_2871__bF_buf3), .C(_2882_), .Y(_66__10_) );
NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(data_159__11_), .B(_2871__bF_buf2), .Y(_2883_) );
AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_2871__bF_buf1), .C(_2883_), .Y(_66__11_) );
NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(data_159__12_), .B(_2871__bF_buf0), .Y(_2884_) );
AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_2871__bF_buf4), .C(_2884_), .Y(_66__12_) );
NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(data_159__13_), .B(_2871__bF_buf3), .Y(_2885_) );
AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_2871__bF_buf2), .C(_2885_), .Y(_66__13_) );
NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(data_159__14_), .B(_2871__bF_buf1), .Y(_2886_) );
AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_2871__bF_buf0), .C(_2886_), .Y(_66__14_) );
NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(data_159__15_), .B(_2871__bF_buf4), .Y(_2887_) );
AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_2871__bF_buf3), .C(_2887_), .Y(_66__15_) );
INVX1 INVX1_1464 ( .gnd(gnd), .vdd(vdd), .A(data_158__0_), .Y(_2888_) );
OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15066__bF_buf0), .C(_2888_), .Y(_2889_) );
NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_14941_), .C(_15793__bF_buf4), .Y(_2890_) );
AND2X2 AND2X2_653 ( .gnd(gnd), .vdd(vdd), .A(_2889_), .B(_2890_), .Y(_65__0_) );
NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_14941_), .B(_15793__bF_buf3), .Y(_2891_) );
INVX1 INVX1_1465 ( .gnd(gnd), .vdd(vdd), .A(data_158__1_), .Y(_2892_) );
OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15066__bF_buf3), .C(_2892_), .Y(_2893_) );
OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf0), .B(_2891_), .C(_2893_), .Y(_2894_) );
INVX1 INVX1_1466 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .Y(_65__1_) );
INVX1 INVX1_1467 ( .gnd(gnd), .vdd(vdd), .A(data_158__2_), .Y(_2895_) );
OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15066__bF_buf2), .C(_2895_), .Y(_2896_) );
NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_14941_), .C(_15793__bF_buf2), .Y(_2897_) );
AND2X2 AND2X2_654 ( .gnd(gnd), .vdd(vdd), .A(_2896_), .B(_2897_), .Y(_65__2_) );
INVX1 INVX1_1468 ( .gnd(gnd), .vdd(vdd), .A(data_158__3_), .Y(_2898_) );
OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15066__bF_buf1), .C(_2898_), .Y(_2899_) );
OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf3), .B(_2891_), .C(_2899_), .Y(_2900_) );
INVX1 INVX1_1469 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .Y(_65__3_) );
NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf0), .B(_15788__bF_buf9), .Y(_2901_) );
NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(data_158__4_), .B(_2901_), .Y(_2902_) );
NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf1), .B(_2891_), .Y(_2903_) );
NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2903_), .B(_2902_), .Y(_65__4_) );
INVX1 INVX1_1470 ( .gnd(gnd), .vdd(vdd), .A(data_158__5_), .Y(_2904_) );
OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15066__bF_buf3), .C(_2904_), .Y(_2905_) );
OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf0), .B(_2891_), .C(_2905_), .Y(_2906_) );
INVX1 INVX1_1471 ( .gnd(gnd), .vdd(vdd), .A(_2906_), .Y(_65__5_) );
INVX1 INVX1_1472 ( .gnd(gnd), .vdd(vdd), .A(data_158__6_), .Y(_2907_) );
OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15066__bF_buf2), .C(_2907_), .Y(_2908_) );
NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_14941_), .C(_15793__bF_buf1), .Y(_2909_) );
AND2X2 AND2X2_655 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_2909_), .Y(_65__6_) );
INVX1 INVX1_1473 ( .gnd(gnd), .vdd(vdd), .A(data_158__7_), .Y(_2910_) );
OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15066__bF_buf1), .C(_2910_), .Y(_2911_) );
OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf4), .B(_2891_), .C(_2911_), .Y(_2912_) );
INVX1 INVX1_1474 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .Y(_65__7_) );
INVX1 INVX1_1475 ( .gnd(gnd), .vdd(vdd), .A(data_158__8_), .Y(_2913_) );
OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15066__bF_buf0), .C(_2913_), .Y(_2914_) );
NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_2901_), .Y(_2915_) );
AND2X2 AND2X2_656 ( .gnd(gnd), .vdd(vdd), .A(_2915_), .B(_2914_), .Y(_65__8_) );
NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(data_158__9_), .B(_2901_), .Y(_2916_) );
AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_2901_), .C(_2916_), .Y(_65__9_) );
INVX1 INVX1_1476 ( .gnd(gnd), .vdd(vdd), .A(data_158__10_), .Y(_2917_) );
OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15066__bF_buf3), .C(_2917_), .Y(_2918_) );
NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_2901_), .Y(_2919_) );
AND2X2 AND2X2_657 ( .gnd(gnd), .vdd(vdd), .A(_2919_), .B(_2918_), .Y(_65__10_) );
NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(data_158__11_), .B(_2901_), .Y(_2920_) );
NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf4), .B(_2891_), .Y(_2921_) );
NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2921_), .B(_2920_), .Y(_65__11_) );
INVX1 INVX1_1477 ( .gnd(gnd), .vdd(vdd), .A(data_158__12_), .Y(_2922_) );
OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15066__bF_buf2), .C(_2922_), .Y(_2923_) );
OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf0), .B(_2891_), .C(_2923_), .Y(_2924_) );
INVX1 INVX1_1478 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .Y(_65__12_) );
INVX1 INVX1_1479 ( .gnd(gnd), .vdd(vdd), .A(data_158__13_), .Y(_2925_) );
OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15066__bF_buf1), .C(_2925_), .Y(_2926_) );
OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf1), .B(_2891_), .C(_2926_), .Y(_2927_) );
INVX1 INVX1_1480 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .Y(_65__13_) );
NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(data_158__14_), .B(_2901_), .Y(_2928_) );
NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf0), .B(_2891_), .Y(_2929_) );
NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2929_), .B(_2928_), .Y(_65__14_) );
INVX1 INVX1_1481 ( .gnd(gnd), .vdd(vdd), .A(data_158__15_), .Y(_2930_) );
OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15066__bF_buf0), .C(_2930_), .Y(_2931_) );
OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf4), .B(_2891_), .C(_2931_), .Y(_2932_) );
INVX1 INVX1_1482 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .Y(_65__15_) );
INVX1 INVX1_1483 ( .gnd(gnd), .vdd(vdd), .A(data_157__0_), .Y(_2933_) );
OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf3), .B(_15835_), .C(_2866_), .Y(_2934_) );
NOR3X1 NOR3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_2679_), .B(_2934_), .C(_2621__bF_buf4), .Y(_2935_) );
OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf3), .B(_2868_), .C(_2935_), .Y(_2936_) );
MUX2X1 MUX2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2933_), .B(_14932__bF_buf5), .S(_2936_), .Y(_64__0_) );
INVX1 INVX1_1484 ( .gnd(gnd), .vdd(vdd), .A(data_157__1_), .Y(_2937_) );
MUX2X1 MUX2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .B(_14894__bF_buf5), .S(_2936_), .Y(_64__1_) );
INVX1 INVX1_1485 ( .gnd(gnd), .vdd(vdd), .A(data_157__2_), .Y(_2938_) );
MUX2X1 MUX2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2938_), .B(_14897__bF_buf1), .S(_2936_), .Y(_64__2_) );
AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2869_), .B(_2935_), .C(data_157__3_), .Y(_2939_) );
NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2678_), .C(_2671_), .Y(_2940_) );
INVX1 INVX1_1486 ( .gnd(gnd), .vdd(vdd), .A(_2934_), .Y(_2941_) );
OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf2), .B(_2868_), .C(_2941_), .Y(_2942_) );
NOR3X1 NOR3X1_108 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf2), .B(_2940_), .C(_2942_), .Y(_2943_) );
NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2943_), .B(_2939_), .Y(_64__3_) );
INVX1 INVX1_1487 ( .gnd(gnd), .vdd(vdd), .A(data_157__4_), .Y(_2944_) );
MUX2X1 MUX2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2944_), .B(_14902__bF_buf12), .S(_2936_), .Y(_64__4_) );
INVX1 INVX1_1488 ( .gnd(gnd), .vdd(vdd), .A(data_157__5_), .Y(_2945_) );
MUX2X1 MUX2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2945_), .B(_14903__bF_buf13), .S(_2936_), .Y(_64__5_) );
INVX1 INVX1_1489 ( .gnd(gnd), .vdd(vdd), .A(data_157__6_), .Y(_2946_) );
MUX2X1 MUX2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2946_), .B(_15049__bF_buf1), .S(_2936_), .Y(_64__6_) );
INVX1 INVX1_1490 ( .gnd(gnd), .vdd(vdd), .A(data_157__7_), .Y(_2947_) );
MUX2X1 MUX2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_2947_), .B(_14908__bF_buf12), .S(_2936_), .Y(_64__7_) );
INVX1 INVX1_1491 ( .gnd(gnd), .vdd(vdd), .A(data_157__8_), .Y(_2948_) );
MUX2X1 MUX2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2948_), .B(_15052__bF_buf12), .S(_2936_), .Y(_64__8_) );
INVX1 INVX1_1492 ( .gnd(gnd), .vdd(vdd), .A(data_157__9_), .Y(_2949_) );
MUX2X1 MUX2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2949_), .B(_14913__bF_buf1), .S(_2936_), .Y(_64__9_) );
INVX1 INVX1_1493 ( .gnd(gnd), .vdd(vdd), .A(data_157__10_), .Y(_2950_) );
MUX2X1 MUX2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_2950_), .B(_15055__bF_buf12), .S(_2936_), .Y(_64__10_) );
INVX1 INVX1_1494 ( .gnd(gnd), .vdd(vdd), .A(data_157__11_), .Y(_2951_) );
MUX2X1 MUX2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2951_), .B(_14918__bF_buf0), .S(_2936_), .Y(_64__11_) );
INVX1 INVX1_1495 ( .gnd(gnd), .vdd(vdd), .A(data_157__12_), .Y(_2952_) );
MUX2X1 MUX2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2952_), .B(_14920__bF_buf13), .S(_2936_), .Y(_64__12_) );
INVX1 INVX1_1496 ( .gnd(gnd), .vdd(vdd), .A(data_157__13_), .Y(_2953_) );
MUX2X1 MUX2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2953_), .B(_14924__bF_buf12), .S(_2936_), .Y(_64__13_) );
INVX1 INVX1_1497 ( .gnd(gnd), .vdd(vdd), .A(data_157__14_), .Y(_2954_) );
MUX2X1 MUX2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2954_), .B(_15060__bF_buf5), .S(_2936_), .Y(_64__14_) );
INVX1 INVX1_1498 ( .gnd(gnd), .vdd(vdd), .A(data_157__15_), .Y(_2955_) );
MUX2X1 MUX2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2955_), .B(_15062__bF_buf12), .S(_2936_), .Y(_64__15_) );
OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf2), .B(_15174_), .C(_2866_), .Y(_2956_) );
INVX1 INVX1_1499 ( .gnd(gnd), .vdd(vdd), .A(_2956_), .Y(_2957_) );
OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_2621__bF_buf1), .B(_2868_), .C(_2957_), .Y(_2958_) );
NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2940_), .B(_2958__bF_buf7), .Y(_2959_) );
NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(data_156__0_), .B(_2959__bF_buf4), .Y(_2960_) );
AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_2959__bF_buf3), .C(_2960_), .Y(_63__0_) );
NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(data_156__1_), .B(_2959__bF_buf2), .Y(_2961_) );
AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_2959__bF_buf1), .C(_2961_), .Y(_63__1_) );
NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(data_156__2_), .B(_2959__bF_buf0), .Y(_2962_) );
AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_2959__bF_buf4), .C(_2962_), .Y(_63__2_) );
NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(data_156__3_), .B(_2959__bF_buf3), .Y(_2963_) );
AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_2959__bF_buf2), .C(_2963_), .Y(_63__3_) );
NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(data_156__4_), .B(_2959__bF_buf1), .Y(_2964_) );
AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_2959__bF_buf0), .C(_2964_), .Y(_63__4_) );
NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(data_156__5_), .B(_2959__bF_buf4), .Y(_2965_) );
AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_2959__bF_buf3), .C(_2965_), .Y(_63__5_) );
NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(data_156__6_), .B(_2959__bF_buf2), .Y(_2966_) );
AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf0), .B(_2959__bF_buf1), .C(_2966_), .Y(_63__6_) );
NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(data_156__7_), .B(_2959__bF_buf0), .Y(_2967_) );
AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_2959__bF_buf4), .C(_2967_), .Y(_63__7_) );
NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(data_156__8_), .B(_2959__bF_buf3), .Y(_2968_) );
AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_2959__bF_buf2), .C(_2968_), .Y(_63__8_) );
NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(data_156__9_), .B(_2959__bF_buf1), .Y(_2969_) );
AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_2959__bF_buf0), .C(_2969_), .Y(_63__9_) );
NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(data_156__10_), .B(_2959__bF_buf4), .Y(_2970_) );
AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_2959__bF_buf3), .C(_2970_), .Y(_63__10_) );
NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(data_156__11_), .B(_2959__bF_buf2), .Y(_2971_) );
AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_2959__bF_buf1), .C(_2971_), .Y(_63__11_) );
NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(data_156__12_), .B(_2959__bF_buf0), .Y(_2972_) );
AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_2959__bF_buf4), .C(_2972_), .Y(_63__12_) );
NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(data_156__13_), .B(_2959__bF_buf3), .Y(_2973_) );
AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_2959__bF_buf2), .C(_2973_), .Y(_63__13_) );
NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(data_156__14_), .B(_2959__bF_buf1), .Y(_2974_) );
AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_2959__bF_buf0), .C(_2974_), .Y(_63__14_) );
NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(data_156__15_), .B(_2959__bF_buf4), .Y(_2975_) );
AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_2959__bF_buf3), .C(_2975_), .Y(_63__15_) );
INVX1 INVX1_1500 ( .gnd(gnd), .vdd(vdd), .A(data_155__0_), .Y(_2976_) );
NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_2113_), .Y(_2977_) );
NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_2977_), .B(_2621__bF_buf0), .Y(_2978_) );
OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_15951_), .B(_15161_), .C(_14941_), .Y(_2979_) );
NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_2979_), .B(_15739_), .Y(_2980_) );
INVX1 INVX1_1501 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .Y(_2981_) );
NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_2981_), .B(_2978_), .Y(_2982_) );
OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf6), .C(_2976_), .Y(_2983_) );
INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(_2958__bF_buf5), .Y(_2984_) );
NOR3X1 NOR3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_2977_), .B(_2980_), .C(_2621__bF_buf7), .Y(_2985_) );
NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_2985_), .C(_2984__bF_buf6), .Y(_2986_) );
AND2X2 AND2X2_658 ( .gnd(gnd), .vdd(vdd), .A(_2983_), .B(_2986_), .Y(_62__0_) );
INVX1 INVX1_1502 ( .gnd(gnd), .vdd(vdd), .A(data_155__1_), .Y(_2987_) );
OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf4), .C(_2987_), .Y(_2988_) );
NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_2985_), .C(_2984__bF_buf5), .Y(_2989_) );
AND2X2 AND2X2_659 ( .gnd(gnd), .vdd(vdd), .A(_2988_), .B(_2989_), .Y(_62__1_) );
INVX1 INVX1_1503 ( .gnd(gnd), .vdd(vdd), .A(data_155__2_), .Y(_2990_) );
OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf3), .C(_2990_), .Y(_2991_) );
NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_2985_), .C(_2984__bF_buf4), .Y(_2992_) );
AND2X2 AND2X2_660 ( .gnd(gnd), .vdd(vdd), .A(_2991_), .B(_2992_), .Y(_62__2_) );
INVX1 INVX1_1504 ( .gnd(gnd), .vdd(vdd), .A(data_155__3_), .Y(_2993_) );
OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf2), .C(_2993_), .Y(_2994_) );
NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_2985_), .C(_2984__bF_buf3), .Y(_2995_) );
AND2X2 AND2X2_661 ( .gnd(gnd), .vdd(vdd), .A(_2994_), .B(_2995_), .Y(_62__3_) );
INVX1 INVX1_1505 ( .gnd(gnd), .vdd(vdd), .A(data_155__4_), .Y(_2996_) );
OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf1), .C(_2996_), .Y(_2997_) );
NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_2985_), .C(_2984__bF_buf2), .Y(_2998_) );
AND2X2 AND2X2_662 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_2998_), .Y(_62__4_) );
INVX1 INVX1_1506 ( .gnd(gnd), .vdd(vdd), .A(data_155__5_), .Y(_2999_) );
OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf0), .C(_2999_), .Y(_3000_) );
NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_2985_), .C(_2984__bF_buf1), .Y(_3001_) );
AND2X2 AND2X2_663 ( .gnd(gnd), .vdd(vdd), .A(_3000_), .B(_3001_), .Y(_62__5_) );
INVX1 INVX1_1507 ( .gnd(gnd), .vdd(vdd), .A(data_155__6_), .Y(_3002_) );
OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf7), .C(_3002_), .Y(_3003_) );
NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_2985_), .C(_2984__bF_buf0), .Y(_3004_) );
AND2X2 AND2X2_664 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(_3004_), .Y(_62__6_) );
INVX1 INVX1_1508 ( .gnd(gnd), .vdd(vdd), .A(data_155__7_), .Y(_3005_) );
OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf6), .C(_3005_), .Y(_3006_) );
NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_2985_), .C(_2984__bF_buf6), .Y(_3007_) );
AND2X2 AND2X2_665 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .B(_3007_), .Y(_62__7_) );
INVX1 INVX1_1509 ( .gnd(gnd), .vdd(vdd), .A(data_155__8_), .Y(_3008_) );
OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf5), .C(_3008_), .Y(_3009_) );
NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_2985_), .C(_2984__bF_buf5), .Y(_3010_) );
AND2X2 AND2X2_666 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_3010_), .Y(_62__8_) );
INVX1 INVX1_1510 ( .gnd(gnd), .vdd(vdd), .A(data_155__9_), .Y(_3011_) );
OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf4), .C(_3011_), .Y(_3012_) );
NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf14), .B(_2985_), .C(_2984__bF_buf4), .Y(_3013_) );
AND2X2 AND2X2_667 ( .gnd(gnd), .vdd(vdd), .A(_3012_), .B(_3013_), .Y(_62__9_) );
INVX1 INVX1_1511 ( .gnd(gnd), .vdd(vdd), .A(data_155__10_), .Y(_3014_) );
OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf3), .C(_3014_), .Y(_3015_) );
NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_2985_), .C(_2984__bF_buf3), .Y(_3016_) );
AND2X2 AND2X2_668 ( .gnd(gnd), .vdd(vdd), .A(_3015_), .B(_3016_), .Y(_62__10_) );
INVX1 INVX1_1512 ( .gnd(gnd), .vdd(vdd), .A(data_155__11_), .Y(_3017_) );
OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf2), .C(_3017_), .Y(_3018_) );
NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_2985_), .C(_2984__bF_buf2), .Y(_3019_) );
AND2X2 AND2X2_669 ( .gnd(gnd), .vdd(vdd), .A(_3018_), .B(_3019_), .Y(_62__11_) );
INVX1 INVX1_1513 ( .gnd(gnd), .vdd(vdd), .A(data_155__12_), .Y(_3020_) );
OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf1), .C(_3020_), .Y(_3021_) );
NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_2985_), .C(_2984__bF_buf1), .Y(_3022_) );
AND2X2 AND2X2_670 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_3022_), .Y(_62__12_) );
INVX1 INVX1_1514 ( .gnd(gnd), .vdd(vdd), .A(data_155__13_), .Y(_3023_) );
OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf0), .C(_3023_), .Y(_3024_) );
NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_2985_), .C(_2984__bF_buf0), .Y(_3025_) );
AND2X2 AND2X2_671 ( .gnd(gnd), .vdd(vdd), .A(_3024_), .B(_3025_), .Y(_62__13_) );
INVX1 INVX1_1515 ( .gnd(gnd), .vdd(vdd), .A(data_155__14_), .Y(_3026_) );
OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf7), .C(_3026_), .Y(_3027_) );
NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_2985_), .C(_2984__bF_buf6), .Y(_3028_) );
AND2X2 AND2X2_672 ( .gnd(gnd), .vdd(vdd), .A(_3027_), .B(_3028_), .Y(_62__14_) );
INVX1 INVX1_1516 ( .gnd(gnd), .vdd(vdd), .A(data_155__15_), .Y(_3029_) );
OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2958__bF_buf6), .C(_3029_), .Y(_3030_) );
NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf10), .B(_2985_), .C(_2984__bF_buf5), .Y(_3031_) );
AND2X2 AND2X2_673 ( .gnd(gnd), .vdd(vdd), .A(_3030_), .B(_3031_), .Y(_62__15_) );
INVX1 INVX1_1517 ( .gnd(gnd), .vdd(vdd), .A(data_154__0_), .Y(_3032_) );
OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_14938_), .B(_14940_), .C(IDATA_PROG_write_bF_buf2), .Y(_3033_) );
INVX4 INVX4_11 ( .gnd(gnd), .vdd(vdd), .A(_3033_), .Y(_3034_) );
OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14952__bF_buf1), .C(_14941_), .Y(_3035_) );
OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_3034_), .C(_3035_), .Y(_3036_) );
NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .B(_2671_), .Y(_3037_) );
NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_3036_), .B(_3037_), .Y(_3038_) );
NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_3038_), .B(_2984__bF_buf4), .Y(_3039_) );
NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_3032_), .B(_3039__bF_buf4), .Y(_3040_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf3), .B(IDATA_PROG_data_0_bF_buf4), .Y(_3041_) );
AND2X2 AND2X2_674 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3040_), .Y(_61__0_) );
INVX1 INVX1_1518 ( .gnd(gnd), .vdd(vdd), .A(data_154__1_), .Y(_3042_) );
NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .B(_3039__bF_buf2), .Y(_3043_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf1), .B(IDATA_PROG_data_1_bF_buf4), .Y(_3044_) );
AND2X2 AND2X2_675 ( .gnd(gnd), .vdd(vdd), .A(_3044_), .B(_3043_), .Y(_61__1_) );
INVX1 INVX1_1519 ( .gnd(gnd), .vdd(vdd), .A(data_154__2_), .Y(_3045_) );
NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3045_), .B(_3039__bF_buf0), .Y(_3046_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf4), .B(IDATA_PROG_data_2_bF_buf0), .Y(_3047_) );
AND2X2 AND2X2_676 ( .gnd(gnd), .vdd(vdd), .A(_3047_), .B(_3046_), .Y(_61__2_) );
INVX1 INVX1_1520 ( .gnd(gnd), .vdd(vdd), .A(data_154__3_), .Y(_3048_) );
NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3039__bF_buf3), .Y(_3049_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf2), .B(IDATA_PROG_data_3_bF_buf1), .Y(_3050_) );
AND2X2 AND2X2_677 ( .gnd(gnd), .vdd(vdd), .A(_3050_), .B(_3049_), .Y(_61__3_) );
INVX1 INVX1_1521 ( .gnd(gnd), .vdd(vdd), .A(data_154__4_), .Y(_3051_) );
NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_3039__bF_buf1), .Y(_3052_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf0), .B(IDATA_PROG_data_4_bF_buf0), .Y(_3053_) );
AND2X2 AND2X2_678 ( .gnd(gnd), .vdd(vdd), .A(_3053_), .B(_3052_), .Y(_61__4_) );
INVX1 INVX1_1522 ( .gnd(gnd), .vdd(vdd), .A(data_154__5_), .Y(_3054_) );
NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_3054_), .B(_3039__bF_buf4), .Y(_3055_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf3), .B(IDATA_PROG_data_5_bF_buf4), .Y(_3056_) );
AND2X2 AND2X2_679 ( .gnd(gnd), .vdd(vdd), .A(_3056_), .B(_3055_), .Y(_61__5_) );
INVX1 INVX1_1523 ( .gnd(gnd), .vdd(vdd), .A(data_154__6_), .Y(_3057_) );
NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .B(_3039__bF_buf2), .Y(_3058_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf1), .B(IDATA_PROG_data_6_bF_buf3), .Y(_3059_) );
AND2X2 AND2X2_680 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .B(_3058_), .Y(_61__6_) );
INVX1 INVX1_1524 ( .gnd(gnd), .vdd(vdd), .A(data_154__7_), .Y(_3060_) );
NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(_3060_), .B(_3039__bF_buf0), .Y(_3061_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf4), .B(IDATA_PROG_data_7_bF_buf3), .Y(_3062_) );
AND2X2 AND2X2_681 ( .gnd(gnd), .vdd(vdd), .A(_3062_), .B(_3061_), .Y(_61__7_) );
INVX1 INVX1_1525 ( .gnd(gnd), .vdd(vdd), .A(data_154__8_), .Y(_3063_) );
NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_3063_), .B(_3039__bF_buf3), .Y(_3064_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf2), .B(IDATA_PROG_data_8_bF_buf0), .Y(_3065_) );
AND2X2 AND2X2_682 ( .gnd(gnd), .vdd(vdd), .A(_3065_), .B(_3064_), .Y(_61__8_) );
INVX1 INVX1_1526 ( .gnd(gnd), .vdd(vdd), .A(data_154__9_), .Y(_3066_) );
NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3066_), .B(_3039__bF_buf1), .Y(_3067_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf0), .B(IDATA_PROG_data_9_bF_buf3), .Y(_3068_) );
AND2X2 AND2X2_683 ( .gnd(gnd), .vdd(vdd), .A(_3068_), .B(_3067_), .Y(_61__9_) );
INVX1 INVX1_1527 ( .gnd(gnd), .vdd(vdd), .A(data_154__10_), .Y(_3069_) );
NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_3069_), .B(_3039__bF_buf4), .Y(_3070_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf3), .B(IDATA_PROG_data_10_bF_buf0), .Y(_3071_) );
AND2X2 AND2X2_684 ( .gnd(gnd), .vdd(vdd), .A(_3071_), .B(_3070_), .Y(_61__10_) );
INVX1 INVX1_1528 ( .gnd(gnd), .vdd(vdd), .A(data_154__11_), .Y(_3072_) );
NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_3072_), .B(_3039__bF_buf2), .Y(_3073_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf1), .B(IDATA_PROG_data_11_bF_buf3), .Y(_3074_) );
AND2X2 AND2X2_685 ( .gnd(gnd), .vdd(vdd), .A(_3074_), .B(_3073_), .Y(_61__11_) );
INVX1 INVX1_1529 ( .gnd(gnd), .vdd(vdd), .A(data_154__12_), .Y(_3075_) );
NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_3075_), .B(_3039__bF_buf0), .Y(_3076_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf4), .B(IDATA_PROG_data_12_bF_buf4), .Y(_3077_) );
AND2X2 AND2X2_686 ( .gnd(gnd), .vdd(vdd), .A(_3077_), .B(_3076_), .Y(_61__12_) );
INVX1 INVX1_1530 ( .gnd(gnd), .vdd(vdd), .A(data_154__13_), .Y(_3078_) );
NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3039__bF_buf3), .Y(_3079_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf2), .B(IDATA_PROG_data_13_bF_buf0), .Y(_3080_) );
AND2X2 AND2X2_687 ( .gnd(gnd), .vdd(vdd), .A(_3080_), .B(_3079_), .Y(_61__13_) );
INVX1 INVX1_1531 ( .gnd(gnd), .vdd(vdd), .A(data_154__14_), .Y(_3081_) );
NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_3081_), .B(_3039__bF_buf1), .Y(_3082_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf0), .B(IDATA_PROG_data_14_bF_buf4), .Y(_3083_) );
AND2X2 AND2X2_688 ( .gnd(gnd), .vdd(vdd), .A(_3083_), .B(_3082_), .Y(_61__14_) );
INVX1 INVX1_1532 ( .gnd(gnd), .vdd(vdd), .A(data_154__15_), .Y(_3084_) );
NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(_3084_), .B(_3039__bF_buf4), .Y(_3085_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_3039__bF_buf3), .B(IDATA_PROG_data_15_bF_buf3), .Y(_3086_) );
AND2X2 AND2X2_689 ( .gnd(gnd), .vdd(vdd), .A(_3086_), .B(_3085_), .Y(_61__15_) );
NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .B(_2621__bF_buf6), .Y(_3087_) );
OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_3034_), .C(_3087_), .Y(_3088_) );
NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2958__bF_buf5), .B(_3088_), .Y(_3089_) );
NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(data_153__0_), .B(_3089__bF_buf3), .Y(_3090_) );
AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_3089__bF_buf2), .C(_3090_), .Y(_60__0_) );
INVX1 INVX1_1533 ( .gnd(gnd), .vdd(vdd), .A(data_153__1_), .Y(_3091_) );
OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf4), .C(_3091_), .Y(_3092_) );
AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_3033_), .C(_3037_), .Y(_3093_) );
NAND3X1 NAND3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_3093_), .C(_2984__bF_buf3), .Y(_3094_) );
AND2X2 AND2X2_690 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3094_), .Y(_60__1_) );
INVX1 INVX1_1534 ( .gnd(gnd), .vdd(vdd), .A(data_153__2_), .Y(_3095_) );
OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf3), .C(_3095_), .Y(_3096_) );
NAND3X1 NAND3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf13), .B(_3093_), .C(_2984__bF_buf2), .Y(_3097_) );
AND2X2 AND2X2_691 ( .gnd(gnd), .vdd(vdd), .A(_3096_), .B(_3097_), .Y(_60__2_) );
INVX1 INVX1_1535 ( .gnd(gnd), .vdd(vdd), .A(data_153__3_), .Y(_3098_) );
OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf2), .C(_3098_), .Y(_3099_) );
NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_3089__bF_buf1), .Y(_3100_) );
AND2X2 AND2X2_692 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3099_), .Y(_60__3_) );
INVX1 INVX1_1536 ( .gnd(gnd), .vdd(vdd), .A(data_153__4_), .Y(_3101_) );
OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf1), .C(_3101_), .Y(_3102_) );
NAND3X1 NAND3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_3093_), .C(_2984__bF_buf1), .Y(_3103_) );
AND2X2 AND2X2_693 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .B(_3103_), .Y(_60__4_) );
NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(data_153__5_), .B(_3089__bF_buf0), .Y(_3104_) );
AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_3089__bF_buf3), .C(_3104_), .Y(_60__5_) );
NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(data_153__6_), .B(_3089__bF_buf2), .Y(_3105_) );
AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_3089__bF_buf1), .C(_3105_), .Y(_60__6_) );
NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(data_153__7_), .B(_3089__bF_buf0), .Y(_3106_) );
AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_3089__bF_buf3), .C(_3106_), .Y(_60__7_) );
NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(data_153__8_), .B(_3089__bF_buf2), .Y(_3107_) );
AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_3089__bF_buf1), .C(_3107_), .Y(_60__8_) );
INVX1 INVX1_1537 ( .gnd(gnd), .vdd(vdd), .A(data_153__9_), .Y(_3108_) );
OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf0), .C(_3108_), .Y(_3109_) );
NAND3X1 NAND3X1_376 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_3093_), .C(_2984__bF_buf0), .Y(_3110_) );
AND2X2 AND2X2_694 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .B(_3110_), .Y(_60__9_) );
NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(data_153__10_), .B(_3089__bF_buf0), .Y(_3111_) );
AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_3089__bF_buf3), .C(_3111_), .Y(_60__10_) );
INVX1 INVX1_1538 ( .gnd(gnd), .vdd(vdd), .A(data_153__11_), .Y(_3112_) );
OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf7), .C(_3112_), .Y(_3113_) );
NAND3X1 NAND3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_3093_), .C(_2984__bF_buf6), .Y(_3114_) );
AND2X2 AND2X2_695 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .B(_3114_), .Y(_60__11_) );
NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(data_153__12_), .B(_3089__bF_buf2), .Y(_3115_) );
AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_3089__bF_buf1), .C(_3115_), .Y(_60__12_) );
NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(data_153__13_), .B(_3089__bF_buf0), .Y(_3116_) );
AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_3089__bF_buf3), .C(_3116_), .Y(_60__13_) );
INVX1 INVX1_1539 ( .gnd(gnd), .vdd(vdd), .A(data_153__14_), .Y(_3117_) );
OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_2958__bF_buf6), .C(_3117_), .Y(_3118_) );
NAND3X1 NAND3X1_378 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_3093_), .C(_2984__bF_buf5), .Y(_3119_) );
AND2X2 AND2X2_696 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_3119_), .Y(_60__14_) );
NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(data_153__15_), .B(_3089__bF_buf2), .Y(_3120_) );
AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_3089__bF_buf1), .C(_3120_), .Y(_60__15_) );
INVX1 INVX1_1540 ( .gnd(gnd), .vdd(vdd), .A(data_152__0_), .Y(_3121_) );
OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_14965__bF_buf2), .B(_14952__bF_buf0), .C(_14941_), .Y(_3122_) );
NAND3X1 NAND3X1_379 ( .gnd(gnd), .vdd(vdd), .A(_15739_), .B(_3122_), .C(_2978_), .Y(_3123_) );
NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_2958__bF_buf5), .B(_3123_), .Y(_3124_) );
MUX2X1 MUX2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_3121_), .S(_3124_), .Y(_59__0_) );
INVX1 INVX1_1541 ( .gnd(gnd), .vdd(vdd), .A(data_152__1_), .Y(_3125_) );
MUX2X1 MUX2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_3125_), .S(_3124_), .Y(_59__1_) );
INVX1 INVX1_1542 ( .gnd(gnd), .vdd(vdd), .A(data_152__2_), .Y(_3126_) );
MUX2X1 MUX2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf12), .B(_3126_), .S(_3124_), .Y(_59__2_) );
INVX1 INVX1_1543 ( .gnd(gnd), .vdd(vdd), .A(data_152__3_), .Y(_3127_) );
OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_3123_), .B(_2958__bF_buf4), .C(_3127_), .Y(_3128_) );
NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_3124_), .Y(_3129_) );
AND2X2 AND2X2_697 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .B(_3128_), .Y(_59__3_) );
INVX1 INVX1_1544 ( .gnd(gnd), .vdd(vdd), .A(data_152__4_), .Y(_3130_) );
MUX2X1 MUX2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_3130_), .S(_3124_), .Y(_59__4_) );
INVX1 INVX1_1545 ( .gnd(gnd), .vdd(vdd), .A(data_152__5_), .Y(_3131_) );
MUX2X1 MUX2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_3131_), .S(_3124_), .Y(_59__5_) );
INVX1 INVX1_1546 ( .gnd(gnd), .vdd(vdd), .A(data_152__6_), .Y(_3132_) );
MUX2X1 MUX2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_3132_), .S(_3124_), .Y(_59__6_) );
INVX1 INVX1_1547 ( .gnd(gnd), .vdd(vdd), .A(data_152__7_), .Y(_3133_) );
MUX2X1 MUX2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_3133_), .S(_3124_), .Y(_59__7_) );
INVX1 INVX1_1548 ( .gnd(gnd), .vdd(vdd), .A(data_152__8_), .Y(_3134_) );
MUX2X1 MUX2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_3134_), .S(_3124_), .Y(_59__8_) );
INVX1 INVX1_1549 ( .gnd(gnd), .vdd(vdd), .A(data_152__9_), .Y(_3135_) );
MUX2X1 MUX2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_3135_), .S(_3124_), .Y(_59__9_) );
INVX1 INVX1_1550 ( .gnd(gnd), .vdd(vdd), .A(data_152__10_), .Y(_3136_) );
MUX2X1 MUX2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_3136_), .S(_3124_), .Y(_59__10_) );
INVX1 INVX1_1551 ( .gnd(gnd), .vdd(vdd), .A(data_152__11_), .Y(_3137_) );
MUX2X1 MUX2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_3137_), .S(_3124_), .Y(_59__11_) );
INVX1 INVX1_1552 ( .gnd(gnd), .vdd(vdd), .A(data_152__12_), .Y(_3138_) );
MUX2X1 MUX2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_3138_), .S(_3124_), .Y(_59__12_) );
INVX1 INVX1_1553 ( .gnd(gnd), .vdd(vdd), .A(data_152__13_), .Y(_3139_) );
MUX2X1 MUX2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_3139_), .S(_3124_), .Y(_59__13_) );
INVX1 INVX1_1554 ( .gnd(gnd), .vdd(vdd), .A(data_152__14_), .Y(_3140_) );
MUX2X1 MUX2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_3140_), .S(_3124_), .Y(_59__14_) );
INVX1 INVX1_1555 ( .gnd(gnd), .vdd(vdd), .A(data_152__15_), .Y(_3141_) );
MUX2X1 MUX2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_3141_), .S(_3124_), .Y(_59__15_) );
INVX1 INVX1_1556 ( .gnd(gnd), .vdd(vdd), .A(data_151__0_), .Y(_3142_) );
OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_3034_), .C(_3087_), .Y(_3143_) );
NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2958__bF_buf3), .B(_3143_), .Y(_3144_) );
MUX2X1 MUX2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_3142_), .S(_3144_), .Y(_58__0_) );
INVX1 INVX1_1557 ( .gnd(gnd), .vdd(vdd), .A(data_151__1_), .Y(_3145_) );
OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_2958__bF_buf2), .C(_3145_), .Y(_3146_) );
AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_3033_), .C(_3037_), .Y(_3147_) );
NAND3X1 NAND3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_3147_), .C(_2984__bF_buf4), .Y(_3148_) );
AND2X2 AND2X2_698 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_3148_), .Y(_58__1_) );
INVX1 INVX1_1558 ( .gnd(gnd), .vdd(vdd), .A(data_151__2_), .Y(_3149_) );
OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_2958__bF_buf1), .C(_3149_), .Y(_3150_) );
NAND3X1 NAND3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_3147_), .C(_2984__bF_buf3), .Y(_3151_) );
AND2X2 AND2X2_699 ( .gnd(gnd), .vdd(vdd), .A(_3150_), .B(_3151_), .Y(_58__2_) );
NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(data_151__3_), .B(_3144_), .Y(_3152_) );
AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_3144_), .C(_3152_), .Y(_58__3_) );
INVX1 INVX1_1559 ( .gnd(gnd), .vdd(vdd), .A(data_151__4_), .Y(_3153_) );
OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_2958__bF_buf0), .C(_3153_), .Y(_3154_) );
NAND3X1 NAND3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_3147_), .C(_2984__bF_buf2), .Y(_3155_) );
AND2X2 AND2X2_700 ( .gnd(gnd), .vdd(vdd), .A(_3154_), .B(_3155_), .Y(_58__4_) );
INVX1 INVX1_1560 ( .gnd(gnd), .vdd(vdd), .A(data_151__5_), .Y(_3156_) );
MUX2X1 MUX2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_3156_), .S(_3144_), .Y(_58__5_) );
INVX1 INVX1_1561 ( .gnd(gnd), .vdd(vdd), .A(data_151__6_), .Y(_3157_) );
MUX2X1 MUX2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_3157_), .S(_3144_), .Y(_58__6_) );
INVX1 INVX1_1562 ( .gnd(gnd), .vdd(vdd), .A(data_151__7_), .Y(_3158_) );
MUX2X1 MUX2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_3158_), .S(_3144_), .Y(_58__7_) );
INVX1 INVX1_1563 ( .gnd(gnd), .vdd(vdd), .A(data_151__8_), .Y(_3159_) );
MUX2X1 MUX2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_3159_), .S(_3144_), .Y(_58__8_) );
INVX1 INVX1_1564 ( .gnd(gnd), .vdd(vdd), .A(data_151__9_), .Y(_3160_) );
OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_2958__bF_buf7), .C(_3160_), .Y(_3161_) );
NAND3X1 NAND3X1_383 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_3147_), .C(_2984__bF_buf1), .Y(_3162_) );
AND2X2 AND2X2_701 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .B(_3162_), .Y(_58__9_) );
INVX1 INVX1_1565 ( .gnd(gnd), .vdd(vdd), .A(data_151__10_), .Y(_3163_) );
MUX2X1 MUX2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_3163_), .S(_3144_), .Y(_58__10_) );
INVX1 INVX1_1566 ( .gnd(gnd), .vdd(vdd), .A(data_151__11_), .Y(_3164_) );
OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_2958__bF_buf6), .C(_3164_), .Y(_3165_) );
NAND3X1 NAND3X1_384 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_3147_), .C(_2984__bF_buf0), .Y(_3166_) );
AND2X2 AND2X2_702 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3166_), .Y(_58__11_) );
INVX1 INVX1_1567 ( .gnd(gnd), .vdd(vdd), .A(data_151__12_), .Y(_3167_) );
MUX2X1 MUX2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_3167_), .S(_3144_), .Y(_58__12_) );
INVX1 INVX1_1568 ( .gnd(gnd), .vdd(vdd), .A(data_151__13_), .Y(_3168_) );
MUX2X1 MUX2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_3168_), .S(_3144_), .Y(_58__13_) );
INVX1 INVX1_1569 ( .gnd(gnd), .vdd(vdd), .A(data_151__14_), .Y(_3169_) );
OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_2958__bF_buf5), .C(_3169_), .Y(_3170_) );
NAND3X1 NAND3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_3147_), .C(_2984__bF_buf6), .Y(_3171_) );
AND2X2 AND2X2_703 ( .gnd(gnd), .vdd(vdd), .A(_3170_), .B(_3171_), .Y(_58__14_) );
INVX1 INVX1_1570 ( .gnd(gnd), .vdd(vdd), .A(data_151__15_), .Y(_3172_) );
MUX2X1 MUX2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_3172_), .S(_3144_), .Y(_58__15_) );
INVX1 INVX1_1571 ( .gnd(gnd), .vdd(vdd), .A(data_150__0_), .Y(_3173_) );
OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_1989_), .B(_16204_), .C(_3033_), .Y(_3174_) );
NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .B(_3087_), .Y(_3175_) );
OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf4), .C(_3173_), .Y(_3176_) );
INVX1 INVX1_1572 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .Y(_3177_) );
NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3037_), .Y(_3178_) );
NAND3X1 NAND3X1_386 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_3178_), .C(_2984__bF_buf5), .Y(_3179_) );
AND2X2 AND2X2_704 ( .gnd(gnd), .vdd(vdd), .A(_3176_), .B(_3179_), .Y(_57__0_) );
INVX1 INVX1_1573 ( .gnd(gnd), .vdd(vdd), .A(data_150__1_), .Y(_3180_) );
NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2958__bF_buf3), .B(_3175_), .Y(_3181_) );
MUX2X1 MUX2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_3180_), .S(_3181_), .Y(_57__1_) );
INVX1 INVX1_1574 ( .gnd(gnd), .vdd(vdd), .A(data_150__2_), .Y(_3182_) );
MUX2X1 MUX2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_3182_), .S(_3181_), .Y(_57__2_) );
NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(data_150__3_), .B(_3181_), .Y(_3183_) );
AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_3181_), .C(_3183_), .Y(_57__3_) );
INVX1 INVX1_1575 ( .gnd(gnd), .vdd(vdd), .A(data_150__4_), .Y(_3184_) );
MUX2X1 MUX2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_3184_), .S(_3181_), .Y(_57__4_) );
INVX1 INVX1_1576 ( .gnd(gnd), .vdd(vdd), .A(data_150__5_), .Y(_3185_) );
OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf2), .C(_3185_), .Y(_3186_) );
NAND3X1 NAND3X1_387 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_3178_), .C(_2984__bF_buf4), .Y(_3187_) );
AND2X2 AND2X2_705 ( .gnd(gnd), .vdd(vdd), .A(_3186_), .B(_3187_), .Y(_57__5_) );
INVX1 INVX1_1577 ( .gnd(gnd), .vdd(vdd), .A(data_150__6_), .Y(_3188_) );
OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf1), .C(_3188_), .Y(_3189_) );
NAND3X1 NAND3X1_388 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_3178_), .C(_2984__bF_buf3), .Y(_3190_) );
AND2X2 AND2X2_706 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_3190_), .Y(_57__6_) );
INVX1 INVX1_1578 ( .gnd(gnd), .vdd(vdd), .A(data_150__7_), .Y(_3191_) );
OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf0), .C(_3191_), .Y(_3192_) );
NAND3X1 NAND3X1_389 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_3178_), .C(_2984__bF_buf2), .Y(_3193_) );
AND2X2 AND2X2_707 ( .gnd(gnd), .vdd(vdd), .A(_3192_), .B(_3193_), .Y(_57__7_) );
INVX1 INVX1_1579 ( .gnd(gnd), .vdd(vdd), .A(data_150__8_), .Y(_3194_) );
OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf7), .C(_3194_), .Y(_3195_) );
NAND3X1 NAND3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_3178_), .C(_2984__bF_buf1), .Y(_3196_) );
AND2X2 AND2X2_708 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3196_), .Y(_57__8_) );
INVX1 INVX1_1580 ( .gnd(gnd), .vdd(vdd), .A(data_150__9_), .Y(_3197_) );
MUX2X1 MUX2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_3197_), .S(_3181_), .Y(_57__9_) );
INVX1 INVX1_1581 ( .gnd(gnd), .vdd(vdd), .A(data_150__10_), .Y(_3198_) );
OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf6), .C(_3198_), .Y(_3199_) );
NAND3X1 NAND3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_3178_), .C(_2984__bF_buf0), .Y(_3200_) );
AND2X2 AND2X2_709 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .B(_3200_), .Y(_57__10_) );
INVX1 INVX1_1582 ( .gnd(gnd), .vdd(vdd), .A(data_150__11_), .Y(_3201_) );
MUX2X1 MUX2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_3201_), .S(_3181_), .Y(_57__11_) );
INVX1 INVX1_1583 ( .gnd(gnd), .vdd(vdd), .A(data_150__12_), .Y(_3202_) );
OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf5), .C(_3202_), .Y(_3203_) );
NAND3X1 NAND3X1_392 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_3178_), .C(_2984__bF_buf6), .Y(_3204_) );
AND2X2 AND2X2_710 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .B(_3204_), .Y(_57__12_) );
INVX1 INVX1_1584 ( .gnd(gnd), .vdd(vdd), .A(data_150__13_), .Y(_3205_) );
OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf4), .C(_3205_), .Y(_3206_) );
NAND3X1 NAND3X1_393 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_3178_), .C(_2984__bF_buf5), .Y(_3207_) );
AND2X2 AND2X2_711 ( .gnd(gnd), .vdd(vdd), .A(_3206_), .B(_3207_), .Y(_57__13_) );
INVX1 INVX1_1585 ( .gnd(gnd), .vdd(vdd), .A(data_150__14_), .Y(_3208_) );
MUX2X1 MUX2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf14), .B(_3208_), .S(_3181_), .Y(_57__14_) );
INVX1 INVX1_1586 ( .gnd(gnd), .vdd(vdd), .A(data_150__15_), .Y(_3209_) );
OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_3175_), .B(_2958__bF_buf3), .C(_3209_), .Y(_3210_) );
NAND3X1 NAND3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_3178_), .C(_2984__bF_buf4), .Y(_3211_) );
AND2X2 AND2X2_712 ( .gnd(gnd), .vdd(vdd), .A(_3210_), .B(_3211_), .Y(_57__15_) );
INVX1 INVX1_1587 ( .gnd(gnd), .vdd(vdd), .A(data_149__0_), .Y(_3212_) );
OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .B(_3034_), .C(_3087_), .Y(_3213_) );
OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf2), .C(_3212_), .Y(_3214_) );
NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_3034_), .B(_2030_), .Y(_3215_) );
NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3037_), .Y(_3216_) );
NAND3X1 NAND3X1_395 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_3216_), .C(_2984__bF_buf3), .Y(_3217_) );
AND2X2 AND2X2_713 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_3217_), .Y(_55__0_) );
INVX1 INVX1_1588 ( .gnd(gnd), .vdd(vdd), .A(data_149__1_), .Y(_3218_) );
NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2958__bF_buf1), .B(_3213_), .Y(_3219_) );
MUX2X1 MUX2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_3218_), .S(_3219_), .Y(_55__1_) );
INVX1 INVX1_1589 ( .gnd(gnd), .vdd(vdd), .A(data_149__2_), .Y(_3220_) );
MUX2X1 MUX2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_3220_), .S(_3219_), .Y(_55__2_) );
NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_3219_), .Y(_3221_) );
OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(data_149__3_), .B(_3219_), .C(_3221_), .Y(_3222_) );
INVX1 INVX1_1590 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .Y(_55__3_) );
INVX1 INVX1_1591 ( .gnd(gnd), .vdd(vdd), .A(data_149__4_), .Y(_3223_) );
MUX2X1 MUX2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_3223_), .S(_3219_), .Y(_55__4_) );
INVX1 INVX1_1592 ( .gnd(gnd), .vdd(vdd), .A(data_149__5_), .Y(_3224_) );
OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf0), .C(_3224_), .Y(_3225_) );
NAND3X1 NAND3X1_396 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_3216_), .C(_2984__bF_buf2), .Y(_3226_) );
AND2X2 AND2X2_714 ( .gnd(gnd), .vdd(vdd), .A(_3225_), .B(_3226_), .Y(_55__5_) );
INVX1 INVX1_1593 ( .gnd(gnd), .vdd(vdd), .A(data_149__6_), .Y(_3227_) );
OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf7), .C(_3227_), .Y(_3228_) );
NAND3X1 NAND3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_3216_), .C(_2984__bF_buf1), .Y(_3229_) );
AND2X2 AND2X2_715 ( .gnd(gnd), .vdd(vdd), .A(_3228_), .B(_3229_), .Y(_55__6_) );
INVX1 INVX1_1594 ( .gnd(gnd), .vdd(vdd), .A(data_149__7_), .Y(_3230_) );
OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf6), .C(_3230_), .Y(_3231_) );
NAND3X1 NAND3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_3216_), .C(_2984__bF_buf0), .Y(_3232_) );
AND2X2 AND2X2_716 ( .gnd(gnd), .vdd(vdd), .A(_3231_), .B(_3232_), .Y(_55__7_) );
INVX1 INVX1_1595 ( .gnd(gnd), .vdd(vdd), .A(data_149__8_), .Y(_3233_) );
OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf5), .C(_3233_), .Y(_3234_) );
NAND3X1 NAND3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_3216_), .C(_2984__bF_buf6), .Y(_3235_) );
AND2X2 AND2X2_717 ( .gnd(gnd), .vdd(vdd), .A(_3234_), .B(_3235_), .Y(_55__8_) );
INVX1 INVX1_1596 ( .gnd(gnd), .vdd(vdd), .A(data_149__9_), .Y(_3236_) );
MUX2X1 MUX2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_3236_), .S(_3219_), .Y(_55__9_) );
INVX1 INVX1_1597 ( .gnd(gnd), .vdd(vdd), .A(data_149__10_), .Y(_3237_) );
OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf4), .C(_3237_), .Y(_3238_) );
NAND3X1 NAND3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_3216_), .C(_2984__bF_buf5), .Y(_3239_) );
AND2X2 AND2X2_718 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_3239_), .Y(_55__10_) );
INVX1 INVX1_1598 ( .gnd(gnd), .vdd(vdd), .A(data_149__11_), .Y(_3240_) );
MUX2X1 MUX2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_3240_), .S(_3219_), .Y(_55__11_) );
INVX1 INVX1_1599 ( .gnd(gnd), .vdd(vdd), .A(data_149__12_), .Y(_3241_) );
OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf3), .C(_3241_), .Y(_3242_) );
NAND3X1 NAND3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_3216_), .C(_2984__bF_buf4), .Y(_3243_) );
AND2X2 AND2X2_719 ( .gnd(gnd), .vdd(vdd), .A(_3242_), .B(_3243_), .Y(_55__12_) );
INVX1 INVX1_1600 ( .gnd(gnd), .vdd(vdd), .A(data_149__13_), .Y(_3244_) );
OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf2), .C(_3244_), .Y(_3245_) );
NAND3X1 NAND3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_3216_), .C(_2984__bF_buf3), .Y(_3246_) );
AND2X2 AND2X2_720 ( .gnd(gnd), .vdd(vdd), .A(_3245_), .B(_3246_), .Y(_55__13_) );
INVX1 INVX1_1601 ( .gnd(gnd), .vdd(vdd), .A(data_149__14_), .Y(_3247_) );
MUX2X1 MUX2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_3247_), .S(_3219_), .Y(_55__14_) );
INVX1 INVX1_1602 ( .gnd(gnd), .vdd(vdd), .A(data_149__15_), .Y(_3248_) );
OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_2958__bF_buf1), .C(_3248_), .Y(_3249_) );
NAND3X1 NAND3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_3216_), .C(_2984__bF_buf2), .Y(_3250_) );
AND2X2 AND2X2_721 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .B(_3250_), .Y(_55__15_) );
INVX1 INVX1_1603 ( .gnd(gnd), .vdd(vdd), .A(data_148__0_), .Y(_3251_) );
OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_14959_), .B(_14965__bF_buf1), .C(_14941_), .Y(_3252_) );
NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(_3252_), .B(_15739_), .Y(_3253_) );
INVX1 INVX1_1604 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .Y(_3254_) );
NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_3254_), .B(_2978_), .Y(_3255_) );
OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf0), .C(_3251_), .Y(_3256_) );
NOR3X1 NOR3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_2977_), .B(_3253_), .C(_2621__bF_buf5), .Y(_3257_) );
NAND3X1 NAND3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_3257_), .C(_2984__bF_buf1), .Y(_3258_) );
AND2X2 AND2X2_722 ( .gnd(gnd), .vdd(vdd), .A(_3256_), .B(_3258_), .Y(_54__0_) );
INVX1 INVX1_1605 ( .gnd(gnd), .vdd(vdd), .A(data_148__1_), .Y(_3259_) );
OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf7), .C(_3259_), .Y(_3260_) );
NAND3X1 NAND3X1_405 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_3257_), .C(_2984__bF_buf0), .Y(_3261_) );
AND2X2 AND2X2_723 ( .gnd(gnd), .vdd(vdd), .A(_3260_), .B(_3261_), .Y(_54__1_) );
INVX1 INVX1_1606 ( .gnd(gnd), .vdd(vdd), .A(data_148__2_), .Y(_3262_) );
OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf6), .C(_3262_), .Y(_3263_) );
NAND3X1 NAND3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_3257_), .C(_2984__bF_buf6), .Y(_3264_) );
AND2X2 AND2X2_724 ( .gnd(gnd), .vdd(vdd), .A(_3263_), .B(_3264_), .Y(_54__2_) );
INVX1 INVX1_1607 ( .gnd(gnd), .vdd(vdd), .A(data_148__3_), .Y(_3265_) );
NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3257_), .B(_2984__bF_buf5), .Y(_3266_) );
MUX2X1 MUX2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3265_), .B(_14899__bF_buf10), .S(_3266_), .Y(_54__3_) );
INVX1 INVX1_1608 ( .gnd(gnd), .vdd(vdd), .A(data_148__4_), .Y(_3267_) );
OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf5), .C(_3267_), .Y(_3268_) );
NAND3X1 NAND3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_3257_), .C(_2984__bF_buf4), .Y(_3269_) );
AND2X2 AND2X2_725 ( .gnd(gnd), .vdd(vdd), .A(_3268_), .B(_3269_), .Y(_54__4_) );
INVX1 INVX1_1609 ( .gnd(gnd), .vdd(vdd), .A(data_148__5_), .Y(_3270_) );
OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf4), .C(_3270_), .Y(_3271_) );
NAND3X1 NAND3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_3257_), .C(_2984__bF_buf3), .Y(_3272_) );
AND2X2 AND2X2_726 ( .gnd(gnd), .vdd(vdd), .A(_3271_), .B(_3272_), .Y(_54__5_) );
INVX1 INVX1_1610 ( .gnd(gnd), .vdd(vdd), .A(data_148__6_), .Y(_3273_) );
OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf3), .C(_3273_), .Y(_3274_) );
NAND3X1 NAND3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_3257_), .C(_2984__bF_buf2), .Y(_3275_) );
AND2X2 AND2X2_727 ( .gnd(gnd), .vdd(vdd), .A(_3274_), .B(_3275_), .Y(_54__6_) );
INVX1 INVX1_1611 ( .gnd(gnd), .vdd(vdd), .A(data_148__7_), .Y(_3276_) );
OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf2), .C(_3276_), .Y(_3277_) );
NAND3X1 NAND3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_3257_), .C(_2984__bF_buf1), .Y(_3278_) );
AND2X2 AND2X2_728 ( .gnd(gnd), .vdd(vdd), .A(_3277_), .B(_3278_), .Y(_54__7_) );
INVX1 INVX1_1612 ( .gnd(gnd), .vdd(vdd), .A(data_148__8_), .Y(_3279_) );
OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf1), .C(_3279_), .Y(_3280_) );
NAND3X1 NAND3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_3257_), .C(_2984__bF_buf0), .Y(_3281_) );
AND2X2 AND2X2_729 ( .gnd(gnd), .vdd(vdd), .A(_3280_), .B(_3281_), .Y(_54__8_) );
INVX1 INVX1_1613 ( .gnd(gnd), .vdd(vdd), .A(data_148__9_), .Y(_3282_) );
OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf0), .C(_3282_), .Y(_3283_) );
NAND3X1 NAND3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_3257_), .C(_2984__bF_buf6), .Y(_3284_) );
AND2X2 AND2X2_730 ( .gnd(gnd), .vdd(vdd), .A(_3283_), .B(_3284_), .Y(_54__9_) );
INVX1 INVX1_1614 ( .gnd(gnd), .vdd(vdd), .A(data_148__10_), .Y(_3285_) );
OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf7), .C(_3285_), .Y(_3286_) );
NAND3X1 NAND3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_3257_), .C(_2984__bF_buf5), .Y(_3287_) );
AND2X2 AND2X2_731 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_3287_), .Y(_54__10_) );
INVX1 INVX1_1615 ( .gnd(gnd), .vdd(vdd), .A(data_148__11_), .Y(_3288_) );
OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf6), .C(_3288_), .Y(_3289_) );
NAND3X1 NAND3X1_414 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_3257_), .C(_2984__bF_buf4), .Y(_3290_) );
AND2X2 AND2X2_732 ( .gnd(gnd), .vdd(vdd), .A(_3289_), .B(_3290_), .Y(_54__11_) );
INVX1 INVX1_1616 ( .gnd(gnd), .vdd(vdd), .A(data_148__12_), .Y(_3291_) );
OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf5), .C(_3291_), .Y(_3292_) );
NAND3X1 NAND3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_3257_), .C(_2984__bF_buf3), .Y(_3293_) );
AND2X2 AND2X2_733 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_3293_), .Y(_54__12_) );
INVX1 INVX1_1617 ( .gnd(gnd), .vdd(vdd), .A(data_148__13_), .Y(_3294_) );
OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf4), .C(_3294_), .Y(_3295_) );
NAND3X1 NAND3X1_416 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_3257_), .C(_2984__bF_buf2), .Y(_3296_) );
AND2X2 AND2X2_734 ( .gnd(gnd), .vdd(vdd), .A(_3295_), .B(_3296_), .Y(_54__13_) );
INVX1 INVX1_1618 ( .gnd(gnd), .vdd(vdd), .A(data_148__14_), .Y(_3297_) );
OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf3), .C(_3297_), .Y(_3298_) );
NAND3X1 NAND3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_3257_), .C(_2984__bF_buf1), .Y(_3299_) );
AND2X2 AND2X2_735 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3299_), .Y(_54__14_) );
INVX1 INVX1_1619 ( .gnd(gnd), .vdd(vdd), .A(data_148__15_), .Y(_3300_) );
OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_2958__bF_buf2), .C(_3300_), .Y(_3301_) );
NAND3X1 NAND3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_3257_), .C(_2984__bF_buf0), .Y(_3302_) );
AND2X2 AND2X2_736 ( .gnd(gnd), .vdd(vdd), .A(_3301_), .B(_3302_), .Y(_54__15_) );
INVX1 INVX1_1620 ( .gnd(gnd), .vdd(vdd), .A(data_147__0_), .Y(_3303_) );
NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(_14885__bF_buf2), .B(_15036_), .Y(_3304_) );
NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_15039_), .B(_15018_), .Y(_3305_) );
OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_15074__bF_buf1), .B(_3305_), .C(_3304_), .Y(_3306_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf0), .B(_15011__bF_buf2), .C(_15035_), .D(_14885__bF_buf1), .Y(_3307_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .Y(_3308_) );
NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_15008_), .B(_15028_), .Y(_3309_) );
OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_14943_), .C(_14942__bF_buf3), .Y(_3310_) );
OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf2), .B(_15011__bF_buf1), .C(_3310_), .Y(_3311_) );
NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .B(_3309_), .Y(_3312_) );
NOR3X1 NOR3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_3312_), .C(_3306__bF_buf6), .Y(_3313_) );
NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_14936__bF_buf2), .Y(_3314_) );
NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_15066__bF_buf1), .Y(_3315_) );
NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3314_), .B(_3315_), .Y(_3316_) );
OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf0), .B(_15171_), .C(_3316_), .Y(_3317_) );
NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_15072_), .B(_3317_), .Y(_3318_) );
OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf1), .B(_15508_), .C(_3318_), .Y(_3319_) );
NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_15020_), .B(_14970_), .Y(_3320_) );
NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_15171_), .B(_3320_), .Y(_3321_) );
NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_14933_), .B(_14970_), .Y(_3322_) );
NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[6]), .B(_14934_), .Y(_3323_) );
NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_3323_), .Y(_3324_) );
NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_14986_), .B(_3324_), .Y(_3325_) );
OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_3322_), .C(_3325_), .Y(_3326_) );
AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_14953_), .C(_3320_), .Y(_3327_) );
NOR3X1 NOR3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(_3327_), .C(_3326_), .Y(_3328_) );
NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_15171_), .B(_3322_), .Y(_3329_) );
NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf2), .B(_14998__bF_buf2), .Y(_3330_) );
OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_3322_), .C(_3330_), .Y(_3331_) );
NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_15064_), .Y(_3332_) );
OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf1), .B(_14994_), .C(_3332_), .Y(_3333_) );
INVX1 INVX1_1621 ( .gnd(gnd), .vdd(vdd), .A(_3333_), .Y(_3334_) );
NOR3X1 NOR3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3331_), .C(_3334_), .Y(_3335_) );
NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_14962_), .B(_14958_), .Y(_3336_) );
NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_15174_), .B(_14964_), .Y(_3337_) );
OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3337_), .C(_3332_), .Y(_3338_) );
NAND3X1 NAND3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .B(_3328_), .C(_3335_), .Y(_3339_) );
OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3337_), .C(_3324_), .Y(_3340_) );
OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3337_), .C(_14998__bF_buf1), .Y(_3341_) );
MUX2X1 MUX2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf1), .B(_14946__bF_buf1), .S(_14974_), .Y(_3342_) );
INVX1 INVX1_1622 ( .gnd(gnd), .vdd(vdd), .A(_3342_), .Y(_3343_) );
NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf0), .B(_14975_), .Y(_3344_) );
NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf3), .B(_14986_), .Y(_3345_) );
NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf0), .B(_16157_), .Y(_3346_) );
NAND3X1 NAND3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_3344_), .C(_3346_), .Y(_3347_) );
NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_15010_), .B(_14968_), .Y(_3348_) );
NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf2), .B(_14978__bF_buf0), .Y(_3349_) );
OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_14953_), .B(_3348_), .C(_3349_), .Y(_3350_) );
NOR3X1 NOR3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3350_), .B(_3343_), .C(_3347_), .Y(_3351_) );
NAND3X1 NAND3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_3340_), .B(_3341_), .C(_3351_), .Y(_3352_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .B(_3339_), .Y(_3353_) );
NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .B(_3323_), .Y(_3354_) );
NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_3354__bF_buf3), .B(_14975_), .Y(_3355_) );
NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_3320_), .Y(_3356_) );
NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_14969_), .B(_14970_), .Y(_3357_) );
NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_3357_), .Y(_3358_) );
NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_3356_), .B(_3358_), .Y(_3359_) );
OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf4), .B(_14994_), .C(_3354__bF_buf2), .Y(_3360_) );
NAND3X1 NAND3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3355_), .B(_3360_), .C(_3359_), .Y(_3361_) );
INVX4 INVX4_12 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .Y(_3362_) );
OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_15565_), .B(_14991_), .C(_3354__bF_buf1), .Y(_3363_) );
OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3357_), .C(_3363_), .Y(_3364_) );
NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_3364_), .B(_3361_), .Y(_3365_) );
NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(_14968_), .B(_14970_), .Y(_3366_) );
NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_15171_), .B(_3366_), .Y(_3367_) );
INVX1 INVX1_1623 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .Y(_3368_) );
NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf1), .B(_3354__bF_buf0), .Y(_3369_) );
NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_14884_), .B(_3323_), .Y(_3370_) );
NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_14986_), .B(_3370_), .Y(_3371_) );
AND2X2 AND2X2_737 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_3371_), .Y(_3372_) );
OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf3), .B(_14994_), .C(_3370_), .Y(_3373_) );
NAND3X1 NAND3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_3368_), .B(_3373_), .C(_3372_), .Y(_3374_) );
OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_15565_), .B(_14991_), .C(_3370_), .Y(_3375_) );
OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3366_), .C(_3375_), .Y(_3376_) );
NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .B(_3374_), .Y(_3377_) );
OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf2), .B(_14994_), .C(_15065__bF_buf2), .Y(_3378_) );
NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf0), .B(_3370_), .Y(_3379_) );
OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf1), .B(_15030_), .C(_3379_), .Y(_3380_) );
AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf1), .B(_14975_), .C(_3380_), .Y(_3381_) );
NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3378_), .B(_3381_), .Y(_3382_) );
OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3337_), .C(_15065__bF_buf0), .Y(_3383_) );
INVX1 INVX1_1624 ( .gnd(gnd), .vdd(vdd), .A(_3383_), .Y(_3384_) );
NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_3382_), .Y(_3385_) );
NAND3X1 NAND3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_3377_), .C(_3385_), .Y(_3386_) );
NOR3X1 NOR3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf4), .B(_3319_), .C(_3386_), .Y(_3387_) );
NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(_3313__bF_buf91), .Y(_3388_) );
OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf13_bF_buf3), .C(_3303_), .Y(_3389_) );
INVX1 INVX1_1625 ( .gnd(gnd), .vdd(vdd), .A(_3304_), .Y(_3390_) );
AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_15040_), .B(_15183__bF_buf4), .C(_3390_), .Y(_3391_) );
INVX1 INVX1_1626 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .Y(_3392_) );
NAND3X1 NAND3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_3392_), .C(_3391__bF_buf6), .Y(_3393_) );
INVX1 INVX1_1627 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .Y(_3394_) );
NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .B(_3352_), .Y(_3395_) );
NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3377_), .B(_3365_), .Y(_3396_) );
AND2X2 AND2X2_738 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3378_), .Y(_3397_) );
NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_3383_), .B(_3397_), .Y(_3398_) );
NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_3398_), .B(_3396_), .Y(_3399_) );
NAND3X1 NAND3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3394_), .B(_3395__bF_buf3), .C(_3399_), .Y(_3400_) );
NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_3393__bF_buf69), .Y(_3401_) );
NAND3X1 NAND3X1_427 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(IDATA_PROG_write_bF_buf1), .C(_3401_), .Y(_3402_) );
AND2X2 AND2X2_739 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .B(_3389_), .Y(_53__0_) );
INVX1 INVX1_1628 ( .gnd(gnd), .vdd(vdd), .A(data_147__1_), .Y(_3403_) );
OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf12), .C(_3403_), .Y(_3404_) );
NAND3X1 NAND3X1_428 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf0), .B(_14894__bF_buf11), .C(_3401_), .Y(_3405_) );
AND2X2 AND2X2_740 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .B(_3404_), .Y(_53__1_) );
INVX1 INVX1_1629 ( .gnd(gnd), .vdd(vdd), .A(data_147__2_), .Y(_3406_) );
OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf11), .C(_3406_), .Y(_3407_) );
NAND3X1 NAND3X1_429 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .B(_14897__bF_buf7), .C(_3401_), .Y(_3408_) );
AND2X2 AND2X2_741 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3407_), .Y(_53__2_) );
INVX1 INVX1_1630 ( .gnd(gnd), .vdd(vdd), .A(data_147__3_), .Y(_3409_) );
OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf10), .C(_3409_), .Y(_3410_) );
NAND3X1 NAND3X1_430 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_14899__bF_buf9), .C(_3401_), .Y(_3411_) );
AND2X2 AND2X2_742 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .B(_3410_), .Y(_53__3_) );
INVX1 INVX1_1631 ( .gnd(gnd), .vdd(vdd), .A(data_147__4_), .Y(_3412_) );
OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf9), .C(_3412_), .Y(_3413_) );
NAND3X1 NAND3X1_431 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_14902__bF_buf3), .C(_3401_), .Y(_3414_) );
AND2X2 AND2X2_743 ( .gnd(gnd), .vdd(vdd), .A(_3414_), .B(_3413_), .Y(_53__4_) );
INVX1 INVX1_1632 ( .gnd(gnd), .vdd(vdd), .A(data_147__5_), .Y(_3415_) );
OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf8), .C(_3415_), .Y(_3416_) );
NAND3X1 NAND3X1_432 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf5), .B(_14903__bF_buf4), .C(_3401_), .Y(_3417_) );
AND2X2 AND2X2_744 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_3416_), .Y(_53__5_) );
INVX1 INVX1_1633 ( .gnd(gnd), .vdd(vdd), .A(data_147__6_), .Y(_3418_) );
OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf7), .C(_3418_), .Y(_3419_) );
NAND3X1 NAND3X1_433 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_15049__bF_buf7), .C(_3401_), .Y(_3420_) );
AND2X2 AND2X2_745 ( .gnd(gnd), .vdd(vdd), .A(_3420_), .B(_3419_), .Y(_53__6_) );
INVX1 INVX1_1634 ( .gnd(gnd), .vdd(vdd), .A(data_147__7_), .Y(_3421_) );
OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf6), .C(_3421_), .Y(_3422_) );
NAND3X1 NAND3X1_434 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf3), .B(_14908__bF_buf3), .C(_3401_), .Y(_3423_) );
AND2X2 AND2X2_746 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(_3422_), .Y(_53__7_) );
INVX1 INVX1_1635 ( .gnd(gnd), .vdd(vdd), .A(data_147__8_), .Y(_3424_) );
OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf5), .C(_3424_), .Y(_3425_) );
NAND3X1 NAND3X1_435 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_15052__bF_buf3), .C(_3401_), .Y(_3426_) );
AND2X2 AND2X2_747 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_3425_), .Y(_53__8_) );
INVX1 INVX1_1636 ( .gnd(gnd), .vdd(vdd), .A(data_147__9_), .Y(_3427_) );
OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf4), .C(_3427_), .Y(_3428_) );
NAND3X1 NAND3X1_436 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_14913__bF_buf7), .C(_3401_), .Y(_3429_) );
AND2X2 AND2X2_748 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(_3428_), .Y(_53__9_) );
INVX1 INVX1_1637 ( .gnd(gnd), .vdd(vdd), .A(data_147__10_), .Y(_3430_) );
OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf3), .C(_3430_), .Y(_3431_) );
NAND3X1 NAND3X1_437 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf0), .B(_15055__bF_buf3), .C(_3401_), .Y(_3432_) );
AND2X2 AND2X2_749 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .B(_3431_), .Y(_53__10_) );
INVX1 INVX1_1638 ( .gnd(gnd), .vdd(vdd), .A(data_147__11_), .Y(_3433_) );
OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf2), .C(_3433_), .Y(_3434_) );
NAND3X1 NAND3X1_438 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .B(_14918__bF_buf5), .C(_3401_), .Y(_3435_) );
AND2X2 AND2X2_750 ( .gnd(gnd), .vdd(vdd), .A(_3435_), .B(_3434_), .Y(_53__11_) );
INVX1 INVX1_1639 ( .gnd(gnd), .vdd(vdd), .A(data_147__12_), .Y(_3436_) );
OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf1), .C(_3436_), .Y(_3437_) );
NAND3X1 NAND3X1_439 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_14920__bF_buf4), .C(_3401_), .Y(_3438_) );
AND2X2 AND2X2_751 ( .gnd(gnd), .vdd(vdd), .A(_3438_), .B(_3437_), .Y(_53__12_) );
INVX1 INVX1_1640 ( .gnd(gnd), .vdd(vdd), .A(data_147__13_), .Y(_3439_) );
OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf0), .C(_3439_), .Y(_3440_) );
NAND3X1 NAND3X1_440 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_14924__bF_buf3), .C(_3401_), .Y(_3441_) );
AND2X2 AND2X2_752 ( .gnd(gnd), .vdd(vdd), .A(_3441_), .B(_3440_), .Y(_53__13_) );
INVX1 INVX1_1641 ( .gnd(gnd), .vdd(vdd), .A(data_147__14_), .Y(_3442_) );
OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf15_bF_buf2), .C(_3442_), .Y(_3443_) );
NAND3X1 NAND3X1_441 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf5), .B(_15060__bF_buf11), .C(_3401_), .Y(_3444_) );
AND2X2 AND2X2_753 ( .gnd(gnd), .vdd(vdd), .A(_3444_), .B(_3443_), .Y(_53__14_) );
INVX1 INVX1_1642 ( .gnd(gnd), .vdd(vdd), .A(data_147__15_), .Y(_3445_) );
OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_14882__bF_buf14_bF_buf2), .C(_3445_), .Y(_3446_) );
NAND3X1 NAND3X1_442 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_15062__bF_buf3), .C(_3401_), .Y(_3447_) );
AND2X2 AND2X2_754 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .B(_3446_), .Y(_53__15_) );
INVX1 INVX1_1643 ( .gnd(gnd), .vdd(vdd), .A(data_146__0_), .Y(_3448_) );
OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf0), .B(_15508_), .C(_14966_), .Y(_3449_) );
NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf1), .B(_14954_), .Y(_3450_) );
OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_14980_), .C(_3450_), .Y(_3451_) );
INVX1 INVX1_1644 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3452_) );
AND2X2 AND2X2_755 ( .gnd(gnd), .vdd(vdd), .A(_3316_), .B(IDATA_PROG_write_bF_buf3), .Y(_3453_) );
OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf3), .B(_3452_), .C(_3453_), .Y(_3454_) );
NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3454_), .Y(_3455_) );
NAND3X1 NAND3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3455_), .B(_3395__bF_buf2), .C(_3399_), .Y(_3456_) );
OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_3456_), .C(_3448_), .Y(_3457_) );
INVX1 INVX1_1645 ( .gnd(gnd), .vdd(vdd), .A(_3455_), .Y(_3458_) );
NOR3X1 NOR3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .B(_3353__bF_buf3), .C(_3458_), .Y(_3459_) );
NAND3X1 NAND3X1_444 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_3459_), .C(_3313__bF_buf90), .Y(_3460_) );
AND2X2 AND2X2_756 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_3460_), .Y(_52__0_) );
INVX1 INVX1_1646 ( .gnd(gnd), .vdd(vdd), .A(data_146__1_), .Y(_3461_) );
OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_3456_), .C(_3461_), .Y(_3462_) );
NAND3X1 NAND3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_3459_), .C(_3313__bF_buf89), .Y(_3463_) );
AND2X2 AND2X2_757 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3463_), .Y(_52__1_) );
INVX1 INVX1_1647 ( .gnd(gnd), .vdd(vdd), .A(data_146__2_), .Y(_3464_) );
NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .B(_3313__bF_buf88), .Y(_3465_) );
MUX2X1 MUX2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3464_), .B(_14897__bF_buf6), .S(_3465_), .Y(_52__2_) );
INVX1 INVX1_1648 ( .gnd(gnd), .vdd(vdd), .A(data_146__3_), .Y(_3466_) );
OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_3456_), .C(_3466_), .Y(_3467_) );
NAND3X1 NAND3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_3459_), .C(_3313__bF_buf87), .Y(_3468_) );
AND2X2 AND2X2_758 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3468_), .Y(_52__3_) );
INVX1 INVX1_1649 ( .gnd(gnd), .vdd(vdd), .A(data_146__4_), .Y(_3469_) );
OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_3456_), .C(_3469_), .Y(_3470_) );
NAND3X1 NAND3X1_447 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_3459_), .C(_3313__bF_buf86), .Y(_3471_) );
AND2X2 AND2X2_759 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3471_), .Y(_52__4_) );
INVX1 INVX1_1650 ( .gnd(gnd), .vdd(vdd), .A(data_146__5_), .Y(_3472_) );
OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_3456_), .C(_3472_), .Y(_3473_) );
NAND3X1 NAND3X1_448 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_3459_), .C(_3313__bF_buf85), .Y(_3474_) );
AND2X2 AND2X2_760 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_3474_), .Y(_52__5_) );
INVX1 INVX1_1651 ( .gnd(gnd), .vdd(vdd), .A(data_146__6_), .Y(_3475_) );
MUX2X1 MUX2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_3475_), .B(_15049__bF_buf6), .S(_3465_), .Y(_52__6_) );
INVX1 INVX1_1652 ( .gnd(gnd), .vdd(vdd), .A(data_146__7_), .Y(_3476_) );
OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_3456_), .C(_3476_), .Y(_3477_) );
NAND3X1 NAND3X1_449 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_3459_), .C(_3313__bF_buf84), .Y(_3478_) );
AND2X2 AND2X2_761 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .B(_3478_), .Y(_52__7_) );
INVX1 INVX1_1653 ( .gnd(gnd), .vdd(vdd), .A(data_146__8_), .Y(_3479_) );
MUX2X1 MUX2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_3479_), .B(_15052__bF_buf2), .S(_3465_), .Y(_52__8_) );
INVX1 INVX1_1654 ( .gnd(gnd), .vdd(vdd), .A(data_146__9_), .Y(_3480_) );
MUX2X1 MUX2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_3480_), .B(_14913__bF_buf6), .S(_3465_), .Y(_52__9_) );
INVX1 INVX1_1655 ( .gnd(gnd), .vdd(vdd), .A(data_146__10_), .Y(_3481_) );
MUX2X1 MUX2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3481_), .B(_15055__bF_buf2), .S(_3465_), .Y(_52__10_) );
INVX1 INVX1_1656 ( .gnd(gnd), .vdd(vdd), .A(data_146__11_), .Y(_3482_) );
OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_3456_), .C(_3482_), .Y(_3483_) );
NAND3X1 NAND3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_3459_), .C(_3313__bF_buf83), .Y(_3484_) );
AND2X2 AND2X2_762 ( .gnd(gnd), .vdd(vdd), .A(_3483_), .B(_3484_), .Y(_52__11_) );
INVX1 INVX1_1657 ( .gnd(gnd), .vdd(vdd), .A(data_146__12_), .Y(_3485_) );
OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_3456_), .C(_3485_), .Y(_3486_) );
NAND3X1 NAND3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_3459_), .C(_3313__bF_buf82), .Y(_3487_) );
AND2X2 AND2X2_763 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .B(_3487_), .Y(_52__12_) );
INVX1 INVX1_1658 ( .gnd(gnd), .vdd(vdd), .A(data_146__13_), .Y(_3488_) );
MUX2X1 MUX2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3488_), .B(_14924__bF_buf2), .S(_3465_), .Y(_52__13_) );
INVX1 INVX1_1659 ( .gnd(gnd), .vdd(vdd), .A(data_146__14_), .Y(_3489_) );
MUX2X1 MUX2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(_15060__bF_buf10), .S(_3465_), .Y(_52__14_) );
INVX1 INVX1_1660 ( .gnd(gnd), .vdd(vdd), .A(data_146__15_), .Y(_3490_) );
MUX2X1 MUX2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .B(_15062__bF_buf2), .S(_3465_), .Y(_52__15_) );
INVX1 INVX1_1661 ( .gnd(gnd), .vdd(vdd), .A(data_145__0_), .Y(_3491_) );
OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_14950_), .B(_14954_), .C(_14942__bF_buf0), .Y(_3492_) );
OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_15066__bF_buf2), .B(_3492_), .C(_3453_), .Y(_3493_) );
NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3493_), .Y(_3494_) );
NAND3X1 NAND3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3494_), .B(_3395__bF_buf1), .C(_3399_), .Y(_3495_) );
OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_3495_), .C(_3491_), .Y(_3496_) );
INVX1 INVX1_1662 ( .gnd(gnd), .vdd(vdd), .A(_3494_), .Y(_3497_) );
NOR3X1 NOR3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .B(_3353__bF_buf2), .C(_3497_), .Y(_3498_) );
NAND3X1 NAND3X1_453 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_3498_), .C(_3313__bF_buf81), .Y(_3499_) );
AND2X2 AND2X2_764 ( .gnd(gnd), .vdd(vdd), .A(_3496_), .B(_3499_), .Y(_51__0_) );
INVX1 INVX1_1663 ( .gnd(gnd), .vdd(vdd), .A(data_145__1_), .Y(_3500_) );
OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_3495_), .C(_3500_), .Y(_3501_) );
NAND3X1 NAND3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_3498_), .C(_3313__bF_buf80), .Y(_3502_) );
AND2X2 AND2X2_765 ( .gnd(gnd), .vdd(vdd), .A(_3501_), .B(_3502_), .Y(_51__1_) );
INVX1 INVX1_1664 ( .gnd(gnd), .vdd(vdd), .A(data_145__2_), .Y(_3503_) );
NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3313__bF_buf79), .Y(_3504_) );
MUX2X1 MUX2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3503_), .B(_14897__bF_buf5), .S(_3504_), .Y(_51__2_) );
INVX1 INVX1_1665 ( .gnd(gnd), .vdd(vdd), .A(data_145__3_), .Y(_3505_) );
OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_3495_), .C(_3505_), .Y(_3506_) );
NAND3X1 NAND3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_3498_), .C(_3313__bF_buf78), .Y(_3507_) );
AND2X2 AND2X2_766 ( .gnd(gnd), .vdd(vdd), .A(_3506_), .B(_3507_), .Y(_51__3_) );
INVX1 INVX1_1666 ( .gnd(gnd), .vdd(vdd), .A(data_145__4_), .Y(_3508_) );
OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_3495_), .C(_3508_), .Y(_3509_) );
NAND3X1 NAND3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_3498_), .C(_3313__bF_buf77), .Y(_3510_) );
AND2X2 AND2X2_767 ( .gnd(gnd), .vdd(vdd), .A(_3509_), .B(_3510_), .Y(_51__4_) );
INVX1 INVX1_1667 ( .gnd(gnd), .vdd(vdd), .A(data_145__5_), .Y(_3511_) );
OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_3495_), .C(_3511_), .Y(_3512_) );
NAND3X1 NAND3X1_457 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_3498_), .C(_3313__bF_buf76), .Y(_3513_) );
AND2X2 AND2X2_768 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .B(_3513_), .Y(_51__5_) );
INVX1 INVX1_1668 ( .gnd(gnd), .vdd(vdd), .A(data_145__6_), .Y(_3514_) );
MUX2X1 MUX2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_3514_), .B(_15049__bF_buf5), .S(_3504_), .Y(_51__6_) );
INVX1 INVX1_1669 ( .gnd(gnd), .vdd(vdd), .A(data_145__7_), .Y(_3515_) );
OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_3495_), .C(_3515_), .Y(_3516_) );
NAND3X1 NAND3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_3498_), .C(_3313__bF_buf75), .Y(_3517_) );
AND2X2 AND2X2_769 ( .gnd(gnd), .vdd(vdd), .A(_3516_), .B(_3517_), .Y(_51__7_) );
INVX1 INVX1_1670 ( .gnd(gnd), .vdd(vdd), .A(data_145__8_), .Y(_3518_) );
MUX2X1 MUX2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_3518_), .B(_15052__bF_buf1), .S(_3504_), .Y(_51__8_) );
INVX1 INVX1_1671 ( .gnd(gnd), .vdd(vdd), .A(data_145__9_), .Y(_3519_) );
MUX2X1 MUX2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(_14913__bF_buf5), .S(_3504_), .Y(_51__9_) );
INVX1 INVX1_1672 ( .gnd(gnd), .vdd(vdd), .A(data_145__10_), .Y(_3520_) );
MUX2X1 MUX2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_15055__bF_buf1), .S(_3504_), .Y(_51__10_) );
INVX1 INVX1_1673 ( .gnd(gnd), .vdd(vdd), .A(data_145__11_), .Y(_3521_) );
OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_3495_), .C(_3521_), .Y(_3522_) );
NAND3X1 NAND3X1_459 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_3498_), .C(_3313__bF_buf74), .Y(_3523_) );
AND2X2 AND2X2_770 ( .gnd(gnd), .vdd(vdd), .A(_3522_), .B(_3523_), .Y(_51__11_) );
INVX1 INVX1_1674 ( .gnd(gnd), .vdd(vdd), .A(data_145__12_), .Y(_3524_) );
OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_3495_), .C(_3524_), .Y(_3525_) );
NAND3X1 NAND3X1_460 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_3498_), .C(_3313__bF_buf73), .Y(_3526_) );
AND2X2 AND2X2_771 ( .gnd(gnd), .vdd(vdd), .A(_3525_), .B(_3526_), .Y(_51__12_) );
INVX1 INVX1_1675 ( .gnd(gnd), .vdd(vdd), .A(data_145__13_), .Y(_3527_) );
MUX2X1 MUX2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_3527_), .B(_14924__bF_buf1), .S(_3504_), .Y(_51__13_) );
INVX1 INVX1_1676 ( .gnd(gnd), .vdd(vdd), .A(data_145__14_), .Y(_3528_) );
MUX2X1 MUX2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_3528_), .B(_15060__bF_buf9), .S(_3504_), .Y(_51__14_) );
INVX1 INVX1_1677 ( .gnd(gnd), .vdd(vdd), .A(data_145__15_), .Y(_3529_) );
MUX2X1 MUX2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_3529_), .B(_15062__bF_buf1), .S(_3504_), .Y(_51__15_) );
NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_3315_), .Y(_3530_) );
INVX1 INVX1_1678 ( .gnd(gnd), .vdd(vdd), .A(data_144__0_), .Y(_3531_) );
NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_14986_), .B(_14941_), .Y(_3532_) );
OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf13_bF_buf2), .C(_3531_), .Y(_3533_) );
OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_0_bF_buf3), .C(_3533_), .Y(_3534_) );
INVX1 INVX1_1679 ( .gnd(gnd), .vdd(vdd), .A(_3534_), .Y(_50__0_) );
INVX1 INVX1_1680 ( .gnd(gnd), .vdd(vdd), .A(data_144__1_), .Y(_3535_) );
OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf12), .C(_3535_), .Y(_3536_) );
OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_1_bF_buf3), .C(_3536_), .Y(_3537_) );
INVX1 INVX1_1681 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .Y(_50__1_) );
INVX1 INVX1_1682 ( .gnd(gnd), .vdd(vdd), .A(data_144__2_), .Y(_3538_) );
MUX2X1 MUX2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_3538_), .B(_14897__bF_buf4), .S(_3530_), .Y(_50__2_) );
INVX1 INVX1_1683 ( .gnd(gnd), .vdd(vdd), .A(data_144__3_), .Y(_3539_) );
OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf11), .C(_3539_), .Y(_3540_) );
OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_3_bF_buf0), .C(_3540_), .Y(_3541_) );
INVX1 INVX1_1684 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .Y(_50__3_) );
INVX1 INVX1_1685 ( .gnd(gnd), .vdd(vdd), .A(data_144__4_), .Y(_3542_) );
OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf10), .C(_3542_), .Y(_3543_) );
OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_4_bF_buf4), .C(_3543_), .Y(_3544_) );
INVX1 INVX1_1686 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .Y(_50__4_) );
INVX1 INVX1_1687 ( .gnd(gnd), .vdd(vdd), .A(data_144__5_), .Y(_3545_) );
OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf9), .C(_3545_), .Y(_3546_) );
OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_5_bF_buf3), .C(_3546_), .Y(_3547_) );
INVX1 INVX1_1688 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .Y(_50__5_) );
INVX1 INVX1_1689 ( .gnd(gnd), .vdd(vdd), .A(data_144__6_), .Y(_3548_) );
OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf8), .C(_3548_), .Y(_3549_) );
OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_6_bF_buf2), .C(_3549_), .Y(_3550_) );
INVX1 INVX1_1690 ( .gnd(gnd), .vdd(vdd), .A(_3550_), .Y(_50__6_) );
INVX1 INVX1_1691 ( .gnd(gnd), .vdd(vdd), .A(data_144__7_), .Y(_3551_) );
OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf7), .C(_3551_), .Y(_3552_) );
OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_7_bF_buf2), .C(_3552_), .Y(_3553_) );
INVX1 INVX1_1692 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .Y(_50__7_) );
INVX1 INVX1_1693 ( .gnd(gnd), .vdd(vdd), .A(data_144__8_), .Y(_3554_) );
OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf6), .C(_3554_), .Y(_3555_) );
OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_8_bF_buf4), .C(_3555_), .Y(_3556_) );
INVX1 INVX1_1694 ( .gnd(gnd), .vdd(vdd), .A(_3556_), .Y(_50__8_) );
INVX1 INVX1_1695 ( .gnd(gnd), .vdd(vdd), .A(data_144__9_), .Y(_3557_) );
OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf5), .C(_3557_), .Y(_3558_) );
OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_9_bF_buf2), .C(_3558_), .Y(_3559_) );
INVX1 INVX1_1696 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .Y(_50__9_) );
INVX1 INVX1_1697 ( .gnd(gnd), .vdd(vdd), .A(data_144__10_), .Y(_3560_) );
OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf4), .C(_3560_), .Y(_3561_) );
OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_10_bF_buf4), .C(_3561_), .Y(_3562_) );
INVX1 INVX1_1698 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .Y(_50__10_) );
INVX1 INVX1_1699 ( .gnd(gnd), .vdd(vdd), .A(data_144__11_), .Y(_3563_) );
OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf3), .C(_3563_), .Y(_3564_) );
OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_11_bF_buf2), .C(_3564_), .Y(_3565_) );
INVX1 INVX1_1700 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .Y(_50__11_) );
INVX1 INVX1_1701 ( .gnd(gnd), .vdd(vdd), .A(data_144__12_), .Y(_3566_) );
OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf2), .C(_3566_), .Y(_3567_) );
OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_12_bF_buf3), .C(_3567_), .Y(_3568_) );
INVX1 INVX1_1702 ( .gnd(gnd), .vdd(vdd), .A(_3568_), .Y(_50__12_) );
INVX1 INVX1_1703 ( .gnd(gnd), .vdd(vdd), .A(data_144__13_), .Y(_3569_) );
OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf1), .C(_3569_), .Y(_3570_) );
OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_13_bF_buf4), .C(_3570_), .Y(_3571_) );
INVX1 INVX1_1704 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .Y(_50__13_) );
INVX1 INVX1_1705 ( .gnd(gnd), .vdd(vdd), .A(data_144__14_), .Y(_3572_) );
OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf0), .C(_3572_), .Y(_3573_) );
OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_14_bF_buf3), .C(_3573_), .Y(_3574_) );
INVX1 INVX1_1706 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .Y(_50__14_) );
INVX1 INVX1_1707 ( .gnd(gnd), .vdd(vdd), .A(data_144__15_), .Y(_3575_) );
OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_3532_), .B(_14882__bF_buf15_bF_buf1), .C(_3575_), .Y(_3576_) );
OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_3530_), .B(IDATA_PROG_data_15_bF_buf2), .C(_3576_), .Y(_3577_) );
INVX1 INVX1_1708 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .Y(_50__15_) );
NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_3314_), .Y(_3578_) );
INVX1 INVX1_1709 ( .gnd(gnd), .vdd(vdd), .A(data_143__0_), .Y(_3579_) );
NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf3), .B(_15065__bF_buf3), .Y(_3580_) );
OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf14_bF_buf1), .C(_3579_), .Y(_3581_) );
OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_0_bF_buf2), .C(_3581_), .Y(_3582_) );
INVX1 INVX1_1710 ( .gnd(gnd), .vdd(vdd), .A(_3582_), .Y(_49__0_) );
INVX1 INVX1_1711 ( .gnd(gnd), .vdd(vdd), .A(data_143__1_), .Y(_3583_) );
OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf13_bF_buf1), .C(_3583_), .Y(_3584_) );
NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf12), .B(_3580_), .Y(_3585_) );
NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_3585_), .Y(_3586_) );
AND2X2 AND2X2_772 ( .gnd(gnd), .vdd(vdd), .A(_3586_), .B(_3584_), .Y(_49__1_) );
NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(data_143__2_), .B(_3585_), .Y(_3587_) );
AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_3585_), .C(_3587_), .Y(_49__2_) );
INVX1 INVX1_1712 ( .gnd(gnd), .vdd(vdd), .A(data_143__3_), .Y(_3588_) );
OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf11), .C(_3588_), .Y(_3589_) );
OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_3_bF_buf4), .C(_3589_), .Y(_3590_) );
INVX1 INVX1_1713 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .Y(_49__3_) );
INVX1 INVX1_1714 ( .gnd(gnd), .vdd(vdd), .A(data_143__4_), .Y(_3591_) );
OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf10), .C(_3591_), .Y(_3592_) );
NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_3585_), .Y(_3593_) );
AND2X2 AND2X2_773 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(_3592_), .Y(_49__4_) );
INVX1 INVX1_1715 ( .gnd(gnd), .vdd(vdd), .A(data_143__5_), .Y(_3594_) );
OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf9), .C(_3594_), .Y(_3595_) );
OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_5_bF_buf2), .C(_3595_), .Y(_3596_) );
INVX1 INVX1_1716 ( .gnd(gnd), .vdd(vdd), .A(_3596_), .Y(_49__5_) );
INVX1 INVX1_1717 ( .gnd(gnd), .vdd(vdd), .A(data_143__6_), .Y(_3597_) );
OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf8), .C(_3597_), .Y(_3598_) );
OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_6_bF_buf1), .C(_3598_), .Y(_3599_) );
INVX1 INVX1_1718 ( .gnd(gnd), .vdd(vdd), .A(_3599_), .Y(_49__6_) );
INVX1 INVX1_1719 ( .gnd(gnd), .vdd(vdd), .A(data_143__7_), .Y(_3600_) );
OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf7), .C(_3600_), .Y(_3601_) );
OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_7_bF_buf1), .C(_3601_), .Y(_3602_) );
INVX1 INVX1_1720 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .Y(_49__7_) );
INVX1 INVX1_1721 ( .gnd(gnd), .vdd(vdd), .A(data_143__8_), .Y(_3603_) );
OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf6), .C(_3603_), .Y(_3604_) );
NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_3585_), .Y(_3605_) );
AND2X2 AND2X2_774 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3604_), .Y(_49__8_) );
NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(data_143__9_), .B(_3585_), .Y(_3606_) );
AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_3585_), .C(_3606_), .Y(_49__9_) );
INVX1 INVX1_1722 ( .gnd(gnd), .vdd(vdd), .A(data_143__10_), .Y(_3607_) );
OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf5), .C(_3607_), .Y(_3608_) );
OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_10_bF_buf3), .C(_3608_), .Y(_3609_) );
INVX1 INVX1_1723 ( .gnd(gnd), .vdd(vdd), .A(_3609_), .Y(_49__10_) );
INVX1 INVX1_1724 ( .gnd(gnd), .vdd(vdd), .A(data_143__11_), .Y(_3610_) );
OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf4), .C(_3610_), .Y(_3611_) );
NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_3585_), .Y(_3612_) );
AND2X2 AND2X2_775 ( .gnd(gnd), .vdd(vdd), .A(_3612_), .B(_3611_), .Y(_49__11_) );
INVX1 INVX1_1725 ( .gnd(gnd), .vdd(vdd), .A(data_143__12_), .Y(_3613_) );
OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf3), .C(_3613_), .Y(_3614_) );
OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_12_bF_buf2), .C(_3614_), .Y(_3615_) );
INVX1 INVX1_1726 ( .gnd(gnd), .vdd(vdd), .A(_3615_), .Y(_49__12_) );
INVX1 INVX1_1727 ( .gnd(gnd), .vdd(vdd), .A(data_143__13_), .Y(_3616_) );
OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf2), .C(_3616_), .Y(_3617_) );
NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_3585_), .Y(_3618_) );
AND2X2 AND2X2_776 ( .gnd(gnd), .vdd(vdd), .A(_3618_), .B(_3617_), .Y(_49__13_) );
INVX1 INVX1_1728 ( .gnd(gnd), .vdd(vdd), .A(data_143__14_), .Y(_3619_) );
OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf1), .C(_3619_), .Y(_3620_) );
OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_14_bF_buf2), .C(_3620_), .Y(_3621_) );
INVX1 INVX1_1729 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .Y(_49__14_) );
INVX1 INVX1_1730 ( .gnd(gnd), .vdd(vdd), .A(data_143__15_), .Y(_3622_) );
OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .B(_14882__bF_buf0), .C(_3622_), .Y(_3623_) );
OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(IDATA_PROG_data_15_bF_buf1), .C(_3623_), .Y(_3624_) );
INVX1 INVX1_1731 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .Y(_49__15_) );
INVX1 INVX1_1732 ( .gnd(gnd), .vdd(vdd), .A(data_142__0_), .Y(_3625_) );
NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_14986_), .B(_3354__bF_buf3), .Y(_3626_) );
OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_3320_), .C(_3626_), .Y(_3627_) );
AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_3354__bF_buf2), .B(_14975_), .C(_3627_), .Y(_3628_) );
OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_14990_), .C(_3354__bF_buf1), .Y(_3629_) );
AND2X2 AND2X2_777 ( .gnd(gnd), .vdd(vdd), .A(_3363_), .B(_3629_), .Y(_3630_) );
NAND3X1 NAND3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3360_), .B(_3630_), .C(_3628_), .Y(_3631_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_3376_), .Y(_3632_) );
NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_3632_), .Y(_3633_) );
NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_14966_), .B(_14960_), .Y(_3634_) );
OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14954_), .C(_14963__bF_buf3), .Y(_3635_) );
NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf0), .B(_3635_), .Y(_3636_) );
INVX1 INVX1_1733 ( .gnd(gnd), .vdd(vdd), .A(_3636_), .Y(_3637_) );
OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_14936__bF_buf3), .C(IDATA_PROG_write_bF_buf0), .Y(_3638_) );
AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf2), .B(_3336_), .C(_3638_), .Y(_3639_) );
NAND3X1 NAND3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_3639_), .C(_3397_), .Y(_3640_) );
NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .B(_3640_), .Y(_3641_) );
NAND3X1 NAND3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf0), .B(_3633_), .C(_3641_), .Y(_3642_) );
OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_3642_), .C(_3625_), .Y(_3643_) );
NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_15072_), .B(_15068_), .Y(_3644_) );
NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3636_), .B(_3382_), .Y(_3645_) );
NAND3X1 NAND3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3639_), .C(_3645_), .Y(_3646_) );
NOR3X1 NOR3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf1), .B(_3396_), .C(_3646_), .Y(_3647_) );
NAND3X1 NAND3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_3647_), .C(_3313__bF_buf72), .Y(_3648_) );
AND2X2 AND2X2_778 ( .gnd(gnd), .vdd(vdd), .A(_3643_), .B(_3648_), .Y(_48__0_) );
INVX1 INVX1_1734 ( .gnd(gnd), .vdd(vdd), .A(data_142__1_), .Y(_3649_) );
OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_3642_), .C(_3649_), .Y(_3650_) );
NAND3X1 NAND3X1_466 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_3647_), .C(_3313__bF_buf71), .Y(_3651_) );
AND2X2 AND2X2_779 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_3651_), .Y(_48__1_) );
INVX1 INVX1_1735 ( .gnd(gnd), .vdd(vdd), .A(data_142__2_), .Y(_3652_) );
NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3313__bF_buf70), .Y(_3653_) );
MUX2X1 MUX2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .B(_14897__bF_buf2), .S(_3653_), .Y(_48__2_) );
INVX1 INVX1_1736 ( .gnd(gnd), .vdd(vdd), .A(data_142__3_), .Y(_3654_) );
OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_3642_), .C(_3654_), .Y(_3655_) );
NAND3X1 NAND3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_3647_), .C(_3313__bF_buf69), .Y(_3656_) );
AND2X2 AND2X2_780 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .B(_3656_), .Y(_48__3_) );
INVX1 INVX1_1737 ( .gnd(gnd), .vdd(vdd), .A(data_142__4_), .Y(_3657_) );
OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_3642_), .C(_3657_), .Y(_3658_) );
NAND3X1 NAND3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_3647_), .C(_3313__bF_buf68), .Y(_3659_) );
AND2X2 AND2X2_781 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3659_), .Y(_48__4_) );
INVX1 INVX1_1738 ( .gnd(gnd), .vdd(vdd), .A(data_142__5_), .Y(_3660_) );
OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_3642_), .C(_3660_), .Y(_3661_) );
NAND3X1 NAND3X1_469 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_3647_), .C(_3313__bF_buf67), .Y(_3662_) );
AND2X2 AND2X2_782 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_3662_), .Y(_48__5_) );
INVX1 INVX1_1739 ( .gnd(gnd), .vdd(vdd), .A(data_142__6_), .Y(_3663_) );
MUX2X1 MUX2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_3663_), .B(_15049__bF_buf4), .S(_3653_), .Y(_48__6_) );
INVX1 INVX1_1740 ( .gnd(gnd), .vdd(vdd), .A(data_142__7_), .Y(_3664_) );
OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_3642_), .C(_3664_), .Y(_3665_) );
NAND3X1 NAND3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_3647_), .C(_3313__bF_buf66), .Y(_3666_) );
AND2X2 AND2X2_783 ( .gnd(gnd), .vdd(vdd), .A(_3665_), .B(_3666_), .Y(_48__7_) );
INVX1 INVX1_1741 ( .gnd(gnd), .vdd(vdd), .A(data_142__8_), .Y(_3667_) );
MUX2X1 MUX2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_3667_), .B(_15052__bF_buf13), .S(_3653_), .Y(_48__8_) );
INVX1 INVX1_1742 ( .gnd(gnd), .vdd(vdd), .A(data_142__9_), .Y(_3668_) );
MUX2X1 MUX2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .B(_14913__bF_buf3), .S(_3653_), .Y(_48__9_) );
INVX1 INVX1_1743 ( .gnd(gnd), .vdd(vdd), .A(data_142__10_), .Y(_3669_) );
MUX2X1 MUX2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_3669_), .B(_15055__bF_buf0), .S(_3653_), .Y(_48__10_) );
INVX1 INVX1_1744 ( .gnd(gnd), .vdd(vdd), .A(data_142__11_), .Y(_3670_) );
OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_3642_), .C(_3670_), .Y(_3671_) );
NAND3X1 NAND3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_3647_), .C(_3313__bF_buf65), .Y(_3672_) );
AND2X2 AND2X2_784 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3672_), .Y(_48__11_) );
INVX1 INVX1_1745 ( .gnd(gnd), .vdd(vdd), .A(data_142__12_), .Y(_3673_) );
OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_3642_), .C(_3673_), .Y(_3674_) );
NAND3X1 NAND3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_3647_), .C(_3313__bF_buf64), .Y(_3675_) );
AND2X2 AND2X2_785 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3675_), .Y(_48__12_) );
INVX1 INVX1_1746 ( .gnd(gnd), .vdd(vdd), .A(data_142__13_), .Y(_3676_) );
MUX2X1 MUX2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_3676_), .B(_14924__bF_buf13), .S(_3653_), .Y(_48__13_) );
INVX1 INVX1_1747 ( .gnd(gnd), .vdd(vdd), .A(data_142__14_), .Y(_3677_) );
MUX2X1 MUX2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_3677_), .B(_15060__bF_buf8), .S(_3653_), .Y(_48__14_) );
INVX1 INVX1_1748 ( .gnd(gnd), .vdd(vdd), .A(data_142__15_), .Y(_3678_) );
MUX2X1 MUX2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_3678_), .B(_15062__bF_buf0), .S(_3653_), .Y(_48__15_) );
INVX1 INVX1_1749 ( .gnd(gnd), .vdd(vdd), .A(data_141__0_), .Y(_3679_) );
AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf1), .B(_2672_), .C(_3382_), .Y(_3680_) );
NAND3X1 NAND3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3639_), .C(_3680_), .Y(_3681_) );
NOR3X1 NOR3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf0), .B(_3396_), .C(_3681_), .Y(_3682_) );
NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3313__bF_buf63), .Y(_3683_) );
MUX2X1 MUX2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_3679_), .B(_14932__bF_buf7), .S(_3683_), .Y(_47__0_) );
INVX1 INVX1_1750 ( .gnd(gnd), .vdd(vdd), .A(data_141__1_), .Y(_3684_) );
MUX2X1 MUX2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_3684_), .B(_14894__bF_buf6), .S(_3683_), .Y(_47__1_) );
INVX1 INVX1_1751 ( .gnd(gnd), .vdd(vdd), .A(data_141__2_), .Y(_3685_) );
MUX2X1 MUX2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_3685_), .B(_14897__bF_buf1), .S(_3683_), .Y(_47__2_) );
INVX1 INVX1_1752 ( .gnd(gnd), .vdd(vdd), .A(data_141__3_), .Y(_3686_) );
MUX2X1 MUX2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_3686_), .B(_14899__bF_buf5), .S(_3683_), .Y(_47__3_) );
INVX1 INVX1_1753 ( .gnd(gnd), .vdd(vdd), .A(data_141__4_), .Y(_3687_) );
MUX2X1 MUX2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_3687_), .B(_14902__bF_buf12), .S(_3683_), .Y(_47__4_) );
INVX1 INVX1_1754 ( .gnd(gnd), .vdd(vdd), .A(data_141__5_), .Y(_3688_) );
OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_14936__bF_buf2), .C(IDATA_PROG_write_bF_buf8), .Y(_3689_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(_3689_), .Y(_3690_) );
NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3690_), .Y(_3691_) );
AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf0), .B(_14991_), .C(_3691_), .Y(_3692_) );
OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf1), .B(_2313_), .C(_3397_), .Y(_3693_) );
NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_3396_), .Y(_3694_) );
NAND3X1 NAND3X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf3), .B(_3692_), .C(_3694_), .Y(_3695_) );
OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_3695_), .C(_3688_), .Y(_3696_) );
NAND3X1 NAND3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_3682_), .C(_3313__bF_buf62), .Y(_3697_) );
AND2X2 AND2X2_786 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3697_), .Y(_47__5_) );
INVX1 INVX1_1755 ( .gnd(gnd), .vdd(vdd), .A(data_141__6_), .Y(_3698_) );
MUX2X1 MUX2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_3698_), .B(_15049__bF_buf3), .S(_3683_), .Y(_47__6_) );
INVX1 INVX1_1756 ( .gnd(gnd), .vdd(vdd), .A(data_141__7_), .Y(_3699_) );
OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_3695_), .C(_3699_), .Y(_3700_) );
NAND3X1 NAND3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_3682_), .C(_3313__bF_buf61), .Y(_3701_) );
AND2X2 AND2X2_787 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .B(_3701_), .Y(_47__7_) );
INVX1 INVX1_1757 ( .gnd(gnd), .vdd(vdd), .A(data_141__8_), .Y(_3702_) );
MUX2X1 MUX2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_15052__bF_buf12), .S(_3683_), .Y(_47__8_) );
NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_3695_), .B(_3393__bF_buf42), .Y(_3703_) );
AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3313__bF_buf60), .C(data_141__9_), .Y(_3704_) );
AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_3703_), .C(_3704_), .Y(_47__9_) );
AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3313__bF_buf59), .C(data_141__10_), .Y(_3705_) );
AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_3703_), .C(_3705_), .Y(_47__10_) );
INVX1 INVX1_1758 ( .gnd(gnd), .vdd(vdd), .A(data_141__11_), .Y(_3706_) );
MUX2X1 MUX2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_3706_), .B(_14918__bF_buf0), .S(_3683_), .Y(_47__11_) );
INVX1 INVX1_1759 ( .gnd(gnd), .vdd(vdd), .A(data_141__12_), .Y(_3707_) );
OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_3695_), .C(_3707_), .Y(_3708_) );
NAND3X1 NAND3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_3682_), .C(_3313__bF_buf58), .Y(_3709_) );
AND2X2 AND2X2_788 ( .gnd(gnd), .vdd(vdd), .A(_3708_), .B(_3709_), .Y(_47__12_) );
AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_3682_), .B(_3313__bF_buf57), .C(data_141__13_), .Y(_3710_) );
AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_3703_), .C(_3710_), .Y(_47__13_) );
INVX1 INVX1_1760 ( .gnd(gnd), .vdd(vdd), .A(data_141__14_), .Y(_3711_) );
MUX2X1 MUX2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_3711_), .B(_15060__bF_buf7), .S(_3683_), .Y(_47__14_) );
INVX1 INVX1_1761 ( .gnd(gnd), .vdd(vdd), .A(data_141__15_), .Y(_3712_) );
MUX2X1 MUX2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_3712_), .B(_15062__bF_buf13), .S(_3683_), .Y(_47__15_) );
INVX1 INVX1_1762 ( .gnd(gnd), .vdd(vdd), .A(data_140__0_), .Y(_3713_) );
NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_14954_), .B(_14957_), .Y(_3714_) );
OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf0), .B(_14980_), .C(_3714_), .Y(_3715_) );
AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf3), .B(_3715_), .C(_3689_), .Y(_3716_) );
NAND3X1 NAND3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3716_), .C(_3680_), .Y(_3717_) );
NOR3X1 NOR3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf4), .B(_3396_), .C(_3717_), .Y(_3718_) );
NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3313__bF_buf56), .Y(_3719_) );
MUX2X1 MUX2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_3713_), .B(_14932__bF_buf6), .S(_3719_), .Y(_46__0_) );
INVX1 INVX1_1763 ( .gnd(gnd), .vdd(vdd), .A(data_140__1_), .Y(_3720_) );
MUX2X1 MUX2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_3720_), .B(_14894__bF_buf5), .S(_3719_), .Y(_46__1_) );
INVX1 INVX1_1764 ( .gnd(gnd), .vdd(vdd), .A(data_140__2_), .Y(_3721_) );
MUX2X1 MUX2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .B(_14897__bF_buf0), .S(_3719_), .Y(_46__2_) );
INVX1 INVX1_1765 ( .gnd(gnd), .vdd(vdd), .A(data_140__3_), .Y(_3722_) );
MUX2X1 MUX2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_14899__bF_buf4), .S(_3719_), .Y(_46__3_) );
INVX1 INVX1_1766 ( .gnd(gnd), .vdd(vdd), .A(data_140__4_), .Y(_3723_) );
MUX2X1 MUX2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_14902__bF_buf11), .S(_3719_), .Y(_46__4_) );
INVX1 INVX1_1767 ( .gnd(gnd), .vdd(vdd), .A(data_140__5_), .Y(_3724_) );
NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_14966_), .Y(_3725_) );
NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3336_), .Y(_3726_) );
OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_14936__bF_buf0), .C(_14960_), .Y(_3727_) );
NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_3727_), .Y(_3728_) );
NAND3X1 NAND3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf2), .B(_3728_), .C(_3694_), .Y(_3729_) );
OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_3729_), .C(_3724_), .Y(_3730_) );
NAND3X1 NAND3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_3718_), .C(_3313__bF_buf55), .Y(_3731_) );
AND2X2 AND2X2_789 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3731_), .Y(_46__5_) );
INVX1 INVX1_1768 ( .gnd(gnd), .vdd(vdd), .A(data_140__6_), .Y(_3732_) );
MUX2X1 MUX2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .B(_15049__bF_buf2), .S(_3719_), .Y(_46__6_) );
INVX1 INVX1_1769 ( .gnd(gnd), .vdd(vdd), .A(data_140__7_), .Y(_3733_) );
OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_3729_), .C(_3733_), .Y(_3734_) );
NAND3X1 NAND3X1_481 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_3718_), .C(_3313__bF_buf54), .Y(_3735_) );
AND2X2 AND2X2_790 ( .gnd(gnd), .vdd(vdd), .A(_3734_), .B(_3735_), .Y(_46__7_) );
INVX1 INVX1_1770 ( .gnd(gnd), .vdd(vdd), .A(data_140__8_), .Y(_3736_) );
MUX2X1 MUX2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .B(_15052__bF_buf11), .S(_3719_), .Y(_46__8_) );
NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_3729_), .B(_3393__bF_buf38), .Y(_3737_) );
AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3313__bF_buf53), .C(data_140__9_), .Y(_3738_) );
AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_3737_), .C(_3738_), .Y(_46__9_) );
AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3313__bF_buf52), .C(data_140__10_), .Y(_3739_) );
AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_3737_), .C(_3739_), .Y(_46__10_) );
INVX1 INVX1_1771 ( .gnd(gnd), .vdd(vdd), .A(data_140__11_), .Y(_3740_) );
MUX2X1 MUX2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .B(_14918__bF_buf13), .S(_3719_), .Y(_46__11_) );
INVX1 INVX1_1772 ( .gnd(gnd), .vdd(vdd), .A(data_140__12_), .Y(_3741_) );
OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_3729_), .C(_3741_), .Y(_3742_) );
NAND3X1 NAND3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_3718_), .C(_3313__bF_buf51), .Y(_3743_) );
AND2X2 AND2X2_791 ( .gnd(gnd), .vdd(vdd), .A(_3742_), .B(_3743_), .Y(_46__12_) );
AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3313__bF_buf50), .C(data_140__13_), .Y(_3744_) );
AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_3737_), .C(_3744_), .Y(_46__13_) );
INVX1 INVX1_1773 ( .gnd(gnd), .vdd(vdd), .A(data_140__14_), .Y(_3745_) );
MUX2X1 MUX2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .B(_15060__bF_buf6), .S(_3719_), .Y(_46__14_) );
INVX1 INVX1_1774 ( .gnd(gnd), .vdd(vdd), .A(data_140__15_), .Y(_3746_) );
MUX2X1 MUX2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_3746_), .B(_15062__bF_buf12), .S(_3719_), .Y(_46__15_) );
INVX1 INVX1_1775 ( .gnd(gnd), .vdd(vdd), .A(data_139__0_), .Y(_3747_) );
NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf2), .B(_15065__bF_buf2), .Y(_3748_) );
NAND3X1 NAND3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .B(_3690_), .C(_3644_), .Y(_3749_) );
NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_3749_), .B(_3396_), .Y(_3750_) );
NAND3X1 NAND3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf1), .B(_3397_), .C(_3750_), .Y(_3751_) );
OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_3751_), .C(_3747_), .Y(_3752_) );
AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf1), .B(_15065__bF_buf1), .C(_3382_), .Y(_3753_) );
NAND3X1 NAND3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3690_), .C(_3753_), .Y(_3754_) );
NOR3X1 NOR3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf3), .B(_3396_), .C(_3754_), .Y(_3755_) );
NAND3X1 NAND3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_3755_), .C(_3313__bF_buf49), .Y(_3756_) );
AND2X2 AND2X2_792 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_3756_), .Y(_44__0_) );
INVX1 INVX1_1776 ( .gnd(gnd), .vdd(vdd), .A(data_139__1_), .Y(_3757_) );
OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_3751_), .C(_3757_), .Y(_3758_) );
NAND3X1 NAND3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_3755_), .C(_3313__bF_buf48), .Y(_3759_) );
AND2X2 AND2X2_793 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .B(_3759_), .Y(_44__1_) );
NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_3751_), .B(_3393__bF_buf34), .Y(_3760_) );
AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3313__bF_buf47), .C(data_139__2_), .Y(_3761_) );
AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_3760_), .C(_3761_), .Y(_44__2_) );
INVX1 INVX1_1777 ( .gnd(gnd), .vdd(vdd), .A(data_139__3_), .Y(_3762_) );
OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_3751_), .C(_3762_), .Y(_3763_) );
NAND3X1 NAND3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_3755_), .C(_3313__bF_buf46), .Y(_3764_) );
AND2X2 AND2X2_794 ( .gnd(gnd), .vdd(vdd), .A(_3763_), .B(_3764_), .Y(_44__3_) );
INVX1 INVX1_1778 ( .gnd(gnd), .vdd(vdd), .A(data_139__4_), .Y(_3765_) );
OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_3751_), .C(_3765_), .Y(_3766_) );
NAND3X1 NAND3X1_489 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_3755_), .C(_3313__bF_buf45), .Y(_3767_) );
AND2X2 AND2X2_795 ( .gnd(gnd), .vdd(vdd), .A(_3766_), .B(_3767_), .Y(_44__4_) );
INVX1 INVX1_1779 ( .gnd(gnd), .vdd(vdd), .A(data_139__5_), .Y(_3768_) );
NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3313__bF_buf44), .Y(_3769_) );
MUX2X1 MUX2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_3768_), .B(_14903__bF_buf12), .S(_3769_), .Y(_44__5_) );
AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3313__bF_buf43), .C(data_139__6_), .Y(_3770_) );
AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_3760_), .C(_3770_), .Y(_44__6_) );
INVX1 INVX1_1780 ( .gnd(gnd), .vdd(vdd), .A(data_139__7_), .Y(_3771_) );
MUX2X1 MUX2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(_14908__bF_buf11), .S(_3769_), .Y(_44__7_) );
AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3313__bF_buf42), .C(data_139__8_), .Y(_3772_) );
AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_3760_), .C(_3772_), .Y(_44__8_) );
INVX1 INVX1_1781 ( .gnd(gnd), .vdd(vdd), .A(data_139__9_), .Y(_3773_) );
MUX2X1 MUX2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .B(_14913__bF_buf0), .S(_3769_), .Y(_44__9_) );
INVX1 INVX1_1782 ( .gnd(gnd), .vdd(vdd), .A(data_139__10_), .Y(_3774_) );
MUX2X1 MUX2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_3774_), .B(_15055__bF_buf11), .S(_3769_), .Y(_44__10_) );
INVX1 INVX1_1783 ( .gnd(gnd), .vdd(vdd), .A(data_139__11_), .Y(_3775_) );
OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_3751_), .C(_3775_), .Y(_3776_) );
NAND3X1 NAND3X1_490 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_3755_), .C(_3313__bF_buf41), .Y(_3777_) );
AND2X2 AND2X2_796 ( .gnd(gnd), .vdd(vdd), .A(_3776_), .B(_3777_), .Y(_44__11_) );
INVX1 INVX1_1784 ( .gnd(gnd), .vdd(vdd), .A(data_139__12_), .Y(_3778_) );
MUX2X1 MUX2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_3778_), .B(_14920__bF_buf12), .S(_3769_), .Y(_44__12_) );
INVX1 INVX1_1785 ( .gnd(gnd), .vdd(vdd), .A(data_139__13_), .Y(_3779_) );
MUX2X1 MUX2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .B(_14924__bF_buf10), .S(_3769_), .Y(_44__13_) );
AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3313__bF_buf40), .C(data_139__14_), .Y(_3780_) );
AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf5), .B(_3760_), .C(_3780_), .Y(_44__14_) );
AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3313__bF_buf39), .C(data_139__15_), .Y(_3781_) );
AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_3760_), .C(_3781_), .Y(_44__15_) );
INVX1 INVX1_1786 ( .gnd(gnd), .vdd(vdd), .A(data_138__0_), .Y(_3782_) );
OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14989_), .C(_3714_), .Y(_3783_) );
INVX1 INVX1_1787 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .Y(_3784_) );
OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .B(_14936__bF_buf3), .C(_3748_), .Y(_3785_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3785_), .Y(_3786_) );
AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf0), .B(_14996_), .C(_14882__bF_buf15_bF_buf0), .Y(_3787_) );
NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_3787_), .B(_3644_), .Y(_3788_) );
NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .B(_3786_), .Y(_3789_) );
NAND3X1 NAND3X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf0), .B(_3633_), .C(_3789_), .Y(_3790_) );
OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_3790_), .C(_3782_), .Y(_3791_) );
NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_3785_), .B(_3382_), .Y(_3792_) );
NAND3X1 NAND3X1_492 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3787_), .C(_3792_), .Y(_3793_) );
NOR3X1 NOR3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf2), .B(_3396_), .C(_3793_), .Y(_3794_) );
NAND3X1 NAND3X1_493 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_3794_), .C(_3313__bF_buf38), .Y(_3795_) );
AND2X2 AND2X2_797 ( .gnd(gnd), .vdd(vdd), .A(_3791_), .B(_3795_), .Y(_43__0_) );
INVX1 INVX1_1788 ( .gnd(gnd), .vdd(vdd), .A(data_138__1_), .Y(_3796_) );
OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_3790_), .C(_3796_), .Y(_3797_) );
NAND3X1 NAND3X1_494 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_3794_), .C(_3313__bF_buf37), .Y(_3798_) );
AND2X2 AND2X2_798 ( .gnd(gnd), .vdd(vdd), .A(_3797_), .B(_3798_), .Y(_43__1_) );
INVX1 INVX1_1789 ( .gnd(gnd), .vdd(vdd), .A(data_138__2_), .Y(_3799_) );
NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_3794_), .B(_3313__bF_buf36), .Y(_3800_) );
MUX2X1 MUX2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_3799_), .B(_14897__bF_buf13), .S(_3800_), .Y(_43__2_) );
INVX1 INVX1_1790 ( .gnd(gnd), .vdd(vdd), .A(data_138__3_), .Y(_3801_) );
OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_3790_), .C(_3801_), .Y(_3802_) );
NAND3X1 NAND3X1_495 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_3794_), .C(_3313__bF_buf35), .Y(_3803_) );
AND2X2 AND2X2_799 ( .gnd(gnd), .vdd(vdd), .A(_3802_), .B(_3803_), .Y(_43__3_) );
INVX1 INVX1_1791 ( .gnd(gnd), .vdd(vdd), .A(data_138__4_), .Y(_3804_) );
OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_3790_), .C(_3804_), .Y(_3805_) );
NAND3X1 NAND3X1_496 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_3794_), .C(_3313__bF_buf34), .Y(_3806_) );
AND2X2 AND2X2_800 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_3806_), .Y(_43__4_) );
INVX1 INVX1_1792 ( .gnd(gnd), .vdd(vdd), .A(data_138__5_), .Y(_3807_) );
OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_3790_), .C(_3807_), .Y(_3808_) );
NAND3X1 NAND3X1_497 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_3794_), .C(_3313__bF_buf33), .Y(_3809_) );
AND2X2 AND2X2_801 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(_3809_), .Y(_43__5_) );
INVX1 INVX1_1793 ( .gnd(gnd), .vdd(vdd), .A(data_138__6_), .Y(_3810_) );
MUX2X1 MUX2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_3810_), .B(_15049__bF_buf0), .S(_3800_), .Y(_43__6_) );
INVX1 INVX1_1794 ( .gnd(gnd), .vdd(vdd), .A(data_138__7_), .Y(_3811_) );
OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_3790_), .C(_3811_), .Y(_3812_) );
NAND3X1 NAND3X1_498 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_3794_), .C(_3313__bF_buf32), .Y(_3813_) );
AND2X2 AND2X2_802 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .B(_3813_), .Y(_43__7_) );
INVX1 INVX1_1795 ( .gnd(gnd), .vdd(vdd), .A(data_138__8_), .Y(_3814_) );
MUX2X1 MUX2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_3814_), .B(_15052__bF_buf9), .S(_3800_), .Y(_43__8_) );
INVX1 INVX1_1796 ( .gnd(gnd), .vdd(vdd), .A(data_138__9_), .Y(_3815_) );
MUX2X1 MUX2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_3815_), .B(_14913__bF_buf14), .S(_3800_), .Y(_43__9_) );
INVX1 INVX1_1797 ( .gnd(gnd), .vdd(vdd), .A(data_138__10_), .Y(_3816_) );
MUX2X1 MUX2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_3816_), .B(_15055__bF_buf10), .S(_3800_), .Y(_43__10_) );
INVX1 INVX1_1798 ( .gnd(gnd), .vdd(vdd), .A(data_138__11_), .Y(_3817_) );
OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf24), .B(_3790_), .C(_3817_), .Y(_3818_) );
NAND3X1 NAND3X1_499 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_3794_), .C(_3313__bF_buf31), .Y(_3819_) );
AND2X2 AND2X2_803 ( .gnd(gnd), .vdd(vdd), .A(_3818_), .B(_3819_), .Y(_43__11_) );
INVX1 INVX1_1799 ( .gnd(gnd), .vdd(vdd), .A(data_138__12_), .Y(_3820_) );
OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_3790_), .C(_3820_), .Y(_3821_) );
NAND3X1 NAND3X1_500 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_3794_), .C(_3313__bF_buf30), .Y(_3822_) );
AND2X2 AND2X2_804 ( .gnd(gnd), .vdd(vdd), .A(_3821_), .B(_3822_), .Y(_43__12_) );
INVX1 INVX1_1800 ( .gnd(gnd), .vdd(vdd), .A(data_138__13_), .Y(_3823_) );
MUX2X1 MUX2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_3823_), .B(_14924__bF_buf9), .S(_3800_), .Y(_43__13_) );
INVX1 INVX1_1801 ( .gnd(gnd), .vdd(vdd), .A(data_138__14_), .Y(_3824_) );
MUX2X1 MUX2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_15060__bF_buf4), .S(_3800_), .Y(_43__14_) );
INVX1 INVX1_1802 ( .gnd(gnd), .vdd(vdd), .A(data_138__15_), .Y(_3825_) );
MUX2X1 MUX2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_3825_), .B(_15062__bF_buf10), .S(_3800_), .Y(_43__15_) );
INVX1 INVX1_1803 ( .gnd(gnd), .vdd(vdd), .A(data_137__0_), .Y(_3826_) );
OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_14950_), .B(_14954_), .C(_14957_), .Y(_3827_) );
OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf2), .B(_3827_), .C(_3748_), .Y(_3828_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3828_), .Y(_3829_) );
NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .B(_3829_), .Y(_3830_) );
NAND3X1 NAND3X1_501 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf3), .B(_3633_), .C(_3830_), .Y(_3831_) );
OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_3831_), .C(_3826_), .Y(_3832_) );
NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_3828_), .B(_3382_), .Y(_3833_) );
NAND3X1 NAND3X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3787_), .C(_3833_), .Y(_3834_) );
NOR3X1 NOR3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf1), .B(_3396_), .C(_3834_), .Y(_3835_) );
NAND3X1 NAND3X1_503 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_3835_), .C(_3313__bF_buf29), .Y(_3836_) );
AND2X2 AND2X2_805 ( .gnd(gnd), .vdd(vdd), .A(_3832_), .B(_3836_), .Y(_42__0_) );
INVX1 INVX1_1804 ( .gnd(gnd), .vdd(vdd), .A(data_137__1_), .Y(_3837_) );
OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_3831_), .C(_3837_), .Y(_3838_) );
NAND3X1 NAND3X1_504 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_3835_), .C(_3313__bF_buf28), .Y(_3839_) );
AND2X2 AND2X2_806 ( .gnd(gnd), .vdd(vdd), .A(_3838_), .B(_3839_), .Y(_42__1_) );
NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_3831_), .B(_3393__bF_buf20), .Y(_3840_) );
AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3313__bF_buf27), .C(data_137__2_), .Y(_3841_) );
AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf12), .B(_3840_), .C(_3841_), .Y(_42__2_) );
INVX1 INVX1_1805 ( .gnd(gnd), .vdd(vdd), .A(data_137__3_), .Y(_3842_) );
OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_3831_), .C(_3842_), .Y(_3843_) );
NAND3X1 NAND3X1_505 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_3835_), .C(_3313__bF_buf26), .Y(_3844_) );
AND2X2 AND2X2_807 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(_3844_), .Y(_42__3_) );
INVX1 INVX1_1806 ( .gnd(gnd), .vdd(vdd), .A(data_137__4_), .Y(_3845_) );
OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_3831_), .C(_3845_), .Y(_3846_) );
NAND3X1 NAND3X1_506 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_3835_), .C(_3313__bF_buf25), .Y(_3847_) );
AND2X2 AND2X2_808 ( .gnd(gnd), .vdd(vdd), .A(_3846_), .B(_3847_), .Y(_42__4_) );
INVX1 INVX1_1807 ( .gnd(gnd), .vdd(vdd), .A(data_137__5_), .Y(_3848_) );
NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3313__bF_buf24), .Y(_3849_) );
MUX2X1 MUX2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_3848_), .B(_14903__bF_buf10), .S(_3849_), .Y(_42__5_) );
AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3313__bF_buf23), .C(data_137__6_), .Y(_3850_) );
AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_3840_), .C(_3850_), .Y(_42__6_) );
INVX1 INVX1_1808 ( .gnd(gnd), .vdd(vdd), .A(data_137__7_), .Y(_3851_) );
MUX2X1 MUX2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_3851_), .B(_14908__bF_buf9), .S(_3849_), .Y(_42__7_) );
AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3313__bF_buf22), .C(data_137__8_), .Y(_3852_) );
AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_3840_), .C(_3852_), .Y(_42__8_) );
INVX1 INVX1_1809 ( .gnd(gnd), .vdd(vdd), .A(data_137__9_), .Y(_3853_) );
MUX2X1 MUX2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_14913__bF_buf13), .S(_3849_), .Y(_42__9_) );
INVX1 INVX1_1810 ( .gnd(gnd), .vdd(vdd), .A(data_137__10_), .Y(_3854_) );
MUX2X1 MUX2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_3854_), .B(_15055__bF_buf9), .S(_3849_), .Y(_42__10_) );
INVX1 INVX1_1811 ( .gnd(gnd), .vdd(vdd), .A(data_137__11_), .Y(_3855_) );
OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf17), .B(_3831_), .C(_3855_), .Y(_3856_) );
NAND3X1 NAND3X1_507 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_3835_), .C(_3313__bF_buf21), .Y(_3857_) );
AND2X2 AND2X2_809 ( .gnd(gnd), .vdd(vdd), .A(_3856_), .B(_3857_), .Y(_42__11_) );
INVX1 INVX1_1812 ( .gnd(gnd), .vdd(vdd), .A(data_137__12_), .Y(_3858_) );
MUX2X1 MUX2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_3858_), .B(_14920__bF_buf10), .S(_3849_), .Y(_42__12_) );
INVX1 INVX1_1813 ( .gnd(gnd), .vdd(vdd), .A(data_137__13_), .Y(_3859_) );
MUX2X1 MUX2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(_14924__bF_buf8), .S(_3849_), .Y(_42__13_) );
AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3313__bF_buf20), .C(data_137__14_), .Y(_3860_) );
AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_3840_), .C(_3860_), .Y(_42__14_) );
AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3313__bF_buf19), .C(data_137__15_), .Y(_3861_) );
AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_3840_), .C(_3861_), .Y(_42__15_) );
INVX1 INVX1_1814 ( .gnd(gnd), .vdd(vdd), .A(data_136__0_), .Y(_3862_) );
NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_14887_), .B(_14977__bF_buf0), .Y(_3863_) );
NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14989_), .Y(_3864_) );
NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_3863_), .B(_3864_), .Y(_3865_) );
OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf1), .B(_3865_), .C(_14960_), .Y(_3866_) );
NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_3866_), .Y(_3867_) );
NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_3867_), .B(_3833_), .Y(_3868_) );
INVX1 INVX1_1815 ( .gnd(gnd), .vdd(vdd), .A(_3868_), .Y(_3869_) );
NAND3X1 NAND3X1_508 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf2), .B(_3633_), .C(_3869_), .Y(_3870_) );
OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf16), .B(_3870_), .C(_3862_), .Y(_3871_) );
NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_3633_), .B(_3395__bF_buf1), .Y(_3872_) );
NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_3868_), .B(_3872_), .Y(_3873_) );
NAND3X1 NAND3X1_509 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_3313__bF_buf18), .C(_3873_), .Y(_3874_) );
AND2X2 AND2X2_810 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3874_), .Y(_41__0_) );
INVX1 INVX1_1816 ( .gnd(gnd), .vdd(vdd), .A(data_136__1_), .Y(_3875_) );
OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf15), .B(_3870_), .C(_3875_), .Y(_3876_) );
NAND3X1 NAND3X1_510 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_3313__bF_buf17), .C(_3873_), .Y(_3877_) );
AND2X2 AND2X2_811 ( .gnd(gnd), .vdd(vdd), .A(_3876_), .B(_3877_), .Y(_41__1_) );
INVX1 INVX1_1817 ( .gnd(gnd), .vdd(vdd), .A(data_136__2_), .Y(_3878_) );
NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf16), .B(_3873_), .Y(_3879_) );
MUX2X1 MUX2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_3878_), .B(_14897__bF_buf11), .S(_3879_), .Y(_41__2_) );
INVX1 INVX1_1818 ( .gnd(gnd), .vdd(vdd), .A(data_136__3_), .Y(_3880_) );
OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf14), .B(_3870_), .C(_3880_), .Y(_3881_) );
NAND3X1 NAND3X1_511 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_3313__bF_buf15), .C(_3873_), .Y(_3882_) );
AND2X2 AND2X2_812 ( .gnd(gnd), .vdd(vdd), .A(_3881_), .B(_3882_), .Y(_41__3_) );
INVX1 INVX1_1819 ( .gnd(gnd), .vdd(vdd), .A(data_136__4_), .Y(_3883_) );
OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf13), .B(_3870_), .C(_3883_), .Y(_3884_) );
NAND3X1 NAND3X1_512 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_3313__bF_buf14), .C(_3873_), .Y(_3885_) );
AND2X2 AND2X2_813 ( .gnd(gnd), .vdd(vdd), .A(_3884_), .B(_3885_), .Y(_41__4_) );
INVX1 INVX1_1820 ( .gnd(gnd), .vdd(vdd), .A(data_136__5_), .Y(_3886_) );
OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_3870_), .C(_3886_), .Y(_3887_) );
NAND3X1 NAND3X1_513 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_3313__bF_buf13), .C(_3873_), .Y(_3888_) );
AND2X2 AND2X2_814 ( .gnd(gnd), .vdd(vdd), .A(_3887_), .B(_3888_), .Y(_41__5_) );
INVX1 INVX1_1821 ( .gnd(gnd), .vdd(vdd), .A(data_136__6_), .Y(_3889_) );
MUX2X1 MUX2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_15049__bF_buf13), .S(_3879_), .Y(_41__6_) );
INVX1 INVX1_1822 ( .gnd(gnd), .vdd(vdd), .A(data_136__7_), .Y(_3890_) );
OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_3870_), .C(_3890_), .Y(_3891_) );
NAND3X1 NAND3X1_514 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_3313__bF_buf12), .C(_3873_), .Y(_3892_) );
AND2X2 AND2X2_815 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_3892_), .Y(_41__7_) );
INVX1 INVX1_1823 ( .gnd(gnd), .vdd(vdd), .A(data_136__8_), .Y(_3893_) );
MUX2X1 MUX2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3893_), .B(_15052__bF_buf7), .S(_3879_), .Y(_41__8_) );
INVX1 INVX1_1824 ( .gnd(gnd), .vdd(vdd), .A(data_136__9_), .Y(_3894_) );
MUX2X1 MUX2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_3894_), .B(_14913__bF_buf12), .S(_3879_), .Y(_41__9_) );
INVX1 INVX1_1825 ( .gnd(gnd), .vdd(vdd), .A(data_136__10_), .Y(_3895_) );
MUX2X1 MUX2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_3895_), .B(_15055__bF_buf8), .S(_3879_), .Y(_41__10_) );
INVX1 INVX1_1826 ( .gnd(gnd), .vdd(vdd), .A(data_136__11_), .Y(_3896_) );
OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_3870_), .C(_3896_), .Y(_3897_) );
NAND3X1 NAND3X1_515 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_3313__bF_buf11), .C(_3873_), .Y(_3898_) );
AND2X2 AND2X2_816 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_3898_), .Y(_41__11_) );
INVX1 INVX1_1827 ( .gnd(gnd), .vdd(vdd), .A(data_136__12_), .Y(_3899_) );
OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_3870_), .C(_3899_), .Y(_3900_) );
NAND3X1 NAND3X1_516 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_3313__bF_buf10), .C(_3873_), .Y(_3901_) );
AND2X2 AND2X2_817 ( .gnd(gnd), .vdd(vdd), .A(_3900_), .B(_3901_), .Y(_41__12_) );
INVX1 INVX1_1828 ( .gnd(gnd), .vdd(vdd), .A(data_136__13_), .Y(_3902_) );
MUX2X1 MUX2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_3902_), .B(_14924__bF_buf7), .S(_3879_), .Y(_41__13_) );
INVX1 INVX1_1829 ( .gnd(gnd), .vdd(vdd), .A(data_136__14_), .Y(_3903_) );
MUX2X1 MUX2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_3903_), .B(_15060__bF_buf2), .S(_3879_), .Y(_41__14_) );
INVX1 INVX1_1830 ( .gnd(gnd), .vdd(vdd), .A(data_136__15_), .Y(_3904_) );
MUX2X1 MUX2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_3904_), .B(_15062__bF_buf8), .S(_3879_), .Y(_41__15_) );
INVX1 INVX1_1831 ( .gnd(gnd), .vdd(vdd), .A(data_135__0_), .Y(_3905_) );
NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf14_bF_buf0), .B(_3380_), .Y(_3906_) );
OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf0), .B(_15171_), .C(_3906_), .Y(_3907_) );
OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_14936__bF_buf3), .C(_3378_), .Y(_3908_) );
NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_3908_), .B(_3907_), .Y(_3909_) );
NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3909_), .Y(_3910_) );
INVX1 INVX1_1832 ( .gnd(gnd), .vdd(vdd), .A(_3910_), .Y(_3911_) );
NAND3X1 NAND3X1_517 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf0), .B(_3633_), .C(_3911_), .Y(_3912_) );
OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_3393__bF_buf8), .C(_3905_), .Y(_3913_) );
NOR3X1 NOR3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3910_), .B(_3396_), .C(_3353__bF_buf0), .Y(_3914_) );
NAND3X1 NAND3X1_518 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_3914_), .C(_3313__bF_buf9), .Y(_3915_) );
AND2X2 AND2X2_818 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3915_), .Y(_40__0_) );
INVX1 INVX1_1833 ( .gnd(gnd), .vdd(vdd), .A(data_135__1_), .Y(_3916_) );
OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_3393__bF_buf7), .C(_3916_), .Y(_3917_) );
NAND3X1 NAND3X1_519 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_3914_), .C(_3313__bF_buf8), .Y(_3918_) );
AND2X2 AND2X2_819 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .B(_3918_), .Y(_40__1_) );
NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_3912_), .Y(_3919_) );
AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3313__bF_buf7), .C(data_135__2_), .Y(_3920_) );
AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_3919_), .C(_3920_), .Y(_40__2_) );
INVX1 INVX1_1834 ( .gnd(gnd), .vdd(vdd), .A(data_135__3_), .Y(_3921_) );
OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_3393__bF_buf5), .C(_3921_), .Y(_3922_) );
NAND3X1 NAND3X1_520 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_3914_), .C(_3313__bF_buf6), .Y(_3923_) );
AND2X2 AND2X2_820 ( .gnd(gnd), .vdd(vdd), .A(_3922_), .B(_3923_), .Y(_40__3_) );
INVX1 INVX1_1835 ( .gnd(gnd), .vdd(vdd), .A(data_135__4_), .Y(_3924_) );
OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_3393__bF_buf4), .C(_3924_), .Y(_3925_) );
NAND3X1 NAND3X1_521 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_3914_), .C(_3313__bF_buf5), .Y(_3926_) );
AND2X2 AND2X2_821 ( .gnd(gnd), .vdd(vdd), .A(_3925_), .B(_3926_), .Y(_40__4_) );
INVX1 INVX1_1836 ( .gnd(gnd), .vdd(vdd), .A(data_135__5_), .Y(_3927_) );
NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3313__bF_buf4), .Y(_3928_) );
MUX2X1 MUX2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_3927_), .B(_14903__bF_buf8), .S(_3928_), .Y(_40__5_) );
AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3313__bF_buf3), .C(data_135__6_), .Y(_3929_) );
AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_3919_), .C(_3929_), .Y(_40__6_) );
INVX1 INVX1_1837 ( .gnd(gnd), .vdd(vdd), .A(data_135__7_), .Y(_3930_) );
MUX2X1 MUX2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_3930_), .B(_14908__bF_buf7), .S(_3928_), .Y(_40__7_) );
AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3313__bF_buf2), .C(data_135__8_), .Y(_3931_) );
AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_3919_), .C(_3931_), .Y(_40__8_) );
INVX1 INVX1_1838 ( .gnd(gnd), .vdd(vdd), .A(data_135__9_), .Y(_3932_) );
MUX2X1 MUX2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_3932_), .B(_14913__bF_buf11), .S(_3928_), .Y(_40__9_) );
INVX1 INVX1_1839 ( .gnd(gnd), .vdd(vdd), .A(data_135__10_), .Y(_3933_) );
MUX2X1 MUX2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_3933_), .B(_15055__bF_buf7), .S(_3928_), .Y(_40__10_) );
INVX1 INVX1_1840 ( .gnd(gnd), .vdd(vdd), .A(data_135__11_), .Y(_3934_) );
OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_3912_), .B(_3393__bF_buf3), .C(_3934_), .Y(_3935_) );
NAND3X1 NAND3X1_522 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_3914_), .C(_3313__bF_buf1), .Y(_3936_) );
AND2X2 AND2X2_822 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3936_), .Y(_40__11_) );
INVX1 INVX1_1841 ( .gnd(gnd), .vdd(vdd), .A(data_135__12_), .Y(_3937_) );
MUX2X1 MUX2X1_596 ( .gnd(gnd), .vdd(vdd), .A(_3937_), .B(_14920__bF_buf8), .S(_3928_), .Y(_40__12_) );
INVX1 INVX1_1842 ( .gnd(gnd), .vdd(vdd), .A(data_135__13_), .Y(_3938_) );
MUX2X1 MUX2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_3938_), .B(_14924__bF_buf6), .S(_3928_), .Y(_40__13_) );
AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3313__bF_buf0), .C(data_135__14_), .Y(_3939_) );
AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_3919_), .C(_3939_), .Y(_40__14_) );
AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3313__bF_buf91), .C(data_135__15_), .Y(_3940_) );
AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_3919_), .C(_3940_), .Y(_40__15_) );
AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf3), .B(_14978__bF_buf1), .C(_14882__bF_buf13_bF_buf0), .Y(_3941_) );
NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_14948_), .B(_14952__bF_buf4), .Y(_3942_) );
OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_14887_), .B(_14977__bF_buf3), .C(_3942_), .Y(_3943_) );
OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_3943_), .B(IDATA_PROG_addr_3_bF_buf2), .C(_15065__bF_buf2), .Y(_3944_) );
NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_14936__bF_buf2), .Y(_3945_) );
NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_2313_), .Y(_3946_) );
AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[0]), .B(_3946_), .C(_3945_), .Y(_3947_) );
OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf1), .B(_15171_), .C(_3947_), .Y(_3948_) );
NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .B(_3948_), .Y(_3949_) );
NAND3X1 NAND3X1_523 ( .gnd(gnd), .vdd(vdd), .A(_3941_), .B(_3944_), .C(_3949_), .Y(_3950_) );
NOR3X1 NOR3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_3396_), .B(_3950_), .C(_3353__bF_buf4), .Y(_3951_) );
AND2X2 AND2X2_823 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf90), .B(_3951_), .Y(_3952_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_3952__bF_buf3), .B(data_134__0_), .Y(_3953_) );
NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_3952__bF_buf2), .Y(_3954_) );
AND2X2 AND2X2_824 ( .gnd(gnd), .vdd(vdd), .A(_3953_), .B(_3954_), .Y(_39__0_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_3952__bF_buf1), .B(data_134__1_), .Y(_3955_) );
NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_3952__bF_buf0), .Y(_3956_) );
AND2X2 AND2X2_825 ( .gnd(gnd), .vdd(vdd), .A(_3955_), .B(_3956_), .Y(_39__1_) );
AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf89), .C(data_134__2_), .Y(_3957_) );
AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_3952__bF_buf3), .C(_3957_), .Y(_39__2_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_3952__bF_buf2), .B(data_134__3_), .Y(_3958_) );
NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_3952__bF_buf1), .Y(_3959_) );
AND2X2 AND2X2_826 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(_3959_), .Y(_39__3_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_3952__bF_buf0), .B(data_134__4_), .Y(_3960_) );
NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_3952__bF_buf3), .Y(_3961_) );
AND2X2 AND2X2_827 ( .gnd(gnd), .vdd(vdd), .A(_3960_), .B(_3961_), .Y(_39__4_) );
AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf88), .C(data_134__5_), .Y(_3962_) );
AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_3952__bF_buf2), .C(_3962_), .Y(_39__5_) );
AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf87), .C(data_134__6_), .Y(_3963_) );
AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_3952__bF_buf1), .C(_3963_), .Y(_39__6_) );
AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf86), .C(data_134__7_), .Y(_3964_) );
AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_3952__bF_buf0), .C(_3964_), .Y(_39__7_) );
AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf85), .C(data_134__8_), .Y(_3965_) );
AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_3952__bF_buf3), .C(_3965_), .Y(_39__8_) );
INVX1 INVX1_1843 ( .gnd(gnd), .vdd(vdd), .A(data_134__9_), .Y(_3966_) );
NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf84), .Y(_3967_) );
NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(_3966_), .B(_3967_), .Y(_3968_) );
NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_3952__bF_buf2), .Y(_3969_) );
AND2X2 AND2X2_828 ( .gnd(gnd), .vdd(vdd), .A(_3969_), .B(_3968_), .Y(_39__9_) );
INVX1 INVX1_1844 ( .gnd(gnd), .vdd(vdd), .A(data_134__10_), .Y(_3970_) );
NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_3970_), .B(_3967_), .Y(_3971_) );
NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_3952__bF_buf1), .Y(_3972_) );
AND2X2 AND2X2_829 ( .gnd(gnd), .vdd(vdd), .A(_3972_), .B(_3971_), .Y(_39__10_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_3952__bF_buf0), .B(data_134__11_), .Y(_3973_) );
NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_3952__bF_buf3), .Y(_3974_) );
AND2X2 AND2X2_830 ( .gnd(gnd), .vdd(vdd), .A(_3973_), .B(_3974_), .Y(_39__11_) );
AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf83), .C(data_134__12_), .Y(_3975_) );
AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_3952__bF_buf2), .C(_3975_), .Y(_39__12_) );
INVX1 INVX1_1845 ( .gnd(gnd), .vdd(vdd), .A(data_134__13_), .Y(_3976_) );
NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_3976_), .B(_3967_), .Y(_3977_) );
NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_3952__bF_buf1), .Y(_3978_) );
AND2X2 AND2X2_831 ( .gnd(gnd), .vdd(vdd), .A(_3978_), .B(_3977_), .Y(_39__13_) );
AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf82), .C(data_134__14_), .Y(_3979_) );
AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_3952__bF_buf0), .C(_3979_), .Y(_39__14_) );
AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3313__bF_buf81), .C(data_134__15_), .Y(_3980_) );
AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_3952__bF_buf3), .C(_3980_), .Y(_39__15_) );
INVX1 INVX1_1846 ( .gnd(gnd), .vdd(vdd), .A(data_133__0_), .Y(_3981_) );
OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_14950_), .B(_14954_), .C(_14952__bF_buf3), .Y(_3982_) );
INVX4 INVX4_13 ( .gnd(gnd), .vdd(vdd), .A(_3982_), .Y(_3983_) );
OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(IDATA_PROG_addr_3_bF_buf1), .C(_15065__bF_buf1), .Y(_3984_) );
NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(_3941_), .B(_3984_), .Y(_3985_) );
NOR3X1 NOR3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_3985_), .C(_3632_), .Y(_3986_) );
NAND3X1 NAND3X1_524 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .B(_3395__bF_buf3), .C(_3986_), .Y(_3987_) );
OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_3987_), .C(_3981_), .Y(_3988_) );
NAND3X1 NAND3X1_525 ( .gnd(gnd), .vdd(vdd), .A(_3304_), .B(_3307_), .C(_15041_), .Y(_3989_) );
NOR3X1 NOR3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3987_), .C(_3989__bF_buf4), .Y(_3990_) );
NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_3990_), .Y(_3991_) );
AND2X2 AND2X2_832 ( .gnd(gnd), .vdd(vdd), .A(_3991_), .B(_3988_), .Y(_38__0_) );
INVX1 INVX1_1847 ( .gnd(gnd), .vdd(vdd), .A(data_133__1_), .Y(_3992_) );
OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_3987_), .C(_3992_), .Y(_3993_) );
NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_3990_), .Y(_3994_) );
AND2X2 AND2X2_833 ( .gnd(gnd), .vdd(vdd), .A(_3994_), .B(_3993_), .Y(_38__1_) );
INVX1 INVX1_1848 ( .gnd(gnd), .vdd(vdd), .A(_3949_), .Y(_3995_) );
INVX1 INVX1_1849 ( .gnd(gnd), .vdd(vdd), .A(_3985_), .Y(_3996_) );
NAND3X1 NAND3X1_526 ( .gnd(gnd), .vdd(vdd), .A(_3996_), .B(_3377_), .C(_3365_), .Y(_3997_) );
NOR3X1 NOR3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_3995_), .B(_3997_), .C(_3353__bF_buf3), .Y(_3998_) );
AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf80), .C(data_133__2_), .Y(_3999_) );
AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_3990_), .C(_3999_), .Y(_38__2_) );
INVX1 INVX1_1850 ( .gnd(gnd), .vdd(vdd), .A(data_133__3_), .Y(_4000_) );
OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_3987_), .C(_4000_), .Y(_4001_) );
NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_3990_), .Y(_4002_) );
AND2X2 AND2X2_834 ( .gnd(gnd), .vdd(vdd), .A(_4002_), .B(_4001_), .Y(_38__3_) );
INVX1 INVX1_1851 ( .gnd(gnd), .vdd(vdd), .A(data_133__4_), .Y(_4003_) );
OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_3987_), .C(_4003_), .Y(_4004_) );
NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_3990_), .Y(_4005_) );
AND2X2 AND2X2_835 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(_4004_), .Y(_38__4_) );
AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf79), .C(data_133__5_), .Y(_4006_) );
AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_3990_), .C(_4006_), .Y(_38__5_) );
AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf78), .C(data_133__6_), .Y(_4007_) );
AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_3990_), .C(_4007_), .Y(_38__6_) );
AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf77), .C(data_133__7_), .Y(_4008_) );
AOI21X1 AOI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_3990_), .C(_4008_), .Y(_38__7_) );
AOI21X1 AOI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf76), .C(data_133__8_), .Y(_4009_) );
AOI21X1 AOI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_3990_), .C(_4009_), .Y(_38__8_) );
INVX1 INVX1_1852 ( .gnd(gnd), .vdd(vdd), .A(data_133__9_), .Y(_4010_) );
OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_3987_), .C(_4010_), .Y(_4011_) );
NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_3990_), .Y(_4012_) );
AND2X2 AND2X2_836 ( .gnd(gnd), .vdd(vdd), .A(_4012_), .B(_4011_), .Y(_38__9_) );
INVX1 INVX1_1853 ( .gnd(gnd), .vdd(vdd), .A(data_133__10_), .Y(_4013_) );
OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_3987_), .C(_4013_), .Y(_4014_) );
NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_3990_), .Y(_4015_) );
AND2X2 AND2X2_837 ( .gnd(gnd), .vdd(vdd), .A(_4015_), .B(_4014_), .Y(_38__10_) );
INVX1 INVX1_1854 ( .gnd(gnd), .vdd(vdd), .A(data_133__11_), .Y(_4016_) );
OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_3987_), .C(_4016_), .Y(_4017_) );
NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_3990_), .Y(_4018_) );
AND2X2 AND2X2_838 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .B(_4017_), .Y(_38__11_) );
AOI21X1 AOI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf75), .C(data_133__12_), .Y(_4019_) );
AOI21X1 AOI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_3990_), .C(_4019_), .Y(_38__12_) );
INVX1 INVX1_1855 ( .gnd(gnd), .vdd(vdd), .A(data_133__13_), .Y(_4020_) );
OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_3987_), .C(_4020_), .Y(_4021_) );
NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_3990_), .Y(_4022_) );
AND2X2 AND2X2_839 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(_4021_), .Y(_38__13_) );
AOI21X1 AOI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf74), .C(data_133__14_), .Y(_4023_) );
AOI21X1 AOI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf14), .B(_3990_), .C(_4023_), .Y(_38__14_) );
AOI21X1 AOI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_3998_), .B(_3313__bF_buf73), .C(data_133__15_), .Y(_4024_) );
AOI21X1 AOI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_3990_), .C(_4024_), .Y(_38__15_) );
INVX1 INVX1_1856 ( .gnd(gnd), .vdd(vdd), .A(data_132__0_), .Y(_4025_) );
OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_14980_), .B(_14977__bF_buf2), .C(_3450_), .Y(_4026_) );
INVX1 INVX1_1857 ( .gnd(gnd), .vdd(vdd), .A(_4026_), .Y(_4027_) );
OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_4027_), .B(_14936__bF_buf0), .C(_3984_), .Y(_4028_) );
NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_4028_), .B(_3907_), .Y(_4029_) );
NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_4029_), .Y(_4030_) );
INVX1 INVX1_1858 ( .gnd(gnd), .vdd(vdd), .A(_4030_), .Y(_4031_) );
NAND3X1 NAND3X1_527 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf2), .B(_3633_), .C(_4031_), .Y(_4032_) );
OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf64), .C(_4025_), .Y(_4033_) );
NOR3X1 NOR3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_4030_), .B(_3396_), .C(_3353__bF_buf2), .Y(_4034_) );
NAND3X1 NAND3X1_528 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_4034_), .C(_3313__bF_buf72), .Y(_4035_) );
AND2X2 AND2X2_840 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .B(_4035_), .Y(_37__0_) );
INVX1 INVX1_1859 ( .gnd(gnd), .vdd(vdd), .A(data_132__1_), .Y(_4036_) );
OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf63), .C(_4036_), .Y(_4037_) );
NAND3X1 NAND3X1_529 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_4034_), .C(_3313__bF_buf71), .Y(_4038_) );
AND2X2 AND2X2_841 ( .gnd(gnd), .vdd(vdd), .A(_4037_), .B(_4038_), .Y(_37__1_) );
INVX1 INVX1_1860 ( .gnd(gnd), .vdd(vdd), .A(data_132__2_), .Y(_4039_) );
NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_4034_), .B(_3313__bF_buf70), .Y(_4040_) );
MUX2X1 MUX2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_4039_), .B(_14897__bF_buf7), .S(_4040_), .Y(_37__2_) );
INVX1 INVX1_1861 ( .gnd(gnd), .vdd(vdd), .A(data_132__3_), .Y(_4041_) );
OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf62), .C(_4041_), .Y(_4042_) );
NAND3X1 NAND3X1_530 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_4034_), .C(_3313__bF_buf69), .Y(_4043_) );
AND2X2 AND2X2_842 ( .gnd(gnd), .vdd(vdd), .A(_4042_), .B(_4043_), .Y(_37__3_) );
INVX1 INVX1_1862 ( .gnd(gnd), .vdd(vdd), .A(data_132__4_), .Y(_4044_) );
OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf61), .C(_4044_), .Y(_4045_) );
NAND3X1 NAND3X1_531 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_4034_), .C(_3313__bF_buf68), .Y(_4046_) );
AND2X2 AND2X2_843 ( .gnd(gnd), .vdd(vdd), .A(_4045_), .B(_4046_), .Y(_37__4_) );
INVX1 INVX1_1863 ( .gnd(gnd), .vdd(vdd), .A(data_132__5_), .Y(_4047_) );
OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf60), .C(_4047_), .Y(_4048_) );
NAND3X1 NAND3X1_532 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_4034_), .C(_3313__bF_buf67), .Y(_4049_) );
AND2X2 AND2X2_844 ( .gnd(gnd), .vdd(vdd), .A(_4048_), .B(_4049_), .Y(_37__5_) );
INVX1 INVX1_1864 ( .gnd(gnd), .vdd(vdd), .A(data_132__6_), .Y(_4050_) );
MUX2X1 MUX2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_15049__bF_buf9), .S(_4040_), .Y(_37__6_) );
INVX1 INVX1_1865 ( .gnd(gnd), .vdd(vdd), .A(data_132__7_), .Y(_4051_) );
OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf59), .C(_4051_), .Y(_4052_) );
NAND3X1 NAND3X1_533 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_4034_), .C(_3313__bF_buf66), .Y(_4053_) );
AND2X2 AND2X2_845 ( .gnd(gnd), .vdd(vdd), .A(_4052_), .B(_4053_), .Y(_37__7_) );
INVX1 INVX1_1866 ( .gnd(gnd), .vdd(vdd), .A(data_132__8_), .Y(_4054_) );
MUX2X1 MUX2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_4054_), .B(_15052__bF_buf3), .S(_4040_), .Y(_37__8_) );
INVX1 INVX1_1867 ( .gnd(gnd), .vdd(vdd), .A(data_132__9_), .Y(_4055_) );
MUX2X1 MUX2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_4055_), .B(_14913__bF_buf8), .S(_4040_), .Y(_37__9_) );
INVX1 INVX1_1868 ( .gnd(gnd), .vdd(vdd), .A(data_132__10_), .Y(_4056_) );
MUX2X1 MUX2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_4056_), .B(_15055__bF_buf4), .S(_4040_), .Y(_37__10_) );
INVX1 INVX1_1869 ( .gnd(gnd), .vdd(vdd), .A(data_132__11_), .Y(_4057_) );
OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf58), .C(_4057_), .Y(_4058_) );
NAND3X1 NAND3X1_534 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_4034_), .C(_3313__bF_buf65), .Y(_4059_) );
AND2X2 AND2X2_846 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4059_), .Y(_37__11_) );
INVX1 INVX1_1870 ( .gnd(gnd), .vdd(vdd), .A(data_132__12_), .Y(_4060_) );
OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_4032_), .B(_3393__bF_buf57), .C(_4060_), .Y(_4061_) );
NAND3X1 NAND3X1_535 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_4034_), .C(_3313__bF_buf64), .Y(_4062_) );
AND2X2 AND2X2_847 ( .gnd(gnd), .vdd(vdd), .A(_4061_), .B(_4062_), .Y(_37__12_) );
INVX1 INVX1_1871 ( .gnd(gnd), .vdd(vdd), .A(data_132__13_), .Y(_4063_) );
MUX2X1 MUX2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_4063_), .B(_14924__bF_buf3), .S(_4040_), .Y(_37__13_) );
INVX1 INVX1_1872 ( .gnd(gnd), .vdd(vdd), .A(data_132__14_), .Y(_4064_) );
MUX2X1 MUX2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_4064_), .B(_15060__bF_buf13), .S(_4040_), .Y(_37__14_) );
INVX1 INVX1_1873 ( .gnd(gnd), .vdd(vdd), .A(data_132__15_), .Y(_4065_) );
MUX2X1 MUX2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_4065_), .B(_15062__bF_buf4), .S(_4040_), .Y(_37__15_) );
INVX1 INVX1_1874 ( .gnd(gnd), .vdd(vdd), .A(data_131__0_), .Y(_4066_) );
OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf3), .B(_14942__bF_buf3), .C(_3644_), .Y(_4067_) );
NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_3907_), .B(_4067_), .Y(_4068_) );
NAND3X1 NAND3X1_536 ( .gnd(gnd), .vdd(vdd), .A(_4068_), .B(_3633_), .C(_3395__bF_buf1), .Y(_4069_) );
OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_4069_), .C(_4066_), .Y(_4070_) );
INVX4 INVX4_14 ( .gnd(gnd), .vdd(vdd), .A(_4069_), .Y(_4071_) );
NAND3X1 NAND3X1_537 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_3313__bF_buf63), .C(_4071_), .Y(_4072_) );
AND2X2 AND2X2_848 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(_4072_), .Y(_36__0_) );
INVX1 INVX1_1875 ( .gnd(gnd), .vdd(vdd), .A(data_131__1_), .Y(_4073_) );
OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_4069_), .C(_4073_), .Y(_4074_) );
NAND3X1 NAND3X1_538 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_3313__bF_buf62), .C(_4071_), .Y(_4075_) );
AND2X2 AND2X2_849 ( .gnd(gnd), .vdd(vdd), .A(_4074_), .B(_4075_), .Y(_36__1_) );
INVX1 INVX1_1876 ( .gnd(gnd), .vdd(vdd), .A(data_131__2_), .Y(_4076_) );
NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf61), .B(_4071_), .Y(_4077_) );
MUX2X1 MUX2X1_606 ( .gnd(gnd), .vdd(vdd), .A(_4076_), .B(_14897__bF_buf6), .S(_4077_), .Y(_36__2_) );
INVX1 INVX1_1877 ( .gnd(gnd), .vdd(vdd), .A(data_131__3_), .Y(_4078_) );
OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_4069_), .C(_4078_), .Y(_4079_) );
NAND3X1 NAND3X1_539 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_3313__bF_buf60), .C(_4071_), .Y(_4080_) );
AND2X2 AND2X2_850 ( .gnd(gnd), .vdd(vdd), .A(_4079_), .B(_4080_), .Y(_36__3_) );
INVX1 INVX1_1878 ( .gnd(gnd), .vdd(vdd), .A(data_131__4_), .Y(_4081_) );
OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_4069_), .C(_4081_), .Y(_4082_) );
NAND3X1 NAND3X1_540 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_3313__bF_buf59), .C(_4071_), .Y(_4083_) );
AND2X2 AND2X2_851 ( .gnd(gnd), .vdd(vdd), .A(_4082_), .B(_4083_), .Y(_36__4_) );
INVX1 INVX1_1879 ( .gnd(gnd), .vdd(vdd), .A(data_131__5_), .Y(_4084_) );
OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_4069_), .C(_4084_), .Y(_4085_) );
NAND3X1 NAND3X1_541 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_3313__bF_buf58), .C(_4071_), .Y(_4086_) );
AND2X2 AND2X2_852 ( .gnd(gnd), .vdd(vdd), .A(_4085_), .B(_4086_), .Y(_36__5_) );
INVX1 INVX1_1880 ( .gnd(gnd), .vdd(vdd), .A(data_131__6_), .Y(_4087_) );
MUX2X1 MUX2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_4087_), .B(_15049__bF_buf8), .S(_4077_), .Y(_36__6_) );
INVX1 INVX1_1881 ( .gnd(gnd), .vdd(vdd), .A(data_131__7_), .Y(_4088_) );
OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_4069_), .C(_4088_), .Y(_4089_) );
NAND3X1 NAND3X1_542 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_3313__bF_buf57), .C(_4071_), .Y(_4090_) );
AND2X2 AND2X2_853 ( .gnd(gnd), .vdd(vdd), .A(_4089_), .B(_4090_), .Y(_36__7_) );
INVX1 INVX1_1882 ( .gnd(gnd), .vdd(vdd), .A(data_131__8_), .Y(_4091_) );
MUX2X1 MUX2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_4091_), .B(_15052__bF_buf2), .S(_4077_), .Y(_36__8_) );
INVX1 INVX1_1883 ( .gnd(gnd), .vdd(vdd), .A(data_131__9_), .Y(_4092_) );
MUX2X1 MUX2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_4092_), .B(_14913__bF_buf7), .S(_4077_), .Y(_36__9_) );
INVX1 INVX1_1884 ( .gnd(gnd), .vdd(vdd), .A(data_131__10_), .Y(_4093_) );
MUX2X1 MUX2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_4093_), .B(_15055__bF_buf3), .S(_4077_), .Y(_36__10_) );
INVX1 INVX1_1885 ( .gnd(gnd), .vdd(vdd), .A(data_131__11_), .Y(_4094_) );
OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_4069_), .C(_4094_), .Y(_4095_) );
NAND3X1 NAND3X1_543 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_3313__bF_buf56), .C(_4071_), .Y(_4096_) );
AND2X2 AND2X2_854 ( .gnd(gnd), .vdd(vdd), .A(_4095_), .B(_4096_), .Y(_36__11_) );
INVX1 INVX1_1886 ( .gnd(gnd), .vdd(vdd), .A(data_131__12_), .Y(_4097_) );
OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_4069_), .C(_4097_), .Y(_4098_) );
NAND3X1 NAND3X1_544 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_3313__bF_buf55), .C(_4071_), .Y(_4099_) );
AND2X2 AND2X2_855 ( .gnd(gnd), .vdd(vdd), .A(_4098_), .B(_4099_), .Y(_36__12_) );
INVX1 INVX1_1887 ( .gnd(gnd), .vdd(vdd), .A(data_131__13_), .Y(_4100_) );
MUX2X1 MUX2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_4100_), .B(_14924__bF_buf2), .S(_4077_), .Y(_36__13_) );
INVX1 INVX1_1888 ( .gnd(gnd), .vdd(vdd), .A(data_131__14_), .Y(_4101_) );
MUX2X1 MUX2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_4101_), .B(_15060__bF_buf12), .S(_4077_), .Y(_36__14_) );
INVX1 INVX1_1889 ( .gnd(gnd), .vdd(vdd), .A(data_131__15_), .Y(_4102_) );
MUX2X1 MUX2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_4102_), .B(_15062__bF_buf3), .S(_4077_), .Y(_36__15_) );
INVX1 INVX1_1890 ( .gnd(gnd), .vdd(vdd), .A(data_130__0_), .Y(_4103_) );
NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3644_), .Y(_4104_) );
AOI21X1 AOI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf0), .B(_475_), .C(_4104_), .Y(_4105_) );
NAND3X1 NAND3X1_545 ( .gnd(gnd), .vdd(vdd), .A(_4105_), .B(_3633_), .C(_3395__bF_buf0), .Y(_4106_) );
OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_4106_), .C(_4103_), .Y(_4107_) );
INVX4 INVX4_15 ( .gnd(gnd), .vdd(vdd), .A(_4106_), .Y(_4108_) );
NAND3X1 NAND3X1_546 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_3313__bF_buf54), .C(_4108_), .Y(_4109_) );
AND2X2 AND2X2_856 ( .gnd(gnd), .vdd(vdd), .A(_4107_), .B(_4109_), .Y(_35__0_) );
INVX1 INVX1_1891 ( .gnd(gnd), .vdd(vdd), .A(data_130__1_), .Y(_4110_) );
OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_4106_), .C(_4110_), .Y(_4111_) );
NAND3X1 NAND3X1_547 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_3313__bF_buf53), .C(_4108_), .Y(_4112_) );
AND2X2 AND2X2_857 ( .gnd(gnd), .vdd(vdd), .A(_4111_), .B(_4112_), .Y(_35__1_) );
INVX1 INVX1_1892 ( .gnd(gnd), .vdd(vdd), .A(data_130__2_), .Y(_4113_) );
NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf52), .B(_4108_), .Y(_4114_) );
MUX2X1 MUX2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_4113_), .B(_14897__bF_buf5), .S(_4114_), .Y(_35__2_) );
INVX1 INVX1_1893 ( .gnd(gnd), .vdd(vdd), .A(data_130__3_), .Y(_4115_) );
OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_4106_), .C(_4115_), .Y(_4116_) );
NAND3X1 NAND3X1_548 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_3313__bF_buf51), .C(_4108_), .Y(_4117_) );
AND2X2 AND2X2_858 ( .gnd(gnd), .vdd(vdd), .A(_4116_), .B(_4117_), .Y(_35__3_) );
INVX1 INVX1_1894 ( .gnd(gnd), .vdd(vdd), .A(data_130__4_), .Y(_4118_) );
OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_4106_), .C(_4118_), .Y(_4119_) );
NAND3X1 NAND3X1_549 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_3313__bF_buf50), .C(_4108_), .Y(_4120_) );
AND2X2 AND2X2_859 ( .gnd(gnd), .vdd(vdd), .A(_4119_), .B(_4120_), .Y(_35__4_) );
INVX1 INVX1_1895 ( .gnd(gnd), .vdd(vdd), .A(data_130__5_), .Y(_4121_) );
OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_4106_), .C(_4121_), .Y(_4122_) );
NAND3X1 NAND3X1_550 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_3313__bF_buf49), .C(_4108_), .Y(_4123_) );
AND2X2 AND2X2_860 ( .gnd(gnd), .vdd(vdd), .A(_4122_), .B(_4123_), .Y(_35__5_) );
INVX1 INVX1_1896 ( .gnd(gnd), .vdd(vdd), .A(data_130__6_), .Y(_4124_) );
MUX2X1 MUX2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_4124_), .B(_15049__bF_buf7), .S(_4114_), .Y(_35__6_) );
INVX1 INVX1_1897 ( .gnd(gnd), .vdd(vdd), .A(data_130__7_), .Y(_4125_) );
OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_4106_), .C(_4125_), .Y(_4126_) );
NAND3X1 NAND3X1_551 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_3313__bF_buf48), .C(_4108_), .Y(_4127_) );
AND2X2 AND2X2_861 ( .gnd(gnd), .vdd(vdd), .A(_4126_), .B(_4127_), .Y(_35__7_) );
INVX1 INVX1_1898 ( .gnd(gnd), .vdd(vdd), .A(data_130__8_), .Y(_4128_) );
MUX2X1 MUX2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_4128_), .B(_15052__bF_buf1), .S(_4114_), .Y(_35__8_) );
INVX1 INVX1_1899 ( .gnd(gnd), .vdd(vdd), .A(data_130__9_), .Y(_4129_) );
MUX2X1 MUX2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_4129_), .B(_14913__bF_buf6), .S(_4114_), .Y(_35__9_) );
INVX1 INVX1_1900 ( .gnd(gnd), .vdd(vdd), .A(data_130__10_), .Y(_4130_) );
MUX2X1 MUX2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_4130_), .B(_15055__bF_buf2), .S(_4114_), .Y(_35__10_) );
INVX1 INVX1_1901 ( .gnd(gnd), .vdd(vdd), .A(data_130__11_), .Y(_4131_) );
OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_4106_), .C(_4131_), .Y(_4132_) );
NAND3X1 NAND3X1_552 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_3313__bF_buf47), .C(_4108_), .Y(_4133_) );
AND2X2 AND2X2_862 ( .gnd(gnd), .vdd(vdd), .A(_4132_), .B(_4133_), .Y(_35__11_) );
INVX1 INVX1_1902 ( .gnd(gnd), .vdd(vdd), .A(data_130__12_), .Y(_4134_) );
OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_4106_), .C(_4134_), .Y(_4135_) );
NAND3X1 NAND3X1_553 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_3313__bF_buf46), .C(_4108_), .Y(_4136_) );
AND2X2 AND2X2_863 ( .gnd(gnd), .vdd(vdd), .A(_4135_), .B(_4136_), .Y(_35__12_) );
INVX1 INVX1_1903 ( .gnd(gnd), .vdd(vdd), .A(data_130__13_), .Y(_4137_) );
MUX2X1 MUX2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_4137_), .B(_14924__bF_buf1), .S(_4114_), .Y(_35__13_) );
INVX1 INVX1_1904 ( .gnd(gnd), .vdd(vdd), .A(data_130__14_), .Y(_4138_) );
MUX2X1 MUX2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_4138_), .B(_15060__bF_buf11), .S(_4114_), .Y(_35__14_) );
INVX1 INVX1_1905 ( .gnd(gnd), .vdd(vdd), .A(data_130__15_), .Y(_4139_) );
MUX2X1 MUX2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_4139_), .B(_15062__bF_buf2), .S(_4114_), .Y(_35__15_) );
INVX1 INVX1_1906 ( .gnd(gnd), .vdd(vdd), .A(data_129__0_), .Y(_4140_) );
AOI21X1 AOI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_15065__bF_buf3), .B(_15571_), .C(_4104_), .Y(_4141_) );
NAND3X1 NAND3X1_554 ( .gnd(gnd), .vdd(vdd), .A(_4141_), .B(_3633_), .C(_3395__bF_buf3), .Y(_4142_) );
OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_4142_), .C(_4140_), .Y(_4143_) );
INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(_4142_), .Y(_4144_) );
NAND3X1 NAND3X1_555 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_3313__bF_buf45), .C(_4144_), .Y(_4145_) );
AND2X2 AND2X2_864 ( .gnd(gnd), .vdd(vdd), .A(_4143_), .B(_4145_), .Y(_33__0_) );
INVX1 INVX1_1907 ( .gnd(gnd), .vdd(vdd), .A(data_129__1_), .Y(_4146_) );
OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_4142_), .C(_4146_), .Y(_4147_) );
NAND3X1 NAND3X1_556 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_3313__bF_buf44), .C(_4144_), .Y(_4148_) );
AND2X2 AND2X2_865 ( .gnd(gnd), .vdd(vdd), .A(_4147_), .B(_4148_), .Y(_33__1_) );
NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4142_), .B(_3393__bF_buf38), .Y(_4149_) );
AOI21X1 AOI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf43), .B(_4144_), .C(data_129__2_), .Y(_4150_) );
AOI21X1 AOI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_4149_), .C(_4150_), .Y(_33__2_) );
INVX1 INVX1_1908 ( .gnd(gnd), .vdd(vdd), .A(data_129__3_), .Y(_4151_) );
OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_4142_), .C(_4151_), .Y(_4152_) );
NAND3X1 NAND3X1_557 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_3313__bF_buf42), .C(_4144_), .Y(_4153_) );
AND2X2 AND2X2_866 ( .gnd(gnd), .vdd(vdd), .A(_4152_), .B(_4153_), .Y(_33__3_) );
INVX1 INVX1_1909 ( .gnd(gnd), .vdd(vdd), .A(data_129__4_), .Y(_4154_) );
OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_4142_), .C(_4154_), .Y(_4155_) );
NAND3X1 NAND3X1_558 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_3313__bF_buf41), .C(_4144_), .Y(_4156_) );
AND2X2 AND2X2_867 ( .gnd(gnd), .vdd(vdd), .A(_4155_), .B(_4156_), .Y(_33__4_) );
INVX1 INVX1_1910 ( .gnd(gnd), .vdd(vdd), .A(data_129__5_), .Y(_4157_) );
NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf40), .B(_4144_), .Y(_4158_) );
MUX2X1 MUX2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_4157_), .B(_14903__bF_buf2), .S(_4158_), .Y(_33__5_) );
AOI21X1 AOI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf39), .B(_4144_), .C(data_129__6_), .Y(_4159_) );
AOI21X1 AOI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_4149_), .C(_4159_), .Y(_33__6_) );
INVX1 INVX1_1911 ( .gnd(gnd), .vdd(vdd), .A(data_129__7_), .Y(_4160_) );
MUX2X1 MUX2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_4160_), .B(_14908__bF_buf1), .S(_4158_), .Y(_33__7_) );
AOI21X1 AOI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf38), .B(_4144_), .C(data_129__8_), .Y(_4161_) );
AOI21X1 AOI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_4149_), .C(_4161_), .Y(_33__8_) );
INVX1 INVX1_1912 ( .gnd(gnd), .vdd(vdd), .A(data_129__9_), .Y(_4162_) );
MUX2X1 MUX2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .B(_14913__bF_buf5), .S(_4158_), .Y(_33__9_) );
INVX1 INVX1_1913 ( .gnd(gnd), .vdd(vdd), .A(data_129__10_), .Y(_4163_) );
MUX2X1 MUX2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_4163_), .B(_15055__bF_buf1), .S(_4158_), .Y(_33__10_) );
INVX1 INVX1_1914 ( .gnd(gnd), .vdd(vdd), .A(data_129__11_), .Y(_4164_) );
OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_4142_), .C(_4164_), .Y(_4165_) );
NAND3X1 NAND3X1_559 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_3313__bF_buf37), .C(_4144_), .Y(_4166_) );
AND2X2 AND2X2_868 ( .gnd(gnd), .vdd(vdd), .A(_4165_), .B(_4166_), .Y(_33__11_) );
INVX1 INVX1_1915 ( .gnd(gnd), .vdd(vdd), .A(data_129__12_), .Y(_4167_) );
MUX2X1 MUX2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_4167_), .B(_14920__bF_buf2), .S(_4158_), .Y(_33__12_) );
INVX1 INVX1_1916 ( .gnd(gnd), .vdd(vdd), .A(data_129__13_), .Y(_4168_) );
MUX2X1 MUX2X1_627 ( .gnd(gnd), .vdd(vdd), .A(_4168_), .B(_14924__bF_buf0), .S(_4158_), .Y(_33__13_) );
AOI21X1 AOI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf36), .B(_4144_), .C(data_129__14_), .Y(_4169_) );
AOI21X1 AOI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_4149_), .C(_4169_), .Y(_33__14_) );
AOI21X1 AOI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf35), .B(_4144_), .C(data_129__15_), .Y(_4170_) );
AOI21X1 AOI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_4149_), .C(_4170_), .Y(_33__15_) );
NOR3X1 NOR3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf12), .B(_15030_), .C(_14936__bF_buf2), .Y(_4171_) );
NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_4171__bF_buf4), .Y(_4172_) );
OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(data_128__0_), .B(_4171__bF_buf3), .C(_4172_), .Y(_4173_) );
INVX1 INVX1_1917 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .Y(_32__0_) );
NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_4171__bF_buf2), .Y(_4174_) );
OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(data_128__1_), .B(_4171__bF_buf1), .C(_4174_), .Y(_4175_) );
INVX1 INVX1_1918 ( .gnd(gnd), .vdd(vdd), .A(_4175_), .Y(_32__1_) );
NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(data_128__2_), .B(_4171__bF_buf0), .Y(_4176_) );
AOI21X1 AOI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_4171__bF_buf4), .C(_4176_), .Y(_32__2_) );
NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_4171__bF_buf3), .Y(_4177_) );
OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(data_128__3_), .B(_4171__bF_buf2), .C(_4177_), .Y(_4178_) );
INVX1 INVX1_1919 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .Y(_32__3_) );
NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_4171__bF_buf1), .Y(_4179_) );
OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(data_128__4_), .B(_4171__bF_buf0), .C(_4179_), .Y(_4180_) );
INVX1 INVX1_1920 ( .gnd(gnd), .vdd(vdd), .A(_4180_), .Y(_32__4_) );
NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_4171__bF_buf4), .Y(_4181_) );
OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(data_128__5_), .B(_4171__bF_buf3), .C(_4181_), .Y(_4182_) );
INVX1 INVX1_1921 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .Y(_32__5_) );
NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_4171__bF_buf2), .Y(_4183_) );
OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(data_128__6_), .B(_4171__bF_buf1), .C(_4183_), .Y(_4184_) );
INVX1 INVX1_1922 ( .gnd(gnd), .vdd(vdd), .A(_4184_), .Y(_32__6_) );
NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_4171__bF_buf0), .Y(_4185_) );
OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(data_128__7_), .B(_4171__bF_buf4), .C(_4185_), .Y(_4186_) );
INVX1 INVX1_1923 ( .gnd(gnd), .vdd(vdd), .A(_4186_), .Y(_32__7_) );
NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_4171__bF_buf3), .Y(_4187_) );
OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(data_128__8_), .B(_4171__bF_buf2), .C(_4187_), .Y(_4188_) );
INVX1 INVX1_1924 ( .gnd(gnd), .vdd(vdd), .A(_4188_), .Y(_32__8_) );
NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(data_128__9_), .B(_4171__bF_buf1), .Y(_4189_) );
AOI21X1 AOI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_4171__bF_buf0), .C(_4189_), .Y(_32__9_) );
NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(data_128__10_), .B(_4171__bF_buf4), .Y(_4190_) );
INVX1 INVX1_1925 ( .gnd(gnd), .vdd(vdd), .A(_4171__bF_buf3), .Y(_4191_) );
NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf2), .B(_4191_), .Y(_4192_) );
NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_4190_), .B(_4192_), .Y(_32__10_) );
NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(data_128__11_), .B(_4171__bF_buf2), .Y(_4193_) );
NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf1), .B(_4191_), .Y(_4194_) );
NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_4193_), .B(_4194_), .Y(_32__11_) );
NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_4171__bF_buf1), .Y(_4195_) );
OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(data_128__12_), .B(_4171__bF_buf0), .C(_4195_), .Y(_4196_) );
INVX1 INVX1_1926 ( .gnd(gnd), .vdd(vdd), .A(_4196_), .Y(_32__12_) );
NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_4171__bF_buf4), .Y(_4197_) );
OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(data_128__13_), .B(_4171__bF_buf3), .C(_4197_), .Y(_4198_) );
INVX1 INVX1_1927 ( .gnd(gnd), .vdd(vdd), .A(_4198_), .Y(_32__13_) );
NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(data_128__14_), .B(_4171__bF_buf2), .Y(_4199_) );
AOI21X1 AOI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_4171__bF_buf1), .C(_4199_), .Y(_32__14_) );
NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_4171__bF_buf0), .Y(_4200_) );
OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(data_128__15_), .B(_4171__bF_buf4), .C(_4200_), .Y(_4201_) );
INVX1 INVX1_1928 ( .gnd(gnd), .vdd(vdd), .A(_4201_), .Y(_32__15_) );
NAND3X1 NAND3X1_560 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_14888__bF_buf2), .C(_3370_), .Y(_4202_) );
MUX2X1 MUX2X1_628 ( .gnd(gnd), .vdd(vdd), .A(data_127__0_), .B(IDATA_PROG_data_0_bF_buf1), .S(_4202_), .Y(_4203_) );
INVX1 INVX1_1929 ( .gnd(gnd), .vdd(vdd), .A(_4203_), .Y(_31__0_) );
INVX8 INVX8_27 ( .gnd(gnd), .vdd(vdd), .A(_4202_), .Y(_4204_) );
NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_4204_), .Y(_4205_) );
OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(data_127__1_), .B(_4204_), .C(_4205_), .Y(_4206_) );
INVX1 INVX1_1930 ( .gnd(gnd), .vdd(vdd), .A(_4206_), .Y(_31__1_) );
NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(data_127__2_), .B(_4204_), .Y(_4207_) );
AOI21X1 AOI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_4204_), .C(_4207_), .Y(_31__2_) );
INVX1 INVX1_1931 ( .gnd(gnd), .vdd(vdd), .A(data_127__3_), .Y(_4208_) );
OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf11), .C(_4208_), .Y(_4209_) );
NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_4204_), .Y(_4210_) );
AND2X2 AND2X2_869 ( .gnd(gnd), .vdd(vdd), .A(_4210_), .B(_4209_), .Y(_31__3_) );
INVX1 INVX1_1932 ( .gnd(gnd), .vdd(vdd), .A(data_127__4_), .Y(_4211_) );
OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf10), .C(_4211_), .Y(_4212_) );
OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf3), .B(_4202_), .C(_4212_), .Y(_4213_) );
INVX1 INVX1_1933 ( .gnd(gnd), .vdd(vdd), .A(_4213_), .Y(_31__4_) );
NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_4204_), .Y(_4214_) );
OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(data_127__5_), .B(_4204_), .C(_4214_), .Y(_4215_) );
INVX1 INVX1_1934 ( .gnd(gnd), .vdd(vdd), .A(_4215_), .Y(_31__5_) );
INVX1 INVX1_1935 ( .gnd(gnd), .vdd(vdd), .A(data_127__6_), .Y(_4216_) );
OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf9), .C(_4216_), .Y(_4217_) );
OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf0), .B(_4202_), .C(_4217_), .Y(_4218_) );
INVX1 INVX1_1936 ( .gnd(gnd), .vdd(vdd), .A(_4218_), .Y(_31__6_) );
MUX2X1 MUX2X1_629 ( .gnd(gnd), .vdd(vdd), .A(data_127__7_), .B(IDATA_PROG_data_7_bF_buf0), .S(_4202_), .Y(_4219_) );
INVX1 INVX1_1937 ( .gnd(gnd), .vdd(vdd), .A(_4219_), .Y(_31__7_) );
INVX1 INVX1_1938 ( .gnd(gnd), .vdd(vdd), .A(data_127__8_), .Y(_4220_) );
OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf8), .C(_4220_), .Y(_4221_) );
OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf3), .B(_4202_), .C(_4221_), .Y(_4222_) );
INVX1 INVX1_1939 ( .gnd(gnd), .vdd(vdd), .A(_4222_), .Y(_31__8_) );
INVX1 INVX1_1940 ( .gnd(gnd), .vdd(vdd), .A(data_127__9_), .Y(_4223_) );
OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf7), .C(_4223_), .Y(_4224_) );
OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf1), .B(_4202_), .C(_4224_), .Y(_4225_) );
INVX1 INVX1_1941 ( .gnd(gnd), .vdd(vdd), .A(_4225_), .Y(_31__9_) );
INVX1 INVX1_1942 ( .gnd(gnd), .vdd(vdd), .A(data_127__10_), .Y(_4226_) );
OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf6), .C(_4226_), .Y(_4227_) );
OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf1), .B(_4202_), .C(_4227_), .Y(_4228_) );
INVX1 INVX1_1943 ( .gnd(gnd), .vdd(vdd), .A(_4228_), .Y(_31__10_) );
NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_4204_), .Y(_4229_) );
OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(data_127__11_), .B(_4204_), .C(_4229_), .Y(_4230_) );
INVX1 INVX1_1944 ( .gnd(gnd), .vdd(vdd), .A(_4230_), .Y(_31__11_) );
INVX1 INVX1_1945 ( .gnd(gnd), .vdd(vdd), .A(data_127__12_), .Y(_4231_) );
OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf5), .C(_4231_), .Y(_4232_) );
OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf1), .B(_4202_), .C(_4232_), .Y(_4233_) );
INVX1 INVX1_1946 ( .gnd(gnd), .vdd(vdd), .A(_4233_), .Y(_31__12_) );
INVX1 INVX1_1947 ( .gnd(gnd), .vdd(vdd), .A(data_127__13_), .Y(_4234_) );
OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf4), .C(_4234_), .Y(_4235_) );
OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf3), .B(_4202_), .C(_4235_), .Y(_4236_) );
INVX1 INVX1_1948 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .Y(_31__13_) );
NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_4204_), .Y(_4237_) );
OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(data_127__14_), .B(_4204_), .C(_4237_), .Y(_4238_) );
INVX1 INVX1_1949 ( .gnd(gnd), .vdd(vdd), .A(_4238_), .Y(_31__14_) );
INVX1 INVX1_1950 ( .gnd(gnd), .vdd(vdd), .A(data_127__15_), .Y(_4239_) );
OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .B(_14882__bF_buf3), .C(_4239_), .Y(_4240_) );
OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf0), .B(_4202_), .C(_4240_), .Y(_4241_) );
INVX1 INVX1_1951 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .Y(_31__15_) );
INVX1 INVX1_1952 ( .gnd(gnd), .vdd(vdd), .A(data_126__0_), .Y(_4242_) );
NOR3X1 NOR3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .B(_14967_), .C(_3352_), .Y(_4243_) );
INVX1 INVX1_1953 ( .gnd(gnd), .vdd(vdd), .A(_3635_), .Y(_4244_) );
AOI21X1 AOI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3336_), .C(_14882__bF_buf2), .Y(_4245_) );
OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_3366_), .C(_4245_), .Y(_4246_) );
NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_4246_), .Y(_4247_) );
NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_4247_), .Y(_4248_) );
AOI21X1 AOI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_4244_), .C(_4248_), .Y(_4249_) );
AND2X2 AND2X2_870 ( .gnd(gnd), .vdd(vdd), .A(_4249_), .B(_4243_), .Y(_4250_) );
NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf34), .B(_4250_), .Y(_4251_) );
MUX2X1 MUX2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_4242_), .B(_14932__bF_buf8), .S(_4251_), .Y(_30__0_) );
INVX1 INVX1_1954 ( .gnd(gnd), .vdd(vdd), .A(data_126__1_), .Y(_4252_) );
MUX2X1 MUX2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_4252_), .B(_14894__bF_buf6), .S(_4251_), .Y(_30__1_) );
NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_4243_), .B(_4249_), .Y(_4253_) );
NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4253_), .B(_3393__bF_buf34), .Y(_4254_) );
AOI21X1 AOI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf33), .B(_4250_), .C(data_126__2_), .Y(_4255_) );
AOI21X1 AOI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_4254_), .C(_4255_), .Y(_30__2_) );
INVX1 INVX1_1955 ( .gnd(gnd), .vdd(vdd), .A(data_126__3_), .Y(_4256_) );
MUX2X1 MUX2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_4256_), .B(_14899__bF_buf5), .S(_4251_), .Y(_30__3_) );
INVX1 INVX1_1956 ( .gnd(gnd), .vdd(vdd), .A(data_126__4_), .Y(_4257_) );
MUX2X1 MUX2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_4257_), .B(_14902__bF_buf12), .S(_4251_), .Y(_30__4_) );
AOI21X1 AOI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf32), .B(_4250_), .C(data_126__5_), .Y(_4258_) );
AOI21X1 AOI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_4254_), .C(_4258_), .Y(_30__5_) );
AOI21X1 AOI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf31), .B(_4250_), .C(data_126__6_), .Y(_4259_) );
AOI21X1 AOI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_4254_), .C(_4259_), .Y(_30__6_) );
AOI21X1 AOI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf30), .B(_4250_), .C(data_126__7_), .Y(_4260_) );
AOI21X1 AOI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_4254_), .C(_4260_), .Y(_30__7_) );
AOI21X1 AOI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf29), .B(_4250_), .C(data_126__8_), .Y(_4261_) );
AOI21X1 AOI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_4254_), .C(_4261_), .Y(_30__8_) );
AOI21X1 AOI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf28), .B(_4250_), .C(data_126__9_), .Y(_4262_) );
AOI21X1 AOI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_4254_), .C(_4262_), .Y(_30__9_) );
AOI21X1 AOI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf27), .B(_4250_), .C(data_126__10_), .Y(_4263_) );
AOI21X1 AOI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_4254_), .C(_4263_), .Y(_30__10_) );
INVX1 INVX1_1957 ( .gnd(gnd), .vdd(vdd), .A(data_126__11_), .Y(_4264_) );
MUX2X1 MUX2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_4264_), .B(_14918__bF_buf0), .S(_4251_), .Y(_30__11_) );
AOI21X1 AOI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf26), .B(_4250_), .C(data_126__12_), .Y(_4265_) );
AOI21X1 AOI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_4254_), .C(_4265_), .Y(_30__12_) );
AOI21X1 AOI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf25), .B(_4250_), .C(data_126__13_), .Y(_4266_) );
AOI21X1 AOI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_4254_), .C(_4266_), .Y(_30__13_) );
AOI21X1 AOI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf24), .B(_4250_), .C(data_126__14_), .Y(_4267_) );
AOI21X1 AOI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_4254_), .C(_4267_), .Y(_30__14_) );
AOI21X1 AOI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf23), .B(_4250_), .C(data_126__15_), .Y(_4268_) );
AOI21X1 AOI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_4254_), .C(_4268_), .Y(_30__15_) );
INVX1 INVX1_1958 ( .gnd(gnd), .vdd(vdd), .A(data_125__0_), .Y(_4269_) );
INVX1 INVX1_1959 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .Y(_4270_) );
NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_3322_), .Y(_4271_) );
NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_15030_), .B(_3320_), .Y(_4272_) );
NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_4271_), .B(_4272_), .Y(_4273_) );
INVX1 INVX1_1960 ( .gnd(gnd), .vdd(vdd), .A(_3327_), .Y(_4274_) );
NAND3X1 NAND3X1_561 ( .gnd(gnd), .vdd(vdd), .A(_4270_), .B(_4273_), .C(_4274_), .Y(_4275_) );
NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3331_), .Y(_4276_) );
NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(_3333_), .B(_4276_), .Y(_4277_) );
INVX1 INVX1_1961 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .Y(_4278_) );
NOR3X1 NOR3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_4275_), .B(_4278_), .C(_4277_), .Y(_4279_) );
INVX1 INVX1_1962 ( .gnd(gnd), .vdd(vdd), .A(_3340_), .Y(_4280_) );
INVX1 INVX1_1963 ( .gnd(gnd), .vdd(vdd), .A(_3341_), .Y(_4281_) );
OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf3), .B(_15579_), .C(_3345_), .Y(_4282_) );
AOI21X1 AOI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_14975_), .B(_14998__bF_buf1), .C(_4282_), .Y(_4283_) );
OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf0), .B(_14994_), .C(_14998__bF_buf0), .Y(_4284_) );
NAND3X1 NAND3X1_562 ( .gnd(gnd), .vdd(vdd), .A(_3342_), .B(_4284_), .C(_4283_), .Y(_4285_) );
NOR3X1 NOR3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_4280_), .B(_4281_), .C(_4285_), .Y(_4286_) );
NAND3X1 NAND3X1_563 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_4279_), .C(_4286_), .Y(_4287_) );
NOR3X1 NOR3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_4248_), .C(_4287_), .Y(_4288_) );
NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf22), .B(_4288_), .Y(_4289_) );
MUX2X1 MUX2X1_635 ( .gnd(gnd), .vdd(vdd), .A(_4269_), .B(_14932__bF_buf7), .S(_4289_), .Y(_29__0_) );
INVX1 INVX1_1964 ( .gnd(gnd), .vdd(vdd), .A(data_125__1_), .Y(_4290_) );
MUX2X1 MUX2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_4290_), .B(_14894__bF_buf5), .S(_4289_), .Y(_29__1_) );
AND2X2 AND2X2_871 ( .gnd(gnd), .vdd(vdd), .A(_4288_), .B(_3313__bF_buf21), .Y(_4291_) );
AOI21X1 AOI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf20), .B(_4288_), .C(data_125__2_), .Y(_4292_) );
AOI21X1 AOI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_4291_), .C(_4292_), .Y(_29__2_) );
INVX1 INVX1_1965 ( .gnd(gnd), .vdd(vdd), .A(data_125__3_), .Y(_4293_) );
MUX2X1 MUX2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(_14899__bF_buf4), .S(_4289_), .Y(_29__3_) );
INVX1 INVX1_1966 ( .gnd(gnd), .vdd(vdd), .A(data_125__4_), .Y(_4294_) );
MUX2X1 MUX2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_4294_), .B(_14902__bF_buf11), .S(_4289_), .Y(_29__4_) );
INVX1 INVX1_1967 ( .gnd(gnd), .vdd(vdd), .A(data_125__5_), .Y(_4295_) );
MUX2X1 MUX2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_4295_), .B(_14903__bF_buf12), .S(_4289_), .Y(_29__5_) );
AOI21X1 AOI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf19), .B(_4288_), .C(data_125__6_), .Y(_4296_) );
AOI21X1 AOI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_4291_), .C(_4296_), .Y(_29__6_) );
INVX1 INVX1_1968 ( .gnd(gnd), .vdd(vdd), .A(data_125__7_), .Y(_4297_) );
MUX2X1 MUX2X1_640 ( .gnd(gnd), .vdd(vdd), .A(_4297_), .B(_14908__bF_buf12), .S(_4289_), .Y(_29__7_) );
AOI21X1 AOI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf18), .B(_4288_), .C(data_125__8_), .Y(_4298_) );
AOI21X1 AOI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_4291_), .C(_4298_), .Y(_29__8_) );
AOI21X1 AOI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf17), .B(_4288_), .C(data_125__9_), .Y(_4299_) );
AOI21X1 AOI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_4291_), .C(_4299_), .Y(_29__9_) );
AOI21X1 AOI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf16), .B(_4288_), .C(data_125__10_), .Y(_4300_) );
AOI21X1 AOI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_4291_), .C(_4300_), .Y(_29__10_) );
INVX1 INVX1_1969 ( .gnd(gnd), .vdd(vdd), .A(data_125__11_), .Y(_4301_) );
MUX2X1 MUX2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_4301_), .B(_14918__bF_buf13), .S(_4289_), .Y(_29__11_) );
INVX1 INVX1_1970 ( .gnd(gnd), .vdd(vdd), .A(data_125__12_), .Y(_4302_) );
MUX2X1 MUX2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_4302_), .B(_14920__bF_buf13), .S(_4289_), .Y(_29__12_) );
AOI21X1 AOI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf15), .B(_4288_), .C(data_125__13_), .Y(_4303_) );
AOI21X1 AOI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_4291_), .C(_4303_), .Y(_29__13_) );
AOI21X1 AOI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf14), .B(_4288_), .C(data_125__14_), .Y(_4304_) );
AOI21X1 AOI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_4291_), .C(_4304_), .Y(_29__14_) );
AOI21X1 AOI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf13), .B(_4288_), .C(data_125__15_), .Y(_4305_) );
AOI21X1 AOI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_4291_), .C(_4305_), .Y(_29__15_) );
INVX1 INVX1_1971 ( .gnd(gnd), .vdd(vdd), .A(data_124__0_), .Y(_4306_) );
OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_2672_), .B(_3715_), .C(_3370_), .Y(_4307_) );
NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_4307_), .B(_4245_), .Y(_4308_) );
NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_4308_), .Y(_4309_) );
NAND3X1 NAND3X1_564 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_3365_), .C(_4309_), .Y(_4310_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf1), .B(_4310_), .Y(_4311_) );
OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_4311_), .C(_4306_), .Y(_4312_) );
NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_4310_), .B(_3353__bF_buf0), .Y(_4313_) );
NAND3X1 NAND3X1_565 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_4313_), .C(_3313__bF_buf12), .Y(_4314_) );
AND2X2 AND2X2_872 ( .gnd(gnd), .vdd(vdd), .A(_4312_), .B(_4314_), .Y(_28__0_) );
INVX1 INVX1_1972 ( .gnd(gnd), .vdd(vdd), .A(data_124__1_), .Y(_4315_) );
OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_4311_), .C(_4315_), .Y(_4316_) );
NAND3X1 NAND3X1_566 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_4313_), .C(_3313__bF_buf11), .Y(_4317_) );
AND2X2 AND2X2_873 ( .gnd(gnd), .vdd(vdd), .A(_4316_), .B(_4317_), .Y(_28__1_) );
INVX1 INVX1_1973 ( .gnd(gnd), .vdd(vdd), .A(data_124__2_), .Y(_4318_) );
NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_4313_), .B(_3313__bF_buf10), .Y(_4319_) );
MUX2X1 MUX2X1_643 ( .gnd(gnd), .vdd(vdd), .A(_4318_), .B(_14897__bF_buf14), .S(_4319_), .Y(_28__2_) );
INVX1 INVX1_1974 ( .gnd(gnd), .vdd(vdd), .A(data_124__3_), .Y(_4320_) );
OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_4311_), .C(_4320_), .Y(_4321_) );
NAND3X1 NAND3X1_567 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_4313_), .C(_3313__bF_buf9), .Y(_4322_) );
AND2X2 AND2X2_874 ( .gnd(gnd), .vdd(vdd), .A(_4321_), .B(_4322_), .Y(_28__3_) );
INVX1 INVX1_1975 ( .gnd(gnd), .vdd(vdd), .A(data_124__4_), .Y(_4323_) );
OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_4311_), .C(_4323_), .Y(_4324_) );
NAND3X1 NAND3X1_568 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_4313_), .C(_3313__bF_buf8), .Y(_4325_) );
AND2X2 AND2X2_875 ( .gnd(gnd), .vdd(vdd), .A(_4324_), .B(_4325_), .Y(_28__4_) );
INVX1 INVX1_1976 ( .gnd(gnd), .vdd(vdd), .A(data_124__5_), .Y(_4326_) );
OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_4311_), .C(_4326_), .Y(_4327_) );
NAND3X1 NAND3X1_569 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_4313_), .C(_3313__bF_buf7), .Y(_4328_) );
AND2X2 AND2X2_876 ( .gnd(gnd), .vdd(vdd), .A(_4327_), .B(_4328_), .Y(_28__5_) );
INVX1 INVX1_1977 ( .gnd(gnd), .vdd(vdd), .A(data_124__6_), .Y(_4329_) );
MUX2X1 MUX2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_4329_), .B(_15049__bF_buf2), .S(_4319_), .Y(_28__6_) );
INVX1 INVX1_1978 ( .gnd(gnd), .vdd(vdd), .A(data_124__7_), .Y(_4330_) );
OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_4311_), .C(_4330_), .Y(_4331_) );
NAND3X1 NAND3X1_570 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_4313_), .C(_3313__bF_buf6), .Y(_4332_) );
AND2X2 AND2X2_877 ( .gnd(gnd), .vdd(vdd), .A(_4331_), .B(_4332_), .Y(_28__7_) );
INVX1 INVX1_1979 ( .gnd(gnd), .vdd(vdd), .A(data_124__8_), .Y(_4333_) );
MUX2X1 MUX2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_4333_), .B(_15052__bF_buf10), .S(_4319_), .Y(_28__8_) );
INVX1 INVX1_1980 ( .gnd(gnd), .vdd(vdd), .A(data_124__9_), .Y(_4334_) );
MUX2X1 MUX2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_4334_), .B(_14913__bF_buf1), .S(_4319_), .Y(_28__9_) );
INVX1 INVX1_1981 ( .gnd(gnd), .vdd(vdd), .A(data_124__10_), .Y(_4335_) );
MUX2X1 MUX2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_15055__bF_buf12), .S(_4319_), .Y(_28__10_) );
INVX1 INVX1_1982 ( .gnd(gnd), .vdd(vdd), .A(data_124__11_), .Y(_4336_) );
OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_4311_), .C(_4336_), .Y(_4337_) );
NAND3X1 NAND3X1_571 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_4313_), .C(_3313__bF_buf5), .Y(_4338_) );
AND2X2 AND2X2_878 ( .gnd(gnd), .vdd(vdd), .A(_4337_), .B(_4338_), .Y(_28__11_) );
INVX1 INVX1_1983 ( .gnd(gnd), .vdd(vdd), .A(data_124__12_), .Y(_4339_) );
OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_4311_), .C(_4339_), .Y(_4340_) );
NAND3X1 NAND3X1_572 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_4313_), .C(_3313__bF_buf4), .Y(_4341_) );
AND2X2 AND2X2_879 ( .gnd(gnd), .vdd(vdd), .A(_4340_), .B(_4341_), .Y(_28__12_) );
INVX1 INVX1_1984 ( .gnd(gnd), .vdd(vdd), .A(data_124__13_), .Y(_4342_) );
MUX2X1 MUX2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_4342_), .B(_14924__bF_buf10), .S(_4319_), .Y(_28__13_) );
INVX1 INVX1_1985 ( .gnd(gnd), .vdd(vdd), .A(data_124__14_), .Y(_4343_) );
MUX2X1 MUX2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_15060__bF_buf5), .S(_4319_), .Y(_28__14_) );
INVX1 INVX1_1986 ( .gnd(gnd), .vdd(vdd), .A(data_124__15_), .Y(_4344_) );
MUX2X1 MUX2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_4344_), .B(_15062__bF_buf11), .S(_4319_), .Y(_28__15_) );
INVX1 INVX1_1987 ( .gnd(gnd), .vdd(vdd), .A(data_123__0_), .Y(_4345_) );
INVX1 INVX1_1988 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .Y(_4346_) );
NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf3), .B(_3366_), .Y(_4347_) );
INVX1 INVX1_1989 ( .gnd(gnd), .vdd(vdd), .A(_4347_), .Y(_4348_) );
AND2X2 AND2X2_880 ( .gnd(gnd), .vdd(vdd), .A(_4245_), .B(_4348_), .Y(_4349_) );
NAND3X1 NAND3X1_573 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_4349_), .C(_4346_), .Y(_4350_) );
NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_4350_), .Y(_4351_) );
NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf2), .B(_4351_), .Y(_4352_) );
OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_4352_), .C(_4345_), .Y(_4353_) );
AND2X2 AND2X2_881 ( .gnd(gnd), .vdd(vdd), .A(_4351_), .B(_3395__bF_buf1), .Y(_4354_) );
NAND3X1 NAND3X1_574 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_4354_), .C(_3313__bF_buf3), .Y(_4355_) );
AND2X2 AND2X2_882 ( .gnd(gnd), .vdd(vdd), .A(_4353_), .B(_4355_), .Y(_27__0_) );
INVX1 INVX1_1990 ( .gnd(gnd), .vdd(vdd), .A(data_123__1_), .Y(_4356_) );
OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf24), .B(_4352_), .C(_4356_), .Y(_4357_) );
NAND3X1 NAND3X1_575 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_4354_), .C(_3313__bF_buf2), .Y(_4358_) );
AND2X2 AND2X2_883 ( .gnd(gnd), .vdd(vdd), .A(_4357_), .B(_4358_), .Y(_27__1_) );
INVX1 INVX1_1991 ( .gnd(gnd), .vdd(vdd), .A(data_123__2_), .Y(_4359_) );
NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_3313__bF_buf1), .Y(_4360_) );
MUX2X1 MUX2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_4359_), .B(_14897__bF_buf13), .S(_4360_), .Y(_27__2_) );
INVX1 INVX1_1992 ( .gnd(gnd), .vdd(vdd), .A(data_123__3_), .Y(_4361_) );
OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_4352_), .C(_4361_), .Y(_4362_) );
NAND3X1 NAND3X1_576 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_4354_), .C(_3313__bF_buf0), .Y(_4363_) );
AND2X2 AND2X2_884 ( .gnd(gnd), .vdd(vdd), .A(_4362_), .B(_4363_), .Y(_27__3_) );
INVX1 INVX1_1993 ( .gnd(gnd), .vdd(vdd), .A(data_123__4_), .Y(_4364_) );
OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_4352_), .C(_4364_), .Y(_4365_) );
NAND3X1 NAND3X1_577 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_4354_), .C(_3313__bF_buf91), .Y(_4366_) );
AND2X2 AND2X2_885 ( .gnd(gnd), .vdd(vdd), .A(_4365_), .B(_4366_), .Y(_27__4_) );
INVX1 INVX1_1994 ( .gnd(gnd), .vdd(vdd), .A(data_123__5_), .Y(_4367_) );
OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_4352_), .C(_4367_), .Y(_4368_) );
NAND3X1 NAND3X1_578 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_4354_), .C(_3313__bF_buf90), .Y(_4369_) );
AND2X2 AND2X2_886 ( .gnd(gnd), .vdd(vdd), .A(_4368_), .B(_4369_), .Y(_27__5_) );
INVX1 INVX1_1995 ( .gnd(gnd), .vdd(vdd), .A(data_123__6_), .Y(_4370_) );
MUX2X1 MUX2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_4370_), .B(_15049__bF_buf1), .S(_4360_), .Y(_27__6_) );
INVX1 INVX1_1996 ( .gnd(gnd), .vdd(vdd), .A(data_123__7_), .Y(_4371_) );
OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf20), .B(_4352_), .C(_4371_), .Y(_4372_) );
NAND3X1 NAND3X1_579 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_4354_), .C(_3313__bF_buf89), .Y(_4373_) );
AND2X2 AND2X2_887 ( .gnd(gnd), .vdd(vdd), .A(_4372_), .B(_4373_), .Y(_27__7_) );
INVX1 INVX1_1997 ( .gnd(gnd), .vdd(vdd), .A(data_123__8_), .Y(_4374_) );
MUX2X1 MUX2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_4374_), .B(_15052__bF_buf9), .S(_4360_), .Y(_27__8_) );
INVX1 INVX1_1998 ( .gnd(gnd), .vdd(vdd), .A(data_123__9_), .Y(_4375_) );
MUX2X1 MUX2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_4375_), .B(_14913__bF_buf0), .S(_4360_), .Y(_27__9_) );
INVX1 INVX1_1999 ( .gnd(gnd), .vdd(vdd), .A(data_123__10_), .Y(_4376_) );
MUX2X1 MUX2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_4376_), .B(_15055__bF_buf11), .S(_4360_), .Y(_27__10_) );
INVX1 INVX1_2000 ( .gnd(gnd), .vdd(vdd), .A(data_123__11_), .Y(_4377_) );
OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_4352_), .C(_4377_), .Y(_4378_) );
NAND3X1 NAND3X1_580 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_4354_), .C(_3313__bF_buf88), .Y(_4379_) );
AND2X2 AND2X2_888 ( .gnd(gnd), .vdd(vdd), .A(_4378_), .B(_4379_), .Y(_27__11_) );
INVX1 INVX1_2001 ( .gnd(gnd), .vdd(vdd), .A(data_123__12_), .Y(_4380_) );
OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_4352_), .C(_4380_), .Y(_4381_) );
NAND3X1 NAND3X1_581 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_4354_), .C(_3313__bF_buf87), .Y(_4382_) );
AND2X2 AND2X2_889 ( .gnd(gnd), .vdd(vdd), .A(_4381_), .B(_4382_), .Y(_27__12_) );
INVX1 INVX1_2002 ( .gnd(gnd), .vdd(vdd), .A(data_123__13_), .Y(_4383_) );
MUX2X1 MUX2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_4383_), .B(_14924__bF_buf9), .S(_4360_), .Y(_27__13_) );
INVX1 INVX1_2003 ( .gnd(gnd), .vdd(vdd), .A(data_123__14_), .Y(_4384_) );
MUX2X1 MUX2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(_15060__bF_buf4), .S(_4360_), .Y(_27__14_) );
INVX1 INVX1_2004 ( .gnd(gnd), .vdd(vdd), .A(data_123__15_), .Y(_4385_) );
MUX2X1 MUX2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_15062__bF_buf10), .S(_4360_), .Y(_27__15_) );
INVX1 INVX1_2005 ( .gnd(gnd), .vdd(vdd), .A(data_122__0_), .Y(_4386_) );
OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(_14884_), .C(IDATA_PROG_write_bF_buf5), .Y(_4387_) );
NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_16204_), .Y(_4388_) );
OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf2), .B(_3366_), .C(_4388_), .Y(_4389_) );
AOI21X1 AOI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .B(_4389_), .C(_3374_), .Y(_4390_) );
NAND3X1 NAND3X1_582 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_3365_), .C(_4390_), .Y(_4391_) );
NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_4391_), .B(_3353__bF_buf4), .Y(_4392_) );
INVX4 INVX4_16 ( .gnd(gnd), .vdd(vdd), .A(_4392_), .Y(_4393_) );
OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf17), .C(_4386_), .Y(_4394_) );
NAND3X1 NAND3X1_583 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_4392_), .C(_3313__bF_buf86), .Y(_4395_) );
AND2X2 AND2X2_890 ( .gnd(gnd), .vdd(vdd), .A(_4394_), .B(_4395_), .Y(_26__0_) );
INVX1 INVX1_2006 ( .gnd(gnd), .vdd(vdd), .A(data_122__1_), .Y(_4396_) );
OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf16), .C(_4396_), .Y(_4397_) );
NAND3X1 NAND3X1_584 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_4392_), .C(_3313__bF_buf85), .Y(_4398_) );
AND2X2 AND2X2_891 ( .gnd(gnd), .vdd(vdd), .A(_4397_), .B(_4398_), .Y(_26__1_) );
INVX1 INVX1_2007 ( .gnd(gnd), .vdd(vdd), .A(data_122__2_), .Y(_4399_) );
NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_4392_), .B(_3313__bF_buf84), .Y(_4400_) );
MUX2X1 MUX2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_4399_), .B(_14897__bF_buf12), .S(_4400_), .Y(_26__2_) );
INVX1 INVX1_2008 ( .gnd(gnd), .vdd(vdd), .A(data_122__3_), .Y(_4401_) );
OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf15), .C(_4401_), .Y(_4402_) );
NAND3X1 NAND3X1_585 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_4392_), .C(_3313__bF_buf83), .Y(_4403_) );
AND2X2 AND2X2_892 ( .gnd(gnd), .vdd(vdd), .A(_4402_), .B(_4403_), .Y(_26__3_) );
INVX1 INVX1_2009 ( .gnd(gnd), .vdd(vdd), .A(data_122__4_), .Y(_4404_) );
OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf14), .C(_4404_), .Y(_4405_) );
NAND3X1 NAND3X1_586 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_4392_), .C(_3313__bF_buf82), .Y(_4406_) );
AND2X2 AND2X2_893 ( .gnd(gnd), .vdd(vdd), .A(_4405_), .B(_4406_), .Y(_26__4_) );
INVX1 INVX1_2010 ( .gnd(gnd), .vdd(vdd), .A(data_122__5_), .Y(_4407_) );
OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf13), .C(_4407_), .Y(_4408_) );
NAND3X1 NAND3X1_587 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_4392_), .C(_3313__bF_buf81), .Y(_4409_) );
AND2X2 AND2X2_894 ( .gnd(gnd), .vdd(vdd), .A(_4408_), .B(_4409_), .Y(_26__5_) );
INVX1 INVX1_2011 ( .gnd(gnd), .vdd(vdd), .A(data_122__6_), .Y(_4410_) );
MUX2X1 MUX2X1_660 ( .gnd(gnd), .vdd(vdd), .A(_4410_), .B(_15049__bF_buf0), .S(_4400_), .Y(_26__6_) );
INVX1 INVX1_2012 ( .gnd(gnd), .vdd(vdd), .A(data_122__7_), .Y(_4411_) );
OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf12), .C(_4411_), .Y(_4412_) );
NAND3X1 NAND3X1_588 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_4392_), .C(_3313__bF_buf80), .Y(_4413_) );
AND2X2 AND2X2_895 ( .gnd(gnd), .vdd(vdd), .A(_4412_), .B(_4413_), .Y(_26__7_) );
INVX1 INVX1_2013 ( .gnd(gnd), .vdd(vdd), .A(data_122__8_), .Y(_4414_) );
MUX2X1 MUX2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_4414_), .B(_15052__bF_buf8), .S(_4400_), .Y(_26__8_) );
INVX1 INVX1_2014 ( .gnd(gnd), .vdd(vdd), .A(data_122__9_), .Y(_4415_) );
MUX2X1 MUX2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_4415_), .B(_14913__bF_buf14), .S(_4400_), .Y(_26__9_) );
INVX1 INVX1_2015 ( .gnd(gnd), .vdd(vdd), .A(data_122__10_), .Y(_4416_) );
MUX2X1 MUX2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_4416_), .B(_15055__bF_buf10), .S(_4400_), .Y(_26__10_) );
INVX1 INVX1_2016 ( .gnd(gnd), .vdd(vdd), .A(data_122__11_), .Y(_4417_) );
OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf11), .C(_4417_), .Y(_4418_) );
NAND3X1 NAND3X1_589 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_4392_), .C(_3313__bF_buf79), .Y(_4419_) );
AND2X2 AND2X2_896 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .B(_4419_), .Y(_26__11_) );
INVX1 INVX1_2017 ( .gnd(gnd), .vdd(vdd), .A(data_122__12_), .Y(_4420_) );
OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_3393__bF_buf10), .C(_4420_), .Y(_4421_) );
NAND3X1 NAND3X1_590 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_4392_), .C(_3313__bF_buf78), .Y(_4422_) );
AND2X2 AND2X2_897 ( .gnd(gnd), .vdd(vdd), .A(_4421_), .B(_4422_), .Y(_26__12_) );
INVX1 INVX1_2018 ( .gnd(gnd), .vdd(vdd), .A(data_122__13_), .Y(_4423_) );
MUX2X1 MUX2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .B(_14924__bF_buf8), .S(_4400_), .Y(_26__13_) );
INVX1 INVX1_2019 ( .gnd(gnd), .vdd(vdd), .A(data_122__14_), .Y(_4424_) );
MUX2X1 MUX2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .B(_15060__bF_buf3), .S(_4400_), .Y(_26__14_) );
INVX1 INVX1_2020 ( .gnd(gnd), .vdd(vdd), .A(data_122__15_), .Y(_4425_) );
MUX2X1 MUX2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_4425_), .B(_15062__bF_buf9), .S(_4400_), .Y(_26__15_) );
INVX1 INVX1_2021 ( .gnd(gnd), .vdd(vdd), .A(data_121__0_), .Y(_4426_) );
OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_14989_), .B(_14949_), .C(IDATA_PROG_write_bF_buf4), .Y(_4427_) );
INVX1 INVX1_2022 ( .gnd(gnd), .vdd(vdd), .A(_4427_), .Y(_4428_) );
NAND3X1 NAND3X1_591 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf1), .B(_14958_), .C(_4428_), .Y(_4429_) );
AOI21X1 AOI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .B(_4429_), .C(_3374_), .Y(_4430_) );
NAND3X1 NAND3X1_592 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_4430_), .C(_3365_), .Y(_4431_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf3), .B(_4431_), .Y(_4432_) );
OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_4432_), .C(_4426_), .Y(_4433_) );
NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_4431_), .B(_3353__bF_buf2), .Y(_4434_) );
NAND3X1 NAND3X1_593 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_4434_), .C(_3313__bF_buf77), .Y(_4435_) );
AND2X2 AND2X2_898 ( .gnd(gnd), .vdd(vdd), .A(_4433_), .B(_4435_), .Y(_25__0_) );
INVX1 INVX1_2023 ( .gnd(gnd), .vdd(vdd), .A(data_121__1_), .Y(_4436_) );
OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf8), .B(_4432_), .C(_4436_), .Y(_4437_) );
NAND3X1 NAND3X1_594 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_4434_), .C(_3313__bF_buf76), .Y(_4438_) );
AND2X2 AND2X2_899 ( .gnd(gnd), .vdd(vdd), .A(_4437_), .B(_4438_), .Y(_25__1_) );
INVX1 INVX1_2024 ( .gnd(gnd), .vdd(vdd), .A(data_121__2_), .Y(_4439_) );
NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_3313__bF_buf75), .Y(_4440_) );
MUX2X1 MUX2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_4439_), .B(_14897__bF_buf11), .S(_4440_), .Y(_25__2_) );
INVX1 INVX1_2025 ( .gnd(gnd), .vdd(vdd), .A(data_121__3_), .Y(_4441_) );
OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_4432_), .C(_4441_), .Y(_4442_) );
NAND3X1 NAND3X1_595 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_4434_), .C(_3313__bF_buf74), .Y(_4443_) );
AND2X2 AND2X2_900 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_4443_), .Y(_25__3_) );
INVX1 INVX1_2026 ( .gnd(gnd), .vdd(vdd), .A(data_121__4_), .Y(_4444_) );
OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_4432_), .C(_4444_), .Y(_4445_) );
NAND3X1 NAND3X1_596 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_4434_), .C(_3313__bF_buf73), .Y(_4446_) );
AND2X2 AND2X2_901 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_4446_), .Y(_25__4_) );
INVX1 INVX1_2027 ( .gnd(gnd), .vdd(vdd), .A(data_121__5_), .Y(_4447_) );
OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_4432_), .C(_4447_), .Y(_4448_) );
NAND3X1 NAND3X1_597 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_4434_), .C(_3313__bF_buf72), .Y(_4449_) );
AND2X2 AND2X2_902 ( .gnd(gnd), .vdd(vdd), .A(_4448_), .B(_4449_), .Y(_25__5_) );
INVX1 INVX1_2028 ( .gnd(gnd), .vdd(vdd), .A(data_121__6_), .Y(_4450_) );
MUX2X1 MUX2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_4450_), .B(_15049__bF_buf14), .S(_4440_), .Y(_25__6_) );
INVX1 INVX1_2029 ( .gnd(gnd), .vdd(vdd), .A(data_121__7_), .Y(_4451_) );
OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_4432_), .C(_4451_), .Y(_4452_) );
NAND3X1 NAND3X1_598 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_4434_), .C(_3313__bF_buf71), .Y(_4453_) );
AND2X2 AND2X2_903 ( .gnd(gnd), .vdd(vdd), .A(_4452_), .B(_4453_), .Y(_25__7_) );
INVX1 INVX1_2030 ( .gnd(gnd), .vdd(vdd), .A(data_121__8_), .Y(_4454_) );
MUX2X1 MUX2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_4454_), .B(_15052__bF_buf7), .S(_4440_), .Y(_25__8_) );
INVX1 INVX1_2031 ( .gnd(gnd), .vdd(vdd), .A(data_121__9_), .Y(_4455_) );
MUX2X1 MUX2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_4455_), .B(_14913__bF_buf13), .S(_4440_), .Y(_25__9_) );
INVX1 INVX1_2032 ( .gnd(gnd), .vdd(vdd), .A(data_121__10_), .Y(_4456_) );
MUX2X1 MUX2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_15055__bF_buf9), .S(_4440_), .Y(_25__10_) );
INVX1 INVX1_2033 ( .gnd(gnd), .vdd(vdd), .A(data_121__11_), .Y(_4457_) );
OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf3), .B(_4432_), .C(_4457_), .Y(_4458_) );
NAND3X1 NAND3X1_599 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_4434_), .C(_3313__bF_buf70), .Y(_4459_) );
AND2X2 AND2X2_904 ( .gnd(gnd), .vdd(vdd), .A(_4458_), .B(_4459_), .Y(_25__11_) );
INVX1 INVX1_2034 ( .gnd(gnd), .vdd(vdd), .A(data_121__12_), .Y(_4460_) );
OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_4432_), .C(_4460_), .Y(_4461_) );
NAND3X1 NAND3X1_600 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_4434_), .C(_3313__bF_buf69), .Y(_4462_) );
AND2X2 AND2X2_905 ( .gnd(gnd), .vdd(vdd), .A(_4461_), .B(_4462_), .Y(_25__12_) );
INVX1 INVX1_2035 ( .gnd(gnd), .vdd(vdd), .A(data_121__13_), .Y(_4463_) );
MUX2X1 MUX2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_4463_), .B(_14924__bF_buf7), .S(_4440_), .Y(_25__13_) );
INVX1 INVX1_2036 ( .gnd(gnd), .vdd(vdd), .A(data_121__14_), .Y(_4464_) );
MUX2X1 MUX2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_4464_), .B(_15060__bF_buf2), .S(_4440_), .Y(_25__14_) );
INVX1 INVX1_2037 ( .gnd(gnd), .vdd(vdd), .A(data_121__15_), .Y(_4465_) );
MUX2X1 MUX2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_4465_), .B(_15062__bF_buf8), .S(_4440_), .Y(_25__15_) );
INVX1 INVX1_2038 ( .gnd(gnd), .vdd(vdd), .A(data_120__0_), .Y(_4466_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .Y(_4467_) );
NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_4427_), .B(_4467_), .Y(_4468_) );
OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf0), .B(_3366_), .C(_4468_), .Y(_4469_) );
AOI21X1 AOI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .B(_4469_), .C(_3374_), .Y(_4470_) );
NAND3X1 NAND3X1_601 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_3365_), .C(_4470_), .Y(_4471_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_4471_), .B(_3353__bF_buf1), .Y(_4472_) );
OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_4472_), .C(_4466_), .Y(_4473_) );
NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf0), .B(_4471_), .Y(_4474_) );
NAND3X1 NAND3X1_602 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_4474_), .C(_3313__bF_buf68), .Y(_4475_) );
AND2X2 AND2X2_906 ( .gnd(gnd), .vdd(vdd), .A(_4473_), .B(_4475_), .Y(_24__0_) );
INVX1 INVX1_2039 ( .gnd(gnd), .vdd(vdd), .A(data_120__1_), .Y(_4476_) );
OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_4472_), .C(_4476_), .Y(_4477_) );
NAND3X1 NAND3X1_603 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_4474_), .C(_3313__bF_buf67), .Y(_4478_) );
AND2X2 AND2X2_907 ( .gnd(gnd), .vdd(vdd), .A(_4477_), .B(_4478_), .Y(_24__1_) );
INVX1 INVX1_2040 ( .gnd(gnd), .vdd(vdd), .A(data_120__2_), .Y(_4479_) );
NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_4474_), .B(_3313__bF_buf66), .Y(_4480_) );
MUX2X1 MUX2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_14897__bF_buf10), .S(_4480_), .Y(_24__2_) );
INVX1 INVX1_2041 ( .gnd(gnd), .vdd(vdd), .A(data_120__3_), .Y(_4481_) );
OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_4472_), .C(_4481_), .Y(_4482_) );
NAND3X1 NAND3X1_604 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_4474_), .C(_3313__bF_buf65), .Y(_4483_) );
AND2X2 AND2X2_908 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4483_), .Y(_24__3_) );
INVX1 INVX1_2042 ( .gnd(gnd), .vdd(vdd), .A(data_120__4_), .Y(_4484_) );
OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_4472_), .C(_4484_), .Y(_4485_) );
NAND3X1 NAND3X1_605 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_4474_), .C(_3313__bF_buf64), .Y(_4486_) );
AND2X2 AND2X2_909 ( .gnd(gnd), .vdd(vdd), .A(_4485_), .B(_4486_), .Y(_24__4_) );
INVX1 INVX1_2043 ( .gnd(gnd), .vdd(vdd), .A(data_120__5_), .Y(_4487_) );
OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_4472_), .C(_4487_), .Y(_4488_) );
NAND3X1 NAND3X1_606 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_4474_), .C(_3313__bF_buf63), .Y(_4489_) );
AND2X2 AND2X2_910 ( .gnd(gnd), .vdd(vdd), .A(_4488_), .B(_4489_), .Y(_24__5_) );
INVX1 INVX1_2044 ( .gnd(gnd), .vdd(vdd), .A(data_120__6_), .Y(_4490_) );
MUX2X1 MUX2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_4490_), .B(_15049__bF_buf13), .S(_4480_), .Y(_24__6_) );
INVX1 INVX1_2045 ( .gnd(gnd), .vdd(vdd), .A(data_120__7_), .Y(_4491_) );
OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_4472_), .C(_4491_), .Y(_4492_) );
NAND3X1 NAND3X1_607 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_4474_), .C(_3313__bF_buf62), .Y(_4493_) );
AND2X2 AND2X2_911 ( .gnd(gnd), .vdd(vdd), .A(_4492_), .B(_4493_), .Y(_24__7_) );
INVX1 INVX1_2046 ( .gnd(gnd), .vdd(vdd), .A(data_120__8_), .Y(_4494_) );
MUX2X1 MUX2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_4494_), .B(_15052__bF_buf6), .S(_4480_), .Y(_24__8_) );
INVX1 INVX1_2047 ( .gnd(gnd), .vdd(vdd), .A(data_120__9_), .Y(_4495_) );
MUX2X1 MUX2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_4495_), .B(_14913__bF_buf12), .S(_4480_), .Y(_24__9_) );
INVX1 INVX1_2048 ( .gnd(gnd), .vdd(vdd), .A(data_120__10_), .Y(_4496_) );
MUX2X1 MUX2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_4496_), .B(_15055__bF_buf8), .S(_4480_), .Y(_24__10_) );
INVX1 INVX1_2049 ( .gnd(gnd), .vdd(vdd), .A(data_120__11_), .Y(_4497_) );
OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_4472_), .C(_4497_), .Y(_4498_) );
NAND3X1 NAND3X1_608 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_4474_), .C(_3313__bF_buf61), .Y(_4499_) );
AND2X2 AND2X2_912 ( .gnd(gnd), .vdd(vdd), .A(_4498_), .B(_4499_), .Y(_24__11_) );
INVX1 INVX1_2050 ( .gnd(gnd), .vdd(vdd), .A(data_120__12_), .Y(_4500_) );
OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_4472_), .C(_4500_), .Y(_4501_) );
NAND3X1 NAND3X1_609 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_4474_), .C(_3313__bF_buf60), .Y(_4502_) );
AND2X2 AND2X2_913 ( .gnd(gnd), .vdd(vdd), .A(_4501_), .B(_4502_), .Y(_24__12_) );
INVX1 INVX1_2051 ( .gnd(gnd), .vdd(vdd), .A(data_120__13_), .Y(_4503_) );
MUX2X1 MUX2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_4503_), .B(_14924__bF_buf6), .S(_4480_), .Y(_24__13_) );
INVX1 INVX1_2052 ( .gnd(gnd), .vdd(vdd), .A(data_120__14_), .Y(_4504_) );
MUX2X1 MUX2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_4504_), .B(_15060__bF_buf1), .S(_4480_), .Y(_24__14_) );
INVX1 INVX1_2053 ( .gnd(gnd), .vdd(vdd), .A(data_120__15_), .Y(_4505_) );
MUX2X1 MUX2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_15062__bF_buf7), .S(_4480_), .Y(_24__15_) );
OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_3357_), .C(_3371_), .Y(_4506_) );
OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_14956_), .C(IDATA_PROG_write_bF_buf3), .Y(_4507_) );
NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_4507_), .B(_4506_), .Y(_4508_) );
NAND3X1 NAND3X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3368_), .B(_3373_), .C(_4508_), .Y(_4509_) );
NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .B(_4509_), .Y(_4510_) );
NAND3X1 NAND3X1_611 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_4510_), .C(_3395__bF_buf0), .Y(_4511_) );
NOR3X1 NOR3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_4511_), .C(_3989__bF_buf3), .Y(_4512_) );
NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_4510_), .Y(_4513_) );
NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf4), .B(_4513_), .Y(_4514_) );
AOI21X1 AOI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf59), .C(data_119__0_), .Y(_4515_) );
AOI21X1 AOI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_4512_), .C(_4515_), .Y(_22__0_) );
AOI21X1 AOI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf58), .C(data_119__1_), .Y(_4516_) );
AOI21X1 AOI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_4512_), .C(_4516_), .Y(_22__1_) );
AOI21X1 AOI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf57), .C(data_119__2_), .Y(_4517_) );
AOI21X1 AOI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_4512_), .C(_4517_), .Y(_22__2_) );
AOI21X1 AOI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf56), .C(data_119__3_), .Y(_4518_) );
AOI21X1 AOI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_4512_), .C(_4518_), .Y(_22__3_) );
AOI21X1 AOI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf55), .C(data_119__4_), .Y(_4519_) );
AOI21X1 AOI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_4512_), .C(_4519_), .Y(_22__4_) );
INVX1 INVX1_2054 ( .gnd(gnd), .vdd(vdd), .A(data_119__5_), .Y(_4520_) );
NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf54), .Y(_4521_) );
MUX2X1 MUX2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_4520_), .B(_14903__bF_buf6), .S(_4521_), .Y(_22__5_) );
AOI21X1 AOI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf53), .C(data_119__6_), .Y(_4522_) );
AOI21X1 AOI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_4512_), .C(_4522_), .Y(_22__6_) );
INVX1 INVX1_2055 ( .gnd(gnd), .vdd(vdd), .A(data_119__7_), .Y(_4523_) );
MUX2X1 MUX2X1_684 ( .gnd(gnd), .vdd(vdd), .A(_4523_), .B(_14908__bF_buf6), .S(_4521_), .Y(_22__7_) );
AOI21X1 AOI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf52), .C(data_119__8_), .Y(_4524_) );
AOI21X1 AOI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_4512_), .C(_4524_), .Y(_22__8_) );
AOI21X1 AOI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf51), .C(data_119__9_), .Y(_4525_) );
AOI21X1 AOI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_4512_), .C(_4525_), .Y(_22__9_) );
AOI21X1 AOI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf50), .C(data_119__10_), .Y(_4526_) );
AOI21X1 AOI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_4512_), .C(_4526_), .Y(_22__10_) );
AOI21X1 AOI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf49), .C(data_119__11_), .Y(_4527_) );
AOI21X1 AOI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_4512_), .C(_4527_), .Y(_22__11_) );
INVX1 INVX1_2056 ( .gnd(gnd), .vdd(vdd), .A(data_119__12_), .Y(_4528_) );
MUX2X1 MUX2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_4528_), .B(_14920__bF_buf7), .S(_4521_), .Y(_22__12_) );
AOI21X1 AOI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf48), .C(data_119__13_), .Y(_4529_) );
AOI21X1 AOI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_4512_), .C(_4529_), .Y(_22__13_) );
AOI21X1 AOI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf47), .C(data_119__14_), .Y(_4530_) );
AOI21X1 AOI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_4512_), .C(_4530_), .Y(_22__14_) );
AOI21X1 AOI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_4514_), .B(_3313__bF_buf46), .C(data_119__15_), .Y(_4531_) );
AOI21X1 AOI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_4512_), .C(_4531_), .Y(_22__15_) );
INVX1 INVX1_2057 ( .gnd(gnd), .vdd(vdd), .A(data_118__0_), .Y(_4532_) );
OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_3366_), .C(IDATA_PROG_write_bF_buf2), .Y(_4533_) );
NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .B(_4506_), .Y(_4534_) );
NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf0), .B(_3943_), .Y(_4535_) );
OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_4535_), .C(_4534_), .Y(_4536_) );
NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_4533_), .B(_4536_), .Y(_4537_) );
NAND3X1 NAND3X1_612 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_3365_), .C(_4537_), .Y(_4538_) );
NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf3), .B(_4538_), .Y(_4539_) );
NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_3313__bF_buf45), .Y(_4540_) );
MUX2X1 MUX2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_4532_), .B(_14932__bF_buf0), .S(_4540_), .Y(_21__0_) );
INVX1 INVX1_2058 ( .gnd(gnd), .vdd(vdd), .A(data_118__1_), .Y(_4541_) );
MUX2X1 MUX2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_4541_), .B(_14894__bF_buf13), .S(_4540_), .Y(_21__1_) );
INVX1 INVX1_2059 ( .gnd(gnd), .vdd(vdd), .A(data_118__2_), .Y(_4542_) );
MUX2X1 MUX2X1_688 ( .gnd(gnd), .vdd(vdd), .A(_4542_), .B(_14897__bF_buf8), .S(_4540_), .Y(_21__2_) );
INVX1 INVX1_2060 ( .gnd(gnd), .vdd(vdd), .A(data_118__3_), .Y(_4543_) );
MUX2X1 MUX2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_4543_), .B(_14899__bF_buf12), .S(_4540_), .Y(_21__3_) );
INVX1 INVX1_2061 ( .gnd(gnd), .vdd(vdd), .A(data_118__4_), .Y(_4544_) );
MUX2X1 MUX2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_4544_), .B(_14902__bF_buf4), .S(_4540_), .Y(_21__4_) );
INVX1 INVX1_2062 ( .gnd(gnd), .vdd(vdd), .A(data_118__5_), .Y(_4545_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_4538_), .B(_3353__bF_buf2), .Y(_4546_) );
OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_4546_), .C(_4545_), .Y(_4547_) );
NAND3X1 NAND3X1_613 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_4539_), .C(_3313__bF_buf44), .Y(_4548_) );
AND2X2 AND2X2_914 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .B(_4548_), .Y(_21__5_) );
INVX1 INVX1_2063 ( .gnd(gnd), .vdd(vdd), .A(data_118__6_), .Y(_4549_) );
MUX2X1 MUX2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_4549_), .B(_15049__bF_buf11), .S(_4540_), .Y(_21__6_) );
INVX1 INVX1_2064 ( .gnd(gnd), .vdd(vdd), .A(data_118__7_), .Y(_4550_) );
OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_4546_), .C(_4550_), .Y(_4551_) );
NAND3X1 NAND3X1_614 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_4539_), .C(_3313__bF_buf43), .Y(_4552_) );
AND2X2 AND2X2_915 ( .gnd(gnd), .vdd(vdd), .A(_4551_), .B(_4552_), .Y(_21__7_) );
INVX1 INVX1_2065 ( .gnd(gnd), .vdd(vdd), .A(data_118__8_), .Y(_4553_) );
MUX2X1 MUX2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_4553_), .B(_15052__bF_buf4), .S(_4540_), .Y(_21__8_) );
NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_4546_), .B(_3393__bF_buf61), .Y(_4554_) );
AOI21X1 AOI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_3313__bF_buf42), .C(data_118__9_), .Y(_4555_) );
AOI21X1 AOI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_4554_), .C(_4555_), .Y(_21__9_) );
AOI21X1 AOI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_3313__bF_buf41), .C(data_118__10_), .Y(_4556_) );
AOI21X1 AOI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_4554_), .C(_4556_), .Y(_21__10_) );
INVX1 INVX1_2066 ( .gnd(gnd), .vdd(vdd), .A(data_118__11_), .Y(_4557_) );
MUX2X1 MUX2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_4557_), .B(_14918__bF_buf6), .S(_4540_), .Y(_21__11_) );
INVX1 INVX1_2067 ( .gnd(gnd), .vdd(vdd), .A(data_118__12_), .Y(_4558_) );
OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_4546_), .C(_4558_), .Y(_4559_) );
NAND3X1 NAND3X1_615 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_4539_), .C(_3313__bF_buf40), .Y(_4560_) );
AND2X2 AND2X2_916 ( .gnd(gnd), .vdd(vdd), .A(_4559_), .B(_4560_), .Y(_21__12_) );
AOI21X1 AOI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_3313__bF_buf39), .C(data_118__13_), .Y(_4561_) );
AOI21X1 AOI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_4554_), .C(_4561_), .Y(_21__13_) );
INVX1 INVX1_2068 ( .gnd(gnd), .vdd(vdd), .A(data_118__14_), .Y(_4562_) );
MUX2X1 MUX2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_15060__bF_buf14), .S(_4540_), .Y(_21__14_) );
INVX1 INVX1_2069 ( .gnd(gnd), .vdd(vdd), .A(data_118__15_), .Y(_4563_) );
MUX2X1 MUX2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_4563_), .B(_15062__bF_buf5), .S(_4540_), .Y(_21__15_) );
INVX1 INVX1_2070 ( .gnd(gnd), .vdd(vdd), .A(data_117__0_), .Y(_4564_) );
OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(IDATA_PROG_addr_3_bF_buf3), .C(_3370_), .Y(_4565_) );
NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_4565_), .B(_4534_), .Y(_4566_) );
NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_4533_), .B(_4566_), .Y(_4567_) );
NAND3X1 NAND3X1_616 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_3365_), .C(_4567_), .Y(_4568_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_4568_), .B(_3353__bF_buf1), .Y(_4569_) );
OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_4569_), .C(_4564_), .Y(_4570_) );
NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf0), .B(_4568_), .Y(_4571_) );
NAND3X1 NAND3X1_617 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_4571_), .C(_3313__bF_buf38), .Y(_4572_) );
AND2X2 AND2X2_917 ( .gnd(gnd), .vdd(vdd), .A(_4570_), .B(_4572_), .Y(_20__0_) );
INVX1 INVX1_2071 ( .gnd(gnd), .vdd(vdd), .A(data_117__1_), .Y(_4573_) );
OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_4569_), .C(_4573_), .Y(_4574_) );
NAND3X1 NAND3X1_618 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_4571_), .C(_3313__bF_buf37), .Y(_4575_) );
AND2X2 AND2X2_918 ( .gnd(gnd), .vdd(vdd), .A(_4574_), .B(_4575_), .Y(_20__1_) );
INVX1 INVX1_2072 ( .gnd(gnd), .vdd(vdd), .A(data_117__2_), .Y(_4576_) );
NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_4571_), .B(_3313__bF_buf36), .Y(_4577_) );
MUX2X1 MUX2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_14897__bF_buf7), .S(_4577_), .Y(_20__2_) );
INVX1 INVX1_2073 ( .gnd(gnd), .vdd(vdd), .A(data_117__3_), .Y(_4578_) );
OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_4569_), .C(_4578_), .Y(_4579_) );
NAND3X1 NAND3X1_619 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_4571_), .C(_3313__bF_buf35), .Y(_4580_) );
AND2X2 AND2X2_919 ( .gnd(gnd), .vdd(vdd), .A(_4579_), .B(_4580_), .Y(_20__3_) );
INVX1 INVX1_2074 ( .gnd(gnd), .vdd(vdd), .A(data_117__4_), .Y(_4581_) );
OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_4569_), .C(_4581_), .Y(_4582_) );
NAND3X1 NAND3X1_620 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_4571_), .C(_3313__bF_buf34), .Y(_4583_) );
AND2X2 AND2X2_920 ( .gnd(gnd), .vdd(vdd), .A(_4582_), .B(_4583_), .Y(_20__4_) );
INVX1 INVX1_2075 ( .gnd(gnd), .vdd(vdd), .A(data_117__5_), .Y(_4584_) );
OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_4569_), .C(_4584_), .Y(_4585_) );
NAND3X1 NAND3X1_621 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_4571_), .C(_3313__bF_buf33), .Y(_4586_) );
AND2X2 AND2X2_921 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .B(_4586_), .Y(_20__5_) );
INVX1 INVX1_2076 ( .gnd(gnd), .vdd(vdd), .A(data_117__6_), .Y(_4587_) );
MUX2X1 MUX2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_4587_), .B(_15049__bF_buf10), .S(_4577_), .Y(_20__6_) );
INVX1 INVX1_2077 ( .gnd(gnd), .vdd(vdd), .A(data_117__7_), .Y(_4588_) );
OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_4569_), .C(_4588_), .Y(_4589_) );
NAND3X1 NAND3X1_622 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_4571_), .C(_3313__bF_buf32), .Y(_4590_) );
AND2X2 AND2X2_922 ( .gnd(gnd), .vdd(vdd), .A(_4589_), .B(_4590_), .Y(_20__7_) );
INVX1 INVX1_2078 ( .gnd(gnd), .vdd(vdd), .A(data_117__8_), .Y(_4591_) );
MUX2X1 MUX2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_4591_), .B(_15052__bF_buf3), .S(_4577_), .Y(_20__8_) );
INVX1 INVX1_2079 ( .gnd(gnd), .vdd(vdd), .A(data_117__9_), .Y(_4592_) );
MUX2X1 MUX2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_4592_), .B(_14913__bF_buf9), .S(_4577_), .Y(_20__9_) );
INVX1 INVX1_2080 ( .gnd(gnd), .vdd(vdd), .A(data_117__10_), .Y(_4593_) );
MUX2X1 MUX2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_4593_), .B(_15055__bF_buf5), .S(_4577_), .Y(_20__10_) );
INVX1 INVX1_2081 ( .gnd(gnd), .vdd(vdd), .A(data_117__11_), .Y(_4594_) );
OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_4569_), .C(_4594_), .Y(_4595_) );
NAND3X1 NAND3X1_623 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_4571_), .C(_3313__bF_buf31), .Y(_4596_) );
AND2X2 AND2X2_923 ( .gnd(gnd), .vdd(vdd), .A(_4595_), .B(_4596_), .Y(_20__11_) );
INVX1 INVX1_2082 ( .gnd(gnd), .vdd(vdd), .A(data_117__12_), .Y(_4597_) );
OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_4569_), .C(_4597_), .Y(_4598_) );
NAND3X1 NAND3X1_624 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_4571_), .C(_3313__bF_buf30), .Y(_4599_) );
AND2X2 AND2X2_924 ( .gnd(gnd), .vdd(vdd), .A(_4598_), .B(_4599_), .Y(_20__12_) );
INVX1 INVX1_2083 ( .gnd(gnd), .vdd(vdd), .A(data_117__13_), .Y(_4600_) );
MUX2X1 MUX2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_4600_), .B(_14924__bF_buf3), .S(_4577_), .Y(_20__13_) );
INVX1 INVX1_2084 ( .gnd(gnd), .vdd(vdd), .A(data_117__14_), .Y(_4601_) );
MUX2X1 MUX2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_4601_), .B(_15060__bF_buf13), .S(_4577_), .Y(_20__14_) );
INVX1 INVX1_2085 ( .gnd(gnd), .vdd(vdd), .A(data_117__15_), .Y(_4602_) );
MUX2X1 MUX2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_4602_), .B(_15062__bF_buf4), .S(_4577_), .Y(_20__15_) );
INVX1 INVX1_2086 ( .gnd(gnd), .vdd(vdd), .A(data_116__0_), .Y(_4603_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .Y(_4604_) );
OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_14977__bF_buf1), .B(_14949_), .C(IDATA_PROG_write_bF_buf1), .Y(_4605_) );
NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_4605_), .B(_4026_), .Y(_4606_) );
OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_4604_), .B(_4606_), .C(_4534_), .Y(_4607_) );
AOI21X1 AOI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf2), .B(_3370_), .C(_4607_), .Y(_4608_) );
NAND3X1 NAND3X1_625 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_3365_), .C(_4608_), .Y(_4609_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_4609_), .B(_3353__bF_buf4), .Y(_4610_) );
OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_4610_), .C(_4603_), .Y(_4611_) );
NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf3), .B(_4609_), .Y(_4612_) );
NAND3X1 NAND3X1_626 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_4612_), .C(_3313__bF_buf29), .Y(_4613_) );
AND2X2 AND2X2_925 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_4613_), .Y(_19__0_) );
INVX1 INVX1_2087 ( .gnd(gnd), .vdd(vdd), .A(data_116__1_), .Y(_4614_) );
OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_4610_), .C(_4614_), .Y(_4615_) );
NAND3X1 NAND3X1_627 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_4612_), .C(_3313__bF_buf28), .Y(_4616_) );
AND2X2 AND2X2_926 ( .gnd(gnd), .vdd(vdd), .A(_4615_), .B(_4616_), .Y(_19__1_) );
INVX1 INVX1_2088 ( .gnd(gnd), .vdd(vdd), .A(data_116__2_), .Y(_4617_) );
NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_4612_), .B(_3313__bF_buf27), .Y(_4618_) );
MUX2X1 MUX2X1_704 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_14897__bF_buf6), .S(_4618_), .Y(_19__2_) );
INVX1 INVX1_2089 ( .gnd(gnd), .vdd(vdd), .A(data_116__3_), .Y(_4619_) );
OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_4610_), .C(_4619_), .Y(_4620_) );
NAND3X1 NAND3X1_628 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_4612_), .C(_3313__bF_buf26), .Y(_4621_) );
AND2X2 AND2X2_927 ( .gnd(gnd), .vdd(vdd), .A(_4620_), .B(_4621_), .Y(_19__3_) );
INVX1 INVX1_2090 ( .gnd(gnd), .vdd(vdd), .A(data_116__4_), .Y(_4622_) );
OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_4610_), .C(_4622_), .Y(_4623_) );
NAND3X1 NAND3X1_629 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_4612_), .C(_3313__bF_buf25), .Y(_4624_) );
AND2X2 AND2X2_928 ( .gnd(gnd), .vdd(vdd), .A(_4623_), .B(_4624_), .Y(_19__4_) );
INVX1 INVX1_2091 ( .gnd(gnd), .vdd(vdd), .A(data_116__5_), .Y(_4625_) );
OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_4610_), .C(_4625_), .Y(_4626_) );
NAND3X1 NAND3X1_630 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_4612_), .C(_3313__bF_buf24), .Y(_4627_) );
AND2X2 AND2X2_929 ( .gnd(gnd), .vdd(vdd), .A(_4626_), .B(_4627_), .Y(_19__5_) );
INVX1 INVX1_2092 ( .gnd(gnd), .vdd(vdd), .A(data_116__6_), .Y(_4628_) );
MUX2X1 MUX2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_4628_), .B(_15049__bF_buf9), .S(_4618_), .Y(_19__6_) );
INVX1 INVX1_2093 ( .gnd(gnd), .vdd(vdd), .A(data_116__7_), .Y(_4629_) );
OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_4610_), .C(_4629_), .Y(_4630_) );
NAND3X1 NAND3X1_631 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_4612_), .C(_3313__bF_buf23), .Y(_4631_) );
AND2X2 AND2X2_930 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(_4631_), .Y(_19__7_) );
INVX1 INVX1_2094 ( .gnd(gnd), .vdd(vdd), .A(data_116__8_), .Y(_4632_) );
MUX2X1 MUX2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_4632_), .B(_15052__bF_buf2), .S(_4618_), .Y(_19__8_) );
INVX1 INVX1_2095 ( .gnd(gnd), .vdd(vdd), .A(data_116__9_), .Y(_4633_) );
MUX2X1 MUX2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_4633_), .B(_14913__bF_buf8), .S(_4618_), .Y(_19__9_) );
INVX1 INVX1_2096 ( .gnd(gnd), .vdd(vdd), .A(data_116__10_), .Y(_4634_) );
MUX2X1 MUX2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .B(_15055__bF_buf4), .S(_4618_), .Y(_19__10_) );
INVX1 INVX1_2097 ( .gnd(gnd), .vdd(vdd), .A(data_116__11_), .Y(_4635_) );
OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_4610_), .C(_4635_), .Y(_4636_) );
NAND3X1 NAND3X1_632 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_4612_), .C(_3313__bF_buf22), .Y(_4637_) );
AND2X2 AND2X2_931 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_4637_), .Y(_19__11_) );
INVX1 INVX1_2098 ( .gnd(gnd), .vdd(vdd), .A(data_116__12_), .Y(_4638_) );
OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_4610_), .C(_4638_), .Y(_4639_) );
NAND3X1 NAND3X1_633 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_4612_), .C(_3313__bF_buf21), .Y(_4640_) );
AND2X2 AND2X2_932 ( .gnd(gnd), .vdd(vdd), .A(_4639_), .B(_4640_), .Y(_19__12_) );
INVX1 INVX1_2099 ( .gnd(gnd), .vdd(vdd), .A(data_116__13_), .Y(_4641_) );
MUX2X1 MUX2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_4641_), .B(_14924__bF_buf2), .S(_4618_), .Y(_19__13_) );
INVX1 INVX1_2100 ( .gnd(gnd), .vdd(vdd), .A(data_116__14_), .Y(_4642_) );
MUX2X1 MUX2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_4642_), .B(_15060__bF_buf12), .S(_4618_), .Y(_19__14_) );
INVX1 INVX1_2101 ( .gnd(gnd), .vdd(vdd), .A(data_116__15_), .Y(_4643_) );
MUX2X1 MUX2X1_711 ( .gnd(gnd), .vdd(vdd), .A(_4643_), .B(_15062__bF_buf3), .S(_4618_), .Y(_19__15_) );
INVX1 INVX1_2102 ( .gnd(gnd), .vdd(vdd), .A(data_115__0_), .Y(_4644_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_4506_), .B(_4507_), .Y(_4645_) );
NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_3367_), .B(_4645_), .Y(_4646_) );
AOI21X1 AOI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf2), .B(_3370_), .C(_3631_), .Y(_4647_) );
NAND3X1 NAND3X1_634 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_4646_), .C(_4647_), .Y(_4648_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_4648_), .B(_3353__bF_buf2), .Y(_4649_) );
OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_4649_), .C(_4644_), .Y(_4650_) );
NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf1), .B(_4648_), .Y(_4651_) );
NAND3X1 NAND3X1_635 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_4651_), .C(_3313__bF_buf20), .Y(_4652_) );
AND2X2 AND2X2_933 ( .gnd(gnd), .vdd(vdd), .A(_4650_), .B(_4652_), .Y(_18__0_) );
INVX1 INVX1_2103 ( .gnd(gnd), .vdd(vdd), .A(data_115__1_), .Y(_4653_) );
OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_4649_), .C(_4653_), .Y(_4654_) );
NAND3X1 NAND3X1_636 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_4651_), .C(_3313__bF_buf19), .Y(_4655_) );
AND2X2 AND2X2_934 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4655_), .Y(_18__1_) );
INVX1 INVX1_2104 ( .gnd(gnd), .vdd(vdd), .A(data_115__2_), .Y(_4656_) );
NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_3313__bF_buf18), .Y(_4657_) );
MUX2X1 MUX2X1_712 ( .gnd(gnd), .vdd(vdd), .A(_4656_), .B(_14897__bF_buf5), .S(_4657_), .Y(_18__2_) );
INVX1 INVX1_2105 ( .gnd(gnd), .vdd(vdd), .A(data_115__3_), .Y(_4658_) );
OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_4649_), .C(_4658_), .Y(_4659_) );
NAND3X1 NAND3X1_637 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_4651_), .C(_3313__bF_buf17), .Y(_4660_) );
AND2X2 AND2X2_935 ( .gnd(gnd), .vdd(vdd), .A(_4659_), .B(_4660_), .Y(_18__3_) );
INVX1 INVX1_2106 ( .gnd(gnd), .vdd(vdd), .A(data_115__4_), .Y(_4661_) );
OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_4649_), .C(_4661_), .Y(_4662_) );
NAND3X1 NAND3X1_638 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_4651_), .C(_3313__bF_buf16), .Y(_4663_) );
AND2X2 AND2X2_936 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_4663_), .Y(_18__4_) );
INVX1 INVX1_2107 ( .gnd(gnd), .vdd(vdd), .A(data_115__5_), .Y(_4664_) );
OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_4649_), .C(_4664_), .Y(_4665_) );
NAND3X1 NAND3X1_639 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_4651_), .C(_3313__bF_buf15), .Y(_4666_) );
AND2X2 AND2X2_937 ( .gnd(gnd), .vdd(vdd), .A(_4665_), .B(_4666_), .Y(_18__5_) );
INVX1 INVX1_2108 ( .gnd(gnd), .vdd(vdd), .A(data_115__6_), .Y(_4667_) );
MUX2X1 MUX2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .B(_15049__bF_buf8), .S(_4657_), .Y(_18__6_) );
INVX1 INVX1_2109 ( .gnd(gnd), .vdd(vdd), .A(data_115__7_), .Y(_4668_) );
OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_4649_), .C(_4668_), .Y(_4669_) );
NAND3X1 NAND3X1_640 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_4651_), .C(_3313__bF_buf14), .Y(_4670_) );
AND2X2 AND2X2_938 ( .gnd(gnd), .vdd(vdd), .A(_4669_), .B(_4670_), .Y(_18__7_) );
INVX1 INVX1_2110 ( .gnd(gnd), .vdd(vdd), .A(data_115__8_), .Y(_4671_) );
MUX2X1 MUX2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_4671_), .B(_15052__bF_buf1), .S(_4657_), .Y(_18__8_) );
INVX1 INVX1_2111 ( .gnd(gnd), .vdd(vdd), .A(data_115__9_), .Y(_4672_) );
MUX2X1 MUX2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_4672_), .B(_14913__bF_buf7), .S(_4657_), .Y(_18__9_) );
INVX1 INVX1_2112 ( .gnd(gnd), .vdd(vdd), .A(data_115__10_), .Y(_4673_) );
MUX2X1 MUX2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_4673_), .B(_15055__bF_buf3), .S(_4657_), .Y(_18__10_) );
INVX1 INVX1_2113 ( .gnd(gnd), .vdd(vdd), .A(data_115__11_), .Y(_4674_) );
OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_4649_), .C(_4674_), .Y(_4675_) );
NAND3X1 NAND3X1_641 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_4651_), .C(_3313__bF_buf13), .Y(_4676_) );
AND2X2 AND2X2_939 ( .gnd(gnd), .vdd(vdd), .A(_4675_), .B(_4676_), .Y(_18__11_) );
INVX1 INVX1_2114 ( .gnd(gnd), .vdd(vdd), .A(data_115__12_), .Y(_4677_) );
OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_4649_), .C(_4677_), .Y(_4678_) );
NAND3X1 NAND3X1_642 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_4651_), .C(_3313__bF_buf12), .Y(_4679_) );
AND2X2 AND2X2_940 ( .gnd(gnd), .vdd(vdd), .A(_4678_), .B(_4679_), .Y(_18__12_) );
INVX1 INVX1_2115 ( .gnd(gnd), .vdd(vdd), .A(data_115__13_), .Y(_4680_) );
MUX2X1 MUX2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_4680_), .B(_14924__bF_buf1), .S(_4657_), .Y(_18__13_) );
INVX1 INVX1_2116 ( .gnd(gnd), .vdd(vdd), .A(data_115__14_), .Y(_4681_) );
MUX2X1 MUX2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_4681_), .B(_15060__bF_buf11), .S(_4657_), .Y(_18__14_) );
INVX1 INVX1_2117 ( .gnd(gnd), .vdd(vdd), .A(data_115__15_), .Y(_4682_) );
MUX2X1 MUX2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_4682_), .B(_15062__bF_buf2), .S(_4657_), .Y(_18__15_) );
OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[0]), .B(IDATA_PROG_addr[2]), .C(_14956_), .Y(_4683_) );
OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_4683_), .C(_4508_), .Y(_4684_) );
NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_14967_), .B(_4684_), .Y(_4685_) );
NAND3X1 NAND3X1_643 ( .gnd(gnd), .vdd(vdd), .A(_3365_), .B(_4685_), .C(_3395__bF_buf3), .Y(_4686_) );
NOR3X1 NOR3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_4686_), .C(_3989__bF_buf2), .Y(_4687_) );
INVX8 INVX8_28 ( .gnd(gnd), .vdd(vdd), .A(_4686_), .Y(_4688_) );
AOI21X1 AOI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf11), .B(_4688_), .C(data_114__0_), .Y(_4689_) );
AOI21X1 AOI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_4687_), .C(_4689_), .Y(_17__0_) );
AOI21X1 AOI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf10), .B(_4688_), .C(data_114__1_), .Y(_4690_) );
AOI21X1 AOI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_4687_), .C(_4690_), .Y(_17__1_) );
INVX1 INVX1_2118 ( .gnd(gnd), .vdd(vdd), .A(data_114__2_), .Y(_4691_) );
OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_4686_), .C(_4691_), .Y(_4692_) );
NAND3X1 NAND3X1_644 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_3313__bF_buf9), .C(_4688_), .Y(_4693_) );
AND2X2 AND2X2_941 ( .gnd(gnd), .vdd(vdd), .A(_4692_), .B(_4693_), .Y(_17__2_) );
AOI21X1 AOI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf8), .B(_4688_), .C(data_114__3_), .Y(_4694_) );
AOI21X1 AOI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_4687_), .C(_4694_), .Y(_17__3_) );
AOI21X1 AOI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf7), .B(_4688_), .C(data_114__4_), .Y(_4695_) );
AOI21X1 AOI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_4687_), .C(_4695_), .Y(_17__4_) );
INVX1 INVX1_2119 ( .gnd(gnd), .vdd(vdd), .A(data_114__5_), .Y(_4696_) );
OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf34), .B(_4686_), .C(_4696_), .Y(_4697_) );
NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_4687_), .Y(_4698_) );
AND2X2 AND2X2_942 ( .gnd(gnd), .vdd(vdd), .A(_4698_), .B(_4697_), .Y(_17__5_) );
INVX1 INVX1_2120 ( .gnd(gnd), .vdd(vdd), .A(data_114__6_), .Y(_4699_) );
OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_4686_), .C(_4699_), .Y(_4700_) );
NAND3X1 NAND3X1_645 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_3313__bF_buf6), .C(_4688_), .Y(_4701_) );
AND2X2 AND2X2_943 ( .gnd(gnd), .vdd(vdd), .A(_4700_), .B(_4701_), .Y(_17__6_) );
INVX1 INVX1_2121 ( .gnd(gnd), .vdd(vdd), .A(data_114__7_), .Y(_4702_) );
OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_4686_), .C(_4702_), .Y(_4703_) );
NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_4687_), .Y(_4704_) );
AND2X2 AND2X2_944 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4703_), .Y(_17__7_) );
INVX1 INVX1_2122 ( .gnd(gnd), .vdd(vdd), .A(data_114__8_), .Y(_4705_) );
OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_4686_), .C(_4705_), .Y(_4706_) );
NAND3X1 NAND3X1_646 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_3313__bF_buf5), .C(_4688_), .Y(_4707_) );
AND2X2 AND2X2_945 ( .gnd(gnd), .vdd(vdd), .A(_4706_), .B(_4707_), .Y(_17__8_) );
AOI21X1 AOI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf4), .B(_4688_), .C(data_114__9_), .Y(_4708_) );
AOI21X1 AOI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_4687_), .C(_4708_), .Y(_17__9_) );
AOI21X1 AOI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf3), .B(_4688_), .C(data_114__10_), .Y(_4709_) );
AOI21X1 AOI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_4687_), .C(_4709_), .Y(_17__10_) );
AOI21X1 AOI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf2), .B(_4688_), .C(data_114__11_), .Y(_4710_) );
AOI21X1 AOI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_4687_), .C(_4710_), .Y(_17__11_) );
INVX1 INVX1_2123 ( .gnd(gnd), .vdd(vdd), .A(data_114__12_), .Y(_4711_) );
OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_4686_), .C(_4711_), .Y(_4712_) );
NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_4687_), .Y(_4713_) );
AND2X2 AND2X2_946 ( .gnd(gnd), .vdd(vdd), .A(_4713_), .B(_4712_), .Y(_17__12_) );
AOI21X1 AOI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf1), .B(_4688_), .C(data_114__13_), .Y(_4714_) );
AOI21X1 AOI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_4687_), .C(_4714_), .Y(_17__13_) );
INVX1 INVX1_2124 ( .gnd(gnd), .vdd(vdd), .A(data_114__14_), .Y(_4715_) );
OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_4686_), .C(_4715_), .Y(_4716_) );
NAND3X1 NAND3X1_647 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_3313__bF_buf0), .C(_4688_), .Y(_4717_) );
AND2X2 AND2X2_947 ( .gnd(gnd), .vdd(vdd), .A(_4716_), .B(_4717_), .Y(_17__14_) );
INVX1 INVX1_2125 ( .gnd(gnd), .vdd(vdd), .A(data_114__15_), .Y(_4718_) );
OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_4686_), .C(_4718_), .Y(_4719_) );
NAND3X1 NAND3X1_648 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_3313__bF_buf91), .C(_4688_), .Y(_4720_) );
AND2X2 AND2X2_948 ( .gnd(gnd), .vdd(vdd), .A(_4719_), .B(_4720_), .Y(_17__15_) );
INVX1 INVX1_2126 ( .gnd(gnd), .vdd(vdd), .A(data_113__0_), .Y(_4721_) );
OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr[1]), .B(IDATA_PROG_addr[2]), .C(_14956_), .Y(_4722_) );
INVX1 INVX1_2127 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .Y(_4723_) );
AOI21X1 AOI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_4723_), .C(_4645_), .Y(_4724_) );
NAND3X1 NAND3X1_649 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_4724_), .C(_3365_), .Y(_4725_) );
NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_4725_), .B(_3353__bF_buf0), .Y(_4726_) );
NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf90), .Y(_4727_) );
NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_4721_), .B(_4727_), .Y(_4728_) );
AND2X2 AND2X2_949 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf89), .B(_4726_), .Y(_4729_) );
NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_4729_), .Y(_4730_) );
AND2X2 AND2X2_950 ( .gnd(gnd), .vdd(vdd), .A(_4730_), .B(_4728_), .Y(_16__0_) );
INVX1 INVX1_2128 ( .gnd(gnd), .vdd(vdd), .A(data_113__1_), .Y(_4731_) );
NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_4731_), .B(_4727_), .Y(_4732_) );
NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_4729_), .Y(_4733_) );
AND2X2 AND2X2_951 ( .gnd(gnd), .vdd(vdd), .A(_4733_), .B(_4732_), .Y(_16__1_) );
AOI21X1 AOI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf88), .C(data_113__2_), .Y(_4734_) );
AOI21X1 AOI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_4729_), .C(_4734_), .Y(_16__2_) );
INVX1 INVX1_2129 ( .gnd(gnd), .vdd(vdd), .A(data_113__3_), .Y(_4735_) );
NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_4735_), .B(_4727_), .Y(_4736_) );
NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_4729_), .Y(_4737_) );
AND2X2 AND2X2_952 ( .gnd(gnd), .vdd(vdd), .A(_4737_), .B(_4736_), .Y(_16__3_) );
INVX1 INVX1_2130 ( .gnd(gnd), .vdd(vdd), .A(data_113__4_), .Y(_4738_) );
NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_4738_), .B(_4727_), .Y(_4739_) );
NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_4729_), .Y(_4740_) );
AND2X2 AND2X2_953 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(_4739_), .Y(_16__4_) );
AOI21X1 AOI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf87), .C(data_113__5_), .Y(_4741_) );
AOI21X1 AOI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_4729_), .C(_4741_), .Y(_16__5_) );
AOI21X1 AOI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf86), .C(data_113__6_), .Y(_4742_) );
AOI21X1 AOI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_4729_), .C(_4742_), .Y(_16__6_) );
AOI21X1 AOI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf85), .C(data_113__7_), .Y(_4743_) );
AOI21X1 AOI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_4729_), .C(_4743_), .Y(_16__7_) );
AOI21X1 AOI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf84), .C(data_113__8_), .Y(_4744_) );
AOI21X1 AOI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_4729_), .C(_4744_), .Y(_16__8_) );
INVX1 INVX1_2131 ( .gnd(gnd), .vdd(vdd), .A(data_113__9_), .Y(_4745_) );
NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_4745_), .B(_4727_), .Y(_4746_) );
NAND3X1 NAND3X1_650 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_4726_), .C(_3313__bF_buf83), .Y(_4747_) );
AND2X2 AND2X2_954 ( .gnd(gnd), .vdd(vdd), .A(_4746_), .B(_4747_), .Y(_16__9_) );
INVX1 INVX1_2132 ( .gnd(gnd), .vdd(vdd), .A(data_113__10_), .Y(_4748_) );
NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_4748_), .B(_4727_), .Y(_4749_) );
NAND3X1 NAND3X1_651 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_4726_), .C(_3313__bF_buf82), .Y(_4750_) );
AND2X2 AND2X2_955 ( .gnd(gnd), .vdd(vdd), .A(_4749_), .B(_4750_), .Y(_16__10_) );
INVX1 INVX1_2133 ( .gnd(gnd), .vdd(vdd), .A(data_113__11_), .Y(_4751_) );
NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_4751_), .B(_4727_), .Y(_4752_) );
NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_4729_), .Y(_4753_) );
AND2X2 AND2X2_956 ( .gnd(gnd), .vdd(vdd), .A(_4753_), .B(_4752_), .Y(_16__11_) );
AOI21X1 AOI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf81), .C(data_113__12_), .Y(_4754_) );
AOI21X1 AOI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_4729_), .C(_4754_), .Y(_16__12_) );
INVX1 INVX1_2134 ( .gnd(gnd), .vdd(vdd), .A(data_113__13_), .Y(_4755_) );
NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_4755_), .B(_4727_), .Y(_4756_) );
NAND3X1 NAND3X1_652 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_4726_), .C(_3313__bF_buf80), .Y(_4757_) );
AND2X2 AND2X2_957 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_4757_), .Y(_16__13_) );
AOI21X1 AOI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf79), .C(data_113__14_), .Y(_4758_) );
AOI21X1 AOI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_4729_), .C(_4758_), .Y(_16__14_) );
AOI21X1 AOI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_3313__bF_buf78), .C(data_113__15_), .Y(_4759_) );
AOI21X1 AOI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_4729_), .C(_4759_), .Y(_16__15_) );
INVX1 INVX1_2135 ( .gnd(gnd), .vdd(vdd), .A(data_112__0_), .Y(_4760_) );
OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_14882__bF_buf1), .C(_4760_), .Y(_4761_) );
NAND3X1 NAND3X1_653 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf0), .B(_14986_), .C(_3370_), .Y(_4762_) );
INVX8 INVX8_29 ( .gnd(gnd), .vdd(vdd), .A(_4762_), .Y(_4763_) );
NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_4763__bF_buf3), .Y(_4764_) );
AND2X2 AND2X2_958 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(_4761_), .Y(_15__0_) );
NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(data_112__1_), .B(_4763__bF_buf2), .Y(_4765_) );
AOI21X1 AOI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_4763__bF_buf1), .C(_4765_), .Y(_15__1_) );
NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(data_112__2_), .B(_4763__bF_buf0), .Y(_4766_) );
NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf3), .B(_4762_), .Y(_4767_) );
NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_4767_), .B(_4766_), .Y(_15__2_) );
INVX1 INVX1_2136 ( .gnd(gnd), .vdd(vdd), .A(data_112__3_), .Y(_4768_) );
OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_14882__bF_buf0), .C(_4768_), .Y(_4769_) );
NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_4763__bF_buf3), .Y(_4770_) );
AND2X2 AND2X2_959 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .B(_4769_), .Y(_15__3_) );
INVX1 INVX1_2137 ( .gnd(gnd), .vdd(vdd), .A(data_112__4_), .Y(_4771_) );
OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_14882__bF_buf15_bF_buf3), .C(_4771_), .Y(_4772_) );
OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf2), .B(_4762_), .C(_4772_), .Y(_4773_) );
INVX1 INVX1_2138 ( .gnd(gnd), .vdd(vdd), .A(_4773_), .Y(_15__4_) );
INVX1 INVX1_2139 ( .gnd(gnd), .vdd(vdd), .A(data_112__5_), .Y(_4774_) );
OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_14882__bF_buf14_bF_buf3), .C(_4774_), .Y(_4775_) );
NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_4763__bF_buf2), .Y(_4776_) );
AND2X2 AND2X2_960 ( .gnd(gnd), .vdd(vdd), .A(_4776_), .B(_4775_), .Y(_15__5_) );
INVX1 INVX1_2140 ( .gnd(gnd), .vdd(vdd), .A(data_112__6_), .Y(_4777_) );
OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_14882__bF_buf13_bF_buf3), .C(_4777_), .Y(_4778_) );
NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_4763__bF_buf1), .Y(_4779_) );
AND2X2 AND2X2_961 ( .gnd(gnd), .vdd(vdd), .A(_4779_), .B(_4778_), .Y(_15__6_) );
MUX2X1 MUX2X1_720 ( .gnd(gnd), .vdd(vdd), .A(data_112__7_), .B(IDATA_PROG_data_7_bF_buf5), .S(_4762_), .Y(_4780_) );
INVX1 INVX1_2141 ( .gnd(gnd), .vdd(vdd), .A(_4780_), .Y(_15__7_) );
NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(data_112__8_), .B(_4763__bF_buf0), .Y(_4781_) );
AOI21X1 AOI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_4763__bF_buf3), .C(_4781_), .Y(_15__8_) );
NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_4763__bF_buf2), .Y(_4782_) );
OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(data_112__9_), .B(_4763__bF_buf1), .C(_4782_), .Y(_4783_) );
INVX1 INVX1_2142 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .Y(_15__9_) );
NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(data_112__10_), .B(_4763__bF_buf0), .Y(_4784_) );
NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf0), .B(_4762_), .Y(_4785_) );
NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(_4784_), .Y(_15__10_) );
INVX1 INVX1_2143 ( .gnd(gnd), .vdd(vdd), .A(data_112__11_), .Y(_4786_) );
OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_14882__bF_buf12), .C(_4786_), .Y(_4787_) );
OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf0), .B(_4762_), .C(_4787_), .Y(_4788_) );
INVX1 INVX1_2144 ( .gnd(gnd), .vdd(vdd), .A(_4788_), .Y(_15__11_) );
NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_4763__bF_buf3), .Y(_4789_) );
OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(data_112__12_), .B(_4763__bF_buf2), .C(_4789_), .Y(_4790_) );
INVX1 INVX1_2145 ( .gnd(gnd), .vdd(vdd), .A(_4790_), .Y(_15__12_) );
NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(data_112__13_), .B(_4763__bF_buf1), .Y(_4791_) );
NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf2), .B(_4762_), .Y(_4792_) );
NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_4791_), .Y(_15__13_) );
NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_4763__bF_buf0), .Y(_4793_) );
OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(data_112__14_), .B(_4763__bF_buf3), .C(_4793_), .Y(_4794_) );
INVX1 INVX1_2146 ( .gnd(gnd), .vdd(vdd), .A(_4794_), .Y(_15__14_) );
NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(data_112__15_), .B(_4763__bF_buf2), .Y(_4795_) );
NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf5), .B(_4762_), .Y(_4796_) );
NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_4796_), .B(_4795_), .Y(_15__15_) );
NAND3X1 NAND3X1_654 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .B(_14888__bF_buf1), .C(_3354__bF_buf0), .Y(_4797_) );
INVX1 INVX1_2147 ( .gnd(gnd), .vdd(vdd), .A(data_111__0_), .Y(_4798_) );
OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf11), .C(_4798_), .Y(_4799_) );
OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf0), .B(_4797_), .C(_4799_), .Y(_4800_) );
INVX1 INVX1_2148 ( .gnd(gnd), .vdd(vdd), .A(_4800_), .Y(_14__0_) );
INVX1 INVX1_2149 ( .gnd(gnd), .vdd(vdd), .A(data_111__1_), .Y(_4801_) );
MUX2X1 MUX2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(_14894__bF_buf6), .S(_4797_), .Y(_14__1_) );
INVX1 INVX1_2150 ( .gnd(gnd), .vdd(vdd), .A(data_111__2_), .Y(_4802_) );
MUX2X1 MUX2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_4802_), .B(_14897__bF_buf2), .S(_4797_), .Y(_14__2_) );
INVX1 INVX1_2151 ( .gnd(gnd), .vdd(vdd), .A(data_111__3_), .Y(_4803_) );
OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf10), .C(_4803_), .Y(_4804_) );
OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(IDATA_PROG_data_3_bF_buf3), .C(_4804_), .Y(_4805_) );
INVX1 INVX1_2152 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .Y(_14__3_) );
INVX1 INVX1_2153 ( .gnd(gnd), .vdd(vdd), .A(data_111__4_), .Y(_4806_) );
OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf9), .C(_4806_), .Y(_4807_) );
OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf1), .B(_4797_), .C(_4807_), .Y(_4808_) );
INVX1 INVX1_2154 ( .gnd(gnd), .vdd(vdd), .A(_4808_), .Y(_14__4_) );
INVX1 INVX1_2155 ( .gnd(gnd), .vdd(vdd), .A(data_111__5_), .Y(_4809_) );
MUX2X1 MUX2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(_14903__bF_buf12), .S(_4797_), .Y(_14__5_) );
INVX1 INVX1_2156 ( .gnd(gnd), .vdd(vdd), .A(data_111__6_), .Y(_4810_) );
OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf8), .C(_4810_), .Y(_4811_) );
OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf4), .B(_4797_), .C(_4811_), .Y(_4812_) );
INVX1 INVX1_2157 ( .gnd(gnd), .vdd(vdd), .A(_4812_), .Y(_14__6_) );
MUX2X1 MUX2X1_724 ( .gnd(gnd), .vdd(vdd), .A(data_111__7_), .B(IDATA_PROG_data_7_bF_buf4), .S(_4797_), .Y(_4813_) );
INVX1 INVX1_2158 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .Y(_14__7_) );
INVX1 INVX1_2159 ( .gnd(gnd), .vdd(vdd), .A(data_111__8_), .Y(_4814_) );
OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf7), .C(_4814_), .Y(_4815_) );
OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(IDATA_PROG_data_8_bF_buf2), .C(_4815_), .Y(_4816_) );
INVX1 INVX1_2160 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .Y(_14__8_) );
INVX1 INVX1_2161 ( .gnd(gnd), .vdd(vdd), .A(data_111__9_), .Y(_4817_) );
OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf6), .C(_4817_), .Y(_4818_) );
OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf0), .B(_4797_), .C(_4818_), .Y(_4819_) );
INVX1 INVX1_2162 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .Y(_14__9_) );
INVX1 INVX1_2163 ( .gnd(gnd), .vdd(vdd), .A(data_111__10_), .Y(_4820_) );
OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf5), .C(_4820_), .Y(_4821_) );
OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(IDATA_PROG_data_10_bF_buf4), .C(_4821_), .Y(_4822_) );
INVX1 INVX1_2164 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .Y(_14__10_) );
INVX1 INVX1_2165 ( .gnd(gnd), .vdd(vdd), .A(data_111__11_), .Y(_4823_) );
OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf4), .C(_4823_), .Y(_4824_) );
OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(IDATA_PROG_data_11_bF_buf4), .C(_4824_), .Y(_4825_) );
INVX1 INVX1_2166 ( .gnd(gnd), .vdd(vdd), .A(_4825_), .Y(_14__11_) );
INVX1 INVX1_2167 ( .gnd(gnd), .vdd(vdd), .A(data_111__12_), .Y(_4826_) );
OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf3), .C(_4826_), .Y(_4827_) );
OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(IDATA_PROG_data_12_bF_buf0), .C(_4827_), .Y(_4828_) );
INVX1 INVX1_2168 ( .gnd(gnd), .vdd(vdd), .A(_4828_), .Y(_14__12_) );
INVX1 INVX1_2169 ( .gnd(gnd), .vdd(vdd), .A(data_111__13_), .Y(_4829_) );
OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf2), .C(_4829_), .Y(_4830_) );
OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf1), .B(_4797_), .C(_4830_), .Y(_4831_) );
INVX1 INVX1_2170 ( .gnd(gnd), .vdd(vdd), .A(_4831_), .Y(_14__13_) );
INVX1 INVX1_2171 ( .gnd(gnd), .vdd(vdd), .A(data_111__14_), .Y(_4832_) );
MUX2X1 MUX2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_15060__bF_buf7), .S(_4797_), .Y(_14__14_) );
INVX1 INVX1_2172 ( .gnd(gnd), .vdd(vdd), .A(data_111__15_), .Y(_4833_) );
OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_14882__bF_buf1), .C(_4833_), .Y(_4834_) );
OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(IDATA_PROG_data_15_bF_buf4), .C(_4834_), .Y(_4835_) );
INVX1 INVX1_2173 ( .gnd(gnd), .vdd(vdd), .A(_4835_), .Y(_14__15_) );
INVX1 INVX1_2174 ( .gnd(gnd), .vdd(vdd), .A(data_110__0_), .Y(_4836_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(_3361_), .Y(_4837_) );
OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3362_), .C(_4837_), .Y(_4838_) );
AOI21X1 AOI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_3354__bF_buf3), .B(_14991_), .C(_4387_), .Y(_4839_) );
OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3635_), .C(_4839_), .Y(_4840_) );
NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(_4838_), .Y(_4841_) );
NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_4841_), .B(_4243_), .Y(_4842_) );
OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_4842_), .C(_4836_), .Y(_4843_) );
AND2X2 AND2X2_962 ( .gnd(gnd), .vdd(vdd), .A(_4243_), .B(_4841_), .Y(_4844_) );
NAND3X1 NAND3X1_655 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_4844_), .C(_3313__bF_buf77), .Y(_4845_) );
AND2X2 AND2X2_963 ( .gnd(gnd), .vdd(vdd), .A(_4843_), .B(_4845_), .Y(_13__0_) );
INVX1 INVX1_2175 ( .gnd(gnd), .vdd(vdd), .A(data_110__1_), .Y(_4846_) );
OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_4842_), .C(_4846_), .Y(_4847_) );
NAND3X1 NAND3X1_656 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_4844_), .C(_3313__bF_buf76), .Y(_4848_) );
AND2X2 AND2X2_964 ( .gnd(gnd), .vdd(vdd), .A(_4847_), .B(_4848_), .Y(_13__1_) );
INVX1 INVX1_2176 ( .gnd(gnd), .vdd(vdd), .A(data_110__2_), .Y(_4849_) );
NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_4844_), .B(_3313__bF_buf75), .Y(_4850_) );
MUX2X1 MUX2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_4849_), .B(_14897__bF_buf1), .S(_4850_), .Y(_13__2_) );
INVX1 INVX1_2177 ( .gnd(gnd), .vdd(vdd), .A(data_110__3_), .Y(_4851_) );
OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_4842_), .C(_4851_), .Y(_4852_) );
NAND3X1 NAND3X1_657 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_4844_), .C(_3313__bF_buf74), .Y(_4853_) );
AND2X2 AND2X2_965 ( .gnd(gnd), .vdd(vdd), .A(_4852_), .B(_4853_), .Y(_13__3_) );
INVX1 INVX1_2178 ( .gnd(gnd), .vdd(vdd), .A(data_110__4_), .Y(_4854_) );
OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf24), .B(_4842_), .C(_4854_), .Y(_4855_) );
NAND3X1 NAND3X1_658 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_4844_), .C(_3313__bF_buf73), .Y(_4856_) );
AND2X2 AND2X2_966 ( .gnd(gnd), .vdd(vdd), .A(_4855_), .B(_4856_), .Y(_13__4_) );
INVX1 INVX1_2179 ( .gnd(gnd), .vdd(vdd), .A(data_110__5_), .Y(_4857_) );
OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_4842_), .C(_4857_), .Y(_4858_) );
NAND3X1 NAND3X1_659 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_4844_), .C(_3313__bF_buf72), .Y(_4859_) );
AND2X2 AND2X2_967 ( .gnd(gnd), .vdd(vdd), .A(_4858_), .B(_4859_), .Y(_13__5_) );
INVX1 INVX1_2180 ( .gnd(gnd), .vdd(vdd), .A(data_110__6_), .Y(_4860_) );
MUX2X1 MUX2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_4860_), .B(_15049__bF_buf4), .S(_4850_), .Y(_13__6_) );
INVX1 INVX1_2181 ( .gnd(gnd), .vdd(vdd), .A(data_110__7_), .Y(_4861_) );
OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_4842_), .C(_4861_), .Y(_4862_) );
NAND3X1 NAND3X1_660 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_4844_), .C(_3313__bF_buf71), .Y(_4863_) );
AND2X2 AND2X2_968 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(_4863_), .Y(_13__7_) );
INVX1 INVX1_2182 ( .gnd(gnd), .vdd(vdd), .A(data_110__8_), .Y(_4864_) );
MUX2X1 MUX2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .B(_15052__bF_buf11), .S(_4850_), .Y(_13__8_) );
INVX1 INVX1_2183 ( .gnd(gnd), .vdd(vdd), .A(data_110__9_), .Y(_4865_) );
MUX2X1 MUX2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_4865_), .B(_14913__bF_buf3), .S(_4850_), .Y(_13__9_) );
INVX1 INVX1_2184 ( .gnd(gnd), .vdd(vdd), .A(data_110__10_), .Y(_4866_) );
MUX2X1 MUX2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_4866_), .B(_15055__bF_buf0), .S(_4850_), .Y(_13__10_) );
INVX1 INVX1_2185 ( .gnd(gnd), .vdd(vdd), .A(data_110__11_), .Y(_4867_) );
OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_4842_), .C(_4867_), .Y(_4868_) );
NAND3X1 NAND3X1_661 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_4844_), .C(_3313__bF_buf70), .Y(_4869_) );
AND2X2 AND2X2_969 ( .gnd(gnd), .vdd(vdd), .A(_4868_), .B(_4869_), .Y(_13__11_) );
INVX1 INVX1_2186 ( .gnd(gnd), .vdd(vdd), .A(data_110__12_), .Y(_4870_) );
OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf20), .B(_4842_), .C(_4870_), .Y(_4871_) );
NAND3X1 NAND3X1_662 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_4844_), .C(_3313__bF_buf69), .Y(_4872_) );
AND2X2 AND2X2_970 ( .gnd(gnd), .vdd(vdd), .A(_4871_), .B(_4872_), .Y(_13__12_) );
INVX1 INVX1_2187 ( .gnd(gnd), .vdd(vdd), .A(data_110__13_), .Y(_4873_) );
MUX2X1 MUX2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_4873_), .B(_14924__bF_buf12), .S(_4850_), .Y(_13__13_) );
INVX1 INVX1_2188 ( .gnd(gnd), .vdd(vdd), .A(data_110__14_), .Y(_4874_) );
MUX2X1 MUX2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_4874_), .B(_15060__bF_buf6), .S(_4850_), .Y(_13__14_) );
INVX1 INVX1_2189 ( .gnd(gnd), .vdd(vdd), .A(data_110__15_), .Y(_4875_) );
MUX2X1 MUX2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(_15062__bF_buf13), .S(_4850_), .Y(_13__15_) );
INVX1 INVX1_2190 ( .gnd(gnd), .vdd(vdd), .A(data_109__0_), .Y(_4876_) );
OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_14991_), .C(_3354__bF_buf2), .Y(_4877_) );
OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_2313_), .C(_4604_), .Y(_4878_) );
NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .B(_3361_), .Y(_4879_) );
AND2X2 AND2X2_971 ( .gnd(gnd), .vdd(vdd), .A(_4879_), .B(_4877_), .Y(_4880_) );
NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .B(_4243_), .Y(_4881_) );
OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_4881_), .C(_4876_), .Y(_4882_) );
AND2X2 AND2X2_972 ( .gnd(gnd), .vdd(vdd), .A(_4243_), .B(_4880_), .Y(_4883_) );
NAND3X1 NAND3X1_663 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_4883_), .C(_3313__bF_buf68), .Y(_4884_) );
AND2X2 AND2X2_973 ( .gnd(gnd), .vdd(vdd), .A(_4882_), .B(_4884_), .Y(_11__0_) );
INVX1 INVX1_2191 ( .gnd(gnd), .vdd(vdd), .A(data_109__1_), .Y(_4885_) );
OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_4881_), .C(_4885_), .Y(_4886_) );
NAND3X1 NAND3X1_664 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_4883_), .C(_3313__bF_buf67), .Y(_4887_) );
AND2X2 AND2X2_974 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .B(_4887_), .Y(_11__1_) );
INVX1 INVX1_2192 ( .gnd(gnd), .vdd(vdd), .A(data_109__2_), .Y(_4888_) );
NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_4883_), .B(_3313__bF_buf66), .Y(_4889_) );
MUX2X1 MUX2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_14897__bF_buf0), .S(_4889_), .Y(_11__2_) );
INVX1 INVX1_2193 ( .gnd(gnd), .vdd(vdd), .A(data_109__3_), .Y(_4890_) );
OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf17), .B(_4881_), .C(_4890_), .Y(_4891_) );
NAND3X1 NAND3X1_665 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_4883_), .C(_3313__bF_buf65), .Y(_4892_) );
AND2X2 AND2X2_975 ( .gnd(gnd), .vdd(vdd), .A(_4891_), .B(_4892_), .Y(_11__3_) );
INVX1 INVX1_2194 ( .gnd(gnd), .vdd(vdd), .A(data_109__4_), .Y(_4893_) );
OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf16), .B(_4881_), .C(_4893_), .Y(_4894_) );
NAND3X1 NAND3X1_666 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_4883_), .C(_3313__bF_buf64), .Y(_4895_) );
AND2X2 AND2X2_976 ( .gnd(gnd), .vdd(vdd), .A(_4894_), .B(_4895_), .Y(_11__4_) );
INVX1 INVX1_2195 ( .gnd(gnd), .vdd(vdd), .A(data_109__5_), .Y(_4896_) );
OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf15), .B(_4881_), .C(_4896_), .Y(_4897_) );
NAND3X1 NAND3X1_667 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_4883_), .C(_3313__bF_buf63), .Y(_4898_) );
AND2X2 AND2X2_977 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .B(_4898_), .Y(_11__5_) );
INVX1 INVX1_2196 ( .gnd(gnd), .vdd(vdd), .A(data_109__6_), .Y(_4899_) );
MUX2X1 MUX2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .B(_15049__bF_buf3), .S(_4889_), .Y(_11__6_) );
INVX1 INVX1_2197 ( .gnd(gnd), .vdd(vdd), .A(data_109__7_), .Y(_4900_) );
OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf14), .B(_4881_), .C(_4900_), .Y(_4901_) );
NAND3X1 NAND3X1_668 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_4883_), .C(_3313__bF_buf62), .Y(_4902_) );
AND2X2 AND2X2_978 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(_4902_), .Y(_11__7_) );
INVX1 INVX1_2198 ( .gnd(gnd), .vdd(vdd), .A(data_109__8_), .Y(_4903_) );
MUX2X1 MUX2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .B(_15052__bF_buf10), .S(_4889_), .Y(_11__8_) );
INVX1 INVX1_2199 ( .gnd(gnd), .vdd(vdd), .A(data_109__9_), .Y(_4904_) );
MUX2X1 MUX2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_4904_), .B(_14913__bF_buf2), .S(_4889_), .Y(_11__9_) );
INVX1 INVX1_2200 ( .gnd(gnd), .vdd(vdd), .A(data_109__10_), .Y(_4905_) );
MUX2X1 MUX2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_4905_), .B(_15055__bF_buf13), .S(_4889_), .Y(_11__10_) );
INVX1 INVX1_2201 ( .gnd(gnd), .vdd(vdd), .A(data_109__11_), .Y(_4906_) );
OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf13), .B(_4881_), .C(_4906_), .Y(_4907_) );
NAND3X1 NAND3X1_669 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_4883_), .C(_3313__bF_buf61), .Y(_4908_) );
AND2X2 AND2X2_979 ( .gnd(gnd), .vdd(vdd), .A(_4907_), .B(_4908_), .Y(_11__11_) );
INVX1 INVX1_2202 ( .gnd(gnd), .vdd(vdd), .A(data_109__12_), .Y(_4909_) );
OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_4881_), .C(_4909_), .Y(_4910_) );
NAND3X1 NAND3X1_670 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_4883_), .C(_3313__bF_buf60), .Y(_4911_) );
AND2X2 AND2X2_980 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .B(_4911_), .Y(_11__12_) );
INVX1 INVX1_2203 ( .gnd(gnd), .vdd(vdd), .A(data_109__13_), .Y(_4912_) );
MUX2X1 MUX2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_4912_), .B(_14924__bF_buf11), .S(_4889_), .Y(_11__13_) );
INVX1 INVX1_2204 ( .gnd(gnd), .vdd(vdd), .A(data_109__14_), .Y(_4913_) );
MUX2X1 MUX2X1_740 ( .gnd(gnd), .vdd(vdd), .A(_4913_), .B(_15060__bF_buf5), .S(_4889_), .Y(_11__14_) );
INVX1 INVX1_2205 ( .gnd(gnd), .vdd(vdd), .A(data_109__15_), .Y(_4914_) );
MUX2X1 MUX2X1_741 ( .gnd(gnd), .vdd(vdd), .A(_4914_), .B(_15062__bF_buf12), .S(_4889_), .Y(_11__15_) );
INVX1 INVX1_2206 ( .gnd(gnd), .vdd(vdd), .A(data_108__0_), .Y(_4915_) );
INVX1 INVX1_2207 ( .gnd(gnd), .vdd(vdd), .A(_4878_), .Y(_4916_) );
INVX1 INVX1_2208 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .Y(_4917_) );
AOI21X1 AOI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_3354__bF_buf1), .B(_4917_), .C(_3361_), .Y(_4918_) );
NAND3X1 NAND3X1_671 ( .gnd(gnd), .vdd(vdd), .A(_15073_), .B(_4916_), .C(_4918_), .Y(_4919_) );
NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(_3353__bF_buf4), .Y(_4920_) );
NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_4920_), .B(_3313__bF_buf59), .Y(_4921_) );
MUX2X1 MUX2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_4915_), .B(_14932__bF_buf6), .S(_4921_), .Y(_10__0_) );
INVX1 INVX1_2209 ( .gnd(gnd), .vdd(vdd), .A(data_108__1_), .Y(_4922_) );
MUX2X1 MUX2X1_743 ( .gnd(gnd), .vdd(vdd), .A(_4922_), .B(_14894__bF_buf3), .S(_4921_), .Y(_10__1_) );
INVX1 INVX1_2210 ( .gnd(gnd), .vdd(vdd), .A(data_108__2_), .Y(_4923_) );
NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_4923_), .B(_4921_), .Y(_4924_) );
AND2X2 AND2X2_981 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf58), .B(_4920_), .Y(_4925_) );
NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_4925_), .Y(_4926_) );
AND2X2 AND2X2_982 ( .gnd(gnd), .vdd(vdd), .A(_4926_), .B(_4924_), .Y(_10__2_) );
INVX1 INVX1_2211 ( .gnd(gnd), .vdd(vdd), .A(data_108__3_), .Y(_4927_) );
MUX2X1 MUX2X1_744 ( .gnd(gnd), .vdd(vdd), .A(_4927_), .B(_14899__bF_buf3), .S(_4921_), .Y(_10__3_) );
INVX1 INVX1_2212 ( .gnd(gnd), .vdd(vdd), .A(data_108__4_), .Y(_4928_) );
MUX2X1 MUX2X1_745 ( .gnd(gnd), .vdd(vdd), .A(_4928_), .B(_14902__bF_buf10), .S(_4921_), .Y(_10__4_) );
INVX1 INVX1_2213 ( .gnd(gnd), .vdd(vdd), .A(data_108__5_), .Y(_4929_) );
MUX2X1 MUX2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_4929_), .B(_14903__bF_buf9), .S(_4921_), .Y(_10__5_) );
INVX1 INVX1_2214 ( .gnd(gnd), .vdd(vdd), .A(data_108__6_), .Y(_4930_) );
NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_4930_), .B(_4921_), .Y(_4931_) );
NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_4925_), .Y(_4932_) );
AND2X2 AND2X2_983 ( .gnd(gnd), .vdd(vdd), .A(_4932_), .B(_4931_), .Y(_10__6_) );
INVX1 INVX1_2215 ( .gnd(gnd), .vdd(vdd), .A(data_108__7_), .Y(_4933_) );
MUX2X1 MUX2X1_747 ( .gnd(gnd), .vdd(vdd), .A(_4933_), .B(_14908__bF_buf11), .S(_4921_), .Y(_10__7_) );
AOI21X1 AOI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_4920_), .B(_3313__bF_buf57), .C(data_108__8_), .Y(_4934_) );
AOI21X1 AOI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_4925_), .C(_4934_), .Y(_10__8_) );
INVX1 INVX1_2216 ( .gnd(gnd), .vdd(vdd), .A(data_108__9_), .Y(_4935_) );
MUX2X1 MUX2X1_748 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_14913__bF_buf1), .S(_4921_), .Y(_10__9_) );
INVX1 INVX1_2217 ( .gnd(gnd), .vdd(vdd), .A(data_108__10_), .Y(_4936_) );
MUX2X1 MUX2X1_749 ( .gnd(gnd), .vdd(vdd), .A(_4936_), .B(_15055__bF_buf12), .S(_4921_), .Y(_10__10_) );
INVX1 INVX1_2218 ( .gnd(gnd), .vdd(vdd), .A(data_108__11_), .Y(_4937_) );
MUX2X1 MUX2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_4937_), .B(_14918__bF_buf12), .S(_4921_), .Y(_10__11_) );
INVX1 INVX1_2219 ( .gnd(gnd), .vdd(vdd), .A(data_108__12_), .Y(_4938_) );
MUX2X1 MUX2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(_14920__bF_buf11), .S(_4921_), .Y(_10__12_) );
INVX1 INVX1_2220 ( .gnd(gnd), .vdd(vdd), .A(data_108__13_), .Y(_4939_) );
MUX2X1 MUX2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_4939_), .B(_14924__bF_buf10), .S(_4921_), .Y(_10__13_) );
INVX1 INVX1_2221 ( .gnd(gnd), .vdd(vdd), .A(data_108__14_), .Y(_4940_) );
NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_4940_), .B(_4921_), .Y(_4941_) );
NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_4925_), .Y(_4942_) );
AND2X2 AND2X2_984 ( .gnd(gnd), .vdd(vdd), .A(_4942_), .B(_4941_), .Y(_10__14_) );
INVX1 INVX1_2222 ( .gnd(gnd), .vdd(vdd), .A(data_108__15_), .Y(_4943_) );
NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4921_), .Y(_4944_) );
NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_4925_), .Y(_4945_) );
AND2X2 AND2X2_985 ( .gnd(gnd), .vdd(vdd), .A(_4945_), .B(_4944_), .Y(_10__15_) );
INVX1 INVX1_2223 ( .gnd(gnd), .vdd(vdd), .A(data_107__0_), .Y(_4946_) );
INVX1 INVX1_2224 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .Y(_4947_) );
AOI21X1 AOI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf0), .B(_3354__bF_buf0), .C(_4387_), .Y(_4948_) );
NAND3X1 NAND3X1_672 ( .gnd(gnd), .vdd(vdd), .A(_4947_), .B(_4948_), .C(_4243_), .Y(_4949_) );
OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_4949_), .C(_4946_), .Y(_4950_) );
INVX1 INVX1_2225 ( .gnd(gnd), .vdd(vdd), .A(_4948_), .Y(_4951_) );
NOR3X1 NOR3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .B(_4951_), .C(_4287_), .Y(_4952_) );
NAND3X1 NAND3X1_673 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_3313__bF_buf56), .C(_4952_), .Y(_4953_) );
AND2X2 AND2X2_986 ( .gnd(gnd), .vdd(vdd), .A(_4950_), .B(_4953_), .Y(_9__0_) );
INVX1 INVX1_2226 ( .gnd(gnd), .vdd(vdd), .A(data_107__1_), .Y(_4954_) );
OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_4949_), .C(_4954_), .Y(_4955_) );
NAND3X1 NAND3X1_674 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_3313__bF_buf55), .C(_4952_), .Y(_4956_) );
AND2X2 AND2X2_987 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4956_), .Y(_9__1_) );
INVX1 INVX1_2227 ( .gnd(gnd), .vdd(vdd), .A(data_107__2_), .Y(_4957_) );
NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf54), .B(_4952_), .Y(_4958_) );
MUX2X1 MUX2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_4957_), .B(_14897__bF_buf13), .S(_4958_), .Y(_9__2_) );
INVX1 INVX1_2228 ( .gnd(gnd), .vdd(vdd), .A(data_107__3_), .Y(_4959_) );
OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_4949_), .C(_4959_), .Y(_4960_) );
NAND3X1 NAND3X1_675 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_3313__bF_buf53), .C(_4952_), .Y(_4961_) );
AND2X2 AND2X2_988 ( .gnd(gnd), .vdd(vdd), .A(_4960_), .B(_4961_), .Y(_9__3_) );
INVX1 INVX1_2229 ( .gnd(gnd), .vdd(vdd), .A(data_107__4_), .Y(_4962_) );
OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf8), .B(_4949_), .C(_4962_), .Y(_4963_) );
NAND3X1 NAND3X1_676 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_3313__bF_buf52), .C(_4952_), .Y(_4964_) );
AND2X2 AND2X2_989 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4964_), .Y(_9__4_) );
INVX1 INVX1_2230 ( .gnd(gnd), .vdd(vdd), .A(data_107__5_), .Y(_4965_) );
OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_4949_), .C(_4965_), .Y(_4966_) );
NAND3X1 NAND3X1_677 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_3313__bF_buf51), .C(_4952_), .Y(_4967_) );
AND2X2 AND2X2_990 ( .gnd(gnd), .vdd(vdd), .A(_4966_), .B(_4967_), .Y(_9__5_) );
INVX1 INVX1_2231 ( .gnd(gnd), .vdd(vdd), .A(data_107__6_), .Y(_4968_) );
MUX2X1 MUX2X1_754 ( .gnd(gnd), .vdd(vdd), .A(_4968_), .B(_15049__bF_buf1), .S(_4958_), .Y(_9__6_) );
INVX1 INVX1_2232 ( .gnd(gnd), .vdd(vdd), .A(data_107__7_), .Y(_4969_) );
OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_4949_), .C(_4969_), .Y(_4970_) );
NAND3X1 NAND3X1_678 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_3313__bF_buf50), .C(_4952_), .Y(_4971_) );
AND2X2 AND2X2_991 ( .gnd(gnd), .vdd(vdd), .A(_4970_), .B(_4971_), .Y(_9__7_) );
INVX1 INVX1_2233 ( .gnd(gnd), .vdd(vdd), .A(data_107__8_), .Y(_4972_) );
MUX2X1 MUX2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_4972_), .B(_15052__bF_buf8), .S(_4958_), .Y(_9__8_) );
INVX1 INVX1_2234 ( .gnd(gnd), .vdd(vdd), .A(data_107__9_), .Y(_4973_) );
MUX2X1 MUX2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_4973_), .B(_14913__bF_buf0), .S(_4958_), .Y(_9__9_) );
INVX1 INVX1_2235 ( .gnd(gnd), .vdd(vdd), .A(data_107__10_), .Y(_4974_) );
MUX2X1 MUX2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_4974_), .B(_15055__bF_buf11), .S(_4958_), .Y(_9__10_) );
INVX1 INVX1_2236 ( .gnd(gnd), .vdd(vdd), .A(data_107__11_), .Y(_4975_) );
OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_4949_), .C(_4975_), .Y(_4976_) );
NAND3X1 NAND3X1_679 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_3313__bF_buf49), .C(_4952_), .Y(_4977_) );
AND2X2 AND2X2_992 ( .gnd(gnd), .vdd(vdd), .A(_4976_), .B(_4977_), .Y(_9__11_) );
INVX1 INVX1_2237 ( .gnd(gnd), .vdd(vdd), .A(data_107__12_), .Y(_4978_) );
OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_4949_), .C(_4978_), .Y(_4979_) );
NAND3X1 NAND3X1_680 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_3313__bF_buf48), .C(_4952_), .Y(_4980_) );
AND2X2 AND2X2_993 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(_4980_), .Y(_9__12_) );
INVX1 INVX1_2238 ( .gnd(gnd), .vdd(vdd), .A(data_107__13_), .Y(_4981_) );
MUX2X1 MUX2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_4981_), .B(_14924__bF_buf9), .S(_4958_), .Y(_9__13_) );
INVX1 INVX1_2239 ( .gnd(gnd), .vdd(vdd), .A(data_107__14_), .Y(_4982_) );
MUX2X1 MUX2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_4982_), .B(_15060__bF_buf3), .S(_4958_), .Y(_9__14_) );
INVX1 INVX1_2240 ( .gnd(gnd), .vdd(vdd), .A(data_107__15_), .Y(_4983_) );
MUX2X1 MUX2X1_760 ( .gnd(gnd), .vdd(vdd), .A(_4983_), .B(_15062__bF_buf10), .S(_4958_), .Y(_9__15_) );
INVX1 INVX1_2241 ( .gnd(gnd), .vdd(vdd), .A(data_106__0_), .Y(_4984_) );
OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_14996_), .C(_3354__bF_buf3), .Y(_4985_) );
NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_4985_), .B(_4837_), .Y(_4986_) );
INVX1 INVX1_2242 ( .gnd(gnd), .vdd(vdd), .A(_4986_), .Y(_4987_) );
NAND3X1 NAND3X1_681 ( .gnd(gnd), .vdd(vdd), .A(_4948_), .B(_4987_), .C(_4243_), .Y(_4988_) );
OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf3), .B(_4988_), .C(_4984_), .Y(_4989_) );
NOR3X1 NOR3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_4951_), .B(_4986_), .C(_4287_), .Y(_4990_) );
NAND3X1 NAND3X1_682 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_3313__bF_buf47), .C(_4990_), .Y(_4991_) );
AND2X2 AND2X2_994 ( .gnd(gnd), .vdd(vdd), .A(_4989_), .B(_4991_), .Y(_8__0_) );
INVX1 INVX1_2243 ( .gnd(gnd), .vdd(vdd), .A(data_106__1_), .Y(_4992_) );
OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_4988_), .C(_4992_), .Y(_4993_) );
NAND3X1 NAND3X1_683 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_3313__bF_buf46), .C(_4990_), .Y(_4994_) );
AND2X2 AND2X2_995 ( .gnd(gnd), .vdd(vdd), .A(_4993_), .B(_4994_), .Y(_8__1_) );
INVX1 INVX1_2244 ( .gnd(gnd), .vdd(vdd), .A(data_106__2_), .Y(_4995_) );
NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf45), .B(_4990_), .Y(_4996_) );
MUX2X1 MUX2X1_761 ( .gnd(gnd), .vdd(vdd), .A(_4995_), .B(_14897__bF_buf12), .S(_4996_), .Y(_8__2_) );
INVX1 INVX1_2245 ( .gnd(gnd), .vdd(vdd), .A(data_106__3_), .Y(_4997_) );
OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_4988_), .C(_4997_), .Y(_4998_) );
NAND3X1 NAND3X1_684 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_3313__bF_buf44), .C(_4990_), .Y(_4999_) );
AND2X2 AND2X2_996 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(_4999_), .Y(_8__3_) );
INVX1 INVX1_2246 ( .gnd(gnd), .vdd(vdd), .A(data_106__4_), .Y(_5000_) );
OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_4988_), .C(_5000_), .Y(_5001_) );
NAND3X1 NAND3X1_685 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_3313__bF_buf43), .C(_4990_), .Y(_5002_) );
AND2X2 AND2X2_997 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_5002_), .Y(_8__4_) );
INVX1 INVX1_2247 ( .gnd(gnd), .vdd(vdd), .A(data_106__5_), .Y(_5003_) );
OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_4988_), .C(_5003_), .Y(_5004_) );
NAND3X1 NAND3X1_686 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_3313__bF_buf42), .C(_4990_), .Y(_5005_) );
AND2X2 AND2X2_998 ( .gnd(gnd), .vdd(vdd), .A(_5004_), .B(_5005_), .Y(_8__5_) );
INVX1 INVX1_2248 ( .gnd(gnd), .vdd(vdd), .A(data_106__6_), .Y(_5006_) );
MUX2X1 MUX2X1_762 ( .gnd(gnd), .vdd(vdd), .A(_5006_), .B(_15049__bF_buf0), .S(_4996_), .Y(_8__6_) );
INVX1 INVX1_2249 ( .gnd(gnd), .vdd(vdd), .A(data_106__7_), .Y(_5007_) );
OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_4988_), .C(_5007_), .Y(_5008_) );
NAND3X1 NAND3X1_687 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_3313__bF_buf41), .C(_4990_), .Y(_5009_) );
AND2X2 AND2X2_999 ( .gnd(gnd), .vdd(vdd), .A(_5008_), .B(_5009_), .Y(_8__7_) );
INVX1 INVX1_2250 ( .gnd(gnd), .vdd(vdd), .A(data_106__8_), .Y(_5010_) );
MUX2X1 MUX2X1_763 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(_15052__bF_buf7), .S(_4996_), .Y(_8__8_) );
INVX1 INVX1_2251 ( .gnd(gnd), .vdd(vdd), .A(data_106__9_), .Y(_5011_) );
MUX2X1 MUX2X1_764 ( .gnd(gnd), .vdd(vdd), .A(_5011_), .B(_14913__bF_buf14), .S(_4996_), .Y(_8__9_) );
INVX1 INVX1_2252 ( .gnd(gnd), .vdd(vdd), .A(data_106__10_), .Y(_5012_) );
MUX2X1 MUX2X1_765 ( .gnd(gnd), .vdd(vdd), .A(_5012_), .B(_15055__bF_buf10), .S(_4996_), .Y(_8__10_) );
INVX1 INVX1_2253 ( .gnd(gnd), .vdd(vdd), .A(data_106__11_), .Y(_5013_) );
OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_4988_), .C(_5013_), .Y(_5014_) );
NAND3X1 NAND3X1_688 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_3313__bF_buf40), .C(_4990_), .Y(_5015_) );
AND2X2 AND2X2_1000 ( .gnd(gnd), .vdd(vdd), .A(_5014_), .B(_5015_), .Y(_8__11_) );
INVX1 INVX1_2254 ( .gnd(gnd), .vdd(vdd), .A(data_106__12_), .Y(_5016_) );
OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_4988_), .C(_5016_), .Y(_5017_) );
NAND3X1 NAND3X1_689 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_3313__bF_buf39), .C(_4990_), .Y(_5018_) );
AND2X2 AND2X2_1001 ( .gnd(gnd), .vdd(vdd), .A(_5017_), .B(_5018_), .Y(_8__12_) );
INVX1 INVX1_2255 ( .gnd(gnd), .vdd(vdd), .A(data_106__13_), .Y(_5019_) );
MUX2X1 MUX2X1_766 ( .gnd(gnd), .vdd(vdd), .A(_5019_), .B(_14924__bF_buf8), .S(_4996_), .Y(_8__13_) );
INVX1 INVX1_2256 ( .gnd(gnd), .vdd(vdd), .A(data_106__14_), .Y(_5020_) );
MUX2X1 MUX2X1_767 ( .gnd(gnd), .vdd(vdd), .A(_5020_), .B(_15060__bF_buf2), .S(_4996_), .Y(_8__14_) );
INVX1 INVX1_2257 ( .gnd(gnd), .vdd(vdd), .A(data_106__15_), .Y(_5021_) );
MUX2X1 MUX2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_5021_), .B(_15062__bF_buf9), .S(_4996_), .Y(_8__15_) );
INVX1 INVX1_2258 ( .gnd(gnd), .vdd(vdd), .A(data_105__0_), .Y(_5022_) );
OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3827_), .C(_4948_), .Y(_5023_) );
AOI21X1 AOI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_3354__bF_buf2), .C(_5023_), .Y(_5024_) );
NAND3X1 NAND3X1_690 ( .gnd(gnd), .vdd(vdd), .A(_4837_), .B(_5024_), .C(_4243_), .Y(_5025_) );
OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_5025__bF_buf3), .C(_5022_), .Y(_5026_) );
NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_5025__bF_buf2), .B(_3393__bF_buf64), .Y(_5027_) );
NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_5027_), .Y(_5028_) );
AND2X2 AND2X2_1002 ( .gnd(gnd), .vdd(vdd), .A(_5028_), .B(_5026_), .Y(_7__0_) );
INVX1 INVX1_2259 ( .gnd(gnd), .vdd(vdd), .A(data_105__1_), .Y(_5029_) );
OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_5025__bF_buf1), .C(_5029_), .Y(_5030_) );
NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_5027_), .Y(_5031_) );
AND2X2 AND2X2_1003 ( .gnd(gnd), .vdd(vdd), .A(_5031_), .B(_5030_), .Y(_7__1_) );
INVX1 INVX1_2260 ( .gnd(gnd), .vdd(vdd), .A(data_105__2_), .Y(_5032_) );
OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_5025__bF_buf0), .C(_5032_), .Y(_5033_) );
NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_5027_), .Y(_5034_) );
AND2X2 AND2X2_1004 ( .gnd(gnd), .vdd(vdd), .A(_5034_), .B(_5033_), .Y(_7__2_) );
INVX1 INVX1_2261 ( .gnd(gnd), .vdd(vdd), .A(data_105__3_), .Y(_5035_) );
OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_5025__bF_buf3), .C(_5035_), .Y(_5036_) );
NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_5027_), .Y(_5037_) );
AND2X2 AND2X2_1005 ( .gnd(gnd), .vdd(vdd), .A(_5037_), .B(_5036_), .Y(_7__3_) );
INVX1 INVX1_2262 ( .gnd(gnd), .vdd(vdd), .A(data_105__4_), .Y(_5038_) );
OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_5025__bF_buf2), .C(_5038_), .Y(_5039_) );
NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_5027_), .Y(_5040_) );
AND2X2 AND2X2_1006 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .B(_5039_), .Y(_7__4_) );
INVX1 INVX1_2263 ( .gnd(gnd), .vdd(vdd), .A(data_105__5_), .Y(_5041_) );
OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_5025__bF_buf1), .C(_5041_), .Y(_5042_) );
NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_5027_), .Y(_5043_) );
AND2X2 AND2X2_1007 ( .gnd(gnd), .vdd(vdd), .A(_5043_), .B(_5042_), .Y(_7__5_) );
INVX1 INVX1_2264 ( .gnd(gnd), .vdd(vdd), .A(data_105__6_), .Y(_5044_) );
OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_5025__bF_buf0), .C(_5044_), .Y(_5045_) );
NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_5027_), .Y(_5046_) );
AND2X2 AND2X2_1008 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_5045_), .Y(_7__6_) );
INVX1 INVX1_2265 ( .gnd(gnd), .vdd(vdd), .A(data_105__7_), .Y(_5047_) );
OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_5025__bF_buf3), .C(_5047_), .Y(_5048_) );
NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_5027_), .Y(_5049_) );
AND2X2 AND2X2_1009 ( .gnd(gnd), .vdd(vdd), .A(_5049_), .B(_5048_), .Y(_7__7_) );
INVX1 INVX1_2266 ( .gnd(gnd), .vdd(vdd), .A(data_105__8_), .Y(_5050_) );
OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_5025__bF_buf2), .C(_5050_), .Y(_5051_) );
NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_5027_), .Y(_5052_) );
AND2X2 AND2X2_1010 ( .gnd(gnd), .vdd(vdd), .A(_5052_), .B(_5051_), .Y(_7__8_) );
INVX1 INVX1_2267 ( .gnd(gnd), .vdd(vdd), .A(data_105__9_), .Y(_5053_) );
OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_5025__bF_buf1), .C(_5053_), .Y(_5054_) );
NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_5027_), .Y(_5055_) );
AND2X2 AND2X2_1011 ( .gnd(gnd), .vdd(vdd), .A(_5055_), .B(_5054_), .Y(_7__9_) );
INVX1 INVX1_2268 ( .gnd(gnd), .vdd(vdd), .A(data_105__10_), .Y(_5056_) );
OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_5025__bF_buf0), .C(_5056_), .Y(_5057_) );
NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_5027_), .Y(_5058_) );
AND2X2 AND2X2_1012 ( .gnd(gnd), .vdd(vdd), .A(_5058_), .B(_5057_), .Y(_7__10_) );
INVX1 INVX1_2269 ( .gnd(gnd), .vdd(vdd), .A(data_105__11_), .Y(_5059_) );
OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_5025__bF_buf3), .C(_5059_), .Y(_5060_) );
NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_5027_), .Y(_5061_) );
AND2X2 AND2X2_1013 ( .gnd(gnd), .vdd(vdd), .A(_5061_), .B(_5060_), .Y(_7__11_) );
INVX1 INVX1_2270 ( .gnd(gnd), .vdd(vdd), .A(data_105__12_), .Y(_5062_) );
OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_5025__bF_buf2), .C(_5062_), .Y(_5063_) );
NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_5027_), .Y(_5064_) );
AND2X2 AND2X2_1014 ( .gnd(gnd), .vdd(vdd), .A(_5064_), .B(_5063_), .Y(_7__12_) );
INVX1 INVX1_2271 ( .gnd(gnd), .vdd(vdd), .A(data_105__13_), .Y(_5065_) );
OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_5025__bF_buf1), .C(_5065_), .Y(_5066_) );
NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_5027_), .Y(_5067_) );
AND2X2 AND2X2_1015 ( .gnd(gnd), .vdd(vdd), .A(_5067_), .B(_5066_), .Y(_7__13_) );
INVX1 INVX1_2272 ( .gnd(gnd), .vdd(vdd), .A(data_105__14_), .Y(_5068_) );
OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_5025__bF_buf0), .C(_5068_), .Y(_5069_) );
NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_5027_), .Y(_5070_) );
AND2X2 AND2X2_1016 ( .gnd(gnd), .vdd(vdd), .A(_5070_), .B(_5069_), .Y(_7__14_) );
INVX1 INVX1_2273 ( .gnd(gnd), .vdd(vdd), .A(data_105__15_), .Y(_5071_) );
OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_5025__bF_buf3), .C(_5071_), .Y(_5072_) );
NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_5027_), .Y(_5073_) );
AND2X2 AND2X2_1017 ( .gnd(gnd), .vdd(vdd), .A(_5073_), .B(_5072_), .Y(_7__15_) );
AOI21X1 AOI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_3354__bF_buf1), .B(_4467_), .C(_5023_), .Y(_5074_) );
NAND3X1 NAND3X1_691 ( .gnd(gnd), .vdd(vdd), .A(_4837_), .B(_5074_), .C(_4243_), .Y(_5075_) );
NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .B(_3393__bF_buf48), .Y(_5076_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf3), .B(data_104__0_), .Y(_5077_) );
NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_5076__bF_buf2), .Y(_5078_) );
AND2X2 AND2X2_1018 ( .gnd(gnd), .vdd(vdd), .A(_5077_), .B(_5078_), .Y(_6__0_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf1), .B(data_104__1_), .Y(_5079_) );
NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_5076__bF_buf0), .Y(_5080_) );
AND2X2 AND2X2_1019 ( .gnd(gnd), .vdd(vdd), .A(_5079_), .B(_5080_), .Y(_6__1_) );
INVX1 INVX1_2274 ( .gnd(gnd), .vdd(vdd), .A(data_104__2_), .Y(_5081_) );
OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_5075_), .C(_5081_), .Y(_5082_) );
NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_5076__bF_buf3), .Y(_5083_) );
AND2X2 AND2X2_1020 ( .gnd(gnd), .vdd(vdd), .A(_5083_), .B(_5082_), .Y(_6__2_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf2), .B(data_104__3_), .Y(_5084_) );
NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_5076__bF_buf1), .Y(_5085_) );
AND2X2 AND2X2_1021 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .B(_5085_), .Y(_6__3_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf0), .B(data_104__4_), .Y(_5086_) );
NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_5076__bF_buf3), .Y(_5087_) );
AND2X2 AND2X2_1022 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .B(_5087_), .Y(_6__4_) );
INVX1 INVX1_2275 ( .gnd(gnd), .vdd(vdd), .A(data_104__5_), .Y(_5088_) );
OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_5075_), .C(_5088_), .Y(_5089_) );
NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_5076__bF_buf2), .Y(_5090_) );
AND2X2 AND2X2_1023 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_5089_), .Y(_6__5_) );
INVX1 INVX1_2276 ( .gnd(gnd), .vdd(vdd), .A(data_104__6_), .Y(_5091_) );
OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_5075_), .C(_5091_), .Y(_5092_) );
NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_5076__bF_buf1), .Y(_5093_) );
AND2X2 AND2X2_1024 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .B(_5092_), .Y(_6__6_) );
INVX1 INVX1_2277 ( .gnd(gnd), .vdd(vdd), .A(data_104__7_), .Y(_5094_) );
OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_5075_), .C(_5094_), .Y(_5095_) );
NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_5076__bF_buf0), .Y(_5096_) );
AND2X2 AND2X2_1025 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .B(_5095_), .Y(_6__7_) );
INVX1 INVX1_2278 ( .gnd(gnd), .vdd(vdd), .A(data_104__8_), .Y(_5097_) );
OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_5075_), .C(_5097_), .Y(_5098_) );
NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_5076__bF_buf3), .Y(_5099_) );
AND2X2 AND2X2_1026 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .B(_5098_), .Y(_6__8_) );
INVX1 INVX1_2279 ( .gnd(gnd), .vdd(vdd), .A(data_104__9_), .Y(_5100_) );
OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_5075_), .C(_5100_), .Y(_5101_) );
NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_5076__bF_buf2), .Y(_5102_) );
AND2X2 AND2X2_1027 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_5101_), .Y(_6__9_) );
INVX1 INVX1_2280 ( .gnd(gnd), .vdd(vdd), .A(data_104__10_), .Y(_5103_) );
OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_5075_), .C(_5103_), .Y(_5104_) );
NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_5076__bF_buf1), .Y(_5105_) );
AND2X2 AND2X2_1028 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_5104_), .Y(_6__10_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_5076__bF_buf0), .B(data_104__11_), .Y(_5106_) );
NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_5076__bF_buf3), .Y(_5107_) );
AND2X2 AND2X2_1029 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_5107_), .Y(_6__11_) );
INVX1 INVX1_2281 ( .gnd(gnd), .vdd(vdd), .A(data_104__12_), .Y(_5108_) );
OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_5075_), .C(_5108_), .Y(_5109_) );
NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_5076__bF_buf2), .Y(_5110_) );
AND2X2 AND2X2_1030 ( .gnd(gnd), .vdd(vdd), .A(_5110_), .B(_5109_), .Y(_6__12_) );
INVX1 INVX1_2282 ( .gnd(gnd), .vdd(vdd), .A(data_104__13_), .Y(_5111_) );
OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_5075_), .C(_5111_), .Y(_5112_) );
NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_5076__bF_buf1), .Y(_5113_) );
AND2X2 AND2X2_1031 ( .gnd(gnd), .vdd(vdd), .A(_5113_), .B(_5112_), .Y(_6__13_) );
INVX1 INVX1_2283 ( .gnd(gnd), .vdd(vdd), .A(data_104__14_), .Y(_5114_) );
OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_5075_), .C(_5114_), .Y(_5115_) );
NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_5076__bF_buf0), .Y(_5116_) );
AND2X2 AND2X2_1032 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_5115_), .Y(_6__14_) );
INVX1 INVX1_2284 ( .gnd(gnd), .vdd(vdd), .A(data_104__15_), .Y(_5117_) );
OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_5075_), .C(_5117_), .Y(_5118_) );
NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_5076__bF_buf3), .Y(_5119_) );
AND2X2 AND2X2_1033 ( .gnd(gnd), .vdd(vdd), .A(_5119_), .B(_5118_), .Y(_6__15_) );
INVX1 INVX1_2285 ( .gnd(gnd), .vdd(vdd), .A(data_103__0_), .Y(_5120_) );
OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_15171_), .C(_3359_), .Y(_5121_) );
NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_4387_), .B(_5121_), .Y(_5122_) );
NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_3357_), .Y(_5123_) );
INVX1 INVX1_2286 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .Y(_5124_) );
NAND3X1 NAND3X1_692 ( .gnd(gnd), .vdd(vdd), .A(_3360_), .B(_5124_), .C(_5122_), .Y(_5125_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_5125_), .Y(_5126_) );
OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_5126_), .C(_5120_), .Y(_5127_) );
NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_5125_), .B(_4287_), .Y(_5128_) );
NAND3X1 NAND3X1_693 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_5128_), .C(_3313__bF_buf38), .Y(_5129_) );
AND2X2 AND2X2_1034 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .B(_5129_), .Y(_5__0_) );
INVX1 INVX1_2287 ( .gnd(gnd), .vdd(vdd), .A(data_103__1_), .Y(_5130_) );
OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_5126_), .C(_5130_), .Y(_5131_) );
NAND3X1 NAND3X1_694 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_5128_), .C(_3313__bF_buf37), .Y(_5132_) );
AND2X2 AND2X2_1035 ( .gnd(gnd), .vdd(vdd), .A(_5131_), .B(_5132_), .Y(_5__1_) );
INVX1 INVX1_2288 ( .gnd(gnd), .vdd(vdd), .A(data_103__2_), .Y(_5133_) );
NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_5128_), .B(_3313__bF_buf36), .Y(_5134_) );
MUX2X1 MUX2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_5133_), .B(_14897__bF_buf9), .S(_5134_), .Y(_5__2_) );
INVX1 INVX1_2289 ( .gnd(gnd), .vdd(vdd), .A(data_103__3_), .Y(_5135_) );
OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf34), .B(_5126_), .C(_5135_), .Y(_5136_) );
NAND3X1 NAND3X1_695 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_5128_), .C(_3313__bF_buf35), .Y(_5137_) );
AND2X2 AND2X2_1036 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_5137_), .Y(_5__3_) );
INVX1 INVX1_2290 ( .gnd(gnd), .vdd(vdd), .A(data_103__4_), .Y(_5138_) );
OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_5126_), .C(_5138_), .Y(_5139_) );
NAND3X1 NAND3X1_696 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_5128_), .C(_3313__bF_buf34), .Y(_5140_) );
AND2X2 AND2X2_1037 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .B(_5140_), .Y(_5__4_) );
INVX1 INVX1_2291 ( .gnd(gnd), .vdd(vdd), .A(data_103__5_), .Y(_5141_) );
OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_5126_), .C(_5141_), .Y(_5142_) );
NAND3X1 NAND3X1_697 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_5128_), .C(_3313__bF_buf33), .Y(_5143_) );
AND2X2 AND2X2_1038 ( .gnd(gnd), .vdd(vdd), .A(_5142_), .B(_5143_), .Y(_5__5_) );
INVX1 INVX1_2292 ( .gnd(gnd), .vdd(vdd), .A(data_103__6_), .Y(_5144_) );
MUX2X1 MUX2X1_770 ( .gnd(gnd), .vdd(vdd), .A(_5144_), .B(_15049__bF_buf12), .S(_5134_), .Y(_5__6_) );
INVX1 INVX1_2293 ( .gnd(gnd), .vdd(vdd), .A(data_103__7_), .Y(_5145_) );
OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_5126_), .C(_5145_), .Y(_5146_) );
NAND3X1 NAND3X1_698 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_5128_), .C(_3313__bF_buf32), .Y(_5147_) );
AND2X2 AND2X2_1039 ( .gnd(gnd), .vdd(vdd), .A(_5146_), .B(_5147_), .Y(_5__7_) );
INVX1 INVX1_2294 ( .gnd(gnd), .vdd(vdd), .A(data_103__8_), .Y(_5148_) );
MUX2X1 MUX2X1_771 ( .gnd(gnd), .vdd(vdd), .A(_5148_), .B(_15052__bF_buf4), .S(_5134_), .Y(_5__8_) );
INVX1 INVX1_2295 ( .gnd(gnd), .vdd(vdd), .A(data_103__9_), .Y(_5149_) );
MUX2X1 MUX2X1_772 ( .gnd(gnd), .vdd(vdd), .A(_5149_), .B(_14913__bF_buf11), .S(_5134_), .Y(_5__9_) );
INVX1 INVX1_2296 ( .gnd(gnd), .vdd(vdd), .A(data_103__10_), .Y(_5150_) );
MUX2X1 MUX2X1_773 ( .gnd(gnd), .vdd(vdd), .A(_5150_), .B(_15055__bF_buf7), .S(_5134_), .Y(_5__10_) );
INVX1 INVX1_2297 ( .gnd(gnd), .vdd(vdd), .A(data_103__11_), .Y(_5151_) );
OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_5126_), .C(_5151_), .Y(_5152_) );
NAND3X1 NAND3X1_699 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_5128_), .C(_3313__bF_buf31), .Y(_5153_) );
AND2X2 AND2X2_1040 ( .gnd(gnd), .vdd(vdd), .A(_5152_), .B(_5153_), .Y(_5__11_) );
INVX1 INVX1_2298 ( .gnd(gnd), .vdd(vdd), .A(data_103__12_), .Y(_5154_) );
OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_5126_), .C(_5154_), .Y(_5155_) );
NAND3X1 NAND3X1_700 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_5128_), .C(_3313__bF_buf30), .Y(_5156_) );
AND2X2 AND2X2_1041 ( .gnd(gnd), .vdd(vdd), .A(_5155_), .B(_5156_), .Y(_5__12_) );
INVX1 INVX1_2299 ( .gnd(gnd), .vdd(vdd), .A(data_103__13_), .Y(_5157_) );
MUX2X1 MUX2X1_774 ( .gnd(gnd), .vdd(vdd), .A(_5157_), .B(_14924__bF_buf5), .S(_5134_), .Y(_5__13_) );
INVX1 INVX1_2300 ( .gnd(gnd), .vdd(vdd), .A(data_103__14_), .Y(_5158_) );
MUX2X1 MUX2X1_775 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_15060__bF_buf14), .S(_5134_), .Y(_5__14_) );
INVX1 INVX1_2301 ( .gnd(gnd), .vdd(vdd), .A(data_103__15_), .Y(_5159_) );
MUX2X1 MUX2X1_776 ( .gnd(gnd), .vdd(vdd), .A(_5159_), .B(_15062__bF_buf6), .S(_5134_), .Y(_5__15_) );
INVX1 INVX1_2302 ( .gnd(gnd), .vdd(vdd), .A(data_102__0_), .Y(_5160_) );
OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf4), .B(IDATA_PROG_addr_3_bF_buf1), .C(_3354__bF_buf0), .Y(_5161_) );
OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_16156_), .B(_3863_), .C(_3354__bF_buf3), .Y(_5162_) );
NAND3X1 NAND3X1_701 ( .gnd(gnd), .vdd(vdd), .A(_5161_), .B(_5162_), .C(_5122_), .Y(_5163_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_5163_), .Y(_5164_) );
OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_5164_), .C(_5160_), .Y(_5165_) );
NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_5163_), .B(_4287_), .Y(_5166_) );
NAND3X1 NAND3X1_702 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_5166_), .C(_3313__bF_buf29), .Y(_5167_) );
AND2X2 AND2X2_1042 ( .gnd(gnd), .vdd(vdd), .A(_5165_), .B(_5167_), .Y(_4__0_) );
INVX1 INVX1_2303 ( .gnd(gnd), .vdd(vdd), .A(data_102__1_), .Y(_5168_) );
OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_5164_), .C(_5168_), .Y(_5169_) );
NAND3X1 NAND3X1_703 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_5166_), .C(_3313__bF_buf28), .Y(_5170_) );
AND2X2 AND2X2_1043 ( .gnd(gnd), .vdd(vdd), .A(_5169_), .B(_5170_), .Y(_4__1_) );
INVX1 INVX1_2304 ( .gnd(gnd), .vdd(vdd), .A(data_102__2_), .Y(_5171_) );
NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_5166_), .B(_3313__bF_buf27), .Y(_5172_) );
MUX2X1 MUX2X1_777 ( .gnd(gnd), .vdd(vdd), .A(_5171_), .B(_14897__bF_buf8), .S(_5172_), .Y(_4__2_) );
INVX1 INVX1_2305 ( .gnd(gnd), .vdd(vdd), .A(data_102__3_), .Y(_5173_) );
OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_5164_), .C(_5173_), .Y(_5174_) );
NAND3X1 NAND3X1_704 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_5166_), .C(_3313__bF_buf26), .Y(_5175_) );
AND2X2 AND2X2_1044 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_5175_), .Y(_4__3_) );
INVX1 INVX1_2306 ( .gnd(gnd), .vdd(vdd), .A(data_102__4_), .Y(_5176_) );
OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_5164_), .C(_5176_), .Y(_5177_) );
NAND3X1 NAND3X1_705 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_5166_), .C(_3313__bF_buf25), .Y(_5178_) );
AND2X2 AND2X2_1045 ( .gnd(gnd), .vdd(vdd), .A(_5177_), .B(_5178_), .Y(_4__4_) );
INVX1 INVX1_2307 ( .gnd(gnd), .vdd(vdd), .A(data_102__5_), .Y(_5179_) );
OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf24), .B(_5164_), .C(_5179_), .Y(_5180_) );
NAND3X1 NAND3X1_706 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_5166_), .C(_3313__bF_buf24), .Y(_5181_) );
AND2X2 AND2X2_1046 ( .gnd(gnd), .vdd(vdd), .A(_5180_), .B(_5181_), .Y(_4__5_) );
INVX1 INVX1_2308 ( .gnd(gnd), .vdd(vdd), .A(data_102__6_), .Y(_5182_) );
MUX2X1 MUX2X1_778 ( .gnd(gnd), .vdd(vdd), .A(_5182_), .B(_15049__bF_buf11), .S(_5172_), .Y(_4__6_) );
INVX1 INVX1_2309 ( .gnd(gnd), .vdd(vdd), .A(data_102__7_), .Y(_5183_) );
OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_5164_), .C(_5183_), .Y(_5184_) );
NAND3X1 NAND3X1_707 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_5166_), .C(_3313__bF_buf23), .Y(_5185_) );
AND2X2 AND2X2_1047 ( .gnd(gnd), .vdd(vdd), .A(_5184_), .B(_5185_), .Y(_4__7_) );
INVX1 INVX1_2310 ( .gnd(gnd), .vdd(vdd), .A(data_102__8_), .Y(_5186_) );
MUX2X1 MUX2X1_779 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_15052__bF_buf3), .S(_5172_), .Y(_4__8_) );
INVX1 INVX1_2311 ( .gnd(gnd), .vdd(vdd), .A(data_102__9_), .Y(_5187_) );
MUX2X1 MUX2X1_780 ( .gnd(gnd), .vdd(vdd), .A(_5187_), .B(_14913__bF_buf10), .S(_5172_), .Y(_4__9_) );
INVX1 INVX1_2312 ( .gnd(gnd), .vdd(vdd), .A(data_102__10_), .Y(_5188_) );
MUX2X1 MUX2X1_781 ( .gnd(gnd), .vdd(vdd), .A(_5188_), .B(_15055__bF_buf6), .S(_5172_), .Y(_4__10_) );
INVX1 INVX1_2313 ( .gnd(gnd), .vdd(vdd), .A(data_102__11_), .Y(_5189_) );
OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_5164_), .C(_5189_), .Y(_5190_) );
NAND3X1 NAND3X1_708 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_5166_), .C(_3313__bF_buf22), .Y(_5191_) );
AND2X2 AND2X2_1048 ( .gnd(gnd), .vdd(vdd), .A(_5190_), .B(_5191_), .Y(_4__11_) );
INVX1 INVX1_2314 ( .gnd(gnd), .vdd(vdd), .A(data_102__12_), .Y(_5192_) );
OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_5164_), .C(_5192_), .Y(_5193_) );
NAND3X1 NAND3X1_709 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_5166_), .C(_3313__bF_buf21), .Y(_5194_) );
AND2X2 AND2X2_1049 ( .gnd(gnd), .vdd(vdd), .A(_5193_), .B(_5194_), .Y(_4__12_) );
INVX1 INVX1_2315 ( .gnd(gnd), .vdd(vdd), .A(data_102__13_), .Y(_5195_) );
MUX2X1 MUX2X1_782 ( .gnd(gnd), .vdd(vdd), .A(_5195_), .B(_14924__bF_buf4), .S(_5172_), .Y(_4__13_) );
INVX1 INVX1_2316 ( .gnd(gnd), .vdd(vdd), .A(data_102__14_), .Y(_5196_) );
MUX2X1 MUX2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_5196_), .B(_15060__bF_buf13), .S(_5172_), .Y(_4__14_) );
INVX1 INVX1_2317 ( .gnd(gnd), .vdd(vdd), .A(data_102__15_), .Y(_5197_) );
MUX2X1 MUX2X1_784 ( .gnd(gnd), .vdd(vdd), .A(_5197_), .B(_15062__bF_buf5), .S(_5172_), .Y(_4__15_) );
OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3982_), .C(_4604_), .Y(_5198_) );
NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(_5121_), .Y(_5199_) );
NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_5161_), .B(_5199_), .Y(_5200_) );
NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_5200_), .B(_4287_), .Y(_5201_) );
AND2X2 AND2X2_1050 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf20), .B(_5201_), .Y(_5202_) );
AOI21X1 AOI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf19), .C(data_101__0_), .Y(_5203_) );
AOI21X1 AOI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_5202_), .C(_5203_), .Y(_3__0_) );
AOI21X1 AOI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf18), .C(data_101__1_), .Y(_5204_) );
AOI21X1 AOI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_5202_), .C(_5204_), .Y(_3__1_) );
AOI21X1 AOI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf17), .C(data_101__2_), .Y(_5205_) );
AOI21X1 AOI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_5202_), .C(_5205_), .Y(_3__2_) );
AOI21X1 AOI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf16), .C(data_101__3_), .Y(_5206_) );
AOI21X1 AOI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_5202_), .C(_5206_), .Y(_3__3_) );
AOI21X1 AOI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf15), .C(data_101__4_), .Y(_5207_) );
AOI21X1 AOI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_5202_), .C(_5207_), .Y(_3__4_) );
INVX1 INVX1_2318 ( .gnd(gnd), .vdd(vdd), .A(data_101__5_), .Y(_5208_) );
NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf14), .Y(_5209_) );
MUX2X1 MUX2X1_785 ( .gnd(gnd), .vdd(vdd), .A(_5208_), .B(_14903__bF_buf2), .S(_5209_), .Y(_3__5_) );
AOI21X1 AOI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf13), .C(data_101__6_), .Y(_5210_) );
AOI21X1 AOI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_5202_), .C(_5210_), .Y(_3__6_) );
INVX1 INVX1_2319 ( .gnd(gnd), .vdd(vdd), .A(data_101__7_), .Y(_5211_) );
MUX2X1 MUX2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_5211_), .B(_14908__bF_buf4), .S(_5209_), .Y(_3__7_) );
AOI21X1 AOI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf12), .C(data_101__8_), .Y(_5212_) );
AOI21X1 AOI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_5202_), .C(_5212_), .Y(_3__8_) );
AOI21X1 AOI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf11), .C(data_101__9_), .Y(_5213_) );
AOI21X1 AOI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_5202_), .C(_5213_), .Y(_3__9_) );
AOI21X1 AOI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf10), .C(data_101__10_), .Y(_5214_) );
AOI21X1 AOI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_5202_), .C(_5214_), .Y(_3__10_) );
AOI21X1 AOI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf9), .C(data_101__11_), .Y(_5215_) );
AOI21X1 AOI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_5202_), .C(_5215_), .Y(_3__11_) );
INVX1 INVX1_2320 ( .gnd(gnd), .vdd(vdd), .A(data_101__12_), .Y(_5216_) );
MUX2X1 MUX2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_5216_), .B(_14920__bF_buf4), .S(_5209_), .Y(_3__12_) );
AOI21X1 AOI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf8), .C(data_101__13_), .Y(_5217_) );
AOI21X1 AOI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_5202_), .C(_5217_), .Y(_3__13_) );
AOI21X1 AOI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf7), .C(data_101__14_), .Y(_5218_) );
AOI21X1 AOI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf12), .B(_5202_), .C(_5218_), .Y(_3__14_) );
AOI21X1 AOI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_3313__bF_buf6), .C(data_101__15_), .Y(_5219_) );
AOI21X1 AOI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_5202_), .C(_5219_), .Y(_3__15_) );
OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_4026_), .B(IDATA_PROG_addr_3_bF_buf0), .C(_3354__bF_buf2), .Y(_5220_) );
NAND3X1 NAND3X1_710 ( .gnd(gnd), .vdd(vdd), .A(_5199_), .B(_5220_), .C(_4243_), .Y(_5221_) );
NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_5221_), .B(_3393__bF_buf20), .Y(_5222_) );
INVX1 INVX1_2321 ( .gnd(gnd), .vdd(vdd), .A(_5199_), .Y(_5223_) );
INVX1 INVX1_2322 ( .gnd(gnd), .vdd(vdd), .A(_5220_), .Y(_5224_) );
NOR3X1 NOR3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_5223_), .B(_5224_), .C(_4287_), .Y(_5225_) );
AOI21X1 AOI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf5), .B(_5225_), .C(data_100__0_), .Y(_5226_) );
AOI21X1 AOI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_5222_), .C(_5226_), .Y(_2__0_) );
AOI21X1 AOI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf4), .B(_5225_), .C(data_100__1_), .Y(_5227_) );
AOI21X1 AOI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_5222_), .C(_5227_), .Y(_2__1_) );
NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf3), .B(_5225_), .Y(_5228_) );
INVX1 INVX1_2323 ( .gnd(gnd), .vdd(vdd), .A(data_100__2_), .Y(_5229_) );
OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_5221_), .C(_5229_), .Y(_5230_) );
OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf2), .B(_5228_), .C(_5230_), .Y(_5231_) );
INVX1 INVX1_2324 ( .gnd(gnd), .vdd(vdd), .A(_5231_), .Y(_2__2_) );
AOI21X1 AOI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf2), .B(_5225_), .C(data_100__3_), .Y(_5232_) );
AOI21X1 AOI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_5222_), .C(_5232_), .Y(_2__3_) );
AOI21X1 AOI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf1), .B(_5225_), .C(data_100__4_), .Y(_5233_) );
AOI21X1 AOI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_5222_), .C(_5233_), .Y(_2__4_) );
INVX1 INVX1_2325 ( .gnd(gnd), .vdd(vdd), .A(data_100__5_), .Y(_5234_) );
OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_5221_), .C(_5234_), .Y(_5235_) );
OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf1), .B(_5228_), .C(_5235_), .Y(_5236_) );
INVX1 INVX1_2326 ( .gnd(gnd), .vdd(vdd), .A(_5236_), .Y(_2__5_) );
INVX1 INVX1_2327 ( .gnd(gnd), .vdd(vdd), .A(data_100__6_), .Y(_5237_) );
OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf17), .B(_5221_), .C(_5237_), .Y(_5238_) );
OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf3), .B(_5228_), .C(_5238_), .Y(_5239_) );
INVX1 INVX1_2328 ( .gnd(gnd), .vdd(vdd), .A(_5239_), .Y(_2__6_) );
INVX1 INVX1_2329 ( .gnd(gnd), .vdd(vdd), .A(data_100__7_), .Y(_5240_) );
OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf16), .B(_5221_), .C(_5240_), .Y(_5241_) );
OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf3), .B(_5228_), .C(_5241_), .Y(_5242_) );
INVX1 INVX1_2330 ( .gnd(gnd), .vdd(vdd), .A(_5242_), .Y(_2__7_) );
INVX1 INVX1_2331 ( .gnd(gnd), .vdd(vdd), .A(data_100__8_), .Y(_5243_) );
OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf15), .B(_5221_), .C(_5243_), .Y(_5244_) );
OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf1), .B(_5228_), .C(_5244_), .Y(_5245_) );
INVX1 INVX1_2332 ( .gnd(gnd), .vdd(vdd), .A(_5245_), .Y(_2__8_) );
AOI21X1 AOI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf0), .B(_5225_), .C(data_100__9_), .Y(_5246_) );
AOI21X1 AOI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_5222_), .C(_5246_), .Y(_2__9_) );
AOI21X1 AOI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf91), .B(_5225_), .C(data_100__10_), .Y(_5247_) );
AOI21X1 AOI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_5222_), .C(_5247_), .Y(_2__10_) );
AOI21X1 AOI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf90), .B(_5225_), .C(data_100__11_), .Y(_5248_) );
AOI21X1 AOI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_5222_), .C(_5248_), .Y(_2__11_) );
INVX1 INVX1_2333 ( .gnd(gnd), .vdd(vdd), .A(data_100__12_), .Y(_5249_) );
OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf14), .B(_5221_), .C(_5249_), .Y(_5250_) );
OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf4), .B(_5228_), .C(_5250_), .Y(_5251_) );
INVX1 INVX1_2334 ( .gnd(gnd), .vdd(vdd), .A(_5251_), .Y(_2__12_) );
AOI21X1 AOI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf89), .B(_5225_), .C(data_100__13_), .Y(_5252_) );
AOI21X1 AOI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_5222_), .C(_5252_), .Y(_2__13_) );
INVX1 INVX1_2335 ( .gnd(gnd), .vdd(vdd), .A(data_100__14_), .Y(_5253_) );
OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf13), .B(_5221_), .C(_5253_), .Y(_5254_) );
OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf1), .B(_5228_), .C(_5254_), .Y(_5255_) );
INVX1 INVX1_2336 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .Y(_2__14_) );
INVX1 INVX1_2337 ( .gnd(gnd), .vdd(vdd), .A(data_100__15_), .Y(_5256_) );
OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_5221_), .C(_5256_), .Y(_5257_) );
OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf3), .B(_5228_), .C(_5257_), .Y(_5258_) );
INVX1 INVX1_2338 ( .gnd(gnd), .vdd(vdd), .A(_5258_), .Y(_2__15_) );
INVX1 INVX1_2339 ( .gnd(gnd), .vdd(vdd), .A(data_99__0_), .Y(_5259_) );
OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf2), .B(_3357_), .C(_5122_), .Y(_5260_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_5260_), .Y(_5261_) );
OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_5261_), .C(_5259_), .Y(_5262_) );
NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_5260_), .B(_4287_), .Y(_5263_) );
NAND3X1 NAND3X1_711 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_5263_), .C(_3313__bF_buf88), .Y(_5264_) );
AND2X2 AND2X2_1051 ( .gnd(gnd), .vdd(vdd), .A(_5262_), .B(_5264_), .Y(_255__0_) );
INVX1 INVX1_2340 ( .gnd(gnd), .vdd(vdd), .A(data_99__1_), .Y(_5265_) );
OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_5261_), .C(_5265_), .Y(_5266_) );
NAND3X1 NAND3X1_712 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_5263_), .C(_3313__bF_buf87), .Y(_5267_) );
AND2X2 AND2X2_1052 ( .gnd(gnd), .vdd(vdd), .A(_5266_), .B(_5267_), .Y(_255__1_) );
NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_5261_), .B(_3393__bF_buf9), .Y(_5268_) );
AOI21X1 AOI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_3313__bF_buf86), .C(data_99__2_), .Y(_5269_) );
AOI21X1 AOI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_5268_), .C(_5269_), .Y(_255__2_) );
INVX1 INVX1_2341 ( .gnd(gnd), .vdd(vdd), .A(data_99__3_), .Y(_5270_) );
OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf8), .B(_5261_), .C(_5270_), .Y(_5271_) );
NAND3X1 NAND3X1_713 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_5263_), .C(_3313__bF_buf85), .Y(_5272_) );
AND2X2 AND2X2_1053 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .B(_5272_), .Y(_255__3_) );
INVX1 INVX1_2342 ( .gnd(gnd), .vdd(vdd), .A(data_99__4_), .Y(_5273_) );
OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_5261_), .C(_5273_), .Y(_5274_) );
NAND3X1 NAND3X1_714 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_5263_), .C(_3313__bF_buf84), .Y(_5275_) );
AND2X2 AND2X2_1054 ( .gnd(gnd), .vdd(vdd), .A(_5274_), .B(_5275_), .Y(_255__4_) );
INVX1 INVX1_2343 ( .gnd(gnd), .vdd(vdd), .A(data_99__5_), .Y(_5276_) );
NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_3313__bF_buf83), .Y(_5277_) );
MUX2X1 MUX2X1_788 ( .gnd(gnd), .vdd(vdd), .A(_5276_), .B(_14903__bF_buf1), .S(_5277_), .Y(_255__5_) );
AOI21X1 AOI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_3313__bF_buf82), .C(data_99__6_), .Y(_5278_) );
AOI21X1 AOI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_5268_), .C(_5278_), .Y(_255__6_) );
INVX1 INVX1_2344 ( .gnd(gnd), .vdd(vdd), .A(data_99__7_), .Y(_5279_) );
MUX2X1 MUX2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_5279_), .B(_14908__bF_buf3), .S(_5277_), .Y(_255__7_) );
AOI21X1 AOI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_3313__bF_buf81), .C(data_99__8_), .Y(_5280_) );
AOI21X1 AOI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_5268_), .C(_5280_), .Y(_255__8_) );
INVX1 INVX1_2345 ( .gnd(gnd), .vdd(vdd), .A(data_99__9_), .Y(_5281_) );
MUX2X1 MUX2X1_790 ( .gnd(gnd), .vdd(vdd), .A(_5281_), .B(_14913__bF_buf7), .S(_5277_), .Y(_255__9_) );
INVX1 INVX1_2346 ( .gnd(gnd), .vdd(vdd), .A(data_99__10_), .Y(_5282_) );
MUX2X1 MUX2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_5282_), .B(_15055__bF_buf3), .S(_5277_), .Y(_255__10_) );
INVX1 INVX1_2347 ( .gnd(gnd), .vdd(vdd), .A(data_99__11_), .Y(_5283_) );
OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_5261_), .C(_5283_), .Y(_5284_) );
NAND3X1 NAND3X1_715 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_5263_), .C(_3313__bF_buf80), .Y(_5285_) );
AND2X2 AND2X2_1055 ( .gnd(gnd), .vdd(vdd), .A(_5284_), .B(_5285_), .Y(_255__11_) );
INVX1 INVX1_2348 ( .gnd(gnd), .vdd(vdd), .A(data_99__12_), .Y(_5286_) );
MUX2X1 MUX2X1_792 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .B(_14920__bF_buf3), .S(_5277_), .Y(_255__12_) );
INVX1 INVX1_2349 ( .gnd(gnd), .vdd(vdd), .A(data_99__13_), .Y(_5287_) );
MUX2X1 MUX2X1_793 ( .gnd(gnd), .vdd(vdd), .A(_5287_), .B(_14924__bF_buf1), .S(_5277_), .Y(_255__13_) );
AOI21X1 AOI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_3313__bF_buf79), .C(data_99__14_), .Y(_5288_) );
AOI21X1 AOI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_5268_), .C(_5288_), .Y(_255__14_) );
AOI21X1 AOI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_3313__bF_buf78), .C(data_99__15_), .Y(_5289_) );
AOI21X1 AOI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_5268_), .C(_5289_), .Y(_255__15_) );
INVX1 INVX1_2350 ( .gnd(gnd), .vdd(vdd), .A(data_98__0_), .Y(_5290_) );
NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_4604_), .B(_3359_), .Y(_5291_) );
NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_5123_), .B(_5291_), .Y(_5292_) );
OAI21X1 OAI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .B(_14952__bF_buf1), .C(_3354__bF_buf1), .Y(_5293_) );
NAND3X1 NAND3X1_716 ( .gnd(gnd), .vdd(vdd), .A(_5292_), .B(_5293_), .C(_4243_), .Y(_5294_) );
OAI21X1 OAI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_5294_), .C(_5290_), .Y(_5295_) );
INVX1 INVX1_2351 ( .gnd(gnd), .vdd(vdd), .A(_5292_), .Y(_5296_) );
INVX1 INVX1_2352 ( .gnd(gnd), .vdd(vdd), .A(_5293_), .Y(_5297_) );
NOR3X1 NOR3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_5296_), .B(_5297_), .C(_4287_), .Y(_5298_) );
NAND3X1 NAND3X1_717 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_3313__bF_buf77), .C(_5298_), .Y(_5299_) );
AND2X2 AND2X2_1056 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .B(_5299_), .Y(_254__0_) );
INVX1 INVX1_2353 ( .gnd(gnd), .vdd(vdd), .A(data_98__1_), .Y(_5300_) );
OAI21X1 OAI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_5294_), .C(_5300_), .Y(_5301_) );
NAND3X1 NAND3X1_718 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_3313__bF_buf76), .C(_5298_), .Y(_5302_) );
AND2X2 AND2X2_1057 ( .gnd(gnd), .vdd(vdd), .A(_5301_), .B(_5302_), .Y(_254__1_) );
NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_5294_), .B(_3393__bF_buf3), .Y(_5303_) );
AOI21X1 AOI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf75), .B(_5298_), .C(data_98__2_), .Y(_5304_) );
AOI21X1 AOI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_5303_), .C(_5304_), .Y(_254__2_) );
INVX1 INVX1_2354 ( .gnd(gnd), .vdd(vdd), .A(data_98__3_), .Y(_5305_) );
OAI21X1 OAI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_5294_), .C(_5305_), .Y(_5306_) );
NAND3X1 NAND3X1_719 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_3313__bF_buf74), .C(_5298_), .Y(_5307_) );
AND2X2 AND2X2_1058 ( .gnd(gnd), .vdd(vdd), .A(_5306_), .B(_5307_), .Y(_254__3_) );
INVX1 INVX1_2355 ( .gnd(gnd), .vdd(vdd), .A(data_98__4_), .Y(_5308_) );
OAI21X1 OAI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_5294_), .C(_5308_), .Y(_5309_) );
NAND3X1 NAND3X1_720 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_3313__bF_buf73), .C(_5298_), .Y(_5310_) );
AND2X2 AND2X2_1059 ( .gnd(gnd), .vdd(vdd), .A(_5309_), .B(_5310_), .Y(_254__4_) );
INVX1 INVX1_2356 ( .gnd(gnd), .vdd(vdd), .A(data_98__5_), .Y(_5311_) );
NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf72), .B(_5298_), .Y(_5312_) );
MUX2X1 MUX2X1_794 ( .gnd(gnd), .vdd(vdd), .A(_5311_), .B(_14903__bF_buf0), .S(_5312_), .Y(_254__5_) );
AOI21X1 AOI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf71), .B(_5298_), .C(data_98__6_), .Y(_5313_) );
AOI21X1 AOI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_5303_), .C(_5313_), .Y(_254__6_) );
INVX1 INVX1_2357 ( .gnd(gnd), .vdd(vdd), .A(data_98__7_), .Y(_5314_) );
MUX2X1 MUX2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_5314_), .B(_14908__bF_buf2), .S(_5312_), .Y(_254__7_) );
AOI21X1 AOI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf70), .B(_5298_), .C(data_98__8_), .Y(_5315_) );
AOI21X1 AOI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_5303_), .C(_5315_), .Y(_254__8_) );
INVX1 INVX1_2358 ( .gnd(gnd), .vdd(vdd), .A(data_98__9_), .Y(_5316_) );
MUX2X1 MUX2X1_796 ( .gnd(gnd), .vdd(vdd), .A(_5316_), .B(_14913__bF_buf6), .S(_5312_), .Y(_254__9_) );
INVX1 INVX1_2359 ( .gnd(gnd), .vdd(vdd), .A(data_98__10_), .Y(_5317_) );
MUX2X1 MUX2X1_797 ( .gnd(gnd), .vdd(vdd), .A(_5317_), .B(_15055__bF_buf2), .S(_5312_), .Y(_254__10_) );
INVX1 INVX1_2360 ( .gnd(gnd), .vdd(vdd), .A(data_98__11_), .Y(_5318_) );
OAI21X1 OAI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_5294_), .C(_5318_), .Y(_5319_) );
NAND3X1 NAND3X1_721 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_3313__bF_buf69), .C(_5298_), .Y(_5320_) );
AND2X2 AND2X2_1060 ( .gnd(gnd), .vdd(vdd), .A(_5319_), .B(_5320_), .Y(_254__11_) );
INVX1 INVX1_2361 ( .gnd(gnd), .vdd(vdd), .A(data_98__12_), .Y(_5321_) );
MUX2X1 MUX2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_5321_), .B(_14920__bF_buf2), .S(_5312_), .Y(_254__12_) );
INVX1 INVX1_2362 ( .gnd(gnd), .vdd(vdd), .A(data_98__13_), .Y(_5322_) );
MUX2X1 MUX2X1_799 ( .gnd(gnd), .vdd(vdd), .A(_5322_), .B(_14924__bF_buf0), .S(_5312_), .Y(_254__13_) );
AOI21X1 AOI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf68), .B(_5298_), .C(data_98__14_), .Y(_5323_) );
AOI21X1 AOI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_5303_), .C(_5323_), .Y(_254__14_) );
AOI21X1 AOI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf67), .B(_5298_), .C(data_98__15_), .Y(_5324_) );
AOI21X1 AOI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf2), .B(_5303_), .C(_5324_), .Y(_254__15_) );
INVX1 INVX1_2363 ( .gnd(gnd), .vdd(vdd), .A(data_97__0_), .Y(_5325_) );
INVX1 INVX1_2364 ( .gnd(gnd), .vdd(vdd), .A(_3492_), .Y(_5326_) );
OAI21X1 OAI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_5326_), .B(_14952__bF_buf0), .C(_3354__bF_buf0), .Y(_5327_) );
INVX1 INVX1_2365 ( .gnd(gnd), .vdd(vdd), .A(_5327_), .Y(_5328_) );
NOR3X1 NOR3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_5296_), .B(_5328_), .C(_4287_), .Y(_5329_) );
NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf66), .B(_5329_), .Y(_5330_) );
MUX2X1 MUX2X1_800 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .B(_14932__bF_buf10), .S(_5330_), .Y(_253__0_) );
INVX1 INVX1_2366 ( .gnd(gnd), .vdd(vdd), .A(data_97__1_), .Y(_5331_) );
MUX2X1 MUX2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_5331_), .B(_14894__bF_buf7), .S(_5330_), .Y(_253__1_) );
INVX1 INVX1_2367 ( .gnd(gnd), .vdd(vdd), .A(data_97__2_), .Y(_5332_) );
MUX2X1 MUX2X1_802 ( .gnd(gnd), .vdd(vdd), .A(_5332_), .B(_14897__bF_buf4), .S(_5330_), .Y(_253__2_) );
INVX1 INVX1_2368 ( .gnd(gnd), .vdd(vdd), .A(data_97__3_), .Y(_5333_) );
MUX2X1 MUX2X1_803 ( .gnd(gnd), .vdd(vdd), .A(_5333_), .B(_14899__bF_buf7), .S(_5330_), .Y(_253__3_) );
INVX1 INVX1_2369 ( .gnd(gnd), .vdd(vdd), .A(data_97__4_), .Y(_5334_) );
MUX2X1 MUX2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_5334_), .B(_14902__bF_buf13), .S(_5330_), .Y(_253__4_) );
INVX1 INVX1_2370 ( .gnd(gnd), .vdd(vdd), .A(data_97__5_), .Y(_5335_) );
NAND3X1 NAND3X1_722 ( .gnd(gnd), .vdd(vdd), .A(_5292_), .B(_5327_), .C(_4243_), .Y(_5336_) );
OAI21X1 OAI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_5336_), .C(_5335_), .Y(_5337_) );
NAND3X1 NAND3X1_723 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_3313__bF_buf65), .C(_5329_), .Y(_5338_) );
AND2X2 AND2X2_1061 ( .gnd(gnd), .vdd(vdd), .A(_5337_), .B(_5338_), .Y(_253__5_) );
INVX1 INVX1_2371 ( .gnd(gnd), .vdd(vdd), .A(data_97__6_), .Y(_5339_) );
MUX2X1 MUX2X1_805 ( .gnd(gnd), .vdd(vdd), .A(_5339_), .B(_15049__bF_buf7), .S(_5330_), .Y(_253__6_) );
INVX1 INVX1_2372 ( .gnd(gnd), .vdd(vdd), .A(data_97__7_), .Y(_5340_) );
OAI21X1 OAI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_5336_), .C(_5340_), .Y(_5341_) );
NAND3X1 NAND3X1_724 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_3313__bF_buf64), .C(_5329_), .Y(_5342_) );
AND2X2 AND2X2_1062 ( .gnd(gnd), .vdd(vdd), .A(_5341_), .B(_5342_), .Y(_253__7_) );
INVX1 INVX1_2373 ( .gnd(gnd), .vdd(vdd), .A(data_97__8_), .Y(_5343_) );
MUX2X1 MUX2X1_806 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .B(_15052__bF_buf13), .S(_5330_), .Y(_253__8_) );
NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(_5336_), .B(_3393__bF_buf67), .Y(_5344_) );
AOI21X1 AOI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf63), .B(_5329_), .C(data_97__9_), .Y(_5345_) );
AOI21X1 AOI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_5344_), .C(_5345_), .Y(_253__9_) );
AOI21X1 AOI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf62), .B(_5329_), .C(data_97__10_), .Y(_5346_) );
AOI21X1 AOI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_5344_), .C(_5346_), .Y(_253__10_) );
INVX1 INVX1_2374 ( .gnd(gnd), .vdd(vdd), .A(data_97__11_), .Y(_5347_) );
MUX2X1 MUX2X1_807 ( .gnd(gnd), .vdd(vdd), .A(_5347_), .B(_14918__bF_buf1), .S(_5330_), .Y(_253__11_) );
INVX1 INVX1_2375 ( .gnd(gnd), .vdd(vdd), .A(data_97__12_), .Y(_5348_) );
OAI21X1 OAI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_5336_), .C(_5348_), .Y(_5349_) );
NAND3X1 NAND3X1_725 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_3313__bF_buf61), .C(_5329_), .Y(_5350_) );
AND2X2 AND2X2_1063 ( .gnd(gnd), .vdd(vdd), .A(_5349_), .B(_5350_), .Y(_253__12_) );
AOI21X1 AOI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf60), .B(_5329_), .C(data_97__13_), .Y(_5351_) );
AOI21X1 AOI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_5344_), .C(_5351_), .Y(_253__13_) );
INVX1 INVX1_2376 ( .gnd(gnd), .vdd(vdd), .A(data_97__14_), .Y(_5352_) );
MUX2X1 MUX2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_5352_), .B(_15060__bF_buf9), .S(_5330_), .Y(_253__14_) );
INVX1 INVX1_2377 ( .gnd(gnd), .vdd(vdd), .A(data_97__15_), .Y(_5353_) );
MUX2X1 MUX2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_5353_), .B(_15062__bF_buf1), .S(_5330_), .Y(_253__15_) );
NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf0), .B(_3626_), .Y(_5354_) );
NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(data_96__0_), .B(_5354__bF_buf3), .Y(_5355_) );
AOI21X1 AOI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_5354__bF_buf2), .C(_5355_), .Y(_252__0_) );
INVX1 INVX1_2378 ( .gnd(gnd), .vdd(vdd), .A(data_96__1_), .Y(_5356_) );
MUX2X1 MUX2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_5356_), .S(_5354__bF_buf1), .Y(_252__1_) );
NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(data_96__2_), .B(_5354__bF_buf0), .Y(_5357_) );
NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_3358_), .Y(_5358_) );
NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf1), .B(_5358_), .Y(_5359_) );
NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_5357_), .B(_5359_), .Y(_252__2_) );
NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(data_96__3_), .B(_5354__bF_buf3), .Y(_5360_) );
AOI21X1 AOI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_5354__bF_buf2), .C(_5360_), .Y(_252__3_) );
INVX1 INVX1_2379 ( .gnd(gnd), .vdd(vdd), .A(data_96__4_), .Y(_5361_) );
OAI21X1 OAI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_14882__bF_buf15_bF_buf2), .C(_5361_), .Y(_5362_) );
OAI21X1 OAI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_5358_), .B(IDATA_PROG_data_4_bF_buf0), .C(_5362_), .Y(_5363_) );
INVX1 INVX1_2380 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .Y(_252__4_) );
INVX1 INVX1_2381 ( .gnd(gnd), .vdd(vdd), .A(data_96__5_), .Y(_5364_) );
OAI21X1 OAI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_14882__bF_buf14_bF_buf2), .C(_5364_), .Y(_5365_) );
OAI21X1 OAI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_5358_), .B(IDATA_PROG_data_5_bF_buf0), .C(_5365_), .Y(_5366_) );
INVX1 INVX1_2382 ( .gnd(gnd), .vdd(vdd), .A(_5366_), .Y(_252__5_) );
NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(data_96__6_), .B(_5354__bF_buf1), .Y(_5367_) );
AOI21X1 AOI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_5354__bF_buf0), .C(_5367_), .Y(_252__6_) );
NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_5354__bF_buf3), .Y(_5368_) );
OAI21X1 OAI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(data_96__7_), .B(_5354__bF_buf2), .C(_5368_), .Y(_5369_) );
INVX1 INVX1_2383 ( .gnd(gnd), .vdd(vdd), .A(_5369_), .Y(_252__7_) );
NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(data_96__8_), .B(_5354__bF_buf1), .Y(_5370_) );
AOI21X1 AOI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_5354__bF_buf0), .C(_5370_), .Y(_252__8_) );
MUX2X1 MUX2X1_811 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf4), .B(data_96__9_), .S(_5354__bF_buf3), .Y(_5371_) );
INVX1 INVX1_2384 ( .gnd(gnd), .vdd(vdd), .A(_5371_), .Y(_252__9_) );
INVX1 INVX1_2385 ( .gnd(gnd), .vdd(vdd), .A(data_96__10_), .Y(_5372_) );
OAI21X1 OAI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_14882__bF_buf13_bF_buf2), .C(_5372_), .Y(_5373_) );
OAI21X1 OAI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_5358_), .B(IDATA_PROG_data_10_bF_buf3), .C(_5373_), .Y(_5374_) );
INVX1 INVX1_2386 ( .gnd(gnd), .vdd(vdd), .A(_5374_), .Y(_252__10_) );
INVX1 INVX1_2387 ( .gnd(gnd), .vdd(vdd), .A(data_96__11_), .Y(_5375_) );
MUX2X1 MUX2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_5375_), .S(_5354__bF_buf2), .Y(_252__11_) );
INVX1 INVX1_2388 ( .gnd(gnd), .vdd(vdd), .A(data_96__12_), .Y(_5376_) );
OAI21X1 OAI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_14882__bF_buf12), .C(_5376_), .Y(_5377_) );
OAI21X1 OAI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_5358_), .B(IDATA_PROG_data_12_bF_buf3), .C(_5377_), .Y(_5378_) );
INVX1 INVX1_2389 ( .gnd(gnd), .vdd(vdd), .A(_5378_), .Y(_252__12_) );
NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_5354__bF_buf1), .Y(_5379_) );
OAI21X1 OAI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(data_96__13_), .B(_5354__bF_buf0), .C(_5379_), .Y(_5380_) );
INVX1 INVX1_2390 ( .gnd(gnd), .vdd(vdd), .A(_5380_), .Y(_252__13_) );
NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(data_96__14_), .B(_5354__bF_buf3), .Y(_5381_) );
AOI21X1 AOI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_5354__bF_buf2), .C(_5381_), .Y(_252__14_) );
NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(data_96__15_), .B(_5354__bF_buf1), .Y(_5382_) );
AOI21X1 AOI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_5354__bF_buf0), .C(_5382_), .Y(_252__15_) );
NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf0), .B(_3324_), .Y(_5383_) );
NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf11), .B(_5383_), .Y(_5384_) );
NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(data_95__0_), .B(_5384__bF_buf3), .Y(_5385_) );
AOI21X1 AOI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_5384__bF_buf2), .C(_5385_), .Y(_251__0_) );
NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_3356_), .Y(_5386_) );
INVX1 INVX1_2391 ( .gnd(gnd), .vdd(vdd), .A(data_95__1_), .Y(_5387_) );
OAI21X1 OAI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_14882__bF_buf10), .C(_5387_), .Y(_5388_) );
OAI21X1 OAI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(IDATA_PROG_data_1_bF_buf2), .C(_5388_), .Y(_5389_) );
INVX1 INVX1_2392 ( .gnd(gnd), .vdd(vdd), .A(_5389_), .Y(_251__1_) );
NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(data_95__2_), .B(_5384__bF_buf1), .Y(_5390_) );
AOI21X1 AOI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_5384__bF_buf0), .C(_5390_), .Y(_251__2_) );
NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(data_95__3_), .B(_5384__bF_buf3), .Y(_5391_) );
AOI21X1 AOI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_5384__bF_buf2), .C(_5391_), .Y(_251__3_) );
INVX1 INVX1_2393 ( .gnd(gnd), .vdd(vdd), .A(data_95__4_), .Y(_5392_) );
OAI21X1 OAI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_14882__bF_buf9), .C(_5392_), .Y(_5393_) );
NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_5384__bF_buf1), .Y(_5394_) );
AND2X2 AND2X2_1064 ( .gnd(gnd), .vdd(vdd), .A(_5394_), .B(_5393_), .Y(_251__4_) );
NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_5384__bF_buf0), .Y(_5395_) );
OAI21X1 OAI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(data_95__5_), .B(_5384__bF_buf3), .C(_5395_), .Y(_5396_) );
INVX1 INVX1_2394 ( .gnd(gnd), .vdd(vdd), .A(_5396_), .Y(_251__5_) );
NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(data_95__6_), .B(_5384__bF_buf2), .Y(_5397_) );
AOI21X1 AOI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_5384__bF_buf1), .C(_5397_), .Y(_251__6_) );
INVX1 INVX1_2395 ( .gnd(gnd), .vdd(vdd), .A(data_95__7_), .Y(_5398_) );
OAI21X1 OAI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_14882__bF_buf8), .C(_5398_), .Y(_5399_) );
OAI21X1 OAI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(IDATA_PROG_data_7_bF_buf2), .C(_5399_), .Y(_5400_) );
INVX1 INVX1_2396 ( .gnd(gnd), .vdd(vdd), .A(_5400_), .Y(_251__7_) );
INVX1 INVX1_2397 ( .gnd(gnd), .vdd(vdd), .A(data_95__8_), .Y(_5401_) );
OAI21X1 OAI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_14882__bF_buf7), .C(_5401_), .Y(_5402_) );
OAI21X1 OAI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(IDATA_PROG_data_8_bF_buf0), .C(_5402_), .Y(_5403_) );
INVX1 INVX1_2398 ( .gnd(gnd), .vdd(vdd), .A(_5403_), .Y(_251__8_) );
INVX1 INVX1_2399 ( .gnd(gnd), .vdd(vdd), .A(data_95__9_), .Y(_5404_) );
OAI21X1 OAI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_14882__bF_buf6), .C(_5404_), .Y(_5405_) );
OAI21X1 OAI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(IDATA_PROG_data_9_bF_buf3), .C(_5405_), .Y(_5406_) );
INVX1 INVX1_2400 ( .gnd(gnd), .vdd(vdd), .A(_5406_), .Y(_251__9_) );
NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_5384__bF_buf0), .Y(_5407_) );
OAI21X1 OAI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(data_95__10_), .B(_5384__bF_buf3), .C(_5407_), .Y(_5408_) );
INVX1 INVX1_2401 ( .gnd(gnd), .vdd(vdd), .A(_5408_), .Y(_251__10_) );
NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_5384__bF_buf2), .Y(_5409_) );
OAI21X1 OAI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(data_95__11_), .B(_5384__bF_buf1), .C(_5409_), .Y(_5410_) );
INVX1 INVX1_2402 ( .gnd(gnd), .vdd(vdd), .A(_5410_), .Y(_251__11_) );
INVX1 INVX1_2403 ( .gnd(gnd), .vdd(vdd), .A(data_95__12_), .Y(_5411_) );
OAI21X1 OAI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_5383_), .B(_14882__bF_buf5), .C(_5411_), .Y(_5412_) );
OAI21X1 OAI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_5386_), .B(IDATA_PROG_data_12_bF_buf2), .C(_5412_), .Y(_5413_) );
INVX1 INVX1_2404 ( .gnd(gnd), .vdd(vdd), .A(_5413_), .Y(_251__12_) );
NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_5384__bF_buf0), .Y(_5414_) );
OAI21X1 OAI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(data_95__13_), .B(_5384__bF_buf3), .C(_5414_), .Y(_5415_) );
INVX1 INVX1_2405 ( .gnd(gnd), .vdd(vdd), .A(_5415_), .Y(_251__13_) );
NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(data_95__14_), .B(_5384__bF_buf2), .Y(_5416_) );
AOI21X1 AOI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_5384__bF_buf1), .C(_5416_), .Y(_251__14_) );
NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(data_95__15_), .B(_5384__bF_buf0), .Y(_5417_) );
AOI21X1 AOI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_5384__bF_buf3), .C(_5417_), .Y(_251__15_) );
INVX1 INVX1_2406 ( .gnd(gnd), .vdd(vdd), .A(data_94__0_), .Y(_5418_) );
NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(_4285_), .Y(_5419_) );
NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_5419_), .Y(_5420_) );
OAI21X1 OAI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_14940_), .B(_3323_), .C(IDATA_PROG_write_bF_buf5), .Y(_5421_) );
OAI21X1 OAI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_14947_), .B(_14886__bF_buf3), .C(_3362_), .Y(_5422_) );
OAI21X1 OAI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_5422_), .B(_749_), .C(_5421_), .Y(_5423_) );
NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_5423_), .B(_4279_), .Y(_5424_) );
NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_5420__bF_buf3), .B(_5424_), .Y(_5425_) );
INVX4 INVX4_17 ( .gnd(gnd), .vdd(vdd), .A(_5425_), .Y(_5426_) );
OAI21X1 OAI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_5426_), .C(_5418_), .Y(_5427_) );
NAND3X1 NAND3X1_726 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_5425_), .C(_3313__bF_buf59), .Y(_5428_) );
AND2X2 AND2X2_1065 ( .gnd(gnd), .vdd(vdd), .A(_5427_), .B(_5428_), .Y(_250__0_) );
INVX1 INVX1_2407 ( .gnd(gnd), .vdd(vdd), .A(data_94__1_), .Y(_5429_) );
OAI21X1 OAI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_5426_), .C(_5429_), .Y(_5430_) );
NAND3X1 NAND3X1_727 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_5425_), .C(_3313__bF_buf58), .Y(_5431_) );
AND2X2 AND2X2_1066 ( .gnd(gnd), .vdd(vdd), .A(_5430_), .B(_5431_), .Y(_250__1_) );
INVX1 INVX1_2408 ( .gnd(gnd), .vdd(vdd), .A(data_94__2_), .Y(_5432_) );
NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_5425_), .B(_3313__bF_buf57), .Y(_5433_) );
MUX2X1 MUX2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_5432_), .B(_14897__bF_buf2), .S(_5433_), .Y(_250__2_) );
INVX1 INVX1_2409 ( .gnd(gnd), .vdd(vdd), .A(data_94__3_), .Y(_5434_) );
OAI21X1 OAI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_5426_), .C(_5434_), .Y(_5435_) );
NAND3X1 NAND3X1_728 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_5425_), .C(_3313__bF_buf56), .Y(_5436_) );
AND2X2 AND2X2_1067 ( .gnd(gnd), .vdd(vdd), .A(_5435_), .B(_5436_), .Y(_250__3_) );
INVX1 INVX1_2410 ( .gnd(gnd), .vdd(vdd), .A(data_94__4_), .Y(_5437_) );
OAI21X1 OAI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_5426_), .C(_5437_), .Y(_5438_) );
NAND3X1 NAND3X1_729 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_5425_), .C(_3313__bF_buf55), .Y(_5439_) );
AND2X2 AND2X2_1068 ( .gnd(gnd), .vdd(vdd), .A(_5438_), .B(_5439_), .Y(_250__4_) );
INVX1 INVX1_2411 ( .gnd(gnd), .vdd(vdd), .A(data_94__5_), .Y(_5440_) );
OAI21X1 OAI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_5426_), .C(_5440_), .Y(_5441_) );
NAND3X1 NAND3X1_730 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_5425_), .C(_3313__bF_buf54), .Y(_5442_) );
AND2X2 AND2X2_1069 ( .gnd(gnd), .vdd(vdd), .A(_5441_), .B(_5442_), .Y(_250__5_) );
INVX1 INVX1_2412 ( .gnd(gnd), .vdd(vdd), .A(data_94__6_), .Y(_5443_) );
MUX2X1 MUX2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_5443_), .B(_15049__bF_buf4), .S(_5433_), .Y(_250__6_) );
NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_5426_), .B(_3393__bF_buf60), .Y(_5444_) );
AOI21X1 AOI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_5425_), .B(_3313__bF_buf53), .C(data_94__7_), .Y(_5445_) );
AOI21X1 AOI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_5444_), .C(_5445_), .Y(_250__7_) );
INVX1 INVX1_2413 ( .gnd(gnd), .vdd(vdd), .A(data_94__8_), .Y(_5446_) );
MUX2X1 MUX2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_5446_), .B(_15052__bF_buf11), .S(_5433_), .Y(_250__8_) );
AOI21X1 AOI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_5425_), .B(_3313__bF_buf52), .C(data_94__9_), .Y(_5447_) );
AOI21X1 AOI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_5444_), .C(_5447_), .Y(_250__9_) );
AOI21X1 AOI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_5425_), .B(_3313__bF_buf51), .C(data_94__10_), .Y(_5448_) );
AOI21X1 AOI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_5444_), .C(_5448_), .Y(_250__10_) );
INVX1 INVX1_2414 ( .gnd(gnd), .vdd(vdd), .A(data_94__11_), .Y(_5449_) );
OAI21X1 OAI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_5426_), .C(_5449_), .Y(_5450_) );
NAND3X1 NAND3X1_731 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_5425_), .C(_3313__bF_buf50), .Y(_5451_) );
AND2X2 AND2X2_1070 ( .gnd(gnd), .vdd(vdd), .A(_5450_), .B(_5451_), .Y(_250__11_) );
INVX1 INVX1_2415 ( .gnd(gnd), .vdd(vdd), .A(data_94__12_), .Y(_5452_) );
OAI21X1 OAI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_5426_), .C(_5452_), .Y(_5453_) );
NAND3X1 NAND3X1_732 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_5425_), .C(_3313__bF_buf49), .Y(_5454_) );
AND2X2 AND2X2_1071 ( .gnd(gnd), .vdd(vdd), .A(_5453_), .B(_5454_), .Y(_250__12_) );
INVX1 INVX1_2416 ( .gnd(gnd), .vdd(vdd), .A(data_94__13_), .Y(_5455_) );
MUX2X1 MUX2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_5455_), .B(_14924__bF_buf10), .S(_5433_), .Y(_250__13_) );
INVX1 INVX1_2417 ( .gnd(gnd), .vdd(vdd), .A(data_94__14_), .Y(_5456_) );
MUX2X1 MUX2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_5456_), .B(_15060__bF_buf6), .S(_5433_), .Y(_250__14_) );
INVX1 INVX1_2418 ( .gnd(gnd), .vdd(vdd), .A(data_94__15_), .Y(_5457_) );
MUX2X1 MUX2X1_818 ( .gnd(gnd), .vdd(vdd), .A(_5457_), .B(_15062__bF_buf12), .S(_5433_), .Y(_250__15_) );
INVX1 INVX1_2419 ( .gnd(gnd), .vdd(vdd), .A(data_93__0_), .Y(_5458_) );
NAND3X1 NAND3X1_733 ( .gnd(gnd), .vdd(vdd), .A(_14936__bF_buf1), .B(_14971_), .C(_3644_), .Y(_5459_) );
NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_3341_), .B(_3351_), .Y(_5460_) );
NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_5460_), .B(_5459__bF_buf3), .Y(_5461_) );
OAI21X1 OAI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_14949_), .B(_14886__bF_buf2), .C(_3362_), .Y(_5462_) );
INVX1 INVX1_2420 ( .gnd(gnd), .vdd(vdd), .A(_5462_), .Y(_5463_) );
NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_5463_), .Y(_5464_) );
AOI21X1 AOI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_5421_), .B(_5464_), .C(_3339_), .Y(_5465_) );
NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5465_), .Y(_5466_) );
OAI21X1 OAI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_5466_), .C(_5458_), .Y(_5467_) );
AND2X2 AND2X2_1072 ( .gnd(gnd), .vdd(vdd), .A(_5465_), .B(_5461_), .Y(_5468_) );
NAND3X1 NAND3X1_734 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_5468_), .C(_3313__bF_buf48), .Y(_5469_) );
AND2X2 AND2X2_1073 ( .gnd(gnd), .vdd(vdd), .A(_5467_), .B(_5469_), .Y(_249__0_) );
INVX1 INVX1_2421 ( .gnd(gnd), .vdd(vdd), .A(data_93__1_), .Y(_5470_) );
OAI21X1 OAI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_5466_), .C(_5470_), .Y(_5471_) );
NAND3X1 NAND3X1_735 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_5468_), .C(_3313__bF_buf47), .Y(_5472_) );
AND2X2 AND2X2_1074 ( .gnd(gnd), .vdd(vdd), .A(_5471_), .B(_5472_), .Y(_249__1_) );
INVX1 INVX1_2422 ( .gnd(gnd), .vdd(vdd), .A(data_93__2_), .Y(_5473_) );
NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_5468_), .B(_3313__bF_buf46), .Y(_5474_) );
MUX2X1 MUX2X1_819 ( .gnd(gnd), .vdd(vdd), .A(_5473_), .B(_14897__bF_buf1), .S(_5474_), .Y(_249__2_) );
INVX1 INVX1_2423 ( .gnd(gnd), .vdd(vdd), .A(data_93__3_), .Y(_5475_) );
OAI21X1 OAI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_5466_), .C(_5475_), .Y(_5476_) );
NAND3X1 NAND3X1_736 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_5468_), .C(_3313__bF_buf45), .Y(_5477_) );
AND2X2 AND2X2_1075 ( .gnd(gnd), .vdd(vdd), .A(_5476_), .B(_5477_), .Y(_249__3_) );
INVX1 INVX1_2424 ( .gnd(gnd), .vdd(vdd), .A(data_93__4_), .Y(_5478_) );
OAI21X1 OAI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_5466_), .C(_5478_), .Y(_5479_) );
NAND3X1 NAND3X1_737 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_5468_), .C(_3313__bF_buf44), .Y(_5480_) );
AND2X2 AND2X2_1076 ( .gnd(gnd), .vdd(vdd), .A(_5479_), .B(_5480_), .Y(_249__4_) );
INVX1 INVX1_2425 ( .gnd(gnd), .vdd(vdd), .A(data_93__5_), .Y(_5481_) );
OAI21X1 OAI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_5466_), .C(_5481_), .Y(_5482_) );
NAND3X1 NAND3X1_738 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_5468_), .C(_3313__bF_buf43), .Y(_5483_) );
AND2X2 AND2X2_1077 ( .gnd(gnd), .vdd(vdd), .A(_5482_), .B(_5483_), .Y(_249__5_) );
INVX1 INVX1_2426 ( .gnd(gnd), .vdd(vdd), .A(data_93__6_), .Y(_5484_) );
MUX2X1 MUX2X1_820 ( .gnd(gnd), .vdd(vdd), .A(_5484_), .B(_15049__bF_buf3), .S(_5474_), .Y(_249__6_) );
INVX1 INVX1_2427 ( .gnd(gnd), .vdd(vdd), .A(data_93__7_), .Y(_5485_) );
MUX2X1 MUX2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_5485_), .B(_14908__bF_buf12), .S(_5474_), .Y(_249__7_) );
INVX1 INVX1_2428 ( .gnd(gnd), .vdd(vdd), .A(data_93__8_), .Y(_5486_) );
MUX2X1 MUX2X1_822 ( .gnd(gnd), .vdd(vdd), .A(_5486_), .B(_15052__bF_buf10), .S(_5474_), .Y(_249__8_) );
NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_5466_), .B(_3393__bF_buf52), .Y(_5487_) );
AOI21X1 AOI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_5468_), .B(_3313__bF_buf42), .C(data_93__9_), .Y(_5488_) );
AOI21X1 AOI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_5487_), .C(_5488_), .Y(_249__9_) );
AOI21X1 AOI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_5468_), .B(_3313__bF_buf41), .C(data_93__10_), .Y(_5489_) );
AOI21X1 AOI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_5487_), .C(_5489_), .Y(_249__10_) );
INVX1 INVX1_2429 ( .gnd(gnd), .vdd(vdd), .A(data_93__11_), .Y(_5490_) );
OAI21X1 OAI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_5466_), .C(_5490_), .Y(_5491_) );
NAND3X1 NAND3X1_739 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_5468_), .C(_3313__bF_buf40), .Y(_5492_) );
AND2X2 AND2X2_1078 ( .gnd(gnd), .vdd(vdd), .A(_5491_), .B(_5492_), .Y(_249__11_) );
INVX1 INVX1_2430 ( .gnd(gnd), .vdd(vdd), .A(data_93__12_), .Y(_5493_) );
OAI21X1 OAI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_5466_), .C(_5493_), .Y(_5494_) );
NAND3X1 NAND3X1_740 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_5468_), .C(_3313__bF_buf39), .Y(_5495_) );
AND2X2 AND2X2_1079 ( .gnd(gnd), .vdd(vdd), .A(_5494_), .B(_5495_), .Y(_249__12_) );
INVX1 INVX1_2431 ( .gnd(gnd), .vdd(vdd), .A(data_93__13_), .Y(_5496_) );
MUX2X1 MUX2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_5496_), .B(_14924__bF_buf9), .S(_5474_), .Y(_249__13_) );
INVX1 INVX1_2432 ( .gnd(gnd), .vdd(vdd), .A(data_93__14_), .Y(_5497_) );
MUX2X1 MUX2X1_824 ( .gnd(gnd), .vdd(vdd), .A(_5497_), .B(_15060__bF_buf5), .S(_5474_), .Y(_249__14_) );
AOI21X1 AOI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_5468_), .B(_3313__bF_buf38), .C(data_93__15_), .Y(_5498_) );
AOI21X1 AOI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_5487_), .C(_5498_), .Y(_249__15_) );
INVX1 INVX1_2433 ( .gnd(gnd), .vdd(vdd), .A(data_92__0_), .Y(_5499_) );
NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_3338_), .B(_3335_), .Y(_5500_) );
NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_5500_), .B(_5459__bF_buf2), .Y(_5501_) );
OAI21X1 OAI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_5462_), .B(_3715_), .C(_3324_), .Y(_5502_) );
NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(_3326_), .Y(_5503_) );
NAND3X1 NAND3X1_741 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_4274_), .C(_5503_), .Y(_5504_) );
NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_5504_), .B(_5460_), .Y(_5505_) );
NAND3X1 NAND3X1_742 ( .gnd(gnd), .vdd(vdd), .A(_5502_), .B(_5505_), .C(_5501_), .Y(_5506_) );
OAI21X1 OAI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_5506_), .C(_5499_), .Y(_5507_) );
INVX8 INVX8_30 ( .gnd(gnd), .vdd(vdd), .A(_5506_), .Y(_5508_) );
NAND3X1 NAND3X1_743 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_5508_), .C(_3313__bF_buf37), .Y(_5509_) );
AND2X2 AND2X2_1080 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .B(_5509_), .Y(_248__0_) );
INVX1 INVX1_2434 ( .gnd(gnd), .vdd(vdd), .A(data_92__1_), .Y(_5510_) );
OAI21X1 OAI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_5506_), .C(_5510_), .Y(_5511_) );
NAND3X1 NAND3X1_744 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_5508_), .C(_3313__bF_buf36), .Y(_5512_) );
AND2X2 AND2X2_1081 ( .gnd(gnd), .vdd(vdd), .A(_5511_), .B(_5512_), .Y(_248__1_) );
NOR3X1 NOR3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_5506_), .C(_3989__bF_buf1), .Y(_5513_) );
AOI21X1 AOI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_5508_), .B(_3313__bF_buf35), .C(data_92__2_), .Y(_5514_) );
AOI21X1 AOI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_5513_), .C(_5514_), .Y(_248__2_) );
INVX1 INVX1_2435 ( .gnd(gnd), .vdd(vdd), .A(data_92__3_), .Y(_5515_) );
OAI21X1 OAI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_5506_), .C(_5515_), .Y(_5516_) );
NAND3X1 NAND3X1_745 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_5508_), .C(_3313__bF_buf34), .Y(_5517_) );
AND2X2 AND2X2_1082 ( .gnd(gnd), .vdd(vdd), .A(_5516_), .B(_5517_), .Y(_248__3_) );
INVX1 INVX1_2436 ( .gnd(gnd), .vdd(vdd), .A(data_92__4_), .Y(_5518_) );
OAI21X1 OAI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_5506_), .C(_5518_), .Y(_5519_) );
NAND3X1 NAND3X1_746 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_5508_), .C(_3313__bF_buf33), .Y(_5520_) );
AND2X2 AND2X2_1083 ( .gnd(gnd), .vdd(vdd), .A(_5519_), .B(_5520_), .Y(_248__4_) );
INVX1 INVX1_2437 ( .gnd(gnd), .vdd(vdd), .A(data_92__5_), .Y(_5521_) );
OAI21X1 OAI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_5506_), .C(_5521_), .Y(_5522_) );
NAND3X1 NAND3X1_747 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_5508_), .C(_3313__bF_buf32), .Y(_5523_) );
AND2X2 AND2X2_1084 ( .gnd(gnd), .vdd(vdd), .A(_5522_), .B(_5523_), .Y(_248__5_) );
AOI21X1 AOI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_5508_), .B(_3313__bF_buf31), .C(data_92__6_), .Y(_5524_) );
AOI21X1 AOI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_5513_), .C(_5524_), .Y(_248__6_) );
INVX1 INVX1_2438 ( .gnd(gnd), .vdd(vdd), .A(data_92__7_), .Y(_5525_) );
OAI21X1 OAI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_5506_), .C(_5525_), .Y(_5526_) );
NAND3X1 NAND3X1_748 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_5508_), .C(_3313__bF_buf30), .Y(_5527_) );
AND2X2 AND2X2_1085 ( .gnd(gnd), .vdd(vdd), .A(_5526_), .B(_5527_), .Y(_248__7_) );
AOI21X1 AOI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_5508_), .B(_3313__bF_buf29), .C(data_92__8_), .Y(_5528_) );
AOI21X1 AOI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_5513_), .C(_5528_), .Y(_248__8_) );
INVX1 INVX1_2439 ( .gnd(gnd), .vdd(vdd), .A(data_92__9_), .Y(_5529_) );
NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_5508_), .B(_3313__bF_buf28), .Y(_5530_) );
MUX2X1 MUX2X1_825 ( .gnd(gnd), .vdd(vdd), .A(_5529_), .B(_14913__bF_buf2), .S(_5530_), .Y(_248__9_) );
INVX1 INVX1_2440 ( .gnd(gnd), .vdd(vdd), .A(data_92__10_), .Y(_5531_) );
MUX2X1 MUX2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_5531_), .B(_15055__bF_buf11), .S(_5530_), .Y(_248__10_) );
INVX1 INVX1_2441 ( .gnd(gnd), .vdd(vdd), .A(data_92__11_), .Y(_5532_) );
OAI21X1 OAI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_5506_), .C(_5532_), .Y(_5533_) );
NAND3X1 NAND3X1_749 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_5508_), .C(_3313__bF_buf27), .Y(_5534_) );
AND2X2 AND2X2_1086 ( .gnd(gnd), .vdd(vdd), .A(_5533_), .B(_5534_), .Y(_248__11_) );
INVX1 INVX1_2442 ( .gnd(gnd), .vdd(vdd), .A(data_92__12_), .Y(_5535_) );
OAI21X1 OAI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_5506_), .C(_5535_), .Y(_5536_) );
NAND3X1 NAND3X1_750 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_5508_), .C(_3313__bF_buf26), .Y(_5537_) );
AND2X2 AND2X2_1087 ( .gnd(gnd), .vdd(vdd), .A(_5536_), .B(_5537_), .Y(_248__12_) );
INVX1 INVX1_2443 ( .gnd(gnd), .vdd(vdd), .A(data_92__13_), .Y(_5538_) );
MUX2X1 MUX2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_5538_), .B(_14924__bF_buf8), .S(_5530_), .Y(_248__13_) );
INVX1 INVX1_2444 ( .gnd(gnd), .vdd(vdd), .A(data_92__14_), .Y(_5539_) );
MUX2X1 MUX2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_5539_), .B(_15060__bF_buf4), .S(_5530_), .Y(_248__14_) );
INVX1 INVX1_2445 ( .gnd(gnd), .vdd(vdd), .A(data_92__15_), .Y(_5540_) );
MUX2X1 MUX2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_5540_), .B(_15062__bF_buf10), .S(_5530_), .Y(_248__15_) );
INVX1 INVX1_2446 ( .gnd(gnd), .vdd(vdd), .A(data_91__0_), .Y(_5541_) );
NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(_4278_), .B(_4277_), .Y(_5542_) );
NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_5542_), .B(_14973_), .Y(_5543_) );
OAI21X1 OAI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_14963__bF_buf3), .C(_3324_), .Y(_5544_) );
NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_5544_), .B(_5505_), .Y(_5545_) );
NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_5543_), .B(_5545_), .Y(_5546_) );
NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf25), .Y(_5547_) );
MUX2X1 MUX2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_5541_), .B(_14932__bF_buf4), .S(_5547_), .Y(_247__0_) );
INVX1 INVX1_2447 ( .gnd(gnd), .vdd(vdd), .A(data_91__1_), .Y(_5548_) );
MUX2X1 MUX2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_5548_), .B(_14894__bF_buf2), .S(_5547_), .Y(_247__1_) );
AND2X2 AND2X2_1088 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf24), .B(_5546_), .Y(_5549_) );
AOI21X1 AOI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf23), .C(data_91__2_), .Y(_5550_) );
AOI21X1 AOI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_5549_), .C(_5550_), .Y(_247__2_) );
INVX1 INVX1_2448 ( .gnd(gnd), .vdd(vdd), .A(data_91__3_), .Y(_5551_) );
MUX2X1 MUX2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_5551_), .B(_14899__bF_buf1), .S(_5547_), .Y(_247__3_) );
INVX1 INVX1_2449 ( .gnd(gnd), .vdd(vdd), .A(data_91__4_), .Y(_5552_) );
MUX2X1 MUX2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_5552_), .B(_14902__bF_buf8), .S(_5547_), .Y(_247__4_) );
INVX1 INVX1_2450 ( .gnd(gnd), .vdd(vdd), .A(data_91__5_), .Y(_5553_) );
MUX2X1 MUX2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_5553_), .B(_14903__bF_buf8), .S(_5547_), .Y(_247__5_) );
AOI21X1 AOI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf22), .C(data_91__6_), .Y(_5554_) );
AOI21X1 AOI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_5549_), .C(_5554_), .Y(_247__6_) );
INVX1 INVX1_2451 ( .gnd(gnd), .vdd(vdd), .A(data_91__7_), .Y(_5555_) );
MUX2X1 MUX2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_5555_), .B(_14908__bF_buf10), .S(_5547_), .Y(_247__7_) );
AOI21X1 AOI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf21), .C(data_91__8_), .Y(_5556_) );
AOI21X1 AOI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_5549_), .C(_5556_), .Y(_247__8_) );
AOI21X1 AOI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf20), .C(data_91__9_), .Y(_5557_) );
AOI21X1 AOI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_5549_), .C(_5557_), .Y(_247__9_) );
AOI21X1 AOI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf19), .C(data_91__10_), .Y(_5558_) );
AOI21X1 AOI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_5549_), .C(_5558_), .Y(_247__10_) );
INVX1 INVX1_2452 ( .gnd(gnd), .vdd(vdd), .A(data_91__11_), .Y(_5559_) );
MUX2X1 MUX2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_5559_), .B(_14918__bF_buf9), .S(_5547_), .Y(_247__11_) );
INVX1 INVX1_2453 ( .gnd(gnd), .vdd(vdd), .A(data_91__12_), .Y(_5560_) );
MUX2X1 MUX2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_5560_), .B(_14920__bF_buf11), .S(_5547_), .Y(_247__12_) );
AOI21X1 AOI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf18), .C(data_91__13_), .Y(_5561_) );
AOI21X1 AOI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_5549_), .C(_5561_), .Y(_247__13_) );
AOI21X1 AOI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf17), .C(data_91__14_), .Y(_5562_) );
AOI21X1 AOI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_5549_), .C(_5562_), .Y(_247__14_) );
AOI21X1 AOI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_5546_), .B(_3313__bF_buf16), .C(data_91__15_), .Y(_5563_) );
AOI21X1 AOI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_5549_), .C(_5563_), .Y(_247__15_) );
INVX1 INVX1_2454 ( .gnd(gnd), .vdd(vdd), .A(data_90__0_), .Y(_5564_) );
NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf2), .B(_3324_), .Y(_5565_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(_5421_), .Y(_5566_) );
OAI21X1 OAI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_4388_), .B(_5566_), .C(_5565_), .Y(_5567_) );
NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_5567_), .B(_3339_), .Y(_5568_) );
NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5568_), .Y(_5569_) );
INVX4 INVX4_18 ( .gnd(gnd), .vdd(vdd), .A(_5569_), .Y(_5570_) );
NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_5570_), .B(_3313__bF_buf15), .Y(_5571_) );
MUX2X1 MUX2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_5564_), .B(_14932__bF_buf3), .S(_5571_), .Y(_246__0_) );
INVX1 INVX1_2455 ( .gnd(gnd), .vdd(vdd), .A(data_90__1_), .Y(_5572_) );
MUX2X1 MUX2X1_839 ( .gnd(gnd), .vdd(vdd), .A(_5572_), .B(_14894__bF_buf1), .S(_5571_), .Y(_246__1_) );
INVX1 INVX1_2456 ( .gnd(gnd), .vdd(vdd), .A(data_90__2_), .Y(_5573_) );
MUX2X1 MUX2X1_840 ( .gnd(gnd), .vdd(vdd), .A(_5573_), .B(_14897__bF_buf13), .S(_5571_), .Y(_246__2_) );
INVX1 INVX1_2457 ( .gnd(gnd), .vdd(vdd), .A(data_90__3_), .Y(_5574_) );
MUX2X1 MUX2X1_841 ( .gnd(gnd), .vdd(vdd), .A(_5574_), .B(_14899__bF_buf0), .S(_5571_), .Y(_246__3_) );
INVX1 INVX1_2458 ( .gnd(gnd), .vdd(vdd), .A(data_90__4_), .Y(_5575_) );
MUX2X1 MUX2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_5575_), .B(_14902__bF_buf7), .S(_5571_), .Y(_246__4_) );
INVX1 INVX1_2459 ( .gnd(gnd), .vdd(vdd), .A(data_90__5_), .Y(_5576_) );
OAI21X1 OAI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_5569_), .C(_5576_), .Y(_5577_) );
NAND3X1 NAND3X1_751 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_5570_), .C(_3313__bF_buf14), .Y(_5578_) );
AND2X2 AND2X2_1089 ( .gnd(gnd), .vdd(vdd), .A(_5577_), .B(_5578_), .Y(_246__5_) );
INVX1 INVX1_2460 ( .gnd(gnd), .vdd(vdd), .A(data_90__6_), .Y(_5579_) );
MUX2X1 MUX2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_5579_), .B(_15049__bF_buf0), .S(_5571_), .Y(_246__6_) );
INVX1 INVX1_2461 ( .gnd(gnd), .vdd(vdd), .A(data_90__7_), .Y(_5580_) );
OAI21X1 OAI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_5569_), .C(_5580_), .Y(_5581_) );
NAND3X1 NAND3X1_752 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_5570_), .C(_3313__bF_buf13), .Y(_5582_) );
AND2X2 AND2X2_1090 ( .gnd(gnd), .vdd(vdd), .A(_5581_), .B(_5582_), .Y(_246__7_) );
INVX1 INVX1_2462 ( .gnd(gnd), .vdd(vdd), .A(data_90__8_), .Y(_5583_) );
MUX2X1 MUX2X1_844 ( .gnd(gnd), .vdd(vdd), .A(_5583_), .B(_15052__bF_buf7), .S(_5571_), .Y(_246__8_) );
NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_5569_), .B(_3393__bF_buf39), .Y(_5584_) );
AOI21X1 AOI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_5570_), .B(_3313__bF_buf12), .C(data_90__9_), .Y(_5585_) );
AOI21X1 AOI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_5584_), .C(_5585_), .Y(_246__9_) );
AOI21X1 AOI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_5570_), .B(_3313__bF_buf11), .C(data_90__10_), .Y(_5586_) );
AOI21X1 AOI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_5584_), .C(_5586_), .Y(_246__10_) );
INVX1 INVX1_2463 ( .gnd(gnd), .vdd(vdd), .A(data_90__11_), .Y(_5587_) );
MUX2X1 MUX2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_5587_), .B(_14918__bF_buf8), .S(_5571_), .Y(_246__11_) );
INVX1 INVX1_2464 ( .gnd(gnd), .vdd(vdd), .A(data_90__12_), .Y(_5588_) );
OAI21X1 OAI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_5569_), .C(_5588_), .Y(_5589_) );
NAND3X1 NAND3X1_753 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_5570_), .C(_3313__bF_buf10), .Y(_5590_) );
AND2X2 AND2X2_1091 ( .gnd(gnd), .vdd(vdd), .A(_5589_), .B(_5590_), .Y(_246__12_) );
AOI21X1 AOI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_5570_), .B(_3313__bF_buf9), .C(data_90__13_), .Y(_5591_) );
AOI21X1 AOI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_5584_), .C(_5591_), .Y(_246__13_) );
INVX1 INVX1_2465 ( .gnd(gnd), .vdd(vdd), .A(data_90__14_), .Y(_5592_) );
MUX2X1 MUX2X1_846 ( .gnd(gnd), .vdd(vdd), .A(_5592_), .B(_15060__bF_buf2), .S(_5571_), .Y(_246__14_) );
INVX1 INVX1_2466 ( .gnd(gnd), .vdd(vdd), .A(data_90__15_), .Y(_5593_) );
MUX2X1 MUX2X1_847 ( .gnd(gnd), .vdd(vdd), .A(_5593_), .B(_15062__bF_buf8), .S(_5571_), .Y(_246__15_) );
INVX1 INVX1_2467 ( .gnd(gnd), .vdd(vdd), .A(data_89__0_), .Y(_5594_) );
AOI21X1 AOI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_5421_), .C(_4275_), .Y(_5595_) );
NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_5595_), .B(_5419_), .Y(_5596_) );
NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_5543_), .B(_5596_), .Y(_5597_) );
NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_5597_), .B(_3313__bF_buf8), .Y(_5598_) );
MUX2X1 MUX2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_5594_), .B(_14932__bF_buf2), .S(_5598_), .Y(_244__0_) );
INVX1 INVX1_2468 ( .gnd(gnd), .vdd(vdd), .A(data_89__1_), .Y(_5599_) );
MUX2X1 MUX2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_5599_), .B(_14894__bF_buf0), .S(_5598_), .Y(_244__1_) );
INVX1 INVX1_2469 ( .gnd(gnd), .vdd(vdd), .A(data_89__2_), .Y(_5600_) );
MUX2X1 MUX2X1_850 ( .gnd(gnd), .vdd(vdd), .A(_5600_), .B(_14897__bF_buf12), .S(_5598_), .Y(_244__2_) );
INVX1 INVX1_2470 ( .gnd(gnd), .vdd(vdd), .A(data_89__3_), .Y(_5601_) );
MUX2X1 MUX2X1_851 ( .gnd(gnd), .vdd(vdd), .A(_5601_), .B(_14899__bF_buf14), .S(_5598_), .Y(_244__3_) );
INVX1 INVX1_2471 ( .gnd(gnd), .vdd(vdd), .A(data_89__4_), .Y(_5602_) );
MUX2X1 MUX2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_5602_), .B(_14902__bF_buf6), .S(_5598_), .Y(_244__4_) );
INVX1 INVX1_2472 ( .gnd(gnd), .vdd(vdd), .A(data_89__5_), .Y(_5603_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_5596_), .B(_5543_), .Y(_5604_) );
OAI21X1 OAI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_5604_), .C(_5603_), .Y(_5605_) );
NAND3X1 NAND3X1_754 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_5597_), .C(_3313__bF_buf7), .Y(_5606_) );
AND2X2 AND2X2_1092 ( .gnd(gnd), .vdd(vdd), .A(_5605_), .B(_5606_), .Y(_244__5_) );
INVX1 INVX1_2473 ( .gnd(gnd), .vdd(vdd), .A(data_89__6_), .Y(_5607_) );
MUX2X1 MUX2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_5607_), .B(_15049__bF_buf14), .S(_5598_), .Y(_244__6_) );
INVX1 INVX1_2474 ( .gnd(gnd), .vdd(vdd), .A(data_89__7_), .Y(_5608_) );
OAI21X1 OAI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_5604_), .C(_5608_), .Y(_5609_) );
NAND3X1 NAND3X1_755 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_5597_), .C(_3313__bF_buf6), .Y(_5610_) );
AND2X2 AND2X2_1093 ( .gnd(gnd), .vdd(vdd), .A(_5609_), .B(_5610_), .Y(_244__7_) );
INVX1 INVX1_2475 ( .gnd(gnd), .vdd(vdd), .A(data_89__8_), .Y(_5611_) );
MUX2X1 MUX2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_5611_), .B(_15052__bF_buf6), .S(_5598_), .Y(_244__8_) );
INVX1 INVX1_2476 ( .gnd(gnd), .vdd(vdd), .A(data_89__9_), .Y(_5612_) );
MUX2X1 MUX2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_5612_), .B(_14913__bF_buf14), .S(_5598_), .Y(_244__9_) );
INVX1 INVX1_2477 ( .gnd(gnd), .vdd(vdd), .A(data_89__10_), .Y(_5613_) );
MUX2X1 MUX2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_5613_), .B(_15055__bF_buf8), .S(_5598_), .Y(_244__10_) );
INVX1 INVX1_2478 ( .gnd(gnd), .vdd(vdd), .A(data_89__11_), .Y(_5614_) );
MUX2X1 MUX2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_5614_), .B(_14918__bF_buf7), .S(_5598_), .Y(_244__11_) );
INVX1 INVX1_2479 ( .gnd(gnd), .vdd(vdd), .A(data_89__12_), .Y(_5615_) );
OAI21X1 OAI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_5604_), .C(_5615_), .Y(_5616_) );
NAND3X1 NAND3X1_756 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_5597_), .C(_3313__bF_buf5), .Y(_5617_) );
AND2X2 AND2X2_1094 ( .gnd(gnd), .vdd(vdd), .A(_5616_), .B(_5617_), .Y(_244__12_) );
INVX1 INVX1_2480 ( .gnd(gnd), .vdd(vdd), .A(data_89__13_), .Y(_5618_) );
MUX2X1 MUX2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_5618_), .B(_14924__bF_buf5), .S(_5598_), .Y(_244__13_) );
NOR3X1 NOR3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_5604_), .C(_3989__bF_buf0), .Y(_5619_) );
AOI21X1 AOI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_5597_), .B(_3313__bF_buf4), .C(data_89__14_), .Y(_5620_) );
AOI21X1 AOI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_5619_), .C(_5620_), .Y(_244__14_) );
AOI21X1 AOI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_5597_), .B(_3313__bF_buf3), .C(data_89__15_), .Y(_5621_) );
AOI21X1 AOI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_5619_), .C(_5621_), .Y(_244__15_) );
INVX1 INVX1_2481 ( .gnd(gnd), .vdd(vdd), .A(data_88__0_), .Y(_5622_) );
OAI21X1 OAI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_4468_), .B(_5566_), .C(_5565_), .Y(_5623_) );
NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_5623_), .B(_5460_), .Y(_5624_) );
NAND3X1 NAND3X1_757 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_4279_), .C(_5624_), .Y(_5625_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_5625_), .Y(_5626_) );
NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_5626_), .B(_3313__bF_buf2), .Y(_5627_) );
MUX2X1 MUX2X1_859 ( .gnd(gnd), .vdd(vdd), .A(_5622_), .B(_14932__bF_buf1), .S(_5627_), .Y(_243__0_) );
INVX1 INVX1_2482 ( .gnd(gnd), .vdd(vdd), .A(data_88__1_), .Y(_5628_) );
MUX2X1 MUX2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_5628_), .B(_14894__bF_buf14), .S(_5627_), .Y(_243__1_) );
INVX1 INVX1_2483 ( .gnd(gnd), .vdd(vdd), .A(data_88__2_), .Y(_5629_) );
MUX2X1 MUX2X1_861 ( .gnd(gnd), .vdd(vdd), .A(_5629_), .B(_14897__bF_buf11), .S(_5627_), .Y(_243__2_) );
INVX1 INVX1_2484 ( .gnd(gnd), .vdd(vdd), .A(data_88__3_), .Y(_5630_) );
MUX2X1 MUX2X1_862 ( .gnd(gnd), .vdd(vdd), .A(_5630_), .B(_14899__bF_buf13), .S(_5627_), .Y(_243__3_) );
INVX1 INVX1_2485 ( .gnd(gnd), .vdd(vdd), .A(data_88__4_), .Y(_5631_) );
MUX2X1 MUX2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_5631_), .B(_14902__bF_buf5), .S(_5627_), .Y(_243__4_) );
INVX1 INVX1_2486 ( .gnd(gnd), .vdd(vdd), .A(data_88__5_), .Y(_5632_) );
OAI21X1 OAI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf34), .B(_5625_), .C(_5632_), .Y(_5633_) );
NAND3X1 NAND3X1_758 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_5626_), .C(_3313__bF_buf1), .Y(_5634_) );
AND2X2 AND2X2_1095 ( .gnd(gnd), .vdd(vdd), .A(_5633_), .B(_5634_), .Y(_243__5_) );
INVX1 INVX1_2487 ( .gnd(gnd), .vdd(vdd), .A(data_88__6_), .Y(_5635_) );
MUX2X1 MUX2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_5635_), .B(_15049__bF_buf13), .S(_5627_), .Y(_243__6_) );
INVX1 INVX1_2488 ( .gnd(gnd), .vdd(vdd), .A(data_88__7_), .Y(_5636_) );
OAI21X1 OAI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_5625_), .C(_5636_), .Y(_5637_) );
NAND3X1 NAND3X1_759 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_5626_), .C(_3313__bF_buf0), .Y(_5638_) );
AND2X2 AND2X2_1096 ( .gnd(gnd), .vdd(vdd), .A(_5637_), .B(_5638_), .Y(_243__7_) );
INVX1 INVX1_2489 ( .gnd(gnd), .vdd(vdd), .A(data_88__8_), .Y(_5639_) );
MUX2X1 MUX2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_5639_), .B(_15052__bF_buf5), .S(_5627_), .Y(_243__8_) );
INVX1 INVX1_2490 ( .gnd(gnd), .vdd(vdd), .A(data_88__9_), .Y(_5640_) );
MUX2X1 MUX2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_5640_), .B(_14913__bF_buf13), .S(_5627_), .Y(_243__9_) );
INVX1 INVX1_2491 ( .gnd(gnd), .vdd(vdd), .A(data_88__10_), .Y(_5641_) );
MUX2X1 MUX2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_5641_), .B(_15055__bF_buf7), .S(_5627_), .Y(_243__10_) );
INVX1 INVX1_2492 ( .gnd(gnd), .vdd(vdd), .A(data_88__11_), .Y(_5642_) );
MUX2X1 MUX2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_5642_), .B(_14918__bF_buf6), .S(_5627_), .Y(_243__11_) );
INVX1 INVX1_2493 ( .gnd(gnd), .vdd(vdd), .A(data_88__12_), .Y(_5643_) );
OAI21X1 OAI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_5625_), .C(_5643_), .Y(_5644_) );
NAND3X1 NAND3X1_760 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_5626_), .C(_3313__bF_buf91), .Y(_5645_) );
AND2X2 AND2X2_1097 ( .gnd(gnd), .vdd(vdd), .A(_5644_), .B(_5645_), .Y(_243__12_) );
INVX1 INVX1_2494 ( .gnd(gnd), .vdd(vdd), .A(data_88__13_), .Y(_5646_) );
MUX2X1 MUX2X1_869 ( .gnd(gnd), .vdd(vdd), .A(_5646_), .B(_14924__bF_buf4), .S(_5627_), .Y(_243__13_) );
NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_5625_), .B(_3393__bF_buf31), .Y(_5647_) );
AOI21X1 AOI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_5626_), .B(_3313__bF_buf90), .C(data_88__14_), .Y(_5648_) );
AOI21X1 AOI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_5647_), .C(_5648_), .Y(_243__14_) );
INVX1 INVX1_2495 ( .gnd(gnd), .vdd(vdd), .A(data_88__15_), .Y(_5649_) );
MUX2X1 MUX2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_5649_), .B(_15062__bF_buf6), .S(_5627_), .Y(_243__15_) );
INVX1 INVX1_2496 ( .gnd(gnd), .vdd(vdd), .A(data_87__0_), .Y(_5650_) );
AOI21X1 AOI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf3), .B(_3324_), .C(_5500_), .Y(_5651_) );
NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_5651_), .B(_5505_), .Y(_5652_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_5652_), .B(_5459__bF_buf1), .Y(_5653_) );
OAI21X1 OAI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf30), .C(_5650_), .Y(_5654_) );
NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(_5459__bF_buf0), .B(_5652_), .Y(_5655_) );
NAND3X1 NAND3X1_761 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_5655_), .C(_3313__bF_buf89), .Y(_5656_) );
AND2X2 AND2X2_1098 ( .gnd(gnd), .vdd(vdd), .A(_5654_), .B(_5656_), .Y(_242__0_) );
INVX1 INVX1_2497 ( .gnd(gnd), .vdd(vdd), .A(data_87__1_), .Y(_5657_) );
OAI21X1 OAI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf29), .C(_5657_), .Y(_5658_) );
NAND3X1 NAND3X1_762 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_5655_), .C(_3313__bF_buf88), .Y(_5659_) );
AND2X2 AND2X2_1099 ( .gnd(gnd), .vdd(vdd), .A(_5658_), .B(_5659_), .Y(_242__1_) );
INVX1 INVX1_2498 ( .gnd(gnd), .vdd(vdd), .A(data_87__2_), .Y(_5660_) );
NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_5655_), .B(_3313__bF_buf87), .Y(_5661_) );
MUX2X1 MUX2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_5660_), .B(_14897__bF_buf10), .S(_5661_), .Y(_242__2_) );
INVX1 INVX1_2499 ( .gnd(gnd), .vdd(vdd), .A(data_87__3_), .Y(_5662_) );
OAI21X1 OAI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf28), .C(_5662_), .Y(_5663_) );
NAND3X1 NAND3X1_763 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_5655_), .C(_3313__bF_buf86), .Y(_5664_) );
AND2X2 AND2X2_1100 ( .gnd(gnd), .vdd(vdd), .A(_5663_), .B(_5664_), .Y(_242__3_) );
INVX1 INVX1_2500 ( .gnd(gnd), .vdd(vdd), .A(data_87__4_), .Y(_5665_) );
OAI21X1 OAI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf27), .C(_5665_), .Y(_5666_) );
NAND3X1 NAND3X1_764 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_5655_), .C(_3313__bF_buf85), .Y(_5667_) );
AND2X2 AND2X2_1101 ( .gnd(gnd), .vdd(vdd), .A(_5666_), .B(_5667_), .Y(_242__4_) );
INVX1 INVX1_2501 ( .gnd(gnd), .vdd(vdd), .A(data_87__5_), .Y(_5668_) );
OAI21X1 OAI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf26), .C(_5668_), .Y(_5669_) );
NAND3X1 NAND3X1_765 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_5655_), .C(_3313__bF_buf84), .Y(_5670_) );
AND2X2 AND2X2_1102 ( .gnd(gnd), .vdd(vdd), .A(_5669_), .B(_5670_), .Y(_242__5_) );
INVX1 INVX1_2502 ( .gnd(gnd), .vdd(vdd), .A(data_87__6_), .Y(_5671_) );
MUX2X1 MUX2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_5671_), .B(_15049__bF_buf12), .S(_5661_), .Y(_242__6_) );
INVX1 INVX1_2503 ( .gnd(gnd), .vdd(vdd), .A(data_87__7_), .Y(_5672_) );
OAI21X1 OAI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf25), .C(_5672_), .Y(_5673_) );
NAND3X1 NAND3X1_766 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_5655_), .C(_3313__bF_buf83), .Y(_5674_) );
AND2X2 AND2X2_1103 ( .gnd(gnd), .vdd(vdd), .A(_5673_), .B(_5674_), .Y(_242__7_) );
INVX1 INVX1_2504 ( .gnd(gnd), .vdd(vdd), .A(data_87__8_), .Y(_5675_) );
MUX2X1 MUX2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_5675_), .B(_15052__bF_buf4), .S(_5661_), .Y(_242__8_) );
INVX1 INVX1_2505 ( .gnd(gnd), .vdd(vdd), .A(data_87__9_), .Y(_5676_) );
MUX2X1 MUX2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_5676_), .B(_14913__bF_buf12), .S(_5661_), .Y(_242__9_) );
INVX1 INVX1_2506 ( .gnd(gnd), .vdd(vdd), .A(data_87__10_), .Y(_5677_) );
MUX2X1 MUX2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_5677_), .B(_15055__bF_buf6), .S(_5661_), .Y(_242__10_) );
INVX1 INVX1_2507 ( .gnd(gnd), .vdd(vdd), .A(data_87__11_), .Y(_5678_) );
OAI21X1 OAI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf24), .C(_5678_), .Y(_5679_) );
NAND3X1 NAND3X1_767 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_5655_), .C(_3313__bF_buf82), .Y(_5680_) );
AND2X2 AND2X2_1104 ( .gnd(gnd), .vdd(vdd), .A(_5679_), .B(_5680_), .Y(_242__11_) );
INVX1 INVX1_2508 ( .gnd(gnd), .vdd(vdd), .A(data_87__12_), .Y(_5681_) );
OAI21X1 OAI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_5653_), .B(_3393__bF_buf23), .C(_5681_), .Y(_5682_) );
NAND3X1 NAND3X1_768 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_5655_), .C(_3313__bF_buf81), .Y(_5683_) );
AND2X2 AND2X2_1105 ( .gnd(gnd), .vdd(vdd), .A(_5682_), .B(_5683_), .Y(_242__12_) );
INVX1 INVX1_2509 ( .gnd(gnd), .vdd(vdd), .A(data_87__13_), .Y(_5684_) );
MUX2X1 MUX2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_5684_), .B(_14924__bF_buf3), .S(_5661_), .Y(_242__13_) );
INVX1 INVX1_2510 ( .gnd(gnd), .vdd(vdd), .A(data_87__14_), .Y(_5685_) );
MUX2X1 MUX2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_5685_), .B(_15060__bF_buf14), .S(_5661_), .Y(_242__14_) );
INVX1 INVX1_2511 ( .gnd(gnd), .vdd(vdd), .A(data_87__15_), .Y(_5686_) );
MUX2X1 MUX2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_5686_), .B(_15062__bF_buf5), .S(_5661_), .Y(_242__15_) );
INVX1 INVX1_2512 ( .gnd(gnd), .vdd(vdd), .A(data_86__0_), .Y(_5687_) );
NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_5542_), .B(_5419_), .Y(_5688_) );
INVX1 INVX1_2513 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .Y(_5689_) );
AOI21X1 AOI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_3324_), .B(_14978__bF_buf3), .C(_14882__bF_buf4), .Y(_5690_) );
OAI21X1 OAI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_4535_), .B(_3320_), .C(_5690_), .Y(_5691_) );
NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_5691_), .B(_5689_), .Y(_5692_) );
NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_5692_), .Y(_5693_) );
NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(_5693_), .B(_5688_), .Y(_5694_) );
INVX4 INVX4_19 ( .gnd(gnd), .vdd(vdd), .A(_5694_), .Y(_5695_) );
OAI21X1 OAI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_5695_), .C(_5687_), .Y(_5696_) );
NAND3X1 NAND3X1_769 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_5694_), .C(_3313__bF_buf80), .Y(_5697_) );
AND2X2 AND2X2_1106 ( .gnd(gnd), .vdd(vdd), .A(_5696_), .B(_5697_), .Y(_241__0_) );
INVX1 INVX1_2514 ( .gnd(gnd), .vdd(vdd), .A(data_86__1_), .Y(_5698_) );
OAI21X1 OAI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_5695_), .C(_5698_), .Y(_5699_) );
NAND3X1 NAND3X1_770 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_5694_), .C(_3313__bF_buf79), .Y(_5700_) );
AND2X2 AND2X2_1107 ( .gnd(gnd), .vdd(vdd), .A(_5699_), .B(_5700_), .Y(_241__1_) );
INVX1 INVX1_2515 ( .gnd(gnd), .vdd(vdd), .A(data_86__2_), .Y(_5701_) );
NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_5694_), .B(_3313__bF_buf78), .Y(_5702_) );
MUX2X1 MUX2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_5701_), .B(_14897__bF_buf9), .S(_5702_), .Y(_241__2_) );
INVX1 INVX1_2516 ( .gnd(gnd), .vdd(vdd), .A(data_86__3_), .Y(_5703_) );
OAI21X1 OAI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf20), .B(_5695_), .C(_5703_), .Y(_5704_) );
NAND3X1 NAND3X1_771 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_5694_), .C(_3313__bF_buf77), .Y(_5705_) );
AND2X2 AND2X2_1108 ( .gnd(gnd), .vdd(vdd), .A(_5704_), .B(_5705_), .Y(_241__3_) );
INVX1 INVX1_2517 ( .gnd(gnd), .vdd(vdd), .A(data_86__4_), .Y(_5706_) );
OAI21X1 OAI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_5695_), .C(_5706_), .Y(_5707_) );
NAND3X1 NAND3X1_772 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_5694_), .C(_3313__bF_buf76), .Y(_5708_) );
AND2X2 AND2X2_1109 ( .gnd(gnd), .vdd(vdd), .A(_5707_), .B(_5708_), .Y(_241__4_) );
INVX1 INVX1_2518 ( .gnd(gnd), .vdd(vdd), .A(data_86__5_), .Y(_5709_) );
OAI21X1 OAI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_5695_), .C(_5709_), .Y(_5710_) );
NAND3X1 NAND3X1_773 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_5694_), .C(_3313__bF_buf75), .Y(_5711_) );
AND2X2 AND2X2_1110 ( .gnd(gnd), .vdd(vdd), .A(_5710_), .B(_5711_), .Y(_241__5_) );
INVX1 INVX1_2519 ( .gnd(gnd), .vdd(vdd), .A(data_86__6_), .Y(_5712_) );
MUX2X1 MUX2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_5712_), .B(_15049__bF_buf11), .S(_5702_), .Y(_241__6_) );
INVX1 INVX1_2520 ( .gnd(gnd), .vdd(vdd), .A(data_86__7_), .Y(_5713_) );
OAI21X1 OAI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf17), .B(_5695_), .C(_5713_), .Y(_5714_) );
NAND3X1 NAND3X1_774 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_5694_), .C(_3313__bF_buf74), .Y(_5715_) );
AND2X2 AND2X2_1111 ( .gnd(gnd), .vdd(vdd), .A(_5714_), .B(_5715_), .Y(_241__7_) );
INVX1 INVX1_2521 ( .gnd(gnd), .vdd(vdd), .A(data_86__8_), .Y(_5716_) );
MUX2X1 MUX2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_5716_), .B(_15052__bF_buf3), .S(_5702_), .Y(_241__8_) );
INVX1 INVX1_2522 ( .gnd(gnd), .vdd(vdd), .A(data_86__9_), .Y(_5717_) );
MUX2X1 MUX2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_5717_), .B(_14913__bF_buf11), .S(_5702_), .Y(_241__9_) );
INVX1 INVX1_2523 ( .gnd(gnd), .vdd(vdd), .A(data_86__10_), .Y(_5718_) );
MUX2X1 MUX2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_5718_), .B(_15055__bF_buf5), .S(_5702_), .Y(_241__10_) );
INVX1 INVX1_2524 ( .gnd(gnd), .vdd(vdd), .A(data_86__11_), .Y(_5719_) );
OAI21X1 OAI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf16), .B(_5695_), .C(_5719_), .Y(_5720_) );
NAND3X1 NAND3X1_775 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_5694_), .C(_3313__bF_buf73), .Y(_5721_) );
AND2X2 AND2X2_1112 ( .gnd(gnd), .vdd(vdd), .A(_5720_), .B(_5721_), .Y(_241__11_) );
INVX1 INVX1_2525 ( .gnd(gnd), .vdd(vdd), .A(data_86__12_), .Y(_5722_) );
OAI21X1 OAI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf15), .B(_5695_), .C(_5722_), .Y(_5723_) );
NAND3X1 NAND3X1_776 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_5694_), .C(_3313__bF_buf72), .Y(_5724_) );
AND2X2 AND2X2_1113 ( .gnd(gnd), .vdd(vdd), .A(_5723_), .B(_5724_), .Y(_241__12_) );
INVX1 INVX1_2526 ( .gnd(gnd), .vdd(vdd), .A(data_86__13_), .Y(_5725_) );
MUX2X1 MUX2X1_884 ( .gnd(gnd), .vdd(vdd), .A(_5725_), .B(_14924__bF_buf2), .S(_5702_), .Y(_241__13_) );
INVX1 INVX1_2527 ( .gnd(gnd), .vdd(vdd), .A(data_86__14_), .Y(_5726_) );
MUX2X1 MUX2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_5726_), .B(_15060__bF_buf13), .S(_5702_), .Y(_241__14_) );
INVX1 INVX1_2528 ( .gnd(gnd), .vdd(vdd), .A(data_86__15_), .Y(_5727_) );
MUX2X1 MUX2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_5727_), .B(_15062__bF_buf4), .S(_5702_), .Y(_241__15_) );
INVX1 INVX1_2529 ( .gnd(gnd), .vdd(vdd), .A(data_85__0_), .Y(_5728_) );
OAI21X1 OAI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(IDATA_PROG_addr_3_bF_buf2), .C(_3324_), .Y(_5729_) );
AND2X2 AND2X2_1114 ( .gnd(gnd), .vdd(vdd), .A(_5503_), .B(_5729_), .Y(_5730_) );
NAND3X1 NAND3X1_777 ( .gnd(gnd), .vdd(vdd), .A(_5690_), .B(_5730_), .C(_14973_), .Y(_5731_) );
NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_5688_), .B(_5731_), .Y(_5732_) );
INVX4 INVX4_20 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .Y(_5733_) );
OAI21X1 OAI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf14), .B(_5733_), .C(_5728_), .Y(_5734_) );
NAND3X1 NAND3X1_778 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_5732_), .C(_3313__bF_buf71), .Y(_5735_) );
AND2X2 AND2X2_1115 ( .gnd(gnd), .vdd(vdd), .A(_5734_), .B(_5735_), .Y(_240__0_) );
INVX1 INVX1_2530 ( .gnd(gnd), .vdd(vdd), .A(data_85__1_), .Y(_5736_) );
OAI21X1 OAI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf13), .B(_5733_), .C(_5736_), .Y(_5737_) );
NAND3X1 NAND3X1_779 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_5732_), .C(_3313__bF_buf70), .Y(_5738_) );
AND2X2 AND2X2_1116 ( .gnd(gnd), .vdd(vdd), .A(_5737_), .B(_5738_), .Y(_240__1_) );
INVX1 INVX1_2531 ( .gnd(gnd), .vdd(vdd), .A(data_85__2_), .Y(_5739_) );
NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_5732_), .B(_3313__bF_buf69), .Y(_5740_) );
MUX2X1 MUX2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_5739_), .B(_14897__bF_buf8), .S(_5740_), .Y(_240__2_) );
INVX1 INVX1_2532 ( .gnd(gnd), .vdd(vdd), .A(data_85__3_), .Y(_5741_) );
OAI21X1 OAI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_5733_), .C(_5741_), .Y(_5742_) );
NAND3X1 NAND3X1_780 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_5732_), .C(_3313__bF_buf68), .Y(_5743_) );
AND2X2 AND2X2_1117 ( .gnd(gnd), .vdd(vdd), .A(_5742_), .B(_5743_), .Y(_240__3_) );
INVX1 INVX1_2533 ( .gnd(gnd), .vdd(vdd), .A(data_85__4_), .Y(_5744_) );
OAI21X1 OAI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_5733_), .C(_5744_), .Y(_5745_) );
NAND3X1 NAND3X1_781 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_5732_), .C(_3313__bF_buf67), .Y(_5746_) );
AND2X2 AND2X2_1118 ( .gnd(gnd), .vdd(vdd), .A(_5745_), .B(_5746_), .Y(_240__4_) );
INVX1 INVX1_2534 ( .gnd(gnd), .vdd(vdd), .A(data_85__5_), .Y(_5747_) );
OAI21X1 OAI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_5733_), .C(_5747_), .Y(_5748_) );
NAND3X1 NAND3X1_782 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_5732_), .C(_3313__bF_buf66), .Y(_5749_) );
AND2X2 AND2X2_1119 ( .gnd(gnd), .vdd(vdd), .A(_5748_), .B(_5749_), .Y(_240__5_) );
INVX1 INVX1_2535 ( .gnd(gnd), .vdd(vdd), .A(data_85__6_), .Y(_5750_) );
MUX2X1 MUX2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_5750_), .B(_15049__bF_buf10), .S(_5740_), .Y(_240__6_) );
INVX1 INVX1_2536 ( .gnd(gnd), .vdd(vdd), .A(data_85__7_), .Y(_5751_) );
OAI21X1 OAI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_5733_), .C(_5751_), .Y(_5752_) );
NAND3X1 NAND3X1_783 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_5732_), .C(_3313__bF_buf65), .Y(_5753_) );
AND2X2 AND2X2_1120 ( .gnd(gnd), .vdd(vdd), .A(_5752_), .B(_5753_), .Y(_240__7_) );
INVX1 INVX1_2537 ( .gnd(gnd), .vdd(vdd), .A(data_85__8_), .Y(_5754_) );
MUX2X1 MUX2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_5754_), .B(_15052__bF_buf2), .S(_5740_), .Y(_240__8_) );
INVX1 INVX1_2538 ( .gnd(gnd), .vdd(vdd), .A(data_85__9_), .Y(_5755_) );
MUX2X1 MUX2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_5755_), .B(_14913__bF_buf10), .S(_5740_), .Y(_240__9_) );
INVX1 INVX1_2539 ( .gnd(gnd), .vdd(vdd), .A(data_85__10_), .Y(_5756_) );
MUX2X1 MUX2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_5756_), .B(_15055__bF_buf4), .S(_5740_), .Y(_240__10_) );
INVX1 INVX1_2540 ( .gnd(gnd), .vdd(vdd), .A(data_85__11_), .Y(_5757_) );
OAI21X1 OAI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf8), .B(_5733_), .C(_5757_), .Y(_5758_) );
NAND3X1 NAND3X1_784 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_5732_), .C(_3313__bF_buf64), .Y(_5759_) );
AND2X2 AND2X2_1121 ( .gnd(gnd), .vdd(vdd), .A(_5758_), .B(_5759_), .Y(_240__11_) );
INVX1 INVX1_2541 ( .gnd(gnd), .vdd(vdd), .A(data_85__12_), .Y(_5760_) );
OAI21X1 OAI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_5733_), .C(_5760_), .Y(_5761_) );
NAND3X1 NAND3X1_785 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_5732_), .C(_3313__bF_buf63), .Y(_5762_) );
AND2X2 AND2X2_1122 ( .gnd(gnd), .vdd(vdd), .A(_5761_), .B(_5762_), .Y(_240__12_) );
INVX1 INVX1_2542 ( .gnd(gnd), .vdd(vdd), .A(data_85__13_), .Y(_5763_) );
MUX2X1 MUX2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_5763_), .B(_14924__bF_buf1), .S(_5740_), .Y(_240__13_) );
INVX1 INVX1_2543 ( .gnd(gnd), .vdd(vdd), .A(data_85__14_), .Y(_5764_) );
MUX2X1 MUX2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_5764_), .B(_15060__bF_buf12), .S(_5740_), .Y(_240__14_) );
INVX1 INVX1_2544 ( .gnd(gnd), .vdd(vdd), .A(data_85__15_), .Y(_5765_) );
MUX2X1 MUX2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_5765_), .B(_15062__bF_buf3), .S(_5740_), .Y(_240__15_) );
INVX1 INVX1_2545 ( .gnd(gnd), .vdd(vdd), .A(data_84__0_), .Y(_5766_) );
OAI21X1 OAI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_3320_), .C(_5542_), .Y(_5767_) );
OAI21X1 OAI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .B(_5566_), .C(_5503_), .Y(_5768_) );
NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_5768_), .B(_5767_), .Y(_5769_) );
NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5769_), .Y(_5770_) );
OAI21X1 OAI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_5770_), .C(_5766_), .Y(_5771_) );
NOR3X1 NOR3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_5767_), .B(_5768_), .C(_5420__bF_buf2), .Y(_5772_) );
NAND3X1 NAND3X1_786 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_5772_), .C(_3313__bF_buf62), .Y(_5773_) );
AND2X2 AND2X2_1123 ( .gnd(gnd), .vdd(vdd), .A(_5771_), .B(_5773_), .Y(_239__0_) );
INVX1 INVX1_2546 ( .gnd(gnd), .vdd(vdd), .A(data_84__1_), .Y(_5774_) );
OAI21X1 OAI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_5770_), .C(_5774_), .Y(_5775_) );
NAND3X1 NAND3X1_787 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_5772_), .C(_3313__bF_buf61), .Y(_5776_) );
AND2X2 AND2X2_1124 ( .gnd(gnd), .vdd(vdd), .A(_5775_), .B(_5776_), .Y(_239__1_) );
INVX1 INVX1_2547 ( .gnd(gnd), .vdd(vdd), .A(data_84__2_), .Y(_5777_) );
NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_5772_), .B(_3313__bF_buf60), .Y(_5778_) );
MUX2X1 MUX2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_5777_), .B(_14897__bF_buf7), .S(_5778_), .Y(_239__2_) );
INVX1 INVX1_2548 ( .gnd(gnd), .vdd(vdd), .A(data_84__3_), .Y(_5779_) );
OAI21X1 OAI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_5770_), .C(_5779_), .Y(_5780_) );
NAND3X1 NAND3X1_788 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_5772_), .C(_3313__bF_buf59), .Y(_5781_) );
AND2X2 AND2X2_1125 ( .gnd(gnd), .vdd(vdd), .A(_5780_), .B(_5781_), .Y(_239__3_) );
INVX1 INVX1_2549 ( .gnd(gnd), .vdd(vdd), .A(data_84__4_), .Y(_5782_) );
OAI21X1 OAI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf3), .B(_5770_), .C(_5782_), .Y(_5783_) );
NAND3X1 NAND3X1_789 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_5772_), .C(_3313__bF_buf58), .Y(_5784_) );
AND2X2 AND2X2_1126 ( .gnd(gnd), .vdd(vdd), .A(_5783_), .B(_5784_), .Y(_239__4_) );
INVX1 INVX1_2550 ( .gnd(gnd), .vdd(vdd), .A(data_84__5_), .Y(_5785_) );
OAI21X1 OAI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_5770_), .C(_5785_), .Y(_5786_) );
NAND3X1 NAND3X1_790 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_5772_), .C(_3313__bF_buf57), .Y(_5787_) );
AND2X2 AND2X2_1127 ( .gnd(gnd), .vdd(vdd), .A(_5786_), .B(_5787_), .Y(_239__5_) );
INVX1 INVX1_2551 ( .gnd(gnd), .vdd(vdd), .A(data_84__6_), .Y(_5788_) );
MUX2X1 MUX2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_5788_), .B(_15049__bF_buf9), .S(_5778_), .Y(_239__6_) );
INVX1 INVX1_2552 ( .gnd(gnd), .vdd(vdd), .A(data_84__7_), .Y(_5789_) );
OAI21X1 OAI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_5770_), .C(_5789_), .Y(_5790_) );
NAND3X1 NAND3X1_791 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_5772_), .C(_3313__bF_buf56), .Y(_5791_) );
AND2X2 AND2X2_1128 ( .gnd(gnd), .vdd(vdd), .A(_5790_), .B(_5791_), .Y(_239__7_) );
INVX1 INVX1_2553 ( .gnd(gnd), .vdd(vdd), .A(data_84__8_), .Y(_5792_) );
MUX2X1 MUX2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_5792_), .B(_15052__bF_buf1), .S(_5778_), .Y(_239__8_) );
INVX1 INVX1_2554 ( .gnd(gnd), .vdd(vdd), .A(data_84__9_), .Y(_5793_) );
MUX2X1 MUX2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_5793_), .B(_14913__bF_buf9), .S(_5778_), .Y(_239__9_) );
INVX1 INVX1_2555 ( .gnd(gnd), .vdd(vdd), .A(data_84__10_), .Y(_5794_) );
MUX2X1 MUX2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_5794_), .B(_15055__bF_buf3), .S(_5778_), .Y(_239__10_) );
INVX1 INVX1_2556 ( .gnd(gnd), .vdd(vdd), .A(data_84__11_), .Y(_5795_) );
OAI21X1 OAI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_5770_), .C(_5795_), .Y(_5796_) );
NAND3X1 NAND3X1_792 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_5772_), .C(_3313__bF_buf55), .Y(_5797_) );
AND2X2 AND2X2_1129 ( .gnd(gnd), .vdd(vdd), .A(_5796_), .B(_5797_), .Y(_239__11_) );
INVX1 INVX1_2557 ( .gnd(gnd), .vdd(vdd), .A(data_84__12_), .Y(_5798_) );
OAI21X1 OAI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_5770_), .C(_5798_), .Y(_5799_) );
NAND3X1 NAND3X1_793 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_5772_), .C(_3313__bF_buf54), .Y(_5800_) );
AND2X2 AND2X2_1130 ( .gnd(gnd), .vdd(vdd), .A(_5799_), .B(_5800_), .Y(_239__12_) );
INVX1 INVX1_2558 ( .gnd(gnd), .vdd(vdd), .A(data_84__13_), .Y(_5801_) );
MUX2X1 MUX2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_5801_), .B(_14924__bF_buf0), .S(_5778_), .Y(_239__13_) );
INVX1 INVX1_2559 ( .gnd(gnd), .vdd(vdd), .A(data_84__14_), .Y(_5802_) );
MUX2X1 MUX2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_5802_), .B(_15060__bF_buf11), .S(_5778_), .Y(_239__14_) );
INVX1 INVX1_2560 ( .gnd(gnd), .vdd(vdd), .A(data_84__15_), .Y(_5803_) );
MUX2X1 MUX2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_5803_), .B(_15062__bF_buf2), .S(_5778_), .Y(_239__15_) );
INVX1 INVX1_2561 ( .gnd(gnd), .vdd(vdd), .A(data_83__0_), .Y(_5804_) );
NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf3), .B(_3326_), .Y(_5805_) );
OAI21X1 OAI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_15171_), .B(_3320_), .C(_5805_), .Y(_5806_) );
AOI21X1 AOI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_14974_), .B(_3324_), .C(_5806_), .Y(_5807_) );
NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_5807_), .Y(_5808_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_5808_), .B(_5688_), .Y(_5809_) );
OAI21X1 OAI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_5809_), .C(_5804_), .Y(_5810_) );
NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_5688_), .B(_5808_), .Y(_5811_) );
NAND3X1 NAND3X1_794 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_5811_), .C(_3313__bF_buf53), .Y(_5812_) );
AND2X2 AND2X2_1131 ( .gnd(gnd), .vdd(vdd), .A(_5810_), .B(_5812_), .Y(_238__0_) );
INVX1 INVX1_2562 ( .gnd(gnd), .vdd(vdd), .A(data_83__1_), .Y(_5813_) );
OAI21X1 OAI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_5809_), .C(_5813_), .Y(_5814_) );
NAND3X1 NAND3X1_795 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_5811_), .C(_3313__bF_buf52), .Y(_5815_) );
AND2X2 AND2X2_1132 ( .gnd(gnd), .vdd(vdd), .A(_5814_), .B(_5815_), .Y(_238__1_) );
NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_5809_), .B(_3393__bF_buf66), .Y(_5816_) );
AOI21X1 AOI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_3313__bF_buf51), .C(data_83__2_), .Y(_5817_) );
AOI21X1 AOI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_5816_), .C(_5817_), .Y(_238__2_) );
INVX1 INVX1_2563 ( .gnd(gnd), .vdd(vdd), .A(data_83__3_), .Y(_5818_) );
OAI21X1 OAI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_5809_), .C(_5818_), .Y(_5819_) );
NAND3X1 NAND3X1_796 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_5811_), .C(_3313__bF_buf50), .Y(_5820_) );
AND2X2 AND2X2_1133 ( .gnd(gnd), .vdd(vdd), .A(_5819_), .B(_5820_), .Y(_238__3_) );
INVX1 INVX1_2564 ( .gnd(gnd), .vdd(vdd), .A(data_83__4_), .Y(_5821_) );
OAI21X1 OAI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_5809_), .C(_5821_), .Y(_5822_) );
NAND3X1 NAND3X1_797 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_5811_), .C(_3313__bF_buf49), .Y(_5823_) );
AND2X2 AND2X2_1134 ( .gnd(gnd), .vdd(vdd), .A(_5822_), .B(_5823_), .Y(_238__4_) );
INVX1 INVX1_2565 ( .gnd(gnd), .vdd(vdd), .A(data_83__5_), .Y(_5824_) );
OAI21X1 OAI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_5809_), .C(_5824_), .Y(_5825_) );
NAND3X1 NAND3X1_798 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_5811_), .C(_3313__bF_buf48), .Y(_5826_) );
AND2X2 AND2X2_1135 ( .gnd(gnd), .vdd(vdd), .A(_5825_), .B(_5826_), .Y(_238__5_) );
AOI21X1 AOI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_3313__bF_buf47), .C(data_83__6_), .Y(_5827_) );
AOI21X1 AOI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_5816_), .C(_5827_), .Y(_238__6_) );
INVX1 INVX1_2566 ( .gnd(gnd), .vdd(vdd), .A(data_83__7_), .Y(_5828_) );
OAI21X1 OAI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_5809_), .C(_5828_), .Y(_5829_) );
NAND3X1 NAND3X1_799 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_5811_), .C(_3313__bF_buf46), .Y(_5830_) );
AND2X2 AND2X2_1136 ( .gnd(gnd), .vdd(vdd), .A(_5829_), .B(_5830_), .Y(_238__7_) );
AOI21X1 AOI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_3313__bF_buf45), .C(data_83__8_), .Y(_5831_) );
AOI21X1 AOI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_5816_), .C(_5831_), .Y(_238__8_) );
INVX1 INVX1_2567 ( .gnd(gnd), .vdd(vdd), .A(data_83__9_), .Y(_5832_) );
NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_3313__bF_buf44), .Y(_5833_) );
MUX2X1 MUX2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_5832_), .B(_14913__bF_buf8), .S(_5833_), .Y(_238__9_) );
INVX1 INVX1_2568 ( .gnd(gnd), .vdd(vdd), .A(data_83__10_), .Y(_5834_) );
MUX2X1 MUX2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_5834_), .B(_15055__bF_buf2), .S(_5833_), .Y(_238__10_) );
INVX1 INVX1_2569 ( .gnd(gnd), .vdd(vdd), .A(data_83__11_), .Y(_5835_) );
OAI21X1 OAI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_5809_), .C(_5835_), .Y(_5836_) );
NAND3X1 NAND3X1_800 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_5811_), .C(_3313__bF_buf43), .Y(_5837_) );
AND2X2 AND2X2_1137 ( .gnd(gnd), .vdd(vdd), .A(_5836_), .B(_5837_), .Y(_238__11_) );
INVX1 INVX1_2570 ( .gnd(gnd), .vdd(vdd), .A(data_83__12_), .Y(_5838_) );
OAI21X1 OAI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_5809_), .C(_5838_), .Y(_5839_) );
NAND3X1 NAND3X1_801 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_5811_), .C(_3313__bF_buf42), .Y(_5840_) );
AND2X2 AND2X2_1138 ( .gnd(gnd), .vdd(vdd), .A(_5839_), .B(_5840_), .Y(_238__12_) );
AOI21X1 AOI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_5811_), .B(_3313__bF_buf41), .C(data_83__13_), .Y(_5841_) );
AOI21X1 AOI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_5816_), .C(_5841_), .Y(_238__13_) );
INVX1 INVX1_2571 ( .gnd(gnd), .vdd(vdd), .A(data_83__14_), .Y(_5842_) );
MUX2X1 MUX2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_5842_), .B(_15060__bF_buf10), .S(_5833_), .Y(_238__14_) );
INVX1 INVX1_2572 ( .gnd(gnd), .vdd(vdd), .A(data_83__15_), .Y(_5843_) );
MUX2X1 MUX2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_5843_), .B(_15062__bF_buf1), .S(_5833_), .Y(_238__15_) );
INVX1 INVX1_2573 ( .gnd(gnd), .vdd(vdd), .A(data_82__0_), .Y(_5844_) );
OAI21X1 OAI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_3320_), .B(_4683_), .C(_5805_), .Y(_5845_) );
NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_5845_), .B(_5767_), .Y(_5846_) );
NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5846_), .Y(_5847_) );
OAI21X1 OAI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_5847_), .C(_5844_), .Y(_5848_) );
NOR3X1 NOR3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_5767_), .B(_5845_), .C(_5420__bF_buf1), .Y(_5849_) );
NAND3X1 NAND3X1_802 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_5849_), .C(_3313__bF_buf40), .Y(_5850_) );
AND2X2 AND2X2_1139 ( .gnd(gnd), .vdd(vdd), .A(_5848_), .B(_5850_), .Y(_237__0_) );
INVX1 INVX1_2574 ( .gnd(gnd), .vdd(vdd), .A(data_82__1_), .Y(_5851_) );
OAI21X1 OAI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_5847_), .C(_5851_), .Y(_5852_) );
NAND3X1 NAND3X1_803 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_5849_), .C(_3313__bF_buf39), .Y(_5853_) );
AND2X2 AND2X2_1140 ( .gnd(gnd), .vdd(vdd), .A(_5852_), .B(_5853_), .Y(_237__1_) );
INVX1 INVX1_2575 ( .gnd(gnd), .vdd(vdd), .A(data_82__2_), .Y(_5854_) );
NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .B(_3313__bF_buf38), .Y(_5855_) );
MUX2X1 MUX2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_5854_), .B(_14897__bF_buf5), .S(_5855_), .Y(_237__2_) );
INVX1 INVX1_2576 ( .gnd(gnd), .vdd(vdd), .A(data_82__3_), .Y(_5856_) );
OAI21X1 OAI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_5847_), .C(_5856_), .Y(_5857_) );
NAND3X1 NAND3X1_804 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_5849_), .C(_3313__bF_buf37), .Y(_5858_) );
AND2X2 AND2X2_1141 ( .gnd(gnd), .vdd(vdd), .A(_5857_), .B(_5858_), .Y(_237__3_) );
INVX1 INVX1_2577 ( .gnd(gnd), .vdd(vdd), .A(data_82__4_), .Y(_5859_) );
OAI21X1 OAI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_5847_), .C(_5859_), .Y(_5860_) );
NAND3X1 NAND3X1_805 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_5849_), .C(_3313__bF_buf36), .Y(_5861_) );
AND2X2 AND2X2_1142 ( .gnd(gnd), .vdd(vdd), .A(_5860_), .B(_5861_), .Y(_237__4_) );
NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_5847_), .B(_3393__bF_buf55), .Y(_5862_) );
AOI21X1 AOI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .B(_3313__bF_buf35), .C(data_82__5_), .Y(_5863_) );
AOI21X1 AOI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_5862_), .C(_5863_), .Y(_237__5_) );
INVX1 INVX1_2578 ( .gnd(gnd), .vdd(vdd), .A(data_82__6_), .Y(_5864_) );
MUX2X1 MUX2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_5864_), .B(_15049__bF_buf7), .S(_5855_), .Y(_237__6_) );
INVX1 INVX1_2579 ( .gnd(gnd), .vdd(vdd), .A(data_82__7_), .Y(_5865_) );
OAI21X1 OAI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_5847_), .C(_5865_), .Y(_5866_) );
NAND3X1 NAND3X1_806 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_5849_), .C(_3313__bF_buf34), .Y(_5867_) );
AND2X2 AND2X2_1143 ( .gnd(gnd), .vdd(vdd), .A(_5866_), .B(_5867_), .Y(_237__7_) );
INVX1 INVX1_2580 ( .gnd(gnd), .vdd(vdd), .A(data_82__8_), .Y(_5868_) );
MUX2X1 MUX2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_5868_), .B(_15052__bF_buf13), .S(_5855_), .Y(_237__8_) );
INVX1 INVX1_2581 ( .gnd(gnd), .vdd(vdd), .A(data_82__9_), .Y(_5869_) );
MUX2X1 MUX2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_5869_), .B(_14913__bF_buf7), .S(_5855_), .Y(_237__9_) );
INVX1 INVX1_2582 ( .gnd(gnd), .vdd(vdd), .A(data_82__10_), .Y(_5870_) );
MUX2X1 MUX2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_5870_), .B(_15055__bF_buf1), .S(_5855_), .Y(_237__10_) );
INVX1 INVX1_2583 ( .gnd(gnd), .vdd(vdd), .A(data_82__11_), .Y(_5871_) );
OAI21X1 OAI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_5847_), .C(_5871_), .Y(_5872_) );
NAND3X1 NAND3X1_807 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_5849_), .C(_3313__bF_buf33), .Y(_5873_) );
AND2X2 AND2X2_1144 ( .gnd(gnd), .vdd(vdd), .A(_5872_), .B(_5873_), .Y(_237__11_) );
AOI21X1 AOI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .B(_3313__bF_buf32), .C(data_82__12_), .Y(_5874_) );
AOI21X1 AOI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_5862_), .C(_5874_), .Y(_237__12_) );
AOI21X1 AOI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_5849_), .B(_3313__bF_buf31), .C(data_82__13_), .Y(_5875_) );
AOI21X1 AOI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_5862_), .C(_5875_), .Y(_237__13_) );
INVX1 INVX1_2584 ( .gnd(gnd), .vdd(vdd), .A(data_82__14_), .Y(_5876_) );
MUX2X1 MUX2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_5876_), .B(_15060__bF_buf9), .S(_5855_), .Y(_237__14_) );
INVX1 INVX1_2585 ( .gnd(gnd), .vdd(vdd), .A(data_82__15_), .Y(_5877_) );
MUX2X1 MUX2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_5877_), .B(_15062__bF_buf0), .S(_5855_), .Y(_237__15_) );
INVX1 INVX1_2586 ( .gnd(gnd), .vdd(vdd), .A(data_81__0_), .Y(_5878_) );
OAI21X1 OAI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_3320_), .B(_4722_), .C(_5805_), .Y(_5879_) );
NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_5879_), .B(_5767_), .Y(_5880_) );
NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5880_), .Y(_5881_) );
OAI21X1 OAI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_5881_), .C(_5878_), .Y(_5882_) );
NOR3X1 NOR3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_5767_), .B(_5879_), .C(_5420__bF_buf0), .Y(_5883_) );
NAND3X1 NAND3X1_808 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_5883_), .C(_3313__bF_buf30), .Y(_5884_) );
AND2X2 AND2X2_1145 ( .gnd(gnd), .vdd(vdd), .A(_5882_), .B(_5884_), .Y(_236__0_) );
INVX1 INVX1_2587 ( .gnd(gnd), .vdd(vdd), .A(data_81__1_), .Y(_5885_) );
OAI21X1 OAI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_5881_), .C(_5885_), .Y(_5886_) );
NAND3X1 NAND3X1_809 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_5883_), .C(_3313__bF_buf29), .Y(_5887_) );
AND2X2 AND2X2_1146 ( .gnd(gnd), .vdd(vdd), .A(_5886_), .B(_5887_), .Y(_236__1_) );
INVX1 INVX1_2588 ( .gnd(gnd), .vdd(vdd), .A(data_81__2_), .Y(_5888_) );
NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_5883_), .B(_3313__bF_buf28), .Y(_5889_) );
MUX2X1 MUX2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_5888_), .B(_14897__bF_buf4), .S(_5889_), .Y(_236__2_) );
INVX1 INVX1_2589 ( .gnd(gnd), .vdd(vdd), .A(data_81__3_), .Y(_5890_) );
OAI21X1 OAI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_5881_), .C(_5890_), .Y(_5891_) );
NAND3X1 NAND3X1_810 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_5883_), .C(_3313__bF_buf27), .Y(_5892_) );
AND2X2 AND2X2_1147 ( .gnd(gnd), .vdd(vdd), .A(_5891_), .B(_5892_), .Y(_236__3_) );
INVX1 INVX1_2590 ( .gnd(gnd), .vdd(vdd), .A(data_81__4_), .Y(_5893_) );
OAI21X1 OAI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_5881_), .C(_5893_), .Y(_5894_) );
NAND3X1 NAND3X1_811 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_5883_), .C(_3313__bF_buf26), .Y(_5895_) );
AND2X2 AND2X2_1148 ( .gnd(gnd), .vdd(vdd), .A(_5894_), .B(_5895_), .Y(_236__4_) );
INVX1 INVX1_2591 ( .gnd(gnd), .vdd(vdd), .A(data_81__5_), .Y(_5896_) );
MUX2X1 MUX2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_5896_), .B(_14903__bF_buf12), .S(_5889_), .Y(_236__5_) );
INVX1 INVX1_2592 ( .gnd(gnd), .vdd(vdd), .A(data_81__6_), .Y(_5897_) );
MUX2X1 MUX2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_5897_), .B(_15049__bF_buf6), .S(_5889_), .Y(_236__6_) );
INVX1 INVX1_2593 ( .gnd(gnd), .vdd(vdd), .A(data_81__7_), .Y(_5898_) );
OAI21X1 OAI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_5881_), .C(_5898_), .Y(_5899_) );
NAND3X1 NAND3X1_812 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_5883_), .C(_3313__bF_buf25), .Y(_5900_) );
AND2X2 AND2X2_1149 ( .gnd(gnd), .vdd(vdd), .A(_5899_), .B(_5900_), .Y(_236__7_) );
INVX1 INVX1_2594 ( .gnd(gnd), .vdd(vdd), .A(data_81__8_), .Y(_5901_) );
MUX2X1 MUX2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_5901_), .B(_15052__bF_buf12), .S(_5889_), .Y(_236__8_) );
INVX1 INVX1_2595 ( .gnd(gnd), .vdd(vdd), .A(data_81__9_), .Y(_5902_) );
MUX2X1 MUX2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_5902_), .B(_14913__bF_buf6), .S(_5889_), .Y(_236__9_) );
INVX1 INVX1_2596 ( .gnd(gnd), .vdd(vdd), .A(data_81__10_), .Y(_5903_) );
MUX2X1 MUX2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_5903_), .B(_15055__bF_buf0), .S(_5889_), .Y(_236__10_) );
INVX1 INVX1_2597 ( .gnd(gnd), .vdd(vdd), .A(data_81__11_), .Y(_5904_) );
OAI21X1 OAI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_5881_), .C(_5904_), .Y(_5905_) );
NAND3X1 NAND3X1_813 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_5883_), .C(_3313__bF_buf24), .Y(_5906_) );
AND2X2 AND2X2_1150 ( .gnd(gnd), .vdd(vdd), .A(_5905_), .B(_5906_), .Y(_236__11_) );
INVX1 INVX1_2598 ( .gnd(gnd), .vdd(vdd), .A(data_81__12_), .Y(_5907_) );
MUX2X1 MUX2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_5907_), .B(_14920__bF_buf1), .S(_5889_), .Y(_236__12_) );
INVX1 INVX1_2599 ( .gnd(gnd), .vdd(vdd), .A(data_81__13_), .Y(_5908_) );
MUX2X1 MUX2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_5908_), .B(_14924__bF_buf11), .S(_5889_), .Y(_236__13_) );
INVX1 INVX1_2600 ( .gnd(gnd), .vdd(vdd), .A(data_81__14_), .Y(_5909_) );
MUX2X1 MUX2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_5909_), .B(_15060__bF_buf8), .S(_5889_), .Y(_236__14_) );
INVX1 INVX1_2601 ( .gnd(gnd), .vdd(vdd), .A(data_81__15_), .Y(_5910_) );
MUX2X1 MUX2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_5910_), .B(_15062__bF_buf13), .S(_5889_), .Y(_236__15_) );
NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf2), .B(_3325_), .Y(_5911_) );
NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(data_80__0_), .B(_5911__bF_buf3), .Y(_5912_) );
AOI21X1 AOI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_5911__bF_buf2), .C(_5912_), .Y(_235__0_) );
NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf3), .B(_4272_), .Y(_5913_) );
INVX1 INVX1_2602 ( .gnd(gnd), .vdd(vdd), .A(data_80__1_), .Y(_5914_) );
OAI21X1 OAI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_14882__bF_buf1), .C(_5914_), .Y(_5915_) );
OAI21X1 OAI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(IDATA_PROG_data_1_bF_buf1), .C(_5915_), .Y(_5916_) );
INVX1 INVX1_2603 ( .gnd(gnd), .vdd(vdd), .A(_5916_), .Y(_235__1_) );
NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(data_80__2_), .B(_5911__bF_buf1), .Y(_5917_) );
AOI21X1 AOI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_5911__bF_buf0), .C(_5917_), .Y(_235__2_) );
INVX1 INVX1_2604 ( .gnd(gnd), .vdd(vdd), .A(data_80__3_), .Y(_5918_) );
OAI21X1 OAI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_14882__bF_buf0), .C(_5918_), .Y(_5919_) );
OAI21X1 OAI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(IDATA_PROG_data_3_bF_buf2), .C(_5919_), .Y(_5920_) );
INVX1 INVX1_2605 ( .gnd(gnd), .vdd(vdd), .A(_5920_), .Y(_235__3_) );
NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(data_80__4_), .B(_5911__bF_buf3), .Y(_5921_) );
AOI21X1 AOI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_5911__bF_buf2), .C(_5921_), .Y(_235__4_) );
INVX1 INVX1_2606 ( .gnd(gnd), .vdd(vdd), .A(data_80__5_), .Y(_5922_) );
OAI21X1 OAI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_14882__bF_buf15_bF_buf1), .C(_5922_), .Y(_5923_) );
OAI21X1 OAI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(IDATA_PROG_data_5_bF_buf4), .C(_5923_), .Y(_5924_) );
INVX1 INVX1_2607 ( .gnd(gnd), .vdd(vdd), .A(_5924_), .Y(_235__5_) );
NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(data_80__6_), .B(_5911__bF_buf1), .Y(_5925_) );
AOI21X1 AOI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_5911__bF_buf0), .C(_5925_), .Y(_235__6_) );
NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(data_80__7_), .B(_5911__bF_buf3), .Y(_5926_) );
AOI21X1 AOI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_5911__bF_buf2), .C(_5926_), .Y(_235__7_) );
NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(data_80__8_), .B(_5911__bF_buf1), .Y(_5927_) );
AOI21X1 AOI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_5911__bF_buf0), .C(_5927_), .Y(_235__8_) );
NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(data_80__9_), .B(_5911__bF_buf3), .Y(_5928_) );
AOI21X1 AOI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_5911__bF_buf2), .C(_5928_), .Y(_235__9_) );
NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_5911__bF_buf1), .Y(_5929_) );
OAI21X1 OAI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(data_80__10_), .B(_5911__bF_buf0), .C(_5929_), .Y(_5930_) );
INVX1 INVX1_2608 ( .gnd(gnd), .vdd(vdd), .A(_5930_), .Y(_235__10_) );
INVX1 INVX1_2609 ( .gnd(gnd), .vdd(vdd), .A(data_80__11_), .Y(_5931_) );
OAI21X1 OAI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_14882__bF_buf14_bF_buf1), .C(_5931_), .Y(_5932_) );
OAI21X1 OAI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(IDATA_PROG_data_11_bF_buf3), .C(_5932_), .Y(_5933_) );
INVX1 INVX1_2610 ( .gnd(gnd), .vdd(vdd), .A(_5933_), .Y(_235__11_) );
NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(data_80__12_), .B(_5911__bF_buf3), .Y(_5934_) );
AOI21X1 AOI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_5911__bF_buf2), .C(_5934_), .Y(_235__12_) );
NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(data_80__13_), .B(_5911__bF_buf1), .Y(_5935_) );
NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf0), .B(_5913_), .Y(_5936_) );
NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_5935_), .B(_5936_), .Y(_235__13_) );
NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(data_80__14_), .B(_5911__bF_buf0), .Y(_5937_) );
AOI21X1 AOI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_5911__bF_buf3), .C(_5937_), .Y(_235__14_) );
INVX1 INVX1_2611 ( .gnd(gnd), .vdd(vdd), .A(data_80__15_), .Y(_5938_) );
OAI21X1 OAI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_14882__bF_buf13_bF_buf1), .C(_5938_), .Y(_5939_) );
OAI21X1 OAI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_5913_), .B(IDATA_PROG_data_15_bF_buf2), .C(_5939_), .Y(_5940_) );
INVX1 INVX1_2612 ( .gnd(gnd), .vdd(vdd), .A(_5940_), .Y(_235__15_) );
INVX1 INVX1_2613 ( .gnd(gnd), .vdd(vdd), .A(data_79__0_), .Y(_5941_) );
NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf3), .B(_3332_), .Y(_5942_) );
OAI21X1 OAI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf12), .C(_5941_), .Y(_5943_) );
NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf11), .B(_5942_), .Y(_5944_) );
NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_5944__bF_buf3), .Y(_5945_) );
AND2X2 AND2X2_1151 ( .gnd(gnd), .vdd(vdd), .A(_5945_), .B(_5943_), .Y(_233__0_) );
NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_4271_), .Y(_5946_) );
INVX1 INVX1_2614 ( .gnd(gnd), .vdd(vdd), .A(data_79__1_), .Y(_5947_) );
OAI21X1 OAI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf10), .C(_5947_), .Y(_5948_) );
OAI21X1 OAI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_5946_), .B(IDATA_PROG_data_1_bF_buf0), .C(_5948_), .Y(_5949_) );
INVX1 INVX1_2615 ( .gnd(gnd), .vdd(vdd), .A(_5949_), .Y(_233__1_) );
NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(data_79__2_), .B(_5944__bF_buf2), .Y(_5950_) );
AOI21X1 AOI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_5944__bF_buf1), .C(_5950_), .Y(_233__2_) );
INVX1 INVX1_2616 ( .gnd(gnd), .vdd(vdd), .A(data_79__3_), .Y(_5951_) );
OAI21X1 OAI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf9), .C(_5951_), .Y(_5952_) );
OAI21X1 OAI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_5946_), .B(IDATA_PROG_data_3_bF_buf1), .C(_5952_), .Y(_5953_) );
INVX1 INVX1_2617 ( .gnd(gnd), .vdd(vdd), .A(_5953_), .Y(_233__3_) );
INVX1 INVX1_2618 ( .gnd(gnd), .vdd(vdd), .A(data_79__4_), .Y(_5954_) );
OAI21X1 OAI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf8), .C(_5954_), .Y(_5955_) );
NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_5944__bF_buf0), .Y(_5956_) );
AND2X2 AND2X2_1152 ( .gnd(gnd), .vdd(vdd), .A(_5956_), .B(_5955_), .Y(_233__4_) );
INVX1 INVX1_2619 ( .gnd(gnd), .vdd(vdd), .A(data_79__5_), .Y(_5957_) );
OAI21X1 OAI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf7), .C(_5957_), .Y(_5958_) );
OAI21X1 OAI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_5946_), .B(IDATA_PROG_data_5_bF_buf3), .C(_5958_), .Y(_5959_) );
INVX1 INVX1_2620 ( .gnd(gnd), .vdd(vdd), .A(_5959_), .Y(_233__5_) );
INVX1 INVX1_2621 ( .gnd(gnd), .vdd(vdd), .A(data_79__6_), .Y(_5960_) );
OAI21X1 OAI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf6), .C(_5960_), .Y(_5961_) );
NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_5944__bF_buf3), .Y(_5962_) );
AND2X2 AND2X2_1153 ( .gnd(gnd), .vdd(vdd), .A(_5962_), .B(_5961_), .Y(_233__6_) );
NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(data_79__7_), .B(_5944__bF_buf2), .Y(_5963_) );
AOI21X1 AOI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_5944__bF_buf1), .C(_5963_), .Y(_233__7_) );
INVX1 INVX1_2622 ( .gnd(gnd), .vdd(vdd), .A(data_79__8_), .Y(_5964_) );
OAI21X1 OAI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf5), .C(_5964_), .Y(_5965_) );
NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_5944__bF_buf0), .Y(_5966_) );
AND2X2 AND2X2_1154 ( .gnd(gnd), .vdd(vdd), .A(_5966_), .B(_5965_), .Y(_233__8_) );
MUX2X1 MUX2X1_924 ( .gnd(gnd), .vdd(vdd), .A(data_79__9_), .B(IDATA_PROG_data_9_bF_buf2), .S(_5946_), .Y(_5967_) );
INVX1 INVX1_2623 ( .gnd(gnd), .vdd(vdd), .A(_5967_), .Y(_233__9_) );
NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(data_79__10_), .B(_5944__bF_buf3), .Y(_5968_) );
AOI21X1 AOI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_5944__bF_buf2), .C(_5968_), .Y(_233__10_) );
NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(data_79__11_), .B(_5944__bF_buf1), .Y(_5969_) );
AOI21X1 AOI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_5944__bF_buf0), .C(_5969_), .Y(_233__11_) );
INVX1 INVX1_2624 ( .gnd(gnd), .vdd(vdd), .A(data_79__12_), .Y(_5970_) );
OAI21X1 OAI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_5942_), .B(_14882__bF_buf4), .C(_5970_), .Y(_5971_) );
NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_5944__bF_buf3), .Y(_5972_) );
AND2X2 AND2X2_1155 ( .gnd(gnd), .vdd(vdd), .A(_5972_), .B(_5971_), .Y(_233__12_) );
NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_5944__bF_buf2), .Y(_5973_) );
OAI21X1 OAI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(data_79__13_), .B(_5944__bF_buf1), .C(_5973_), .Y(_5974_) );
INVX1 INVX1_2625 ( .gnd(gnd), .vdd(vdd), .A(_5974_), .Y(_233__13_) );
NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(data_79__14_), .B(_5944__bF_buf0), .Y(_5975_) );
AOI21X1 AOI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_5944__bF_buf3), .C(_5975_), .Y(_233__14_) );
NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(data_79__15_), .B(_5944__bF_buf2), .Y(_5976_) );
AOI21X1 AOI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_5944__bF_buf1), .C(_5976_), .Y(_233__15_) );
INVX1 INVX1_2626 ( .gnd(gnd), .vdd(vdd), .A(data_78__0_), .Y(_5977_) );
OAI21X1 OAI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_4244_), .C(_3332_), .Y(_5978_) );
NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_14964_), .Y(_5979_) );
NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_5421_), .B(_5979_), .Y(_5980_) );
NAND3X1 NAND3X1_814 ( .gnd(gnd), .vdd(vdd), .A(_5978_), .B(_5980_), .C(_3335_), .Y(_5981_) );
NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_5981_), .B(_5420__bF_buf3), .Y(_5982_) );
NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf23), .Y(_5983_) );
MUX2X1 MUX2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_5977_), .B(_14932__bF_buf6), .S(_5983_), .Y(_232__0_) );
INVX1 INVX1_2627 ( .gnd(gnd), .vdd(vdd), .A(data_78__1_), .Y(_5984_) );
MUX2X1 MUX2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_5984_), .B(_14894__bF_buf6), .S(_5983_), .Y(_232__1_) );
AND2X2 AND2X2_1156 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf22), .B(_5982_), .Y(_5985_) );
AOI21X1 AOI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf21), .C(data_78__2_), .Y(_5986_) );
AOI21X1 AOI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_5985_), .C(_5986_), .Y(_232__2_) );
INVX1 INVX1_2628 ( .gnd(gnd), .vdd(vdd), .A(data_78__3_), .Y(_5987_) );
MUX2X1 MUX2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_5987_), .B(_14899__bF_buf5), .S(_5983_), .Y(_232__3_) );
INVX1 INVX1_2629 ( .gnd(gnd), .vdd(vdd), .A(data_78__4_), .Y(_5988_) );
MUX2X1 MUX2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_5988_), .B(_14902__bF_buf9), .S(_5983_), .Y(_232__4_) );
INVX1 INVX1_2630 ( .gnd(gnd), .vdd(vdd), .A(data_78__5_), .Y(_5989_) );
MUX2X1 MUX2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_5989_), .B(_14903__bF_buf11), .S(_5983_), .Y(_232__5_) );
AOI21X1 AOI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf20), .C(data_78__6_), .Y(_5990_) );
AOI21X1 AOI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_5985_), .C(_5990_), .Y(_232__6_) );
INVX1 INVX1_2631 ( .gnd(gnd), .vdd(vdd), .A(data_78__7_), .Y(_5991_) );
MUX2X1 MUX2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_5991_), .B(_14908__bF_buf11), .S(_5983_), .Y(_232__7_) );
AOI21X1 AOI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf19), .C(data_78__8_), .Y(_5992_) );
AOI21X1 AOI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_5985_), .C(_5992_), .Y(_232__8_) );
AOI21X1 AOI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf18), .C(data_78__9_), .Y(_5993_) );
AOI21X1 AOI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_5985_), .C(_5993_), .Y(_232__9_) );
AOI21X1 AOI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf17), .C(data_78__10_), .Y(_5994_) );
AOI21X1 AOI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_5985_), .C(_5994_), .Y(_232__10_) );
INVX1 INVX1_2632 ( .gnd(gnd), .vdd(vdd), .A(data_78__11_), .Y(_5995_) );
MUX2X1 MUX2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_5995_), .B(_14918__bF_buf11), .S(_5983_), .Y(_232__11_) );
INVX1 INVX1_2633 ( .gnd(gnd), .vdd(vdd), .A(data_78__12_), .Y(_5996_) );
MUX2X1 MUX2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_5996_), .B(_14920__bF_buf12), .S(_5983_), .Y(_232__12_) );
AOI21X1 AOI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf16), .C(data_78__13_), .Y(_5997_) );
AOI21X1 AOI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_5985_), .C(_5997_), .Y(_232__13_) );
AOI21X1 AOI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf15), .C(data_78__14_), .Y(_5998_) );
AOI21X1 AOI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf5), .B(_5985_), .C(_5998_), .Y(_232__14_) );
AOI21X1 AOI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_5982_), .B(_3313__bF_buf14), .C(data_78__15_), .Y(_5999_) );
AOI21X1 AOI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_5985_), .C(_5999_), .Y(_232__15_) );
INVX1 INVX1_2634 ( .gnd(gnd), .vdd(vdd), .A(data_77__0_), .Y(_6000_) );
OAI21X1 OAI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_3322_), .C(_5461_), .Y(_6001_) );
AOI21X1 AOI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_3332_), .B(_2672_), .C(_5421_), .Y(_6002_) );
OAI21X1 OAI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3322_), .C(_6002_), .Y(_6003_) );
NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(_6003_), .B(_4277_), .Y(_6004_) );
INVX1 INVX1_2635 ( .gnd(gnd), .vdd(vdd), .A(_6004_), .Y(_6005_) );
NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_6005_), .B(_6001_), .Y(_6006_) );
NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf13), .B(_6006_), .Y(_6007_) );
MUX2X1 MUX2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_6000_), .B(_14932__bF_buf5), .S(_6007_), .Y(_231__0_) );
INVX1 INVX1_2636 ( .gnd(gnd), .vdd(vdd), .A(data_77__1_), .Y(_6008_) );
MUX2X1 MUX2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_6008_), .B(_14894__bF_buf5), .S(_6007_), .Y(_231__1_) );
INVX1 INVX1_2637 ( .gnd(gnd), .vdd(vdd), .A(data_77__2_), .Y(_6009_) );
MUX2X1 MUX2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_6009_), .B(_14897__bF_buf0), .S(_6007_), .Y(_231__2_) );
INVX1 INVX1_2638 ( .gnd(gnd), .vdd(vdd), .A(data_77__3_), .Y(_6010_) );
MUX2X1 MUX2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_6010_), .B(_14899__bF_buf4), .S(_6007_), .Y(_231__3_) );
INVX1 INVX1_2639 ( .gnd(gnd), .vdd(vdd), .A(data_77__4_), .Y(_6011_) );
MUX2X1 MUX2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_6011_), .B(_14902__bF_buf8), .S(_6007_), .Y(_231__4_) );
INVX1 INVX1_2640 ( .gnd(gnd), .vdd(vdd), .A(data_77__5_), .Y(_6012_) );
NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_5979_), .B(_5420__bF_buf2), .Y(_6013_) );
NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_6004_), .B(_6013_), .Y(_6014_) );
OAI21X1 OAI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_3393__bF_buf46), .C(_6012_), .Y(_6015_) );
NAND3X1 NAND3X1_815 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_3313__bF_buf12), .C(_6006_), .Y(_6016_) );
AND2X2 AND2X2_1157 ( .gnd(gnd), .vdd(vdd), .A(_6015_), .B(_6016_), .Y(_231__5_) );
INVX1 INVX1_2641 ( .gnd(gnd), .vdd(vdd), .A(data_77__6_), .Y(_6017_) );
MUX2X1 MUX2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_6017_), .B(_15049__bF_buf2), .S(_6007_), .Y(_231__6_) );
INVX1 INVX1_2642 ( .gnd(gnd), .vdd(vdd), .A(data_77__7_), .Y(_6018_) );
OAI21X1 OAI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_3393__bF_buf45), .C(_6018_), .Y(_6019_) );
NAND3X1 NAND3X1_816 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_3313__bF_buf11), .C(_6006_), .Y(_6020_) );
AND2X2 AND2X2_1158 ( .gnd(gnd), .vdd(vdd), .A(_6019_), .B(_6020_), .Y(_231__7_) );
INVX1 INVX1_2643 ( .gnd(gnd), .vdd(vdd), .A(data_77__8_), .Y(_6021_) );
MUX2X1 MUX2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_6021_), .B(_15052__bF_buf8), .S(_6007_), .Y(_231__8_) );
NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_6014_), .Y(_6022_) );
AOI21X1 AOI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf10), .B(_6006_), .C(data_77__9_), .Y(_6023_) );
AOI21X1 AOI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_6022_), .C(_6023_), .Y(_231__9_) );
AOI21X1 AOI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf9), .B(_6006_), .C(data_77__10_), .Y(_6024_) );
AOI21X1 AOI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf10), .B(_6022_), .C(_6024_), .Y(_231__10_) );
INVX1 INVX1_2644 ( .gnd(gnd), .vdd(vdd), .A(data_77__11_), .Y(_6025_) );
MUX2X1 MUX2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_6025_), .B(_14918__bF_buf10), .S(_6007_), .Y(_231__11_) );
INVX1 INVX1_2645 ( .gnd(gnd), .vdd(vdd), .A(data_77__12_), .Y(_6026_) );
OAI21X1 OAI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_6014_), .B(_3393__bF_buf43), .C(_6026_), .Y(_6027_) );
NAND3X1 NAND3X1_817 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_3313__bF_buf8), .C(_6006_), .Y(_6028_) );
AND2X2 AND2X2_1159 ( .gnd(gnd), .vdd(vdd), .A(_6027_), .B(_6028_), .Y(_231__12_) );
AOI21X1 AOI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf7), .B(_6006_), .C(data_77__13_), .Y(_6029_) );
AOI21X1 AOI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_6022_), .C(_6029_), .Y(_231__13_) );
INVX1 INVX1_2646 ( .gnd(gnd), .vdd(vdd), .A(data_77__14_), .Y(_6030_) );
MUX2X1 MUX2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_6030_), .B(_15060__bF_buf4), .S(_6007_), .Y(_231__14_) );
INVX1 INVX1_2647 ( .gnd(gnd), .vdd(vdd), .A(data_77__15_), .Y(_6031_) );
MUX2X1 MUX2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_6031_), .B(_15062__bF_buf10), .S(_6007_), .Y(_231__15_) );
INVX1 INVX1_2648 ( .gnd(gnd), .vdd(vdd), .A(data_76__0_), .Y(_6032_) );
OAI21X1 OAI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_3322_), .C(_6002_), .Y(_6033_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_6033_), .B(_4277_), .Y(_6034_) );
NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_6034_), .B(_5420__bF_buf1), .Y(_6035_) );
INVX4 INVX4_21 ( .gnd(gnd), .vdd(vdd), .A(_6035_), .Y(_6036_) );
OAI21X1 OAI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_6036_), .C(_6032_), .Y(_6037_) );
NAND3X1 NAND3X1_818 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_6035_), .C(_3313__bF_buf6), .Y(_6038_) );
AND2X2 AND2X2_1160 ( .gnd(gnd), .vdd(vdd), .A(_6037_), .B(_6038_), .Y(_230__0_) );
INVX1 INVX1_2649 ( .gnd(gnd), .vdd(vdd), .A(data_76__1_), .Y(_6039_) );
OAI21X1 OAI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_6036_), .C(_6039_), .Y(_6040_) );
NAND3X1 NAND3X1_819 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_6035_), .C(_3313__bF_buf5), .Y(_6041_) );
AND2X2 AND2X2_1161 ( .gnd(gnd), .vdd(vdd), .A(_6040_), .B(_6041_), .Y(_230__1_) );
INVX1 INVX1_2650 ( .gnd(gnd), .vdd(vdd), .A(data_76__2_), .Y(_6042_) );
NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_6035_), .B(_3313__bF_buf4), .Y(_6043_) );
MUX2X1 MUX2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_6042_), .B(_14897__bF_buf14), .S(_6043_), .Y(_230__2_) );
INVX1 INVX1_2651 ( .gnd(gnd), .vdd(vdd), .A(data_76__3_), .Y(_6044_) );
OAI21X1 OAI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_6036_), .C(_6044_), .Y(_6045_) );
NAND3X1 NAND3X1_820 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_6035_), .C(_3313__bF_buf3), .Y(_6046_) );
AND2X2 AND2X2_1162 ( .gnd(gnd), .vdd(vdd), .A(_6045_), .B(_6046_), .Y(_230__3_) );
INVX1 INVX1_2652 ( .gnd(gnd), .vdd(vdd), .A(data_76__4_), .Y(_6047_) );
OAI21X1 OAI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_6036_), .C(_6047_), .Y(_6048_) );
NAND3X1 NAND3X1_821 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_6035_), .C(_3313__bF_buf2), .Y(_6049_) );
AND2X2 AND2X2_1163 ( .gnd(gnd), .vdd(vdd), .A(_6048_), .B(_6049_), .Y(_230__4_) );
INVX1 INVX1_2653 ( .gnd(gnd), .vdd(vdd), .A(data_76__5_), .Y(_6050_) );
OAI21X1 OAI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_6036_), .C(_6050_), .Y(_6051_) );
NAND3X1 NAND3X1_822 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_6035_), .C(_3313__bF_buf1), .Y(_6052_) );
AND2X2 AND2X2_1164 ( .gnd(gnd), .vdd(vdd), .A(_6051_), .B(_6052_), .Y(_230__5_) );
INVX1 INVX1_2654 ( .gnd(gnd), .vdd(vdd), .A(data_76__6_), .Y(_6053_) );
MUX2X1 MUX2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_6053_), .B(_15049__bF_buf1), .S(_6043_), .Y(_230__6_) );
INVX1 INVX1_2655 ( .gnd(gnd), .vdd(vdd), .A(data_76__7_), .Y(_6054_) );
OAI21X1 OAI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_6036_), .C(_6054_), .Y(_6055_) );
NAND3X1 NAND3X1_823 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_6035_), .C(_3313__bF_buf0), .Y(_6056_) );
AND2X2 AND2X2_1165 ( .gnd(gnd), .vdd(vdd), .A(_6055_), .B(_6056_), .Y(_230__7_) );
INVX1 INVX1_2656 ( .gnd(gnd), .vdd(vdd), .A(data_76__8_), .Y(_6057_) );
MUX2X1 MUX2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_6057_), .B(_15052__bF_buf7), .S(_6043_), .Y(_230__8_) );
INVX1 INVX1_2657 ( .gnd(gnd), .vdd(vdd), .A(data_76__9_), .Y(_6058_) );
MUX2X1 MUX2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_6058_), .B(_14913__bF_buf2), .S(_6043_), .Y(_230__9_) );
INVX1 INVX1_2658 ( .gnd(gnd), .vdd(vdd), .A(data_76__10_), .Y(_6059_) );
MUX2X1 MUX2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_6059_), .B(_15055__bF_buf9), .S(_6043_), .Y(_230__10_) );
INVX1 INVX1_2659 ( .gnd(gnd), .vdd(vdd), .A(data_76__11_), .Y(_6060_) );
OAI21X1 OAI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_6036_), .C(_6060_), .Y(_6061_) );
NAND3X1 NAND3X1_824 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_6035_), .C(_3313__bF_buf91), .Y(_6062_) );
AND2X2 AND2X2_1166 ( .gnd(gnd), .vdd(vdd), .A(_6061_), .B(_6062_), .Y(_230__11_) );
INVX1 INVX1_2660 ( .gnd(gnd), .vdd(vdd), .A(data_76__12_), .Y(_6063_) );
OAI21X1 OAI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_6036_), .C(_6063_), .Y(_6064_) );
NAND3X1 NAND3X1_825 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_6035_), .C(_3313__bF_buf90), .Y(_6065_) );
AND2X2 AND2X2_1167 ( .gnd(gnd), .vdd(vdd), .A(_6064_), .B(_6065_), .Y(_230__12_) );
INVX1 INVX1_2661 ( .gnd(gnd), .vdd(vdd), .A(data_76__13_), .Y(_6066_) );
MUX2X1 MUX2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_6066_), .B(_14924__bF_buf7), .S(_6043_), .Y(_230__13_) );
INVX1 INVX1_2662 ( .gnd(gnd), .vdd(vdd), .A(data_76__14_), .Y(_6067_) );
MUX2X1 MUX2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_6067_), .B(_15060__bF_buf3), .S(_6043_), .Y(_230__14_) );
INVX1 INVX1_2663 ( .gnd(gnd), .vdd(vdd), .A(data_76__15_), .Y(_6068_) );
MUX2X1 MUX2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_6068_), .B(_15062__bF_buf9), .S(_6043_), .Y(_230__15_) );
INVX1 INVX1_2664 ( .gnd(gnd), .vdd(vdd), .A(data_75__0_), .Y(_6069_) );
AOI21X1 AOI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf1), .B(_3332_), .C(_5421_), .Y(_6070_) );
OAI21X1 OAI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(_3322_), .C(_6070_), .Y(_6071_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_4277_), .B(_6071_), .Y(_6072_) );
NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_6072_), .B(_5420__bF_buf0), .Y(_6073_) );
NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_6073_), .B(_3313__bF_buf89), .Y(_6074_) );
MUX2X1 MUX2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_6069_), .B(_14932__bF_buf3), .S(_6074_), .Y(_229__0_) );
INVX1 INVX1_2665 ( .gnd(gnd), .vdd(vdd), .A(data_75__1_), .Y(_6075_) );
MUX2X1 MUX2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_6075_), .B(_14894__bF_buf3), .S(_6074_), .Y(_229__1_) );
INVX1 INVX1_2666 ( .gnd(gnd), .vdd(vdd), .A(data_75__2_), .Y(_6076_) );
MUX2X1 MUX2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_6076_), .B(_14897__bF_buf13), .S(_6074_), .Y(_229__2_) );
INVX1 INVX1_2667 ( .gnd(gnd), .vdd(vdd), .A(data_75__3_), .Y(_6077_) );
MUX2X1 MUX2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_6077_), .B(_14899__bF_buf2), .S(_6074_), .Y(_229__3_) );
INVX1 INVX1_2668 ( .gnd(gnd), .vdd(vdd), .A(data_75__4_), .Y(_6078_) );
MUX2X1 MUX2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_6078_), .B(_14902__bF_buf6), .S(_6074_), .Y(_229__4_) );
INVX1 INVX1_2669 ( .gnd(gnd), .vdd(vdd), .A(data_75__5_), .Y(_6079_) );
MUX2X1 MUX2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_6079_), .B(_14903__bF_buf8), .S(_6074_), .Y(_229__5_) );
INVX1 INVX1_2670 ( .gnd(gnd), .vdd(vdd), .A(data_75__6_), .Y(_6080_) );
MUX2X1 MUX2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_6080_), .B(_15049__bF_buf0), .S(_6074_), .Y(_229__6_) );
INVX1 INVX1_2671 ( .gnd(gnd), .vdd(vdd), .A(data_75__7_), .Y(_6081_) );
MUX2X1 MUX2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_6081_), .B(_14908__bF_buf8), .S(_6074_), .Y(_229__7_) );
INVX1 INVX1_2672 ( .gnd(gnd), .vdd(vdd), .A(data_75__8_), .Y(_6082_) );
MUX2X1 MUX2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_6082_), .B(_15052__bF_buf6), .S(_6074_), .Y(_229__8_) );
INVX1 INVX1_2673 ( .gnd(gnd), .vdd(vdd), .A(data_75__9_), .Y(_6083_) );
MUX2X1 MUX2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_6083_), .B(_14913__bF_buf1), .S(_6074_), .Y(_229__9_) );
INVX1 INVX1_2674 ( .gnd(gnd), .vdd(vdd), .A(data_75__10_), .Y(_6084_) );
MUX2X1 MUX2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_6084_), .B(_15055__bF_buf8), .S(_6074_), .Y(_229__10_) );
INVX1 INVX1_2675 ( .gnd(gnd), .vdd(vdd), .A(data_75__11_), .Y(_6085_) );
MUX2X1 MUX2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_6085_), .B(_14918__bF_buf8), .S(_6074_), .Y(_229__11_) );
INVX1 INVX1_2676 ( .gnd(gnd), .vdd(vdd), .A(data_75__12_), .Y(_6086_) );
MUX2X1 MUX2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_6086_), .B(_14920__bF_buf9), .S(_6074_), .Y(_229__12_) );
INVX1 INVX1_2677 ( .gnd(gnd), .vdd(vdd), .A(data_75__13_), .Y(_6087_) );
MUX2X1 MUX2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_6087_), .B(_14924__bF_buf6), .S(_6074_), .Y(_229__13_) );
INVX1 INVX1_2678 ( .gnd(gnd), .vdd(vdd), .A(data_75__14_), .Y(_6088_) );
MUX2X1 MUX2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_6088_), .B(_15060__bF_buf2), .S(_6074_), .Y(_229__14_) );
INVX1 INVX1_2679 ( .gnd(gnd), .vdd(vdd), .A(data_75__15_), .Y(_6089_) );
MUX2X1 MUX2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_6089_), .B(_15062__bF_buf8), .S(_6074_), .Y(_229__15_) );
INVX1 INVX1_2680 ( .gnd(gnd), .vdd(vdd), .A(data_74__0_), .Y(_6090_) );
OAI21X1 OAI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_3783_), .B(_14996_), .C(_3332_), .Y(_6091_) );
NAND3X1 NAND3X1_826 ( .gnd(gnd), .vdd(vdd), .A(_6070_), .B(_6091_), .C(_3335_), .Y(_6092_) );
NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(_6092_), .B(_5420__bF_buf3), .Y(_6093_) );
INVX4 INVX4_22 ( .gnd(gnd), .vdd(vdd), .A(_6093_), .Y(_6094_) );
OAI21X1 OAI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf34), .B(_6094_), .C(_6090_), .Y(_6095_) );
NAND3X1 NAND3X1_827 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_6093_), .C(_3313__bF_buf88), .Y(_6096_) );
AND2X2 AND2X2_1168 ( .gnd(gnd), .vdd(vdd), .A(_6095_), .B(_6096_), .Y(_228__0_) );
INVX1 INVX1_2681 ( .gnd(gnd), .vdd(vdd), .A(data_74__1_), .Y(_6097_) );
OAI21X1 OAI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_6094_), .C(_6097_), .Y(_6098_) );
NAND3X1 NAND3X1_828 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_6093_), .C(_3313__bF_buf87), .Y(_6099_) );
AND2X2 AND2X2_1169 ( .gnd(gnd), .vdd(vdd), .A(_6098_), .B(_6099_), .Y(_228__1_) );
INVX1 INVX1_2682 ( .gnd(gnd), .vdd(vdd), .A(data_74__2_), .Y(_6100_) );
NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_6093_), .B(_3313__bF_buf86), .Y(_6101_) );
MUX2X1 MUX2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_6100_), .B(_14897__bF_buf12), .S(_6101_), .Y(_228__2_) );
INVX1 INVX1_2683 ( .gnd(gnd), .vdd(vdd), .A(data_74__3_), .Y(_6102_) );
OAI21X1 OAI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_6094_), .C(_6102_), .Y(_6103_) );
NAND3X1 NAND3X1_829 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_6093_), .C(_3313__bF_buf85), .Y(_6104_) );
AND2X2 AND2X2_1170 ( .gnd(gnd), .vdd(vdd), .A(_6103_), .B(_6104_), .Y(_228__3_) );
INVX1 INVX1_2684 ( .gnd(gnd), .vdd(vdd), .A(data_74__4_), .Y(_6105_) );
OAI21X1 OAI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_6094_), .C(_6105_), .Y(_6106_) );
NAND3X1 NAND3X1_830 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_6093_), .C(_3313__bF_buf84), .Y(_6107_) );
AND2X2 AND2X2_1171 ( .gnd(gnd), .vdd(vdd), .A(_6106_), .B(_6107_), .Y(_228__4_) );
INVX1 INVX1_2685 ( .gnd(gnd), .vdd(vdd), .A(data_74__5_), .Y(_6108_) );
OAI21X1 OAI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_6094_), .C(_6108_), .Y(_6109_) );
NAND3X1 NAND3X1_831 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_6093_), .C(_3313__bF_buf83), .Y(_6110_) );
AND2X2 AND2X2_1172 ( .gnd(gnd), .vdd(vdd), .A(_6109_), .B(_6110_), .Y(_228__5_) );
INVX1 INVX1_2686 ( .gnd(gnd), .vdd(vdd), .A(data_74__6_), .Y(_6111_) );
MUX2X1 MUX2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_6111_), .B(_15049__bF_buf14), .S(_6101_), .Y(_228__6_) );
INVX1 INVX1_2687 ( .gnd(gnd), .vdd(vdd), .A(data_74__7_), .Y(_6112_) );
OAI21X1 OAI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_6094_), .C(_6112_), .Y(_6113_) );
NAND3X1 NAND3X1_832 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_6093_), .C(_3313__bF_buf82), .Y(_6114_) );
AND2X2 AND2X2_1173 ( .gnd(gnd), .vdd(vdd), .A(_6113_), .B(_6114_), .Y(_228__7_) );
INVX1 INVX1_2688 ( .gnd(gnd), .vdd(vdd), .A(data_74__8_), .Y(_6115_) );
MUX2X1 MUX2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_6115_), .B(_15052__bF_buf5), .S(_6101_), .Y(_228__8_) );
INVX1 INVX1_2689 ( .gnd(gnd), .vdd(vdd), .A(data_74__9_), .Y(_6116_) );
MUX2X1 MUX2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_6116_), .B(_14913__bF_buf0), .S(_6101_), .Y(_228__9_) );
INVX1 INVX1_2690 ( .gnd(gnd), .vdd(vdd), .A(data_74__10_), .Y(_6117_) );
MUX2X1 MUX2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_6117_), .B(_15055__bF_buf7), .S(_6101_), .Y(_228__10_) );
INVX1 INVX1_2691 ( .gnd(gnd), .vdd(vdd), .A(data_74__11_), .Y(_6118_) );
OAI21X1 OAI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_6094_), .C(_6118_), .Y(_6119_) );
NAND3X1 NAND3X1_833 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_6093_), .C(_3313__bF_buf81), .Y(_6120_) );
AND2X2 AND2X2_1174 ( .gnd(gnd), .vdd(vdd), .A(_6119_), .B(_6120_), .Y(_228__11_) );
INVX1 INVX1_2692 ( .gnd(gnd), .vdd(vdd), .A(data_74__12_), .Y(_6121_) );
OAI21X1 OAI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_6094_), .C(_6121_), .Y(_6122_) );
NAND3X1 NAND3X1_834 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_6093_), .C(_3313__bF_buf80), .Y(_6123_) );
AND2X2 AND2X2_1175 ( .gnd(gnd), .vdd(vdd), .A(_6122_), .B(_6123_), .Y(_228__12_) );
INVX1 INVX1_2693 ( .gnd(gnd), .vdd(vdd), .A(data_74__13_), .Y(_6124_) );
MUX2X1 MUX2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_6124_), .B(_14924__bF_buf5), .S(_6101_), .Y(_228__13_) );
INVX1 INVX1_2694 ( .gnd(gnd), .vdd(vdd), .A(data_74__14_), .Y(_6125_) );
MUX2X1 MUX2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_6125_), .B(_15060__bF_buf1), .S(_6101_), .Y(_228__14_) );
INVX1 INVX1_2695 ( .gnd(gnd), .vdd(vdd), .A(data_74__15_), .Y(_6126_) );
MUX2X1 MUX2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_6126_), .B(_15062__bF_buf7), .S(_6101_), .Y(_228__15_) );
INVX1 INVX1_2696 ( .gnd(gnd), .vdd(vdd), .A(data_73__0_), .Y(_6127_) );
OAI21X1 OAI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_3827_), .C(_6070_), .Y(_6128_) );
AOI21X1 AOI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_3332_), .C(_6128_), .Y(_6129_) );
NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_6129_), .B(_3335_), .Y(_6130_) );
NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_6130_), .B(_5420__bF_buf2), .Y(_6131_) );
NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf79), .Y(_6132_) );
MUX2X1 MUX2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_6127_), .B(_14932__bF_buf1), .S(_6132_), .Y(_227__0_) );
INVX1 INVX1_2697 ( .gnd(gnd), .vdd(vdd), .A(data_73__1_), .Y(_6133_) );
MUX2X1 MUX2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_6133_), .B(_14894__bF_buf1), .S(_6132_), .Y(_227__1_) );
AND2X2 AND2X2_1176 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf78), .B(_6131_), .Y(_6134_) );
AOI21X1 AOI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf77), .C(data_73__2_), .Y(_6135_) );
AOI21X1 AOI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_6134_), .C(_6135_), .Y(_227__2_) );
INVX1 INVX1_2698 ( .gnd(gnd), .vdd(vdd), .A(data_73__3_), .Y(_6136_) );
MUX2X1 MUX2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_6136_), .B(_14899__bF_buf0), .S(_6132_), .Y(_227__3_) );
INVX1 INVX1_2699 ( .gnd(gnd), .vdd(vdd), .A(data_73__4_), .Y(_6137_) );
MUX2X1 MUX2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_6137_), .B(_14902__bF_buf4), .S(_6132_), .Y(_227__4_) );
INVX1 INVX1_2700 ( .gnd(gnd), .vdd(vdd), .A(data_73__5_), .Y(_6138_) );
MUX2X1 MUX2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_6138_), .B(_14903__bF_buf6), .S(_6132_), .Y(_227__5_) );
AOI21X1 AOI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf76), .C(data_73__6_), .Y(_6139_) );
AOI21X1 AOI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_6134_), .C(_6139_), .Y(_227__6_) );
INVX1 INVX1_2701 ( .gnd(gnd), .vdd(vdd), .A(data_73__7_), .Y(_6140_) );
MUX2X1 MUX2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_6140_), .B(_14908__bF_buf6), .S(_6132_), .Y(_227__7_) );
AOI21X1 AOI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf75), .C(data_73__8_), .Y(_6141_) );
AOI21X1 AOI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_6134_), .C(_6141_), .Y(_227__8_) );
AOI21X1 AOI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf74), .C(data_73__9_), .Y(_6142_) );
AOI21X1 AOI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf14), .B(_6134_), .C(_6142_), .Y(_227__9_) );
AOI21X1 AOI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf73), .C(data_73__10_), .Y(_6143_) );
AOI21X1 AOI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_6134_), .C(_6143_), .Y(_227__10_) );
INVX1 INVX1_2702 ( .gnd(gnd), .vdd(vdd), .A(data_73__11_), .Y(_6144_) );
MUX2X1 MUX2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_6144_), .B(_14918__bF_buf6), .S(_6132_), .Y(_227__11_) );
INVX1 INVX1_2703 ( .gnd(gnd), .vdd(vdd), .A(data_73__12_), .Y(_6145_) );
MUX2X1 MUX2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_6145_), .B(_14920__bF_buf7), .S(_6132_), .Y(_227__12_) );
AOI21X1 AOI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf72), .C(data_73__13_), .Y(_6146_) );
AOI21X1 AOI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_6134_), .C(_6146_), .Y(_227__13_) );
AOI21X1 AOI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf71), .C(data_73__14_), .Y(_6147_) );
AOI21X1 AOI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_6134_), .C(_6147_), .Y(_227__14_) );
AOI21X1 AOI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_6131_), .B(_3313__bF_buf70), .C(data_73__15_), .Y(_6148_) );
AOI21X1 AOI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_6134_), .C(_6148_), .Y(_227__15_) );
INVX1 INVX1_2704 ( .gnd(gnd), .vdd(vdd), .A(data_72__0_), .Y(_6149_) );
AOI21X1 AOI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_3332_), .B(_4467_), .C(_6128_), .Y(_6150_) );
NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_6150_), .B(_3335_), .Y(_6151_) );
NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_6151_), .B(_5420__bF_buf1), .Y(_6152_) );
NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(_3313__bF_buf69), .Y(_6153_) );
MUX2X1 MUX2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_6149_), .B(_14932__bF_buf0), .S(_6153_), .Y(_226__0_) );
INVX1 INVX1_2705 ( .gnd(gnd), .vdd(vdd), .A(data_72__1_), .Y(_6154_) );
MUX2X1 MUX2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_6154_), .B(_14894__bF_buf0), .S(_6153_), .Y(_226__1_) );
INVX1 INVX1_2706 ( .gnd(gnd), .vdd(vdd), .A(data_72__2_), .Y(_6155_) );
MUX2X1 MUX2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_6155_), .B(_14897__bF_buf10), .S(_6153_), .Y(_226__2_) );
INVX1 INVX1_2707 ( .gnd(gnd), .vdd(vdd), .A(data_72__3_), .Y(_6156_) );
MUX2X1 MUX2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_6156_), .B(_14899__bF_buf14), .S(_6153_), .Y(_226__3_) );
INVX1 INVX1_2708 ( .gnd(gnd), .vdd(vdd), .A(data_72__4_), .Y(_6157_) );
MUX2X1 MUX2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_6157_), .B(_14902__bF_buf3), .S(_6153_), .Y(_226__4_) );
INVX1 INVX1_2709 ( .gnd(gnd), .vdd(vdd), .A(data_72__5_), .Y(_6158_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .Y(_6159_) );
OAI21X1 OAI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_6159_), .C(_6158_), .Y(_6160_) );
NAND3X1 NAND3X1_835 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_6152_), .C(_3313__bF_buf68), .Y(_6161_) );
AND2X2 AND2X2_1177 ( .gnd(gnd), .vdd(vdd), .A(_6160_), .B(_6161_), .Y(_226__5_) );
INVX1 INVX1_2710 ( .gnd(gnd), .vdd(vdd), .A(data_72__6_), .Y(_6162_) );
MUX2X1 MUX2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_6162_), .B(_15049__bF_buf12), .S(_6153_), .Y(_226__6_) );
INVX1 INVX1_2711 ( .gnd(gnd), .vdd(vdd), .A(data_72__7_), .Y(_6163_) );
OAI21X1 OAI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_6159_), .C(_6163_), .Y(_6164_) );
NAND3X1 NAND3X1_836 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_6152_), .C(_3313__bF_buf67), .Y(_6165_) );
AND2X2 AND2X2_1178 ( .gnd(gnd), .vdd(vdd), .A(_6164_), .B(_6165_), .Y(_226__7_) );
INVX1 INVX1_2712 ( .gnd(gnd), .vdd(vdd), .A(data_72__8_), .Y(_6166_) );
MUX2X1 MUX2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_6166_), .B(_15052__bF_buf3), .S(_6153_), .Y(_226__8_) );
NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_6159_), .B(_3393__bF_buf24), .Y(_6167_) );
AOI21X1 AOI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(_3313__bF_buf66), .C(data_72__9_), .Y(_6168_) );
AOI21X1 AOI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_6167_), .C(_6168_), .Y(_226__9_) );
AOI21X1 AOI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(_3313__bF_buf65), .C(data_72__10_), .Y(_6169_) );
AOI21X1 AOI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_6167_), .C(_6169_), .Y(_226__10_) );
INVX1 INVX1_2713 ( .gnd(gnd), .vdd(vdd), .A(data_72__11_), .Y(_6170_) );
MUX2X1 MUX2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_6170_), .B(_14918__bF_buf5), .S(_6153_), .Y(_226__11_) );
INVX1 INVX1_2714 ( .gnd(gnd), .vdd(vdd), .A(data_72__12_), .Y(_6171_) );
OAI21X1 OAI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_6159_), .C(_6171_), .Y(_6172_) );
NAND3X1 NAND3X1_837 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_6152_), .C(_3313__bF_buf64), .Y(_6173_) );
AND2X2 AND2X2_1179 ( .gnd(gnd), .vdd(vdd), .A(_6172_), .B(_6173_), .Y(_226__12_) );
AOI21X1 AOI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_6152_), .B(_3313__bF_buf63), .C(data_72__13_), .Y(_6174_) );
AOI21X1 AOI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_6167_), .C(_6174_), .Y(_226__13_) );
INVX1 INVX1_2715 ( .gnd(gnd), .vdd(vdd), .A(data_72__14_), .Y(_6175_) );
MUX2X1 MUX2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_6175_), .B(_15060__bF_buf14), .S(_6153_), .Y(_226__14_) );
INVX1 INVX1_2716 ( .gnd(gnd), .vdd(vdd), .A(data_72__15_), .Y(_6176_) );
MUX2X1 MUX2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_6176_), .B(_15062__bF_buf5), .S(_6153_), .Y(_226__15_) );
INVX1 INVX1_2717 ( .gnd(gnd), .vdd(vdd), .A(data_71__0_), .Y(_6177_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_3331_), .B(_5421_), .Y(_6178_) );
NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_6178_), .Y(_6179_) );
AOI21X1 AOI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf1), .B(_3332_), .C(_3334_), .Y(_6180_) );
NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_6180_), .B(_6179_), .Y(_6181_) );
NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_6181_), .B(_5420__bF_buf0), .Y(_6182_) );
INVX4 INVX4_23 ( .gnd(gnd), .vdd(vdd), .A(_6182_), .Y(_6183_) );
OAI21X1 OAI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_6183_), .C(_6177_), .Y(_6184_) );
NAND3X1 NAND3X1_838 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_6182_), .C(_3313__bF_buf62), .Y(_6185_) );
AND2X2 AND2X2_1180 ( .gnd(gnd), .vdd(vdd), .A(_6184_), .B(_6185_), .Y(_225__0_) );
INVX1 INVX1_2718 ( .gnd(gnd), .vdd(vdd), .A(data_71__1_), .Y(_6186_) );
OAI21X1 OAI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_6183_), .C(_6186_), .Y(_6187_) );
NAND3X1 NAND3X1_839 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_6182_), .C(_3313__bF_buf61), .Y(_6188_) );
AND2X2 AND2X2_1181 ( .gnd(gnd), .vdd(vdd), .A(_6187_), .B(_6188_), .Y(_225__1_) );
INVX1 INVX1_2719 ( .gnd(gnd), .vdd(vdd), .A(data_71__2_), .Y(_6189_) );
NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_6182_), .B(_3313__bF_buf60), .Y(_6190_) );
MUX2X1 MUX2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_6189_), .B(_14897__bF_buf9), .S(_6190_), .Y(_225__2_) );
INVX1 INVX1_2720 ( .gnd(gnd), .vdd(vdd), .A(data_71__3_), .Y(_6191_) );
OAI21X1 OAI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf20), .B(_6183_), .C(_6191_), .Y(_6192_) );
NAND3X1 NAND3X1_840 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_6182_), .C(_3313__bF_buf59), .Y(_6193_) );
AND2X2 AND2X2_1182 ( .gnd(gnd), .vdd(vdd), .A(_6192_), .B(_6193_), .Y(_225__3_) );
INVX1 INVX1_2721 ( .gnd(gnd), .vdd(vdd), .A(data_71__4_), .Y(_6194_) );
OAI21X1 OAI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_6183_), .C(_6194_), .Y(_6195_) );
NAND3X1 NAND3X1_841 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_6182_), .C(_3313__bF_buf58), .Y(_6196_) );
AND2X2 AND2X2_1183 ( .gnd(gnd), .vdd(vdd), .A(_6195_), .B(_6196_), .Y(_225__4_) );
INVX1 INVX1_2722 ( .gnd(gnd), .vdd(vdd), .A(data_71__5_), .Y(_6197_) );
OAI21X1 OAI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_6183_), .C(_6197_), .Y(_6198_) );
NAND3X1 NAND3X1_842 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_6182_), .C(_3313__bF_buf57), .Y(_6199_) );
AND2X2 AND2X2_1184 ( .gnd(gnd), .vdd(vdd), .A(_6198_), .B(_6199_), .Y(_225__5_) );
INVX1 INVX1_2723 ( .gnd(gnd), .vdd(vdd), .A(data_71__6_), .Y(_6200_) );
MUX2X1 MUX2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_6200_), .B(_15049__bF_buf11), .S(_6190_), .Y(_225__6_) );
INVX1 INVX1_2724 ( .gnd(gnd), .vdd(vdd), .A(data_71__7_), .Y(_6201_) );
OAI21X1 OAI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf17), .B(_6183_), .C(_6201_), .Y(_6202_) );
NAND3X1 NAND3X1_843 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_6182_), .C(_3313__bF_buf56), .Y(_6203_) );
AND2X2 AND2X2_1185 ( .gnd(gnd), .vdd(vdd), .A(_6202_), .B(_6203_), .Y(_225__7_) );
INVX1 INVX1_2725 ( .gnd(gnd), .vdd(vdd), .A(data_71__8_), .Y(_6204_) );
MUX2X1 MUX2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_6204_), .B(_15052__bF_buf2), .S(_6190_), .Y(_225__8_) );
INVX1 INVX1_2726 ( .gnd(gnd), .vdd(vdd), .A(data_71__9_), .Y(_6205_) );
MUX2X1 MUX2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_6205_), .B(_14913__bF_buf12), .S(_6190_), .Y(_225__9_) );
INVX1 INVX1_2727 ( .gnd(gnd), .vdd(vdd), .A(data_71__10_), .Y(_6206_) );
MUX2X1 MUX2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_6206_), .B(_15055__bF_buf4), .S(_6190_), .Y(_225__10_) );
INVX1 INVX1_2728 ( .gnd(gnd), .vdd(vdd), .A(data_71__11_), .Y(_6207_) );
OAI21X1 OAI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf16), .B(_6183_), .C(_6207_), .Y(_6208_) );
NAND3X1 NAND3X1_844 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_6182_), .C(_3313__bF_buf55), .Y(_6209_) );
AND2X2 AND2X2_1186 ( .gnd(gnd), .vdd(vdd), .A(_6208_), .B(_6209_), .Y(_225__11_) );
INVX1 INVX1_2729 ( .gnd(gnd), .vdd(vdd), .A(data_71__12_), .Y(_6210_) );
OAI21X1 OAI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf15), .B(_6183_), .C(_6210_), .Y(_6211_) );
NAND3X1 NAND3X1_845 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_6182_), .C(_3313__bF_buf54), .Y(_6212_) );
AND2X2 AND2X2_1187 ( .gnd(gnd), .vdd(vdd), .A(_6211_), .B(_6212_), .Y(_225__12_) );
INVX1 INVX1_2730 ( .gnd(gnd), .vdd(vdd), .A(data_71__13_), .Y(_6213_) );
MUX2X1 MUX2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_6213_), .B(_14924__bF_buf2), .S(_6190_), .Y(_225__13_) );
INVX1 INVX1_2731 ( .gnd(gnd), .vdd(vdd), .A(data_71__14_), .Y(_6214_) );
MUX2X1 MUX2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_6214_), .B(_15060__bF_buf13), .S(_6190_), .Y(_225__14_) );
INVX1 INVX1_2732 ( .gnd(gnd), .vdd(vdd), .A(data_71__15_), .Y(_6215_) );
MUX2X1 MUX2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_6215_), .B(_15062__bF_buf4), .S(_6190_), .Y(_225__15_) );
INVX1 INVX1_2733 ( .gnd(gnd), .vdd(vdd), .A(data_70__0_), .Y(_6216_) );
AOI21X1 AOI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_3332_), .B(_14978__bF_buf2), .C(_5421_), .Y(_6217_) );
OAI21X1 OAI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_3943_), .B(IDATA_PROG_addr_3_bF_buf0), .C(_3332_), .Y(_6218_) );
NAND3X1 NAND3X1_846 ( .gnd(gnd), .vdd(vdd), .A(_6217_), .B(_6218_), .C(_4276_), .Y(_6219_) );
NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(_6219_), .B(_5420__bF_buf3), .Y(_6220_) );
INVX4 INVX4_24 ( .gnd(gnd), .vdd(vdd), .A(_6220_), .Y(_6221_) );
OAI21X1 OAI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf14), .B(_6221_), .C(_6216_), .Y(_6222_) );
NAND3X1 NAND3X1_847 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_6220_), .C(_3313__bF_buf53), .Y(_6223_) );
AND2X2 AND2X2_1188 ( .gnd(gnd), .vdd(vdd), .A(_6222_), .B(_6223_), .Y(_224__0_) );
INVX1 INVX1_2734 ( .gnd(gnd), .vdd(vdd), .A(data_70__1_), .Y(_6224_) );
OAI21X1 OAI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf13), .B(_6221_), .C(_6224_), .Y(_6225_) );
NAND3X1 NAND3X1_848 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_6220_), .C(_3313__bF_buf52), .Y(_6226_) );
AND2X2 AND2X2_1189 ( .gnd(gnd), .vdd(vdd), .A(_6225_), .B(_6226_), .Y(_224__1_) );
INVX1 INVX1_2735 ( .gnd(gnd), .vdd(vdd), .A(data_70__2_), .Y(_6227_) );
NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_6220_), .B(_3313__bF_buf51), .Y(_6228_) );
MUX2X1 MUX2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_6227_), .B(_14897__bF_buf8), .S(_6228_), .Y(_224__2_) );
INVX1 INVX1_2736 ( .gnd(gnd), .vdd(vdd), .A(data_70__3_), .Y(_6229_) );
OAI21X1 OAI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_6221_), .C(_6229_), .Y(_6230_) );
NAND3X1 NAND3X1_849 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_6220_), .C(_3313__bF_buf50), .Y(_6231_) );
AND2X2 AND2X2_1190 ( .gnd(gnd), .vdd(vdd), .A(_6230_), .B(_6231_), .Y(_224__3_) );
INVX1 INVX1_2737 ( .gnd(gnd), .vdd(vdd), .A(data_70__4_), .Y(_6232_) );
OAI21X1 OAI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_6221_), .C(_6232_), .Y(_6233_) );
NAND3X1 NAND3X1_850 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_6220_), .C(_3313__bF_buf49), .Y(_6234_) );
AND2X2 AND2X2_1191 ( .gnd(gnd), .vdd(vdd), .A(_6233_), .B(_6234_), .Y(_224__4_) );
INVX1 INVX1_2738 ( .gnd(gnd), .vdd(vdd), .A(data_70__5_), .Y(_6235_) );
OAI21X1 OAI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_6221_), .C(_6235_), .Y(_6236_) );
NAND3X1 NAND3X1_851 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_6220_), .C(_3313__bF_buf48), .Y(_6237_) );
AND2X2 AND2X2_1192 ( .gnd(gnd), .vdd(vdd), .A(_6236_), .B(_6237_), .Y(_224__5_) );
INVX1 INVX1_2739 ( .gnd(gnd), .vdd(vdd), .A(data_70__6_), .Y(_6238_) );
MUX2X1 MUX2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_6238_), .B(_15049__bF_buf10), .S(_6228_), .Y(_224__6_) );
INVX1 INVX1_2740 ( .gnd(gnd), .vdd(vdd), .A(data_70__7_), .Y(_6239_) );
OAI21X1 OAI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_6221_), .C(_6239_), .Y(_6240_) );
NAND3X1 NAND3X1_852 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_6220_), .C(_3313__bF_buf47), .Y(_6241_) );
AND2X2 AND2X2_1193 ( .gnd(gnd), .vdd(vdd), .A(_6240_), .B(_6241_), .Y(_224__7_) );
INVX1 INVX1_2741 ( .gnd(gnd), .vdd(vdd), .A(data_70__8_), .Y(_6242_) );
MUX2X1 MUX2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_6242_), .B(_15052__bF_buf1), .S(_6228_), .Y(_224__8_) );
INVX1 INVX1_2742 ( .gnd(gnd), .vdd(vdd), .A(data_70__9_), .Y(_6243_) );
MUX2X1 MUX2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_6243_), .B(_14913__bF_buf11), .S(_6228_), .Y(_224__9_) );
INVX1 INVX1_2743 ( .gnd(gnd), .vdd(vdd), .A(data_70__10_), .Y(_6244_) );
MUX2X1 MUX2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_6244_), .B(_15055__bF_buf3), .S(_6228_), .Y(_224__10_) );
INVX1 INVX1_2744 ( .gnd(gnd), .vdd(vdd), .A(data_70__11_), .Y(_6245_) );
OAI21X1 OAI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf8), .B(_6221_), .C(_6245_), .Y(_6246_) );
NAND3X1 NAND3X1_853 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_6220_), .C(_3313__bF_buf46), .Y(_6247_) );
AND2X2 AND2X2_1194 ( .gnd(gnd), .vdd(vdd), .A(_6246_), .B(_6247_), .Y(_224__11_) );
INVX1 INVX1_2745 ( .gnd(gnd), .vdd(vdd), .A(data_70__12_), .Y(_6248_) );
OAI21X1 OAI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_6221_), .C(_6248_), .Y(_6249_) );
NAND3X1 NAND3X1_854 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_6220_), .C(_3313__bF_buf45), .Y(_6250_) );
AND2X2 AND2X2_1195 ( .gnd(gnd), .vdd(vdd), .A(_6249_), .B(_6250_), .Y(_224__12_) );
INVX1 INVX1_2746 ( .gnd(gnd), .vdd(vdd), .A(data_70__13_), .Y(_6251_) );
MUX2X1 MUX2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_6251_), .B(_14924__bF_buf1), .S(_6228_), .Y(_224__13_) );
INVX1 INVX1_2747 ( .gnd(gnd), .vdd(vdd), .A(data_70__14_), .Y(_6252_) );
MUX2X1 MUX2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_6252_), .B(_15060__bF_buf12), .S(_6228_), .Y(_224__14_) );
INVX1 INVX1_2748 ( .gnd(gnd), .vdd(vdd), .A(data_70__15_), .Y(_6253_) );
MUX2X1 MUX2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_6253_), .B(_15062__bF_buf3), .S(_6228_), .Y(_224__15_) );
INVX1 INVX1_2749 ( .gnd(gnd), .vdd(vdd), .A(data_69__0_), .Y(_6254_) );
OAI21X1 OAI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(IDATA_PROG_addr_3_bF_buf3), .C(_3332_), .Y(_6255_) );
AND2X2 AND2X2_1196 ( .gnd(gnd), .vdd(vdd), .A(_6179_), .B(_6255_), .Y(_6256_) );
OAI21X1 OAI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_15172_), .B(_3322_), .C(_6256_), .Y(_6257_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_6257_), .B(_5420__bF_buf2), .Y(_6258_) );
OAI21X1 OAI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_6258_), .C(_6254_), .Y(_6259_) );
NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_5420__bF_buf1), .B(_6257_), .Y(_6260_) );
NAND3X1 NAND3X1_855 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_6260_), .C(_3313__bF_buf44), .Y(_6261_) );
AND2X2 AND2X2_1197 ( .gnd(gnd), .vdd(vdd), .A(_6259_), .B(_6261_), .Y(_222__0_) );
INVX1 INVX1_2750 ( .gnd(gnd), .vdd(vdd), .A(data_69__1_), .Y(_6262_) );
OAI21X1 OAI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_6258_), .C(_6262_), .Y(_6263_) );
NAND3X1 NAND3X1_856 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_6260_), .C(_3313__bF_buf43), .Y(_6264_) );
AND2X2 AND2X2_1198 ( .gnd(gnd), .vdd(vdd), .A(_6263_), .B(_6264_), .Y(_222__1_) );
INVX1 INVX1_2751 ( .gnd(gnd), .vdd(vdd), .A(data_69__2_), .Y(_6265_) );
NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_6260_), .B(_3313__bF_buf42), .Y(_6266_) );
MUX2X1 MUX2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_6265_), .B(_14897__bF_buf7), .S(_6266_), .Y(_222__2_) );
INVX1 INVX1_2752 ( .gnd(gnd), .vdd(vdd), .A(data_69__3_), .Y(_6267_) );
OAI21X1 OAI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_6258_), .C(_6267_), .Y(_6268_) );
NAND3X1 NAND3X1_857 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_6260_), .C(_3313__bF_buf41), .Y(_6269_) );
AND2X2 AND2X2_1199 ( .gnd(gnd), .vdd(vdd), .A(_6268_), .B(_6269_), .Y(_222__3_) );
INVX1 INVX1_2753 ( .gnd(gnd), .vdd(vdd), .A(data_69__4_), .Y(_6270_) );
OAI21X1 OAI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf3), .B(_6258_), .C(_6270_), .Y(_6271_) );
NAND3X1 NAND3X1_858 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_6260_), .C(_3313__bF_buf40), .Y(_6272_) );
AND2X2 AND2X2_1200 ( .gnd(gnd), .vdd(vdd), .A(_6271_), .B(_6272_), .Y(_222__4_) );
INVX1 INVX1_2754 ( .gnd(gnd), .vdd(vdd), .A(data_69__5_), .Y(_6273_) );
OAI21X1 OAI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_6258_), .C(_6273_), .Y(_6274_) );
NAND3X1 NAND3X1_859 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_6260_), .C(_3313__bF_buf39), .Y(_6275_) );
AND2X2 AND2X2_1201 ( .gnd(gnd), .vdd(vdd), .A(_6274_), .B(_6275_), .Y(_222__5_) );
INVX1 INVX1_2755 ( .gnd(gnd), .vdd(vdd), .A(data_69__6_), .Y(_6276_) );
MUX2X1 MUX2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_6276_), .B(_15049__bF_buf9), .S(_6266_), .Y(_222__6_) );
INVX1 INVX1_2756 ( .gnd(gnd), .vdd(vdd), .A(data_69__7_), .Y(_6277_) );
OAI21X1 OAI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_6258_), .C(_6277_), .Y(_6278_) );
NAND3X1 NAND3X1_860 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_6260_), .C(_3313__bF_buf38), .Y(_6279_) );
AND2X2 AND2X2_1202 ( .gnd(gnd), .vdd(vdd), .A(_6278_), .B(_6279_), .Y(_222__7_) );
INVX1 INVX1_2757 ( .gnd(gnd), .vdd(vdd), .A(data_69__8_), .Y(_6280_) );
MUX2X1 MUX2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_6280_), .B(_15052__bF_buf0), .S(_6266_), .Y(_222__8_) );
INVX1 INVX1_2758 ( .gnd(gnd), .vdd(vdd), .A(data_69__9_), .Y(_6281_) );
MUX2X1 MUX2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_6281_), .B(_14913__bF_buf10), .S(_6266_), .Y(_222__9_) );
INVX1 INVX1_2759 ( .gnd(gnd), .vdd(vdd), .A(data_69__10_), .Y(_6282_) );
MUX2X1 MUX2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_6282_), .B(_15055__bF_buf2), .S(_6266_), .Y(_222__10_) );
INVX1 INVX1_2760 ( .gnd(gnd), .vdd(vdd), .A(data_69__11_), .Y(_6283_) );
OAI21X1 OAI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_6258_), .C(_6283_), .Y(_6284_) );
NAND3X1 NAND3X1_861 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_6260_), .C(_3313__bF_buf37), .Y(_6285_) );
AND2X2 AND2X2_1203 ( .gnd(gnd), .vdd(vdd), .A(_6284_), .B(_6285_), .Y(_222__11_) );
INVX1 INVX1_2761 ( .gnd(gnd), .vdd(vdd), .A(data_69__12_), .Y(_6286_) );
OAI21X1 OAI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_6258_), .C(_6286_), .Y(_6287_) );
NAND3X1 NAND3X1_862 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_6260_), .C(_3313__bF_buf36), .Y(_6288_) );
AND2X2 AND2X2_1204 ( .gnd(gnd), .vdd(vdd), .A(_6287_), .B(_6288_), .Y(_222__12_) );
INVX1 INVX1_2762 ( .gnd(gnd), .vdd(vdd), .A(data_69__13_), .Y(_6289_) );
MUX2X1 MUX2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_6289_), .B(_14924__bF_buf0), .S(_6266_), .Y(_222__13_) );
INVX1 INVX1_2763 ( .gnd(gnd), .vdd(vdd), .A(data_69__14_), .Y(_6290_) );
MUX2X1 MUX2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_6290_), .B(_15060__bF_buf11), .S(_6266_), .Y(_222__14_) );
INVX1 INVX1_2764 ( .gnd(gnd), .vdd(vdd), .A(data_69__15_), .Y(_6291_) );
MUX2X1 MUX2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_6291_), .B(_15062__bF_buf2), .S(_6266_), .Y(_222__15_) );
INVX1 INVX1_2765 ( .gnd(gnd), .vdd(vdd), .A(data_68__0_), .Y(_6292_) );
OAI21X1 OAI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_3322_), .B(_4027_), .C(_6256_), .Y(_6293_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_6293_), .B(_5420__bF_buf0), .Y(_6294_) );
OAI21X1 OAI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_6294_), .C(_6292_), .Y(_6295_) );
NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_5420__bF_buf3), .B(_6293_), .Y(_6296_) );
NAND3X1 NAND3X1_863 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_6296_), .C(_3313__bF_buf35), .Y(_6297_) );
AND2X2 AND2X2_1205 ( .gnd(gnd), .vdd(vdd), .A(_6295_), .B(_6297_), .Y(_221__0_) );
INVX1 INVX1_2766 ( .gnd(gnd), .vdd(vdd), .A(data_68__1_), .Y(_6298_) );
OAI21X1 OAI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_6294_), .C(_6298_), .Y(_6299_) );
NAND3X1 NAND3X1_864 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_6296_), .C(_3313__bF_buf34), .Y(_6300_) );
AND2X2 AND2X2_1206 ( .gnd(gnd), .vdd(vdd), .A(_6299_), .B(_6300_), .Y(_221__1_) );
INVX1 INVX1_2767 ( .gnd(gnd), .vdd(vdd), .A(data_68__2_), .Y(_6301_) );
NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_6296_), .B(_3313__bF_buf33), .Y(_6302_) );
MUX2X1 MUX2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_6301_), .B(_14897__bF_buf6), .S(_6302_), .Y(_221__2_) );
INVX1 INVX1_2768 ( .gnd(gnd), .vdd(vdd), .A(data_68__3_), .Y(_6303_) );
OAI21X1 OAI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_6294_), .C(_6303_), .Y(_6304_) );
NAND3X1 NAND3X1_865 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_6296_), .C(_3313__bF_buf32), .Y(_6305_) );
AND2X2 AND2X2_1207 ( .gnd(gnd), .vdd(vdd), .A(_6304_), .B(_6305_), .Y(_221__3_) );
INVX1 INVX1_2769 ( .gnd(gnd), .vdd(vdd), .A(data_68__4_), .Y(_6306_) );
OAI21X1 OAI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_6294_), .C(_6306_), .Y(_6307_) );
NAND3X1 NAND3X1_866 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_6296_), .C(_3313__bF_buf31), .Y(_6308_) );
AND2X2 AND2X2_1208 ( .gnd(gnd), .vdd(vdd), .A(_6307_), .B(_6308_), .Y(_221__4_) );
INVX1 INVX1_2770 ( .gnd(gnd), .vdd(vdd), .A(data_68__5_), .Y(_6309_) );
OAI21X1 OAI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_6294_), .C(_6309_), .Y(_6310_) );
NAND3X1 NAND3X1_867 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_6296_), .C(_3313__bF_buf30), .Y(_6311_) );
AND2X2 AND2X2_1209 ( .gnd(gnd), .vdd(vdd), .A(_6310_), .B(_6311_), .Y(_221__5_) );
INVX1 INVX1_2771 ( .gnd(gnd), .vdd(vdd), .A(data_68__6_), .Y(_6312_) );
MUX2X1 MUX2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_6312_), .B(_15049__bF_buf8), .S(_6302_), .Y(_221__6_) );
INVX1 INVX1_2772 ( .gnd(gnd), .vdd(vdd), .A(data_68__7_), .Y(_6313_) );
OAI21X1 OAI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_6294_), .C(_6313_), .Y(_6314_) );
NAND3X1 NAND3X1_868 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_6296_), .C(_3313__bF_buf29), .Y(_6315_) );
AND2X2 AND2X2_1210 ( .gnd(gnd), .vdd(vdd), .A(_6314_), .B(_6315_), .Y(_221__7_) );
INVX1 INVX1_2773 ( .gnd(gnd), .vdd(vdd), .A(data_68__8_), .Y(_6316_) );
MUX2X1 MUX2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_6316_), .B(_15052__bF_buf13), .S(_6302_), .Y(_221__8_) );
INVX1 INVX1_2774 ( .gnd(gnd), .vdd(vdd), .A(data_68__9_), .Y(_6317_) );
MUX2X1 MUX2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_6317_), .B(_14913__bF_buf9), .S(_6302_), .Y(_221__9_) );
INVX1 INVX1_2775 ( .gnd(gnd), .vdd(vdd), .A(data_68__10_), .Y(_6318_) );
MUX2X1 MUX2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_6318_), .B(_15055__bF_buf1), .S(_6302_), .Y(_221__10_) );
INVX1 INVX1_2776 ( .gnd(gnd), .vdd(vdd), .A(data_68__11_), .Y(_6319_) );
OAI21X1 OAI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_6294_), .C(_6319_), .Y(_6320_) );
NAND3X1 NAND3X1_869 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_6296_), .C(_3313__bF_buf28), .Y(_6321_) );
AND2X2 AND2X2_1211 ( .gnd(gnd), .vdd(vdd), .A(_6320_), .B(_6321_), .Y(_221__11_) );
INVX1 INVX1_2777 ( .gnd(gnd), .vdd(vdd), .A(data_68__12_), .Y(_6322_) );
OAI21X1 OAI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_6294_), .C(_6322_), .Y(_6323_) );
NAND3X1 NAND3X1_870 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_6296_), .C(_3313__bF_buf27), .Y(_6324_) );
AND2X2 AND2X2_1212 ( .gnd(gnd), .vdd(vdd), .A(_6323_), .B(_6324_), .Y(_221__12_) );
INVX1 INVX1_2778 ( .gnd(gnd), .vdd(vdd), .A(data_68__13_), .Y(_6325_) );
MUX2X1 MUX2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_6325_), .B(_14924__bF_buf13), .S(_6302_), .Y(_221__13_) );
INVX1 INVX1_2779 ( .gnd(gnd), .vdd(vdd), .A(data_68__14_), .Y(_6326_) );
MUX2X1 MUX2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_6326_), .B(_15060__bF_buf10), .S(_6302_), .Y(_221__14_) );
INVX1 INVX1_2780 ( .gnd(gnd), .vdd(vdd), .A(data_68__15_), .Y(_6327_) );
MUX2X1 MUX2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_6327_), .B(_15062__bF_buf1), .S(_6302_), .Y(_221__15_) );
INVX1 INVX1_2781 ( .gnd(gnd), .vdd(vdd), .A(data_67__0_), .Y(_6328_) );
OAI21X1 OAI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf1), .B(_3322_), .C(_6179_), .Y(_6329_) );
NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_6329_), .B(_5420__bF_buf2), .Y(_6330_) );
INVX4 INVX4_25 ( .gnd(gnd), .vdd(vdd), .A(_6330_), .Y(_6331_) );
OAI21X1 OAI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_6331_), .C(_6328_), .Y(_6332_) );
NAND3X1 NAND3X1_871 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_6330_), .C(_3313__bF_buf26), .Y(_6333_) );
AND2X2 AND2X2_1213 ( .gnd(gnd), .vdd(vdd), .A(_6332_), .B(_6333_), .Y(_220__0_) );
INVX1 INVX1_2782 ( .gnd(gnd), .vdd(vdd), .A(data_67__1_), .Y(_6334_) );
OAI21X1 OAI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_6331_), .C(_6334_), .Y(_6335_) );
NAND3X1 NAND3X1_872 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_6330_), .C(_3313__bF_buf25), .Y(_6336_) );
AND2X2 AND2X2_1214 ( .gnd(gnd), .vdd(vdd), .A(_6335_), .B(_6336_), .Y(_220__1_) );
INVX1 INVX1_2783 ( .gnd(gnd), .vdd(vdd), .A(data_67__2_), .Y(_6337_) );
NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_6330_), .B(_3313__bF_buf24), .Y(_6338_) );
MUX2X1 MUX2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_6337_), .B(_14897__bF_buf5), .S(_6338_), .Y(_220__2_) );
INVX1 INVX1_2784 ( .gnd(gnd), .vdd(vdd), .A(data_67__3_), .Y(_6339_) );
OAI21X1 OAI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_6331_), .C(_6339_), .Y(_6340_) );
NAND3X1 NAND3X1_873 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_6330_), .C(_3313__bF_buf23), .Y(_6341_) );
AND2X2 AND2X2_1215 ( .gnd(gnd), .vdd(vdd), .A(_6340_), .B(_6341_), .Y(_220__3_) );
INVX1 INVX1_2785 ( .gnd(gnd), .vdd(vdd), .A(data_67__4_), .Y(_6342_) );
OAI21X1 OAI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_6331_), .C(_6342_), .Y(_6343_) );
NAND3X1 NAND3X1_874 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_6330_), .C(_3313__bF_buf22), .Y(_6344_) );
AND2X2 AND2X2_1216 ( .gnd(gnd), .vdd(vdd), .A(_6343_), .B(_6344_), .Y(_220__4_) );
INVX1 INVX1_2786 ( .gnd(gnd), .vdd(vdd), .A(data_67__5_), .Y(_6345_) );
OAI21X1 OAI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_6331_), .C(_6345_), .Y(_6346_) );
NAND3X1 NAND3X1_875 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_6330_), .C(_3313__bF_buf21), .Y(_6347_) );
AND2X2 AND2X2_1217 ( .gnd(gnd), .vdd(vdd), .A(_6346_), .B(_6347_), .Y(_220__5_) );
INVX1 INVX1_2787 ( .gnd(gnd), .vdd(vdd), .A(data_67__6_), .Y(_6348_) );
MUX2X1 MUX2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_6348_), .B(_15049__bF_buf7), .S(_6338_), .Y(_220__6_) );
INVX1 INVX1_2788 ( .gnd(gnd), .vdd(vdd), .A(data_67__7_), .Y(_6349_) );
OAI21X1 OAI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_6331_), .C(_6349_), .Y(_6350_) );
NAND3X1 NAND3X1_876 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_6330_), .C(_3313__bF_buf20), .Y(_6351_) );
AND2X2 AND2X2_1218 ( .gnd(gnd), .vdd(vdd), .A(_6350_), .B(_6351_), .Y(_220__7_) );
INVX1 INVX1_2789 ( .gnd(gnd), .vdd(vdd), .A(data_67__8_), .Y(_6352_) );
MUX2X1 MUX2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_6352_), .B(_15052__bF_buf12), .S(_6338_), .Y(_220__8_) );
INVX1 INVX1_2790 ( .gnd(gnd), .vdd(vdd), .A(data_67__9_), .Y(_6353_) );
MUX2X1 MUX2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_6353_), .B(_14913__bF_buf8), .S(_6338_), .Y(_220__9_) );
INVX1 INVX1_2791 ( .gnd(gnd), .vdd(vdd), .A(data_67__10_), .Y(_6354_) );
MUX2X1 MUX2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_6354_), .B(_15055__bF_buf0), .S(_6338_), .Y(_220__10_) );
INVX1 INVX1_2792 ( .gnd(gnd), .vdd(vdd), .A(data_67__11_), .Y(_6355_) );
OAI21X1 OAI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_6331_), .C(_6355_), .Y(_6356_) );
NAND3X1 NAND3X1_877 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_6330_), .C(_3313__bF_buf19), .Y(_6357_) );
AND2X2 AND2X2_1219 ( .gnd(gnd), .vdd(vdd), .A(_6356_), .B(_6357_), .Y(_220__11_) );
INVX1 INVX1_2793 ( .gnd(gnd), .vdd(vdd), .A(data_67__12_), .Y(_6358_) );
OAI21X1 OAI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_6331_), .C(_6358_), .Y(_6359_) );
NAND3X1 NAND3X1_878 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_6330_), .C(_3313__bF_buf18), .Y(_6360_) );
AND2X2 AND2X2_1220 ( .gnd(gnd), .vdd(vdd), .A(_6359_), .B(_6360_), .Y(_220__12_) );
INVX1 INVX1_2794 ( .gnd(gnd), .vdd(vdd), .A(data_67__13_), .Y(_6361_) );
MUX2X1 MUX2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_6361_), .B(_14924__bF_buf12), .S(_6338_), .Y(_220__13_) );
INVX1 INVX1_2795 ( .gnd(gnd), .vdd(vdd), .A(data_67__14_), .Y(_6362_) );
MUX2X1 MUX2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_6362_), .B(_15060__bF_buf9), .S(_6338_), .Y(_220__14_) );
INVX1 INVX1_2796 ( .gnd(gnd), .vdd(vdd), .A(data_67__15_), .Y(_6363_) );
MUX2X1 MUX2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_6363_), .B(_15062__bF_buf0), .S(_6338_), .Y(_220__15_) );
INVX1 INVX1_2797 ( .gnd(gnd), .vdd(vdd), .A(data_66__0_), .Y(_6364_) );
INVX1 INVX1_2798 ( .gnd(gnd), .vdd(vdd), .A(_6178_), .Y(_6365_) );
OAI21X1 OAI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_3322_), .C(_6365_), .Y(_6366_) );
INVX1 INVX1_2799 ( .gnd(gnd), .vdd(vdd), .A(_6366_), .Y(_6367_) );
NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_6367_), .B(_5461_), .Y(_6368_) );
NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_3322_), .Y(_6369_) );
NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_6369_), .B(_6368_), .Y(_6370_) );
NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf17), .B(_6370_), .Y(_6371_) );
MUX2X1 MUX2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_6364_), .B(_14932__bF_buf9), .S(_6371_), .Y(_219__0_) );
INVX1 INVX1_2800 ( .gnd(gnd), .vdd(vdd), .A(data_66__1_), .Y(_6372_) );
MUX2X1 MUX2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_6372_), .B(_14894__bF_buf9), .S(_6371_), .Y(_219__1_) );
AND2X2 AND2X2_1221 ( .gnd(gnd), .vdd(vdd), .A(_6370_), .B(_3313__bF_buf16), .Y(_6373_) );
AOI21X1 AOI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf15), .B(_6370_), .C(data_66__2_), .Y(_6374_) );
AOI21X1 AOI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_6373_), .C(_6374_), .Y(_219__2_) );
INVX1 INVX1_2801 ( .gnd(gnd), .vdd(vdd), .A(data_66__3_), .Y(_6375_) );
MUX2X1 MUX2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_6375_), .B(_14899__bF_buf8), .S(_6371_), .Y(_219__3_) );
INVX1 INVX1_2802 ( .gnd(gnd), .vdd(vdd), .A(data_66__4_), .Y(_6376_) );
MUX2X1 MUX2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_6376_), .B(_14902__bF_buf11), .S(_6371_), .Y(_219__4_) );
INVX1 INVX1_2803 ( .gnd(gnd), .vdd(vdd), .A(data_66__5_), .Y(_6377_) );
MUX2X1 MUX2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_6377_), .B(_14903__bF_buf13), .S(_6371_), .Y(_219__5_) );
AOI21X1 AOI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf14), .B(_6370_), .C(data_66__6_), .Y(_6378_) );
AOI21X1 AOI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_6373_), .C(_6378_), .Y(_219__6_) );
INVX1 INVX1_2804 ( .gnd(gnd), .vdd(vdd), .A(data_66__7_), .Y(_6379_) );
MUX2X1 MUX2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_6379_), .B(_14908__bF_buf13), .S(_6371_), .Y(_219__7_) );
AOI21X1 AOI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf13), .B(_6370_), .C(data_66__8_), .Y(_6380_) );
AOI21X1 AOI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_6373_), .C(_6380_), .Y(_219__8_) );
AOI21X1 AOI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf12), .B(_6370_), .C(data_66__9_), .Y(_6381_) );
AOI21X1 AOI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf7), .B(_6373_), .C(_6381_), .Y(_219__9_) );
AOI21X1 AOI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf11), .B(_6370_), .C(data_66__10_), .Y(_6382_) );
AOI21X1 AOI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf13), .B(_6373_), .C(_6382_), .Y(_219__10_) );
INVX1 INVX1_2805 ( .gnd(gnd), .vdd(vdd), .A(data_66__11_), .Y(_6383_) );
MUX2X1 MUX2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_6383_), .B(_14918__bF_buf13), .S(_6371_), .Y(_219__11_) );
INVX1 INVX1_2806 ( .gnd(gnd), .vdd(vdd), .A(data_66__12_), .Y(_6384_) );
MUX2X1 MUX2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_6384_), .B(_14920__bF_buf0), .S(_6371_), .Y(_219__12_) );
AOI21X1 AOI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf10), .B(_6370_), .C(data_66__13_), .Y(_6385_) );
AOI21X1 AOI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_6373_), .C(_6385_), .Y(_219__13_) );
AOI21X1 AOI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf9), .B(_6370_), .C(data_66__14_), .Y(_6386_) );
AOI21X1 AOI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_6373_), .C(_6386_), .Y(_219__14_) );
AOI21X1 AOI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf8), .B(_6370_), .C(data_66__15_), .Y(_6387_) );
AOI21X1 AOI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_6373_), .C(_6387_), .Y(_219__15_) );
AOI21X1 AOI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_3332_), .B(_4723_), .C(_6368_), .Y(_6388_) );
AND2X2 AND2X2_1222 ( .gnd(gnd), .vdd(vdd), .A(_6388__bF_buf3), .B(_3313__bF_buf7), .Y(_6389_) );
AOI21X1 AOI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf6), .B(_6388__bF_buf2), .C(data_65__0_), .Y(_6390_) );
AOI21X1 AOI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_6389_), .C(_6390_), .Y(_218__0_) );
AOI21X1 AOI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf5), .B(_6388__bF_buf1), .C(data_65__1_), .Y(_6391_) );
AOI21X1 AOI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_6389_), .C(_6391_), .Y(_218__1_) );
AOI21X1 AOI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf4), .B(_6388__bF_buf0), .C(data_65__2_), .Y(_6392_) );
AOI21X1 AOI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_6389_), .C(_6392_), .Y(_218__2_) );
AOI21X1 AOI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf3), .B(_6388__bF_buf3), .C(data_65__3_), .Y(_6393_) );
AOI21X1 AOI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_6389_), .C(_6393_), .Y(_218__3_) );
AOI21X1 AOI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf2), .B(_6388__bF_buf2), .C(data_65__4_), .Y(_6394_) );
AOI21X1 AOI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_6389_), .C(_6394_), .Y(_218__4_) );
AOI21X1 AOI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf1), .B(_6388__bF_buf1), .C(data_65__5_), .Y(_6395_) );
AOI21X1 AOI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_6389_), .C(_6395_), .Y(_218__5_) );
AOI21X1 AOI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf0), .B(_6388__bF_buf0), .C(data_65__6_), .Y(_6396_) );
AOI21X1 AOI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_6389_), .C(_6396_), .Y(_218__6_) );
AOI21X1 AOI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf91), .B(_6388__bF_buf3), .C(data_65__7_), .Y(_6397_) );
AOI21X1 AOI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_6389_), .C(_6397_), .Y(_218__7_) );
AOI21X1 AOI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf90), .B(_6388__bF_buf2), .C(data_65__8_), .Y(_6398_) );
AOI21X1 AOI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_6389_), .C(_6398_), .Y(_218__8_) );
AOI21X1 AOI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf89), .B(_6388__bF_buf1), .C(data_65__9_), .Y(_6399_) );
AOI21X1 AOI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_6389_), .C(_6399_), .Y(_218__9_) );
AOI21X1 AOI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf88), .B(_6388__bF_buf0), .C(data_65__10_), .Y(_6400_) );
AOI21X1 AOI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_6389_), .C(_6400_), .Y(_218__10_) );
AOI21X1 AOI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf87), .B(_6388__bF_buf3), .C(data_65__11_), .Y(_6401_) );
AOI21X1 AOI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_6389_), .C(_6401_), .Y(_218__11_) );
AOI21X1 AOI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf86), .B(_6388__bF_buf2), .C(data_65__12_), .Y(_6402_) );
AOI21X1 AOI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_6389_), .C(_6402_), .Y(_218__12_) );
AOI21X1 AOI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf85), .B(_6388__bF_buf1), .C(data_65__13_), .Y(_6403_) );
AOI21X1 AOI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_6389_), .C(_6403_), .Y(_218__13_) );
AOI21X1 AOI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf84), .B(_6388__bF_buf0), .C(data_65__14_), .Y(_6404_) );
AOI21X1 AOI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_6389_), .C(_6404_), .Y(_218__14_) );
AOI21X1 AOI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf83), .B(_6388__bF_buf3), .C(data_65__15_), .Y(_6405_) );
AOI21X1 AOI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_6389_), .C(_6405_), .Y(_218__15_) );
NOR3X1 NOR3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf3), .B(_15030_), .C(_3322_), .Y(_6406_) );
NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_6406_), .Y(_6407_) );
OAI21X1 OAI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(data_64__0_), .B(_6406_), .C(_6407_), .Y(_6408_) );
INVX1 INVX1_2807 ( .gnd(gnd), .vdd(vdd), .A(_6408_), .Y(_217__0_) );
INVX4 INVX4_26 ( .gnd(gnd), .vdd(vdd), .A(_6406_), .Y(_6409_) );
INVX1 INVX1_2808 ( .gnd(gnd), .vdd(vdd), .A(data_64__1_), .Y(_6410_) );
NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_14986_), .B(_3332_), .Y(_6411_) );
OAI21X1 OAI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf2), .C(_6410_), .Y(_6412_) );
OAI21X1 OAI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_1_bF_buf4), .C(_6412_), .Y(_6413_) );
INVX1 INVX1_2809 ( .gnd(gnd), .vdd(vdd), .A(_6413_), .Y(_217__1_) );
NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(data_64__2_), .B(_6406_), .Y(_6414_) );
AOI21X1 AOI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_6406_), .C(_6414_), .Y(_217__2_) );
INVX1 INVX1_2810 ( .gnd(gnd), .vdd(vdd), .A(data_64__3_), .Y(_6415_) );
OAI21X1 OAI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf1), .C(_6415_), .Y(_6416_) );
OAI21X1 OAI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_3_bF_buf0), .C(_6416_), .Y(_6417_) );
INVX1 INVX1_2811 ( .gnd(gnd), .vdd(vdd), .A(_6417_), .Y(_217__3_) );
INVX1 INVX1_2812 ( .gnd(gnd), .vdd(vdd), .A(data_64__4_), .Y(_6418_) );
OAI21X1 OAI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf0), .C(_6418_), .Y(_6419_) );
OAI21X1 OAI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_4_bF_buf4), .C(_6419_), .Y(_6420_) );
INVX1 INVX1_2813 ( .gnd(gnd), .vdd(vdd), .A(_6420_), .Y(_217__4_) );
INVX1 INVX1_2814 ( .gnd(gnd), .vdd(vdd), .A(data_64__5_), .Y(_6421_) );
OAI21X1 OAI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf15_bF_buf0), .C(_6421_), .Y(_6422_) );
OAI21X1 OAI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_5_bF_buf2), .C(_6422_), .Y(_6423_) );
INVX1 INVX1_2815 ( .gnd(gnd), .vdd(vdd), .A(_6423_), .Y(_217__5_) );
INVX1 INVX1_2816 ( .gnd(gnd), .vdd(vdd), .A(data_64__6_), .Y(_6424_) );
OAI21X1 OAI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf14_bF_buf0), .C(_6424_), .Y(_6425_) );
OAI21X1 OAI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_6_bF_buf2), .C(_6425_), .Y(_6426_) );
INVX1 INVX1_2817 ( .gnd(gnd), .vdd(vdd), .A(_6426_), .Y(_217__6_) );
INVX1 INVX1_2818 ( .gnd(gnd), .vdd(vdd), .A(data_64__7_), .Y(_6427_) );
OAI21X1 OAI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf13_bF_buf0), .C(_6427_), .Y(_6428_) );
OAI21X1 OAI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_7_bF_buf1), .C(_6428_), .Y(_6429_) );
INVX1 INVX1_2819 ( .gnd(gnd), .vdd(vdd), .A(_6429_), .Y(_217__7_) );
INVX1 INVX1_2820 ( .gnd(gnd), .vdd(vdd), .A(data_64__8_), .Y(_6430_) );
OAI21X1 OAI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf12), .C(_6430_), .Y(_6431_) );
OAI21X1 OAI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_8_bF_buf4), .C(_6431_), .Y(_6432_) );
INVX1 INVX1_2821 ( .gnd(gnd), .vdd(vdd), .A(_6432_), .Y(_217__8_) );
NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_6406_), .Y(_6433_) );
OAI21X1 OAI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(data_64__9_), .B(_6406_), .C(_6433_), .Y(_6434_) );
INVX1 INVX1_2822 ( .gnd(gnd), .vdd(vdd), .A(_6434_), .Y(_217__9_) );
NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(data_64__10_), .B(_6406_), .Y(_6435_) );
NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf2), .B(_6409_), .Y(_6436_) );
NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_6435_), .B(_6436_), .Y(_217__10_) );
INVX1 INVX1_2823 ( .gnd(gnd), .vdd(vdd), .A(data_64__11_), .Y(_6437_) );
OAI21X1 OAI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf11), .C(_6437_), .Y(_6438_) );
OAI21X1 OAI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_6409_), .B(IDATA_PROG_data_11_bF_buf2), .C(_6438_), .Y(_6439_) );
INVX1 INVX1_2824 ( .gnd(gnd), .vdd(vdd), .A(_6439_), .Y(_217__11_) );
INVX1 INVX1_2825 ( .gnd(gnd), .vdd(vdd), .A(data_64__12_), .Y(_6440_) );
OAI21X1 OAI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf10), .C(_6440_), .Y(_6441_) );
NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_6406_), .Y(_6442_) );
AND2X2 AND2X2_1223 ( .gnd(gnd), .vdd(vdd), .A(_6442_), .B(_6441_), .Y(_217__12_) );
NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_6406_), .Y(_6443_) );
OAI21X1 OAI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(data_64__13_), .B(_6406_), .C(_6443_), .Y(_6444_) );
INVX1 INVX1_2826 ( .gnd(gnd), .vdd(vdd), .A(_6444_), .Y(_217__13_) );
NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_6406_), .Y(_6445_) );
OAI21X1 OAI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(data_64__14_), .B(_6406_), .C(_6445_), .Y(_6446_) );
INVX1 INVX1_2827 ( .gnd(gnd), .vdd(vdd), .A(_6446_), .Y(_217__14_) );
INVX1 INVX1_2828 ( .gnd(gnd), .vdd(vdd), .A(data_64__15_), .Y(_6447_) );
OAI21X1 OAI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_6411_), .B(_14882__bF_buf9), .C(_6447_), .Y(_6448_) );
NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_6406_), .Y(_6449_) );
AND2X2 AND2X2_1224 ( .gnd(gnd), .vdd(vdd), .A(_6449_), .B(_6448_), .Y(_217__15_) );
INVX1 INVX1_2829 ( .gnd(gnd), .vdd(vdd), .A(data_63__0_), .Y(_6450_) );
NAND3X1 NAND3X1_879 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_14888__bF_buf2), .C(_14998__bF_buf3), .Y(_6451_) );
MUX2X1 MUX2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_6450_), .B(_14932__bF_buf6), .S(_6451_), .Y(_216__0_) );
INVX4 INVX4_27 ( .gnd(gnd), .vdd(vdd), .A(_6451_), .Y(_6452_) );
NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(data_63__1_), .B(_6452_), .Y(_6453_) );
AOI21X1 AOI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_6452_), .C(_6453_), .Y(_216__1_) );
INVX1 INVX1_2830 ( .gnd(gnd), .vdd(vdd), .A(data_63__2_), .Y(_6454_) );
OAI21X1 OAI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf8), .C(_6454_), .Y(_6455_) );
OAI21X1 OAI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf0), .B(_6451_), .C(_6455_), .Y(_6456_) );
INVX1 INVX1_2831 ( .gnd(gnd), .vdd(vdd), .A(_6456_), .Y(_216__2_) );
INVX1 INVX1_2832 ( .gnd(gnd), .vdd(vdd), .A(data_63__3_), .Y(_6457_) );
MUX2X1 MUX2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_6457_), .B(_14899__bF_buf6), .S(_6451_), .Y(_216__3_) );
INVX1 INVX1_2833 ( .gnd(gnd), .vdd(vdd), .A(data_63__4_), .Y(_6458_) );
MUX2X1 MUX2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_6458_), .B(_14902__bF_buf9), .S(_6451_), .Y(_216__4_) );
INVX1 INVX1_2834 ( .gnd(gnd), .vdd(vdd), .A(data_63__5_), .Y(_6459_) );
OAI21X1 OAI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf7), .C(_6459_), .Y(_6460_) );
OAI21X1 OAI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf1), .B(_6451_), .C(_6460_), .Y(_6461_) );
INVX1 INVX1_2835 ( .gnd(gnd), .vdd(vdd), .A(_6461_), .Y(_216__5_) );
INVX1 INVX1_2836 ( .gnd(gnd), .vdd(vdd), .A(data_63__6_), .Y(_6462_) );
OAI21X1 OAI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf6), .C(_6462_), .Y(_6463_) );
OAI21X1 OAI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf1), .B(_6451_), .C(_6463_), .Y(_6464_) );
INVX1 INVX1_2837 ( .gnd(gnd), .vdd(vdd), .A(_6464_), .Y(_216__6_) );
INVX1 INVX1_2838 ( .gnd(gnd), .vdd(vdd), .A(data_63__7_), .Y(_6465_) );
MUX2X1 MUX2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_6465_), .B(_14908__bF_buf11), .S(_6451_), .Y(_216__7_) );
INVX1 INVX1_2839 ( .gnd(gnd), .vdd(vdd), .A(data_63__8_), .Y(_6466_) );
OAI21X1 OAI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf5), .C(_6466_), .Y(_6467_) );
NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_6452_), .Y(_6468_) );
AND2X2 AND2X2_1225 ( .gnd(gnd), .vdd(vdd), .A(_6468_), .B(_6467_), .Y(_216__8_) );
NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(data_63__9_), .B(_6452_), .Y(_6469_) );
AOI21X1 AOI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_6452_), .C(_6469_), .Y(_216__9_) );
INVX1 INVX1_2840 ( .gnd(gnd), .vdd(vdd), .A(data_63__10_), .Y(_6470_) );
MUX2X1 MUX2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_6470_), .B(_15055__bF_buf11), .S(_6451_), .Y(_216__10_) );
INVX1 INVX1_2841 ( .gnd(gnd), .vdd(vdd), .A(data_63__11_), .Y(_6471_) );
MUX2X1 MUX2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_6471_), .B(_14918__bF_buf11), .S(_6451_), .Y(_216__11_) );
INVX1 INVX1_2842 ( .gnd(gnd), .vdd(vdd), .A(data_63__12_), .Y(_6472_) );
OAI21X1 OAI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf4), .C(_6472_), .Y(_6473_) );
OAI21X1 OAI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf1), .B(_6451_), .C(_6473_), .Y(_6474_) );
INVX1 INVX1_2843 ( .gnd(gnd), .vdd(vdd), .A(_6474_), .Y(_216__12_) );
INVX1 INVX1_2844 ( .gnd(gnd), .vdd(vdd), .A(data_63__13_), .Y(_6475_) );
OAI21X1 OAI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf3), .C(_6475_), .Y(_6476_) );
OAI21X1 OAI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf4), .B(_6451_), .C(_6476_), .Y(_6477_) );
INVX1 INVX1_2845 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .Y(_216__13_) );
NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(data_63__14_), .B(_6452_), .Y(_6478_) );
AOI21X1 AOI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf5), .B(_6452_), .C(_6478_), .Y(_216__14_) );
INVX1 INVX1_2846 ( .gnd(gnd), .vdd(vdd), .A(data_63__15_), .Y(_6479_) );
OAI21X1 OAI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_14882__bF_buf2), .C(_6479_), .Y(_6480_) );
OAI21X1 OAI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf1), .B(_6451_), .C(_6480_), .Y(_6481_) );
INVX1 INVX1_2847 ( .gnd(gnd), .vdd(vdd), .A(_6481_), .Y(_216__15_) );
INVX1 INVX1_2848 ( .gnd(gnd), .vdd(vdd), .A(data_62__0_), .Y(_6482_) );
OAI21X1 OAI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_3323_), .B(IDATA_PROG_addr[5]), .C(IDATA_PROG_write_bF_buf0), .Y(_6483_) );
INVX1 INVX1_2849 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .Y(_6484_) );
OAI21X1 OAI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_3348_), .C(_6484_), .Y(_6485_) );
AOI21X1 AOI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf2), .B(_5422_), .C(_6485_), .Y(_6486_) );
NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .B(_6486_), .Y(_6487_) );
NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_5459__bF_buf3), .B(_6487_), .Y(_6488_) );
INVX4 INVX4_28 ( .gnd(gnd), .vdd(vdd), .A(_6488_), .Y(_6489_) );
OAI21X1 OAI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_6489_), .C(_6482_), .Y(_6490_) );
NAND3X1 NAND3X1_880 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_6488_), .C(_3313__bF_buf82), .Y(_6491_) );
AND2X2 AND2X2_1226 ( .gnd(gnd), .vdd(vdd), .A(_6490_), .B(_6491_), .Y(_215__0_) );
INVX1 INVX1_2850 ( .gnd(gnd), .vdd(vdd), .A(data_62__1_), .Y(_6492_) );
OAI21X1 OAI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_6489_), .C(_6492_), .Y(_6493_) );
NAND3X1 NAND3X1_881 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_6488_), .C(_3313__bF_buf81), .Y(_6494_) );
AND2X2 AND2X2_1227 ( .gnd(gnd), .vdd(vdd), .A(_6493_), .B(_6494_), .Y(_215__1_) );
INVX1 INVX1_2851 ( .gnd(gnd), .vdd(vdd), .A(data_62__2_), .Y(_6495_) );
NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_6488_), .B(_3313__bF_buf80), .Y(_6496_) );
MUX2X1 MUX2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_6495_), .B(_14897__bF_buf1), .S(_6496_), .Y(_215__2_) );
INVX1 INVX1_2852 ( .gnd(gnd), .vdd(vdd), .A(data_62__3_), .Y(_6497_) );
OAI21X1 OAI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_6489_), .C(_6497_), .Y(_6498_) );
NAND3X1 NAND3X1_882 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_6488_), .C(_3313__bF_buf79), .Y(_6499_) );
AND2X2 AND2X2_1228 ( .gnd(gnd), .vdd(vdd), .A(_6498_), .B(_6499_), .Y(_215__3_) );
INVX1 INVX1_2853 ( .gnd(gnd), .vdd(vdd), .A(data_62__4_), .Y(_6500_) );
OAI21X1 OAI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_6489_), .C(_6500_), .Y(_6501_) );
NAND3X1 NAND3X1_883 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_6488_), .C(_3313__bF_buf78), .Y(_6502_) );
AND2X2 AND2X2_1229 ( .gnd(gnd), .vdd(vdd), .A(_6501_), .B(_6502_), .Y(_215__4_) );
INVX1 INVX1_2854 ( .gnd(gnd), .vdd(vdd), .A(data_62__5_), .Y(_6503_) );
OAI21X1 OAI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_6489_), .C(_6503_), .Y(_6504_) );
NAND3X1 NAND3X1_884 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_6488_), .C(_3313__bF_buf77), .Y(_6505_) );
AND2X2 AND2X2_1230 ( .gnd(gnd), .vdd(vdd), .A(_6504_), .B(_6505_), .Y(_215__5_) );
INVX1 INVX1_2855 ( .gnd(gnd), .vdd(vdd), .A(data_62__6_), .Y(_6506_) );
MUX2X1 MUX2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_6506_), .B(_15049__bF_buf4), .S(_6496_), .Y(_215__6_) );
INVX1 INVX1_2856 ( .gnd(gnd), .vdd(vdd), .A(data_62__7_), .Y(_6507_) );
OAI21X1 OAI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_6489_), .C(_6507_), .Y(_6508_) );
NAND3X1 NAND3X1_885 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_6488_), .C(_3313__bF_buf76), .Y(_6509_) );
AND2X2 AND2X2_1231 ( .gnd(gnd), .vdd(vdd), .A(_6508_), .B(_6509_), .Y(_215__7_) );
INVX1 INVX1_2857 ( .gnd(gnd), .vdd(vdd), .A(data_62__8_), .Y(_6510_) );
MUX2X1 MUX2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_6510_), .B(_15052__bF_buf8), .S(_6496_), .Y(_215__8_) );
INVX1 INVX1_2858 ( .gnd(gnd), .vdd(vdd), .A(data_62__9_), .Y(_6511_) );
MUX2X1 MUX2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_6511_), .B(_14913__bF_buf3), .S(_6496_), .Y(_215__9_) );
INVX1 INVX1_2859 ( .gnd(gnd), .vdd(vdd), .A(data_62__10_), .Y(_6512_) );
MUX2X1 MUX2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_6512_), .B(_15055__bF_buf10), .S(_6496_), .Y(_215__10_) );
INVX1 INVX1_2860 ( .gnd(gnd), .vdd(vdd), .A(data_62__11_), .Y(_6513_) );
OAI21X1 OAI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_6489_), .C(_6513_), .Y(_6514_) );
NAND3X1 NAND3X1_886 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_6488_), .C(_3313__bF_buf75), .Y(_6515_) );
AND2X2 AND2X2_1232 ( .gnd(gnd), .vdd(vdd), .A(_6514_), .B(_6515_), .Y(_215__11_) );
INVX1 INVX1_2861 ( .gnd(gnd), .vdd(vdd), .A(data_62__12_), .Y(_6516_) );
OAI21X1 OAI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_6489_), .C(_6516_), .Y(_6517_) );
NAND3X1 NAND3X1_887 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_6488_), .C(_3313__bF_buf74), .Y(_6518_) );
AND2X2 AND2X2_1233 ( .gnd(gnd), .vdd(vdd), .A(_6517_), .B(_6518_), .Y(_215__12_) );
INVX1 INVX1_2862 ( .gnd(gnd), .vdd(vdd), .A(data_62__13_), .Y(_6519_) );
MUX2X1 MUX2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_6519_), .B(_14924__bF_buf8), .S(_6496_), .Y(_215__13_) );
INVX1 INVX1_2863 ( .gnd(gnd), .vdd(vdd), .A(data_62__14_), .Y(_6520_) );
MUX2X1 MUX2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_6520_), .B(_15060__bF_buf4), .S(_6496_), .Y(_215__14_) );
INVX1 INVX1_2864 ( .gnd(gnd), .vdd(vdd), .A(data_62__15_), .Y(_6521_) );
MUX2X1 MUX2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_6521_), .B(_15062__bF_buf10), .S(_6496_), .Y(_215__15_) );
INVX1 INVX1_2865 ( .gnd(gnd), .vdd(vdd), .A(data_61__0_), .Y(_6522_) );
OAI21X1 OAI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_5463_), .B(_3348_), .C(_3351_), .Y(_6523_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_5459__bF_buf2), .B(_6523_), .Y(_6524_) );
NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_6485_), .B(_6524_), .Y(_6525_) );
NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_6525_), .B(_3313__bF_buf73), .Y(_6526_) );
MUX2X1 MUX2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_6522_), .B(_14932__bF_buf4), .S(_6526_), .Y(_214__0_) );
INVX1 INVX1_2866 ( .gnd(gnd), .vdd(vdd), .A(data_61__1_), .Y(_6527_) );
MUX2X1 MUX2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_6527_), .B(_14894__bF_buf5), .S(_6526_), .Y(_214__1_) );
INVX1 INVX1_2867 ( .gnd(gnd), .vdd(vdd), .A(data_61__2_), .Y(_6528_) );
MUX2X1 MUX2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_6528_), .B(_14897__bF_buf0), .S(_6526_), .Y(_214__2_) );
INVX1 INVX1_2868 ( .gnd(gnd), .vdd(vdd), .A(data_61__3_), .Y(_6529_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_6524_), .B(_6485_), .Y(_6530_) );
OAI21X1 OAI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_6530_), .C(_6529_), .Y(_6531_) );
NAND3X1 NAND3X1_888 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_6525_), .C(_3313__bF_buf72), .Y(_6532_) );
AND2X2 AND2X2_1234 ( .gnd(gnd), .vdd(vdd), .A(_6531_), .B(_6532_), .Y(_214__3_) );
INVX1 INVX1_2869 ( .gnd(gnd), .vdd(vdd), .A(data_61__4_), .Y(_6533_) );
OAI21X1 OAI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_6530_), .C(_6533_), .Y(_6534_) );
NAND3X1 NAND3X1_889 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_6525_), .C(_3313__bF_buf71), .Y(_6535_) );
AND2X2 AND2X2_1235 ( .gnd(gnd), .vdd(vdd), .A(_6534_), .B(_6535_), .Y(_214__4_) );
INVX1 INVX1_2870 ( .gnd(gnd), .vdd(vdd), .A(data_61__5_), .Y(_6536_) );
OAI21X1 OAI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_6530_), .C(_6536_), .Y(_6537_) );
NAND3X1 NAND3X1_890 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_6525_), .C(_3313__bF_buf70), .Y(_6538_) );
AND2X2 AND2X2_1236 ( .gnd(gnd), .vdd(vdd), .A(_6537_), .B(_6538_), .Y(_214__5_) );
INVX1 INVX1_2871 ( .gnd(gnd), .vdd(vdd), .A(data_61__6_), .Y(_6539_) );
MUX2X1 MUX2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_6539_), .B(_15049__bF_buf3), .S(_6526_), .Y(_214__6_) );
INVX1 INVX1_2872 ( .gnd(gnd), .vdd(vdd), .A(data_61__7_), .Y(_6540_) );
OAI21X1 OAI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_6530_), .C(_6540_), .Y(_6541_) );
NAND3X1 NAND3X1_891 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_6525_), .C(_3313__bF_buf69), .Y(_6542_) );
AND2X2 AND2X2_1237 ( .gnd(gnd), .vdd(vdd), .A(_6541_), .B(_6542_), .Y(_214__7_) );
INVX1 INVX1_2873 ( .gnd(gnd), .vdd(vdd), .A(data_61__8_), .Y(_6543_) );
MUX2X1 MUX2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_6543_), .B(_15052__bF_buf7), .S(_6526_), .Y(_214__8_) );
INVX1 INVX1_2874 ( .gnd(gnd), .vdd(vdd), .A(data_61__9_), .Y(_6544_) );
MUX2X1 MUX2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_6544_), .B(_14913__bF_buf2), .S(_6526_), .Y(_214__9_) );
INVX1 INVX1_2875 ( .gnd(gnd), .vdd(vdd), .A(data_61__10_), .Y(_6545_) );
MUX2X1 MUX2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_6545_), .B(_15055__bF_buf9), .S(_6526_), .Y(_214__10_) );
INVX1 INVX1_2876 ( .gnd(gnd), .vdd(vdd), .A(data_61__11_), .Y(_6546_) );
OAI21X1 OAI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_6530_), .C(_6546_), .Y(_6547_) );
NAND3X1 NAND3X1_892 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_6525_), .C(_3313__bF_buf68), .Y(_6548_) );
AND2X2 AND2X2_1238 ( .gnd(gnd), .vdd(vdd), .A(_6547_), .B(_6548_), .Y(_214__11_) );
INVX1 INVX1_2877 ( .gnd(gnd), .vdd(vdd), .A(data_61__12_), .Y(_6549_) );
OAI21X1 OAI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_6530_), .C(_6549_), .Y(_6550_) );
NAND3X1 NAND3X1_893 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_6525_), .C(_3313__bF_buf67), .Y(_6551_) );
AND2X2 AND2X2_1239 ( .gnd(gnd), .vdd(vdd), .A(_6550_), .B(_6551_), .Y(_214__12_) );
INVX1 INVX1_2878 ( .gnd(gnd), .vdd(vdd), .A(data_61__13_), .Y(_6552_) );
MUX2X1 MUX2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_6552_), .B(_14924__bF_buf7), .S(_6526_), .Y(_214__13_) );
INVX1 INVX1_2879 ( .gnd(gnd), .vdd(vdd), .A(data_61__14_), .Y(_6553_) );
MUX2X1 MUX2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_6553_), .B(_15060__bF_buf3), .S(_6526_), .Y(_214__14_) );
INVX1 INVX1_2880 ( .gnd(gnd), .vdd(vdd), .A(data_61__15_), .Y(_6554_) );
MUX2X1 MUX2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_6554_), .B(_15062__bF_buf9), .S(_6526_), .Y(_214__15_) );
INVX1 INVX1_2881 ( .gnd(gnd), .vdd(vdd), .A(data_60__0_), .Y(_6555_) );
NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_5459__bF_buf1), .B(_6523_), .Y(_6556_) );
AOI21X1 AOI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf1), .B(_3715_), .C(_6483_), .Y(_6557_) );
NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_6557_), .B(_6556_), .Y(_6558_) );
OAI21X1 OAI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_6558_), .C(_6555_), .Y(_6559_) );
AND2X2 AND2X2_1240 ( .gnd(gnd), .vdd(vdd), .A(_6556_), .B(_6557_), .Y(_6560_) );
NAND3X1 NAND3X1_894 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_6560_), .C(_3313__bF_buf66), .Y(_6561_) );
AND2X2 AND2X2_1241 ( .gnd(gnd), .vdd(vdd), .A(_6559_), .B(_6561_), .Y(_213__0_) );
INVX1 INVX1_2882 ( .gnd(gnd), .vdd(vdd), .A(data_60__1_), .Y(_6562_) );
OAI21X1 OAI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_6558_), .C(_6562_), .Y(_6563_) );
NAND3X1 NAND3X1_895 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_6560_), .C(_3313__bF_buf65), .Y(_6564_) );
AND2X2 AND2X2_1242 ( .gnd(gnd), .vdd(vdd), .A(_6563_), .B(_6564_), .Y(_213__1_) );
INVX1 INVX1_2883 ( .gnd(gnd), .vdd(vdd), .A(data_60__2_), .Y(_6565_) );
NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(_3313__bF_buf64), .Y(_6566_) );
MUX2X1 MUX2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_6565_), .B(_14897__bF_buf14), .S(_6566_), .Y(_213__2_) );
INVX1 INVX1_2884 ( .gnd(gnd), .vdd(vdd), .A(data_60__3_), .Y(_6567_) );
MUX2X1 MUX2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_6567_), .B(_14899__bF_buf3), .S(_6566_), .Y(_213__3_) );
INVX1 INVX1_2885 ( .gnd(gnd), .vdd(vdd), .A(data_60__4_), .Y(_6568_) );
MUX2X1 MUX2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_6568_), .B(_14902__bF_buf6), .S(_6566_), .Y(_213__4_) );
INVX1 INVX1_2886 ( .gnd(gnd), .vdd(vdd), .A(data_60__5_), .Y(_6569_) );
OAI21X1 OAI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_6558_), .C(_6569_), .Y(_6570_) );
NAND3X1 NAND3X1_896 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_6560_), .C(_3313__bF_buf63), .Y(_6571_) );
AND2X2 AND2X2_1243 ( .gnd(gnd), .vdd(vdd), .A(_6570_), .B(_6571_), .Y(_213__5_) );
INVX1 INVX1_2887 ( .gnd(gnd), .vdd(vdd), .A(data_60__6_), .Y(_6572_) );
MUX2X1 MUX2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_6572_), .B(_15049__bF_buf2), .S(_6566_), .Y(_213__6_) );
INVX1 INVX1_2888 ( .gnd(gnd), .vdd(vdd), .A(data_60__7_), .Y(_6573_) );
OAI21X1 OAI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_6558_), .C(_6573_), .Y(_6574_) );
NAND3X1 NAND3X1_897 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_6560_), .C(_3313__bF_buf62), .Y(_6575_) );
AND2X2 AND2X2_1244 ( .gnd(gnd), .vdd(vdd), .A(_6574_), .B(_6575_), .Y(_213__7_) );
NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_6558_), .B(_3393__bF_buf34), .Y(_6576_) );
AOI21X1 AOI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(_3313__bF_buf61), .C(data_60__8_), .Y(_6577_) );
AOI21X1 AOI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_6576_), .C(_6577_), .Y(_213__8_) );
AOI21X1 AOI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(_3313__bF_buf60), .C(data_60__9_), .Y(_6578_) );
AOI21X1 AOI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_6576_), .C(_6578_), .Y(_213__9_) );
AOI21X1 AOI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(_3313__bF_buf59), .C(data_60__10_), .Y(_6579_) );
AOI21X1 AOI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_6576_), .C(_6579_), .Y(_213__10_) );
INVX1 INVX1_2889 ( .gnd(gnd), .vdd(vdd), .A(data_60__11_), .Y(_6580_) );
MUX2X1 MUX2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_6580_), .B(_14918__bF_buf8), .S(_6566_), .Y(_213__11_) );
INVX1 INVX1_2890 ( .gnd(gnd), .vdd(vdd), .A(data_60__12_), .Y(_6581_) );
OAI21X1 OAI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_6558_), .C(_6581_), .Y(_6582_) );
NAND3X1 NAND3X1_898 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_6560_), .C(_3313__bF_buf58), .Y(_6583_) );
AND2X2 AND2X2_1245 ( .gnd(gnd), .vdd(vdd), .A(_6582_), .B(_6583_), .Y(_213__12_) );
AOI21X1 AOI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_6560_), .B(_3313__bF_buf57), .C(data_60__13_), .Y(_6584_) );
AOI21X1 AOI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_6576_), .C(_6584_), .Y(_213__13_) );
INVX1 INVX1_2891 ( .gnd(gnd), .vdd(vdd), .A(data_60__14_), .Y(_6585_) );
MUX2X1 MUX2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_6585_), .B(_15060__bF_buf2), .S(_6566_), .Y(_213__14_) );
INVX1 INVX1_2892 ( .gnd(gnd), .vdd(vdd), .A(data_60__15_), .Y(_6586_) );
MUX2X1 MUX2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_6586_), .B(_15062__bF_buf8), .S(_6566_), .Y(_213__15_) );
INVX1 INVX1_2893 ( .gnd(gnd), .vdd(vdd), .A(data_59__0_), .Y(_6587_) );
OAI21X1 OAI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_14990_), .C(_14998__bF_buf0), .Y(_6588_) );
AOI21X1 AOI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf0), .B(_14998__bF_buf3), .C(_6483_), .Y(_6589_) );
NAND3X1 NAND3X1_899 ( .gnd(gnd), .vdd(vdd), .A(_6588_), .B(_6589_), .C(_3351_), .Y(_6590_) );
NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_5459__bF_buf0), .B(_6590_), .Y(_6591_) );
INVX4 INVX4_29 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .Y(_6592_) );
OAI21X1 OAI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_6592_), .C(_6587_), .Y(_6593_) );
NAND3X1 NAND3X1_900 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_6591_), .C(_3313__bF_buf56), .Y(_6594_) );
AND2X2 AND2X2_1246 ( .gnd(gnd), .vdd(vdd), .A(_6593_), .B(_6594_), .Y(_211__0_) );
INVX1 INVX1_2894 ( .gnd(gnd), .vdd(vdd), .A(data_59__1_), .Y(_6595_) );
OAI21X1 OAI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_6592_), .C(_6595_), .Y(_6596_) );
NAND3X1 NAND3X1_901 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_6591_), .C(_3313__bF_buf55), .Y(_6597_) );
AND2X2 AND2X2_1247 ( .gnd(gnd), .vdd(vdd), .A(_6596_), .B(_6597_), .Y(_211__1_) );
INVX1 INVX1_2895 ( .gnd(gnd), .vdd(vdd), .A(data_59__2_), .Y(_6598_) );
NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_6591_), .B(_3313__bF_buf54), .Y(_6599_) );
MUX2X1 MUX2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_6598_), .B(_14897__bF_buf13), .S(_6599_), .Y(_211__2_) );
INVX1 INVX1_2896 ( .gnd(gnd), .vdd(vdd), .A(data_59__3_), .Y(_6600_) );
OAI21X1 OAI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_6592_), .C(_6600_), .Y(_6601_) );
NAND3X1 NAND3X1_902 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_6591_), .C(_3313__bF_buf53), .Y(_6602_) );
AND2X2 AND2X2_1248 ( .gnd(gnd), .vdd(vdd), .A(_6601_), .B(_6602_), .Y(_211__3_) );
INVX1 INVX1_2897 ( .gnd(gnd), .vdd(vdd), .A(data_59__4_), .Y(_6603_) );
OAI21X1 OAI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_6592_), .C(_6603_), .Y(_6604_) );
NAND3X1 NAND3X1_903 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_6591_), .C(_3313__bF_buf52), .Y(_6605_) );
AND2X2 AND2X2_1249 ( .gnd(gnd), .vdd(vdd), .A(_6604_), .B(_6605_), .Y(_211__4_) );
INVX1 INVX1_2898 ( .gnd(gnd), .vdd(vdd), .A(data_59__5_), .Y(_6606_) );
OAI21X1 OAI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_6592_), .C(_6606_), .Y(_6607_) );
NAND3X1 NAND3X1_904 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_6591_), .C(_3313__bF_buf51), .Y(_6608_) );
AND2X2 AND2X2_1250 ( .gnd(gnd), .vdd(vdd), .A(_6607_), .B(_6608_), .Y(_211__5_) );
INVX1 INVX1_2899 ( .gnd(gnd), .vdd(vdd), .A(data_59__6_), .Y(_6609_) );
MUX2X1 MUX2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_6609_), .B(_15049__bF_buf1), .S(_6599_), .Y(_211__6_) );
INVX1 INVX1_2900 ( .gnd(gnd), .vdd(vdd), .A(data_59__7_), .Y(_6610_) );
OAI21X1 OAI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_6592_), .C(_6610_), .Y(_6611_) );
NAND3X1 NAND3X1_905 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_6591_), .C(_3313__bF_buf50), .Y(_6612_) );
AND2X2 AND2X2_1251 ( .gnd(gnd), .vdd(vdd), .A(_6611_), .B(_6612_), .Y(_211__7_) );
INVX1 INVX1_2901 ( .gnd(gnd), .vdd(vdd), .A(data_59__8_), .Y(_6613_) );
MUX2X1 MUX2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_6613_), .B(_15052__bF_buf5), .S(_6599_), .Y(_211__8_) );
INVX1 INVX1_2902 ( .gnd(gnd), .vdd(vdd), .A(data_59__9_), .Y(_6614_) );
MUX2X1 MUX2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_6614_), .B(_14913__bF_buf0), .S(_6599_), .Y(_211__9_) );
INVX1 INVX1_2903 ( .gnd(gnd), .vdd(vdd), .A(data_59__10_), .Y(_6615_) );
MUX2X1 MUX2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_6615_), .B(_15055__bF_buf7), .S(_6599_), .Y(_211__10_) );
INVX1 INVX1_2904 ( .gnd(gnd), .vdd(vdd), .A(data_59__11_), .Y(_6616_) );
OAI21X1 OAI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_6592_), .C(_6616_), .Y(_6617_) );
NAND3X1 NAND3X1_906 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_6591_), .C(_3313__bF_buf49), .Y(_6618_) );
AND2X2 AND2X2_1252 ( .gnd(gnd), .vdd(vdd), .A(_6617_), .B(_6618_), .Y(_211__11_) );
INVX1 INVX1_2905 ( .gnd(gnd), .vdd(vdd), .A(data_59__12_), .Y(_6619_) );
OAI21X1 OAI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_6592_), .C(_6619_), .Y(_6620_) );
NAND3X1 NAND3X1_907 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_6591_), .C(_3313__bF_buf48), .Y(_6621_) );
AND2X2 AND2X2_1253 ( .gnd(gnd), .vdd(vdd), .A(_6620_), .B(_6621_), .Y(_211__12_) );
INVX1 INVX1_2906 ( .gnd(gnd), .vdd(vdd), .A(data_59__13_), .Y(_6622_) );
MUX2X1 MUX2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_6622_), .B(_14924__bF_buf5), .S(_6599_), .Y(_211__13_) );
INVX1 INVX1_2907 ( .gnd(gnd), .vdd(vdd), .A(data_59__14_), .Y(_6623_) );
MUX2X1 MUX2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_6623_), .B(_15060__bF_buf1), .S(_6599_), .Y(_211__14_) );
INVX1 INVX1_2908 ( .gnd(gnd), .vdd(vdd), .A(data_59__15_), .Y(_6624_) );
MUX2X1 MUX2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_6624_), .B(_15062__bF_buf7), .S(_6599_), .Y(_211__15_) );
INVX1 INVX1_2909 ( .gnd(gnd), .vdd(vdd), .A(data_58__0_), .Y(_6625_) );
NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf2), .B(_14996_), .Y(_6626_) );
INVX1 INVX1_2910 ( .gnd(gnd), .vdd(vdd), .A(_6626_), .Y(_6627_) );
OAI21X1 OAI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_3784_), .B(_3348_), .C(_6589_), .Y(_6628_) );
NOR2X1 NOR2X1_722 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .B(_6628_), .Y(_6629_) );
AND2X2 AND2X2_1254 ( .gnd(gnd), .vdd(vdd), .A(_6629_), .B(_3351_), .Y(_6630_) );
NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_6630_), .Y(_6631_) );
OAI21X1 OAI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf24), .B(_6631_), .C(_6625_), .Y(_6632_) );
INVX4 INVX4_30 ( .gnd(gnd), .vdd(vdd), .A(_6631_), .Y(_6633_) );
NAND3X1 NAND3X1_908 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_6633_), .C(_3313__bF_buf47), .Y(_6634_) );
AND2X2 AND2X2_1255 ( .gnd(gnd), .vdd(vdd), .A(_6632_), .B(_6634_), .Y(_210__0_) );
INVX1 INVX1_2911 ( .gnd(gnd), .vdd(vdd), .A(data_58__1_), .Y(_6635_) );
OAI21X1 OAI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_6631_), .C(_6635_), .Y(_6636_) );
NAND3X1 NAND3X1_909 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_6633_), .C(_3313__bF_buf46), .Y(_6637_) );
AND2X2 AND2X2_1256 ( .gnd(gnd), .vdd(vdd), .A(_6636_), .B(_6637_), .Y(_210__1_) );
INVX1 INVX1_2912 ( .gnd(gnd), .vdd(vdd), .A(data_58__2_), .Y(_6638_) );
NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_6633_), .B(_3313__bF_buf45), .Y(_6639_) );
MUX2X1 MUX2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_6638_), .B(_14897__bF_buf12), .S(_6639_), .Y(_210__2_) );
INVX1 INVX1_2913 ( .gnd(gnd), .vdd(vdd), .A(data_58__3_), .Y(_6640_) );
OAI21X1 OAI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_6631_), .C(_6640_), .Y(_6641_) );
NAND3X1 NAND3X1_910 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_6633_), .C(_3313__bF_buf44), .Y(_6642_) );
AND2X2 AND2X2_1257 ( .gnd(gnd), .vdd(vdd), .A(_6641_), .B(_6642_), .Y(_210__3_) );
INVX1 INVX1_2914 ( .gnd(gnd), .vdd(vdd), .A(data_58__4_), .Y(_6643_) );
OAI21X1 OAI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_6631_), .C(_6643_), .Y(_6644_) );
NAND3X1 NAND3X1_911 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_6633_), .C(_3313__bF_buf43), .Y(_6645_) );
AND2X2 AND2X2_1258 ( .gnd(gnd), .vdd(vdd), .A(_6644_), .B(_6645_), .Y(_210__4_) );
INVX1 INVX1_2915 ( .gnd(gnd), .vdd(vdd), .A(data_58__5_), .Y(_6646_) );
OAI21X1 OAI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf20), .B(_6631_), .C(_6646_), .Y(_6647_) );
NAND3X1 NAND3X1_912 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_6633_), .C(_3313__bF_buf42), .Y(_6648_) );
AND2X2 AND2X2_1259 ( .gnd(gnd), .vdd(vdd), .A(_6647_), .B(_6648_), .Y(_210__5_) );
INVX1 INVX1_2916 ( .gnd(gnd), .vdd(vdd), .A(data_58__6_), .Y(_6649_) );
MUX2X1 MUX2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_6649_), .B(_15049__bF_buf0), .S(_6639_), .Y(_210__6_) );
INVX1 INVX1_2917 ( .gnd(gnd), .vdd(vdd), .A(data_58__7_), .Y(_6650_) );
OAI21X1 OAI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf19), .B(_6631_), .C(_6650_), .Y(_6651_) );
NAND3X1 NAND3X1_913 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_6633_), .C(_3313__bF_buf41), .Y(_6652_) );
AND2X2 AND2X2_1260 ( .gnd(gnd), .vdd(vdd), .A(_6651_), .B(_6652_), .Y(_210__7_) );
INVX1 INVX1_2918 ( .gnd(gnd), .vdd(vdd), .A(data_58__8_), .Y(_6653_) );
MUX2X1 MUX2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_6653_), .B(_15052__bF_buf4), .S(_6639_), .Y(_210__8_) );
INVX1 INVX1_2919 ( .gnd(gnd), .vdd(vdd), .A(data_58__9_), .Y(_6654_) );
MUX2X1 MUX2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_6654_), .B(_14913__bF_buf14), .S(_6639_), .Y(_210__9_) );
INVX1 INVX1_2920 ( .gnd(gnd), .vdd(vdd), .A(data_58__10_), .Y(_6655_) );
MUX2X1 MUX2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_6655_), .B(_15055__bF_buf6), .S(_6639_), .Y(_210__10_) );
INVX1 INVX1_2921 ( .gnd(gnd), .vdd(vdd), .A(data_58__11_), .Y(_6656_) );
OAI21X1 OAI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf18), .B(_6631_), .C(_6656_), .Y(_6657_) );
NAND3X1 NAND3X1_914 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_6633_), .C(_3313__bF_buf40), .Y(_6658_) );
AND2X2 AND2X2_1261 ( .gnd(gnd), .vdd(vdd), .A(_6657_), .B(_6658_), .Y(_210__11_) );
INVX1 INVX1_2922 ( .gnd(gnd), .vdd(vdd), .A(data_58__12_), .Y(_6659_) );
OAI21X1 OAI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf17), .B(_6631_), .C(_6659_), .Y(_6660_) );
NAND3X1 NAND3X1_915 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_6633_), .C(_3313__bF_buf39), .Y(_6661_) );
AND2X2 AND2X2_1262 ( .gnd(gnd), .vdd(vdd), .A(_6660_), .B(_6661_), .Y(_210__12_) );
INVX1 INVX1_2923 ( .gnd(gnd), .vdd(vdd), .A(data_58__13_), .Y(_6662_) );
MUX2X1 MUX2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_6662_), .B(_14924__bF_buf4), .S(_6639_), .Y(_210__13_) );
INVX1 INVX1_2924 ( .gnd(gnd), .vdd(vdd), .A(data_58__14_), .Y(_6663_) );
MUX2X1 MUX2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_6663_), .B(_15060__bF_buf0), .S(_6639_), .Y(_210__14_) );
INVX1 INVX1_2925 ( .gnd(gnd), .vdd(vdd), .A(data_58__15_), .Y(_6664_) );
MUX2X1 MUX2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_6664_), .B(_15062__bF_buf6), .S(_6639_), .Y(_210__15_) );
INVX1 INVX1_2926 ( .gnd(gnd), .vdd(vdd), .A(data_57__0_), .Y(_6665_) );
AOI21X1 AOI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_14886__bF_buf1), .B(_3827_), .C(_3348_), .Y(_6666_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_6666_), .B(_6483_), .Y(_6667_) );
NOR2X1 NOR2X1_723 ( .gnd(gnd), .vdd(vdd), .A(_6627_), .B(_6667_), .Y(_6668_) );
NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_3351_), .B(_6668_), .Y(_6669_) );
NOR2X1 NOR2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_5459__bF_buf3), .B(_6669_), .Y(_6670_) );
INVX4 INVX4_31 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .Y(_6671_) );
OAI21X1 OAI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf16), .B(_6671_), .C(_6665_), .Y(_6672_) );
NAND3X1 NAND3X1_916 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_6670_), .C(_3313__bF_buf38), .Y(_6673_) );
AND2X2 AND2X2_1263 ( .gnd(gnd), .vdd(vdd), .A(_6672_), .B(_6673_), .Y(_209__0_) );
INVX1 INVX1_2927 ( .gnd(gnd), .vdd(vdd), .A(data_57__1_), .Y(_6674_) );
OAI21X1 OAI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf15), .B(_6671_), .C(_6674_), .Y(_6675_) );
NAND3X1 NAND3X1_917 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_6670_), .C(_3313__bF_buf37), .Y(_6676_) );
AND2X2 AND2X2_1264 ( .gnd(gnd), .vdd(vdd), .A(_6675_), .B(_6676_), .Y(_209__1_) );
NOR2X1 NOR2X1_725 ( .gnd(gnd), .vdd(vdd), .A(_6671_), .B(_3393__bF_buf14), .Y(_6677_) );
AOI21X1 AOI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .B(_3313__bF_buf36), .C(data_57__2_), .Y(_6678_) );
AOI21X1 AOI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_6677_), .C(_6678_), .Y(_209__2_) );
INVX1 INVX1_2928 ( .gnd(gnd), .vdd(vdd), .A(data_57__3_), .Y(_6679_) );
OAI21X1 OAI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf13), .B(_6671_), .C(_6679_), .Y(_6680_) );
NAND3X1 NAND3X1_918 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_6670_), .C(_3313__bF_buf35), .Y(_6681_) );
AND2X2 AND2X2_1265 ( .gnd(gnd), .vdd(vdd), .A(_6680_), .B(_6681_), .Y(_209__3_) );
INVX1 INVX1_2929 ( .gnd(gnd), .vdd(vdd), .A(data_57__4_), .Y(_6682_) );
OAI21X1 OAI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_6671_), .C(_6682_), .Y(_6683_) );
NAND3X1 NAND3X1_919 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_6670_), .C(_3313__bF_buf34), .Y(_6684_) );
AND2X2 AND2X2_1266 ( .gnd(gnd), .vdd(vdd), .A(_6683_), .B(_6684_), .Y(_209__4_) );
INVX1 INVX1_2930 ( .gnd(gnd), .vdd(vdd), .A(data_57__5_), .Y(_6685_) );
NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .B(_3313__bF_buf33), .Y(_6686_) );
MUX2X1 MUX2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_6685_), .B(_14903__bF_buf6), .S(_6686_), .Y(_209__5_) );
AOI21X1 AOI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .B(_3313__bF_buf32), .C(data_57__6_), .Y(_6687_) );
AOI21X1 AOI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_6677_), .C(_6687_), .Y(_209__6_) );
INVX1 INVX1_2931 ( .gnd(gnd), .vdd(vdd), .A(data_57__7_), .Y(_6688_) );
MUX2X1 MUX2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_6688_), .B(_14908__bF_buf5), .S(_6686_), .Y(_209__7_) );
AOI21X1 AOI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .B(_3313__bF_buf31), .C(data_57__8_), .Y(_6689_) );
AOI21X1 AOI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_6677_), .C(_6689_), .Y(_209__8_) );
INVX1 INVX1_2932 ( .gnd(gnd), .vdd(vdd), .A(data_57__9_), .Y(_6690_) );
MUX2X1 MUX2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_6690_), .B(_14913__bF_buf13), .S(_6686_), .Y(_209__9_) );
INVX1 INVX1_2933 ( .gnd(gnd), .vdd(vdd), .A(data_57__10_), .Y(_6691_) );
MUX2X1 MUX2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_6691_), .B(_15055__bF_buf5), .S(_6686_), .Y(_209__10_) );
INVX1 INVX1_2934 ( .gnd(gnd), .vdd(vdd), .A(data_57__11_), .Y(_6692_) );
OAI21X1 OAI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_6671_), .C(_6692_), .Y(_6693_) );
NAND3X1 NAND3X1_920 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_6670_), .C(_3313__bF_buf30), .Y(_6694_) );
AND2X2 AND2X2_1267 ( .gnd(gnd), .vdd(vdd), .A(_6693_), .B(_6694_), .Y(_209__11_) );
INVX1 INVX1_2935 ( .gnd(gnd), .vdd(vdd), .A(data_57__12_), .Y(_6695_) );
MUX2X1 MUX2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_6695_), .B(_14920__bF_buf6), .S(_6686_), .Y(_209__12_) );
INVX1 INVX1_2936 ( .gnd(gnd), .vdd(vdd), .A(data_57__13_), .Y(_6696_) );
MUX2X1 MUX2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_6696_), .B(_14924__bF_buf3), .S(_6686_), .Y(_209__13_) );
AOI21X1 AOI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .B(_3313__bF_buf29), .C(data_57__14_), .Y(_6697_) );
AOI21X1 AOI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf14), .B(_6677_), .C(_6697_), .Y(_209__14_) );
AOI21X1 AOI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_6670_), .B(_3313__bF_buf28), .C(data_57__15_), .Y(_6698_) );
AOI21X1 AOI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_6677_), .C(_6698_), .Y(_209__15_) );
INVX1 INVX1_2937 ( .gnd(gnd), .vdd(vdd), .A(data_56__0_), .Y(_6699_) );
AOI21X1 AOI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf1), .B(_4467_), .C(_6667_), .Y(_6700_) );
AND2X2 AND2X2_1268 ( .gnd(gnd), .vdd(vdd), .A(_6700_), .B(_3351_), .Y(_6701_) );
NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_14973_), .B(_6701_), .Y(_6702_) );
OAI21X1 OAI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_6702_), .C(_6699_), .Y(_6703_) );
INVX8 INVX8_31 ( .gnd(gnd), .vdd(vdd), .A(_6702_), .Y(_6704_) );
NAND3X1 NAND3X1_921 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_6704_), .C(_3313__bF_buf27), .Y(_6705_) );
AND2X2 AND2X2_1269 ( .gnd(gnd), .vdd(vdd), .A(_6703_), .B(_6705_), .Y(_208__0_) );
INVX1 INVX1_2938 ( .gnd(gnd), .vdd(vdd), .A(data_56__1_), .Y(_6706_) );
OAI21X1 OAI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_6702_), .C(_6706_), .Y(_6707_) );
NAND3X1 NAND3X1_922 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_6704_), .C(_3313__bF_buf26), .Y(_6708_) );
AND2X2 AND2X2_1270 ( .gnd(gnd), .vdd(vdd), .A(_6707_), .B(_6708_), .Y(_208__1_) );
NOR2X1 NOR2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_6702_), .B(_3393__bF_buf8), .Y(_6709_) );
AOI21X1 AOI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(_3313__bF_buf25), .C(data_56__2_), .Y(_6710_) );
AOI21X1 AOI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_6709_), .C(_6710_), .Y(_208__2_) );
INVX1 INVX1_2939 ( .gnd(gnd), .vdd(vdd), .A(data_56__3_), .Y(_6711_) );
OAI21X1 OAI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_6702_), .C(_6711_), .Y(_6712_) );
NAND3X1 NAND3X1_923 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_6704_), .C(_3313__bF_buf24), .Y(_6713_) );
AND2X2 AND2X2_1271 ( .gnd(gnd), .vdd(vdd), .A(_6712_), .B(_6713_), .Y(_208__3_) );
INVX1 INVX1_2940 ( .gnd(gnd), .vdd(vdd), .A(data_56__4_), .Y(_6714_) );
OAI21X1 OAI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_6702_), .C(_6714_), .Y(_6715_) );
NAND3X1 NAND3X1_924 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_6704_), .C(_3313__bF_buf23), .Y(_6716_) );
AND2X2 AND2X2_1272 ( .gnd(gnd), .vdd(vdd), .A(_6715_), .B(_6716_), .Y(_208__4_) );
INVX1 INVX1_2941 ( .gnd(gnd), .vdd(vdd), .A(data_56__5_), .Y(_6717_) );
NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(_3313__bF_buf22), .Y(_6718_) );
MUX2X1 MUX2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_6717_), .B(_14903__bF_buf5), .S(_6718_), .Y(_208__5_) );
AOI21X1 AOI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(_3313__bF_buf21), .C(data_56__6_), .Y(_6719_) );
AOI21X1 AOI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_6709_), .C(_6719_), .Y(_208__6_) );
INVX1 INVX1_2942 ( .gnd(gnd), .vdd(vdd), .A(data_56__7_), .Y(_6720_) );
MUX2X1 MUX2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_6720_), .B(_14908__bF_buf4), .S(_6718_), .Y(_208__7_) );
AOI21X1 AOI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(_3313__bF_buf20), .C(data_56__8_), .Y(_6721_) );
AOI21X1 AOI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_6709_), .C(_6721_), .Y(_208__8_) );
INVX1 INVX1_2943 ( .gnd(gnd), .vdd(vdd), .A(data_56__9_), .Y(_6722_) );
MUX2X1 MUX2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_6722_), .B(_14913__bF_buf12), .S(_6718_), .Y(_208__9_) );
INVX1 INVX1_2944 ( .gnd(gnd), .vdd(vdd), .A(data_56__10_), .Y(_6723_) );
MUX2X1 MUX2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_6723_), .B(_15055__bF_buf4), .S(_6718_), .Y(_208__10_) );
INVX1 INVX1_2945 ( .gnd(gnd), .vdd(vdd), .A(data_56__11_), .Y(_6724_) );
OAI21X1 OAI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_6702_), .C(_6724_), .Y(_6725_) );
NAND3X1 NAND3X1_925 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_6704_), .C(_3313__bF_buf19), .Y(_6726_) );
AND2X2 AND2X2_1273 ( .gnd(gnd), .vdd(vdd), .A(_6725_), .B(_6726_), .Y(_208__11_) );
INVX1 INVX1_2946 ( .gnd(gnd), .vdd(vdd), .A(data_56__12_), .Y(_6727_) );
MUX2X1 MUX2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_6727_), .B(_14920__bF_buf5), .S(_6718_), .Y(_208__12_) );
INVX1 INVX1_2947 ( .gnd(gnd), .vdd(vdd), .A(data_56__13_), .Y(_6728_) );
MUX2X1 MUX2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_6728_), .B(_14924__bF_buf2), .S(_6718_), .Y(_208__13_) );
AOI21X1 AOI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(_3313__bF_buf18), .C(data_56__14_), .Y(_6729_) );
AOI21X1 AOI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf13), .B(_6709_), .C(_6729_), .Y(_208__14_) );
AOI21X1 AOI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_6704_), .B(_3313__bF_buf17), .C(data_56__15_), .Y(_6730_) );
AOI21X1 AOI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_6709_), .C(_6730_), .Y(_208__15_) );
INVX1 INVX1_2948 ( .gnd(gnd), .vdd(vdd), .A(data_55__0_), .Y(_6731_) );
OAI21X1 OAI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_14956_), .B(_3348_), .C(_3342_), .Y(_6732_) );
NOR2X1 NOR2X1_727 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .B(_6732_), .Y(_6733_) );
NAND3X1 NAND3X1_926 ( .gnd(gnd), .vdd(vdd), .A(_4283_), .B(_4284_), .C(_6733_), .Y(_6734_) );
NOR2X1 NOR2X1_728 ( .gnd(gnd), .vdd(vdd), .A(_6734_), .B(_5459__bF_buf2), .Y(_6735_) );
INVX4 INVX4_32 ( .gnd(gnd), .vdd(vdd), .A(_6735_), .Y(_6736_) );
OAI21X1 OAI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_6736_), .C(_6731_), .Y(_6737_) );
NAND3X1 NAND3X1_927 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_6735_), .C(_3313__bF_buf16), .Y(_6738_) );
AND2X2 AND2X2_1274 ( .gnd(gnd), .vdd(vdd), .A(_6737_), .B(_6738_), .Y(_207__0_) );
INVX1 INVX1_2949 ( .gnd(gnd), .vdd(vdd), .A(data_55__1_), .Y(_6739_) );
OAI21X1 OAI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf3), .B(_6736_), .C(_6739_), .Y(_6740_) );
NAND3X1 NAND3X1_928 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_6735_), .C(_3313__bF_buf15), .Y(_6741_) );
AND2X2 AND2X2_1275 ( .gnd(gnd), .vdd(vdd), .A(_6740_), .B(_6741_), .Y(_207__1_) );
INVX1 INVX1_2950 ( .gnd(gnd), .vdd(vdd), .A(data_55__2_), .Y(_6742_) );
NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_6735_), .B(_3313__bF_buf14), .Y(_6743_) );
MUX2X1 MUX2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_6742_), .B(_14897__bF_buf9), .S(_6743_), .Y(_207__2_) );
INVX1 INVX1_2951 ( .gnd(gnd), .vdd(vdd), .A(data_55__3_), .Y(_6744_) );
OAI21X1 OAI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_6736_), .C(_6744_), .Y(_6745_) );
NAND3X1 NAND3X1_929 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_6735_), .C(_3313__bF_buf13), .Y(_6746_) );
AND2X2 AND2X2_1276 ( .gnd(gnd), .vdd(vdd), .A(_6745_), .B(_6746_), .Y(_207__3_) );
INVX1 INVX1_2952 ( .gnd(gnd), .vdd(vdd), .A(data_55__4_), .Y(_6747_) );
OAI21X1 OAI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_6736_), .C(_6747_), .Y(_6748_) );
NAND3X1 NAND3X1_930 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf1), .B(_6735_), .C(_3313__bF_buf12), .Y(_6749_) );
AND2X2 AND2X2_1277 ( .gnd(gnd), .vdd(vdd), .A(_6748_), .B(_6749_), .Y(_207__4_) );
INVX1 INVX1_2953 ( .gnd(gnd), .vdd(vdd), .A(data_55__5_), .Y(_6750_) );
OAI21X1 OAI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_6736_), .C(_6750_), .Y(_6751_) );
NAND3X1 NAND3X1_931 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_6735_), .C(_3313__bF_buf11), .Y(_6752_) );
AND2X2 AND2X2_1278 ( .gnd(gnd), .vdd(vdd), .A(_6751_), .B(_6752_), .Y(_207__5_) );
INVX1 INVX1_2954 ( .gnd(gnd), .vdd(vdd), .A(data_55__6_), .Y(_6753_) );
MUX2X1 MUX2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_6753_), .B(_15049__bF_buf12), .S(_6743_), .Y(_207__6_) );
INVX1 INVX1_2955 ( .gnd(gnd), .vdd(vdd), .A(data_55__7_), .Y(_6754_) );
OAI21X1 OAI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_6736_), .C(_6754_), .Y(_6755_) );
NAND3X1 NAND3X1_932 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_6735_), .C(_3313__bF_buf10), .Y(_6756_) );
AND2X2 AND2X2_1279 ( .gnd(gnd), .vdd(vdd), .A(_6755_), .B(_6756_), .Y(_207__7_) );
INVX1 INVX1_2956 ( .gnd(gnd), .vdd(vdd), .A(data_55__8_), .Y(_6757_) );
MUX2X1 MUX2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_6757_), .B(_15052__bF_buf1), .S(_6743_), .Y(_207__8_) );
INVX1 INVX1_2957 ( .gnd(gnd), .vdd(vdd), .A(data_55__9_), .Y(_6758_) );
MUX2X1 MUX2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_6758_), .B(_14913__bF_buf11), .S(_6743_), .Y(_207__9_) );
INVX1 INVX1_2958 ( .gnd(gnd), .vdd(vdd), .A(data_55__10_), .Y(_6759_) );
MUX2X1 MUX2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_6759_), .B(_15055__bF_buf3), .S(_6743_), .Y(_207__10_) );
INVX1 INVX1_2959 ( .gnd(gnd), .vdd(vdd), .A(data_55__11_), .Y(_6760_) );
OAI21X1 OAI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_6736_), .C(_6760_), .Y(_6761_) );
NAND3X1 NAND3X1_933 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_6735_), .C(_3313__bF_buf9), .Y(_6762_) );
AND2X2 AND2X2_1280 ( .gnd(gnd), .vdd(vdd), .A(_6761_), .B(_6762_), .Y(_207__11_) );
INVX1 INVX1_2960 ( .gnd(gnd), .vdd(vdd), .A(data_55__12_), .Y(_6763_) );
OAI21X1 OAI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_6736_), .C(_6763_), .Y(_6764_) );
NAND3X1 NAND3X1_934 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_6735_), .C(_3313__bF_buf8), .Y(_6765_) );
AND2X2 AND2X2_1281 ( .gnd(gnd), .vdd(vdd), .A(_6764_), .B(_6765_), .Y(_207__12_) );
INVX1 INVX1_2961 ( .gnd(gnd), .vdd(vdd), .A(data_55__13_), .Y(_6766_) );
MUX2X1 MUX2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_6766_), .B(_14924__bF_buf1), .S(_6743_), .Y(_207__13_) );
INVX1 INVX1_2962 ( .gnd(gnd), .vdd(vdd), .A(data_55__14_), .Y(_6767_) );
MUX2X1 MUX2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_6767_), .B(_15060__bF_buf12), .S(_6743_), .Y(_207__14_) );
INVX1 INVX1_2963 ( .gnd(gnd), .vdd(vdd), .A(data_55__15_), .Y(_6768_) );
MUX2X1 MUX2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_6768_), .B(_15062__bF_buf3), .S(_6743_), .Y(_207__15_) );
INVX1 INVX1_2964 ( .gnd(gnd), .vdd(vdd), .A(data_54__0_), .Y(_6769_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(_6732_), .Y(_6770_) );
NAND3X1 NAND3X1_935 ( .gnd(gnd), .vdd(vdd), .A(_4283_), .B(_6770_), .C(_14973_), .Y(_6771_) );
OAI21X1 OAI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_16156_), .B(_3863_), .C(_14998__bF_buf0), .Y(_6772_) );
NAND3X1 NAND3X1_936 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .B(_6484_), .C(_6772_), .Y(_6773_) );
NOR2X1 NOR2X1_729 ( .gnd(gnd), .vdd(vdd), .A(_6773_), .B(_6771_), .Y(_6774_) );
INVX4 INVX4_33 ( .gnd(gnd), .vdd(vdd), .A(_6774_), .Y(_6775_) );
OAI21X1 OAI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_6775_), .C(_6769_), .Y(_6776_) );
NAND3X1 NAND3X1_937 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf12), .B(_6774_), .C(_3313__bF_buf7), .Y(_6777_) );
AND2X2 AND2X2_1282 ( .gnd(gnd), .vdd(vdd), .A(_6776_), .B(_6777_), .Y(_206__0_) );
INVX1 INVX1_2965 ( .gnd(gnd), .vdd(vdd), .A(data_54__1_), .Y(_6778_) );
OAI21X1 OAI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_6775_), .C(_6778_), .Y(_6779_) );
NAND3X1 NAND3X1_938 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_6774_), .C(_3313__bF_buf6), .Y(_6780_) );
AND2X2 AND2X2_1283 ( .gnd(gnd), .vdd(vdd), .A(_6779_), .B(_6780_), .Y(_206__1_) );
INVX1 INVX1_2966 ( .gnd(gnd), .vdd(vdd), .A(data_54__2_), .Y(_6781_) );
NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_6774_), .B(_3313__bF_buf5), .Y(_6782_) );
MUX2X1 MUX2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_6781_), .B(_14897__bF_buf8), .S(_6782_), .Y(_206__2_) );
INVX1 INVX1_2967 ( .gnd(gnd), .vdd(vdd), .A(data_54__3_), .Y(_6783_) );
OAI21X1 OAI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_6775_), .C(_6783_), .Y(_6784_) );
NAND3X1 NAND3X1_939 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_6774_), .C(_3313__bF_buf4), .Y(_6785_) );
AND2X2 AND2X2_1284 ( .gnd(gnd), .vdd(vdd), .A(_6784_), .B(_6785_), .Y(_206__3_) );
INVX1 INVX1_2968 ( .gnd(gnd), .vdd(vdd), .A(data_54__4_), .Y(_6786_) );
OAI21X1 OAI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_6775_), .C(_6786_), .Y(_6787_) );
NAND3X1 NAND3X1_940 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_6774_), .C(_3313__bF_buf3), .Y(_6788_) );
AND2X2 AND2X2_1285 ( .gnd(gnd), .vdd(vdd), .A(_6787_), .B(_6788_), .Y(_206__4_) );
INVX1 INVX1_2969 ( .gnd(gnd), .vdd(vdd), .A(data_54__5_), .Y(_6789_) );
OAI21X1 OAI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_6775_), .C(_6789_), .Y(_6790_) );
NAND3X1 NAND3X1_941 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_6774_), .C(_3313__bF_buf2), .Y(_6791_) );
AND2X2 AND2X2_1286 ( .gnd(gnd), .vdd(vdd), .A(_6790_), .B(_6791_), .Y(_206__5_) );
INVX1 INVX1_2970 ( .gnd(gnd), .vdd(vdd), .A(data_54__6_), .Y(_6792_) );
MUX2X1 MUX2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_6792_), .B(_15049__bF_buf11), .S(_6782_), .Y(_206__6_) );
INVX1 INVX1_2971 ( .gnd(gnd), .vdd(vdd), .A(data_54__7_), .Y(_6793_) );
OAI21X1 OAI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_6775_), .C(_6793_), .Y(_6794_) );
NAND3X1 NAND3X1_942 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_6774_), .C(_3313__bF_buf1), .Y(_6795_) );
AND2X2 AND2X2_1287 ( .gnd(gnd), .vdd(vdd), .A(_6794_), .B(_6795_), .Y(_206__7_) );
INVX1 INVX1_2972 ( .gnd(gnd), .vdd(vdd), .A(data_54__8_), .Y(_6796_) );
MUX2X1 MUX2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_6796_), .B(_15052__bF_buf0), .S(_6782_), .Y(_206__8_) );
INVX1 INVX1_2973 ( .gnd(gnd), .vdd(vdd), .A(data_54__9_), .Y(_6797_) );
MUX2X1 MUX2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_6797_), .B(_14913__bF_buf10), .S(_6782_), .Y(_206__9_) );
INVX1 INVX1_2974 ( .gnd(gnd), .vdd(vdd), .A(data_54__10_), .Y(_6798_) );
MUX2X1 MUX2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_6798_), .B(_15055__bF_buf2), .S(_6782_), .Y(_206__10_) );
INVX1 INVX1_2975 ( .gnd(gnd), .vdd(vdd), .A(data_54__11_), .Y(_6799_) );
OAI21X1 OAI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_6775_), .C(_6799_), .Y(_6800_) );
NAND3X1 NAND3X1_943 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_6774_), .C(_3313__bF_buf0), .Y(_6801_) );
AND2X2 AND2X2_1288 ( .gnd(gnd), .vdd(vdd), .A(_6800_), .B(_6801_), .Y(_206__11_) );
INVX1 INVX1_2976 ( .gnd(gnd), .vdd(vdd), .A(data_54__12_), .Y(_6802_) );
OAI21X1 OAI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_6775_), .C(_6802_), .Y(_6803_) );
NAND3X1 NAND3X1_944 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_6774_), .C(_3313__bF_buf91), .Y(_6804_) );
AND2X2 AND2X2_1289 ( .gnd(gnd), .vdd(vdd), .A(_6803_), .B(_6804_), .Y(_206__12_) );
INVX1 INVX1_2977 ( .gnd(gnd), .vdd(vdd), .A(data_54__13_), .Y(_6805_) );
MUX2X1 MUX2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_6805_), .B(_14924__bF_buf0), .S(_6782_), .Y(_206__13_) );
INVX1 INVX1_2978 ( .gnd(gnd), .vdd(vdd), .A(data_54__14_), .Y(_6806_) );
MUX2X1 MUX2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_6806_), .B(_15060__bF_buf11), .S(_6782_), .Y(_206__14_) );
INVX1 INVX1_2979 ( .gnd(gnd), .vdd(vdd), .A(data_54__15_), .Y(_6807_) );
MUX2X1 MUX2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_6807_), .B(_15062__bF_buf2), .S(_6782_), .Y(_206__15_) );
AOI21X1 AOI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf3), .B(_3983_), .C(_6483_), .Y(_6808_) );
NAND3X1 NAND3X1_945 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .B(_6808_), .C(_4283_), .Y(_6809_) );
NOR2X1 NOR2X1_730 ( .gnd(gnd), .vdd(vdd), .A(_6809_), .B(_5459__bF_buf1), .Y(_6810_) );
AND2X2 AND2X2_1290 ( .gnd(gnd), .vdd(vdd), .A(_6810_), .B(_6770_), .Y(_6811_) );
AND2X2 AND2X2_1291 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf90), .B(_6811_), .Y(_6812_) );
AOI21X1 AOI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf89), .C(data_53__0_), .Y(_6813_) );
AOI21X1 AOI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_6812_), .C(_6813_), .Y(_205__0_) );
AOI21X1 AOI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf88), .C(data_53__1_), .Y(_6814_) );
AOI21X1 AOI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_6812_), .C(_6814_), .Y(_205__1_) );
INVX1 INVX1_2980 ( .gnd(gnd), .vdd(vdd), .A(data_53__2_), .Y(_6815_) );
NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf87), .Y(_6816_) );
NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_6815_), .B(_6816_), .Y(_6817_) );
NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_6812_), .Y(_6818_) );
AND2X2 AND2X2_1292 ( .gnd(gnd), .vdd(vdd), .A(_6818_), .B(_6817_), .Y(_205__2_) );
AOI21X1 AOI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf86), .C(data_53__3_), .Y(_6819_) );
AOI21X1 AOI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_6812_), .C(_6819_), .Y(_205__3_) );
AOI21X1 AOI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf85), .C(data_53__4_), .Y(_6820_) );
AOI21X1 AOI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_6812_), .C(_6820_), .Y(_205__4_) );
INVX1 INVX1_2981 ( .gnd(gnd), .vdd(vdd), .A(data_53__5_), .Y(_6821_) );
MUX2X1 MUX2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_6821_), .B(_14903__bF_buf2), .S(_6816_), .Y(_205__5_) );
INVX1 INVX1_2982 ( .gnd(gnd), .vdd(vdd), .A(data_53__6_), .Y(_6822_) );
NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_6822_), .B(_6816_), .Y(_6823_) );
NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf10), .B(_6812_), .Y(_6824_) );
AND2X2 AND2X2_1293 ( .gnd(gnd), .vdd(vdd), .A(_6824_), .B(_6823_), .Y(_205__6_) );
INVX1 INVX1_2983 ( .gnd(gnd), .vdd(vdd), .A(data_53__7_), .Y(_6825_) );
MUX2X1 MUX2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_6825_), .B(_14908__bF_buf1), .S(_6816_), .Y(_205__7_) );
INVX1 INVX1_2984 ( .gnd(gnd), .vdd(vdd), .A(data_53__8_), .Y(_6826_) );
MUX2X1 MUX2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_6826_), .B(_15052__bF_buf13), .S(_6816_), .Y(_205__8_) );
AOI21X1 AOI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf84), .C(data_53__9_), .Y(_6827_) );
AOI21X1 AOI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_6812_), .C(_6827_), .Y(_205__9_) );
AOI21X1 AOI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf83), .C(data_53__10_), .Y(_6828_) );
AOI21X1 AOI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_6812_), .C(_6828_), .Y(_205__10_) );
AOI21X1 AOI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf82), .C(data_53__11_), .Y(_6829_) );
AOI21X1 AOI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_6812_), .C(_6829_), .Y(_205__11_) );
INVX1 INVX1_2985 ( .gnd(gnd), .vdd(vdd), .A(data_53__12_), .Y(_6830_) );
MUX2X1 MUX2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_6830_), .B(_14920__bF_buf2), .S(_6816_), .Y(_205__12_) );
AOI21X1 AOI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_6811_), .B(_3313__bF_buf81), .C(data_53__13_), .Y(_6831_) );
AOI21X1 AOI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf13), .B(_6812_), .C(_6831_), .Y(_205__13_) );
INVX1 INVX1_2986 ( .gnd(gnd), .vdd(vdd), .A(data_53__14_), .Y(_6832_) );
NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_6832_), .B(_6816_), .Y(_6833_) );
NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_6812_), .Y(_6834_) );
AND2X2 AND2X2_1294 ( .gnd(gnd), .vdd(vdd), .A(_6834_), .B(_6833_), .Y(_205__14_) );
INVX1 INVX1_2987 ( .gnd(gnd), .vdd(vdd), .A(data_53__15_), .Y(_6835_) );
NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_6835_), .B(_6816_), .Y(_6836_) );
NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_6812_), .Y(_6837_) );
AND2X2 AND2X2_1295 ( .gnd(gnd), .vdd(vdd), .A(_6837_), .B(_6836_), .Y(_205__15_) );
AOI21X1 AOI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf2), .B(_4026_), .C(_3347_), .Y(_6838_) );
NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_6808_), .B(_6838_), .Y(_6839_) );
NOR2X1 NOR2X1_731 ( .gnd(gnd), .vdd(vdd), .A(_6839_), .B(_5459__bF_buf0), .Y(_6840_) );
AND2X2 AND2X2_1296 ( .gnd(gnd), .vdd(vdd), .A(_6840_), .B(_6770_), .Y(_6841_) );
AND2X2 AND2X2_1297 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf80), .B(_6841_), .Y(_6842_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_6842__bF_buf3), .B(data_52__0_), .Y(_6843_) );
NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_6842__bF_buf2), .Y(_6844_) );
AND2X2 AND2X2_1298 ( .gnd(gnd), .vdd(vdd), .A(_6843_), .B(_6844_), .Y(_204__0_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_6842__bF_buf1), .B(data_52__1_), .Y(_6845_) );
NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_6842__bF_buf0), .Y(_6846_) );
AND2X2 AND2X2_1299 ( .gnd(gnd), .vdd(vdd), .A(_6845_), .B(_6846_), .Y(_204__1_) );
AOI21X1 AOI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(_3313__bF_buf79), .C(data_52__2_), .Y(_6847_) );
AOI21X1 AOI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_6842__bF_buf3), .C(_6847_), .Y(_204__2_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_6842__bF_buf2), .B(data_52__3_), .Y(_6848_) );
NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_6842__bF_buf1), .Y(_6849_) );
AND2X2 AND2X2_1300 ( .gnd(gnd), .vdd(vdd), .A(_6848_), .B(_6849_), .Y(_204__3_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_6842__bF_buf0), .B(data_52__4_), .Y(_6850_) );
NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_6842__bF_buf3), .Y(_6851_) );
AND2X2 AND2X2_1301 ( .gnd(gnd), .vdd(vdd), .A(_6850_), .B(_6851_), .Y(_204__4_) );
INVX1 INVX1_2988 ( .gnd(gnd), .vdd(vdd), .A(data_52__5_), .Y(_6852_) );
NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(_3313__bF_buf78), .Y(_6853_) );
MUX2X1 MUX2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_6852_), .B(_14903__bF_buf1), .S(_6853_), .Y(_204__5_) );
AOI21X1 AOI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(_3313__bF_buf77), .C(data_52__6_), .Y(_6854_) );
AOI21X1 AOI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_6842__bF_buf2), .C(_6854_), .Y(_204__6_) );
INVX1 INVX1_2989 ( .gnd(gnd), .vdd(vdd), .A(data_52__7_), .Y(_6855_) );
MUX2X1 MUX2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_6855_), .B(_14908__bF_buf0), .S(_6853_), .Y(_204__7_) );
INVX1 INVX1_2990 ( .gnd(gnd), .vdd(vdd), .A(data_52__8_), .Y(_6856_) );
NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_6856_), .B(_6853_), .Y(_6857_) );
NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_6842__bF_buf1), .Y(_6858_) );
AND2X2 AND2X2_1302 ( .gnd(gnd), .vdd(vdd), .A(_6858_), .B(_6857_), .Y(_204__8_) );
INVX1 INVX1_2991 ( .gnd(gnd), .vdd(vdd), .A(data_52__9_), .Y(_6859_) );
NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_6859_), .B(_6853_), .Y(_6860_) );
NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_6842__bF_buf0), .Y(_6861_) );
AND2X2 AND2X2_1303 ( .gnd(gnd), .vdd(vdd), .A(_6861_), .B(_6860_), .Y(_204__9_) );
INVX1 INVX1_2992 ( .gnd(gnd), .vdd(vdd), .A(data_52__10_), .Y(_6862_) );
NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_6862_), .B(_6853_), .Y(_6863_) );
NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_6842__bF_buf3), .Y(_6864_) );
AND2X2 AND2X2_1304 ( .gnd(gnd), .vdd(vdd), .A(_6864_), .B(_6863_), .Y(_204__10_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_6842__bF_buf2), .B(data_52__11_), .Y(_6865_) );
NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_6842__bF_buf1), .Y(_6866_) );
AND2X2 AND2X2_1305 ( .gnd(gnd), .vdd(vdd), .A(_6865_), .B(_6866_), .Y(_204__11_) );
INVX1 INVX1_2993 ( .gnd(gnd), .vdd(vdd), .A(data_52__12_), .Y(_6867_) );
MUX2X1 MUX2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_6867_), .B(_14920__bF_buf1), .S(_6853_), .Y(_204__12_) );
INVX1 INVX1_2994 ( .gnd(gnd), .vdd(vdd), .A(data_52__13_), .Y(_6868_) );
NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_6868_), .B(_6853_), .Y(_6869_) );
NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_6842__bF_buf0), .Y(_6870_) );
AND2X2 AND2X2_1306 ( .gnd(gnd), .vdd(vdd), .A(_6870_), .B(_6869_), .Y(_204__13_) );
AOI21X1 AOI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(_3313__bF_buf76), .C(data_52__14_), .Y(_6871_) );
AOI21X1 AOI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf9), .B(_6842__bF_buf3), .C(_6871_), .Y(_204__14_) );
AOI21X1 AOI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_6841_), .B(_3313__bF_buf75), .C(data_52__15_), .Y(_6872_) );
AOI21X1 AOI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_6842__bF_buf2), .C(_6872_), .Y(_204__15_) );
INVX1 INVX1_2995 ( .gnd(gnd), .vdd(vdd), .A(data_51__0_), .Y(_6873_) );
AOI21X1 AOI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_14952__bF_buf4), .B(_14998__bF_buf1), .C(_3347_), .Y(_6874_) );
NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_6874_), .B(_6733_), .Y(_6875_) );
NOR2X1 NOR2X1_732 ( .gnd(gnd), .vdd(vdd), .A(_6875_), .B(_5459__bF_buf3), .Y(_6876_) );
INVX4 INVX4_34 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .Y(_6877_) );
OAI21X1 OAI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_6877_), .C(_6873_), .Y(_6878_) );
NAND3X1 NAND3X1_946 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_6876_), .C(_3313__bF_buf74), .Y(_6879_) );
AND2X2 AND2X2_1307 ( .gnd(gnd), .vdd(vdd), .A(_6878_), .B(_6879_), .Y(_203__0_) );
INVX1 INVX1_2996 ( .gnd(gnd), .vdd(vdd), .A(data_51__1_), .Y(_6880_) );
OAI21X1 OAI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_6877_), .C(_6880_), .Y(_6881_) );
NAND3X1 NAND3X1_947 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf10), .B(_6876_), .C(_3313__bF_buf73), .Y(_6882_) );
AND2X2 AND2X2_1308 ( .gnd(gnd), .vdd(vdd), .A(_6881_), .B(_6882_), .Y(_203__1_) );
NOR2X1 NOR2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_6877_), .B(_3393__bF_buf56), .Y(_6883_) );
AOI21X1 AOI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_3313__bF_buf72), .C(data_51__2_), .Y(_6884_) );
AOI21X1 AOI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_6883_), .C(_6884_), .Y(_203__2_) );
INVX1 INVX1_2997 ( .gnd(gnd), .vdd(vdd), .A(data_51__3_), .Y(_6885_) );
OAI21X1 OAI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_6877_), .C(_6885_), .Y(_6886_) );
NAND3X1 NAND3X1_948 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_6876_), .C(_3313__bF_buf71), .Y(_6887_) );
AND2X2 AND2X2_1309 ( .gnd(gnd), .vdd(vdd), .A(_6886_), .B(_6887_), .Y(_203__3_) );
INVX1 INVX1_2998 ( .gnd(gnd), .vdd(vdd), .A(data_51__4_), .Y(_6888_) );
OAI21X1 OAI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_6877_), .C(_6888_), .Y(_6889_) );
NAND3X1 NAND3X1_949 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_6876_), .C(_3313__bF_buf70), .Y(_6890_) );
AND2X2 AND2X2_1310 ( .gnd(gnd), .vdd(vdd), .A(_6889_), .B(_6890_), .Y(_203__4_) );
INVX1 INVX1_2999 ( .gnd(gnd), .vdd(vdd), .A(data_51__5_), .Y(_6891_) );
NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_3313__bF_buf69), .Y(_6892_) );
MUX2X1 MUX2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_6891_), .B(_14903__bF_buf0), .S(_6892_), .Y(_203__5_) );
AOI21X1 AOI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_3313__bF_buf68), .C(data_51__6_), .Y(_6893_) );
AOI21X1 AOI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_6883_), .C(_6893_), .Y(_203__6_) );
INVX1 INVX1_3000 ( .gnd(gnd), .vdd(vdd), .A(data_51__7_), .Y(_6894_) );
MUX2X1 MUX2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_6894_), .B(_14908__bF_buf13), .S(_6892_), .Y(_203__7_) );
INVX1 INVX1_3001 ( .gnd(gnd), .vdd(vdd), .A(data_51__8_), .Y(_6895_) );
MUX2X1 MUX2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_6895_), .B(_15052__bF_buf11), .S(_6892_), .Y(_203__8_) );
INVX1 INVX1_3002 ( .gnd(gnd), .vdd(vdd), .A(data_51__9_), .Y(_6896_) );
MUX2X1 MUX2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_6896_), .B(_14913__bF_buf7), .S(_6892_), .Y(_203__9_) );
INVX1 INVX1_3003 ( .gnd(gnd), .vdd(vdd), .A(data_51__10_), .Y(_6897_) );
MUX2X1 MUX2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_6897_), .B(_15055__bF_buf13), .S(_6892_), .Y(_203__10_) );
INVX1 INVX1_3004 ( .gnd(gnd), .vdd(vdd), .A(data_51__11_), .Y(_6898_) );
OAI21X1 OAI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_6877_), .C(_6898_), .Y(_6899_) );
NAND3X1 NAND3X1_950 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_6876_), .C(_3313__bF_buf67), .Y(_6900_) );
AND2X2 AND2X2_1311 ( .gnd(gnd), .vdd(vdd), .A(_6899_), .B(_6900_), .Y(_203__11_) );
INVX1 INVX1_3005 ( .gnd(gnd), .vdd(vdd), .A(data_51__12_), .Y(_6901_) );
MUX2X1 MUX2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_6901_), .B(_14920__bF_buf0), .S(_6892_), .Y(_203__12_) );
INVX1 INVX1_3006 ( .gnd(gnd), .vdd(vdd), .A(data_51__13_), .Y(_6902_) );
MUX2X1 MUX2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_6902_), .B(_14924__bF_buf11), .S(_6892_), .Y(_203__13_) );
AOI21X1 AOI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_3313__bF_buf66), .C(data_51__14_), .Y(_6903_) );
AOI21X1 AOI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_6883_), .C(_6903_), .Y(_203__14_) );
AOI21X1 AOI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_6876_), .B(_3313__bF_buf65), .C(data_51__15_), .Y(_6904_) );
AOI21X1 AOI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf13), .B(_6883_), .C(_6904_), .Y(_203__15_) );
INVX1 INVX1_3007 ( .gnd(gnd), .vdd(vdd), .A(data_50__0_), .Y(_6905_) );
NOR2X1 NOR2X1_734 ( .gnd(gnd), .vdd(vdd), .A(_6483_), .B(_4282_), .Y(_6906_) );
OAI21X1 OAI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_4683_), .C(_6906_), .Y(_6907_) );
NOR2X1 NOR2X1_735 ( .gnd(gnd), .vdd(vdd), .A(_6907_), .B(_5459__bF_buf2), .Y(_6908_) );
AND2X2 AND2X2_1312 ( .gnd(gnd), .vdd(vdd), .A(_6908_), .B(_6770_), .Y(_6909_) );
NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_6909_), .B(_3313__bF_buf64), .Y(_6910_) );
NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_6905_), .B(_6910_), .Y(_6911_) );
AND2X2 AND2X2_1313 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf63), .B(_6909_), .Y(_6912_) );
NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_6912__bF_buf3), .Y(_6913_) );
AND2X2 AND2X2_1314 ( .gnd(gnd), .vdd(vdd), .A(_6913_), .B(_6911_), .Y(_202__0_) );
INVX1 INVX1_3008 ( .gnd(gnd), .vdd(vdd), .A(data_50__1_), .Y(_6914_) );
NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_6914_), .B(_6910_), .Y(_6915_) );
NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_6912__bF_buf2), .Y(_6916_) );
AND2X2 AND2X2_1315 ( .gnd(gnd), .vdd(vdd), .A(_6916_), .B(_6915_), .Y(_202__1_) );
INVX1 INVX1_3009 ( .gnd(gnd), .vdd(vdd), .A(data_50__2_), .Y(_6917_) );
NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_6917_), .B(_6910_), .Y(_6918_) );
NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_6912__bF_buf1), .Y(_6919_) );
AND2X2 AND2X2_1316 ( .gnd(gnd), .vdd(vdd), .A(_6919_), .B(_6918_), .Y(_202__2_) );
INVX1 INVX1_3010 ( .gnd(gnd), .vdd(vdd), .A(data_50__3_), .Y(_6920_) );
NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_6920_), .B(_6910_), .Y(_6921_) );
NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_6912__bF_buf0), .Y(_6922_) );
AND2X2 AND2X2_1317 ( .gnd(gnd), .vdd(vdd), .A(_6922_), .B(_6921_), .Y(_202__3_) );
INVX1 INVX1_3011 ( .gnd(gnd), .vdd(vdd), .A(data_50__4_), .Y(_6923_) );
NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_6923_), .B(_6910_), .Y(_6924_) );
NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_6912__bF_buf3), .Y(_6925_) );
AND2X2 AND2X2_1318 ( .gnd(gnd), .vdd(vdd), .A(_6925_), .B(_6924_), .Y(_202__4_) );
OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_6912__bF_buf2), .B(data_50__5_), .Y(_6926_) );
NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_6912__bF_buf1), .Y(_6927_) );
AND2X2 AND2X2_1319 ( .gnd(gnd), .vdd(vdd), .A(_6926_), .B(_6927_), .Y(_202__5_) );
INVX1 INVX1_3012 ( .gnd(gnd), .vdd(vdd), .A(data_50__6_), .Y(_6928_) );
NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_6928_), .B(_6910_), .Y(_6929_) );
NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf7), .B(_6912__bF_buf0), .Y(_6930_) );
AND2X2 AND2X2_1320 ( .gnd(gnd), .vdd(vdd), .A(_6930_), .B(_6929_), .Y(_202__6_) );
OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_6912__bF_buf3), .B(data_50__7_), .Y(_6931_) );
NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_6912__bF_buf2), .Y(_6932_) );
AND2X2 AND2X2_1321 ( .gnd(gnd), .vdd(vdd), .A(_6931_), .B(_6932_), .Y(_202__7_) );
INVX1 INVX1_3013 ( .gnd(gnd), .vdd(vdd), .A(data_50__8_), .Y(_6933_) );
NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_6933_), .B(_6910_), .Y(_6934_) );
NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_6912__bF_buf1), .Y(_6935_) );
AND2X2 AND2X2_1322 ( .gnd(gnd), .vdd(vdd), .A(_6935_), .B(_6934_), .Y(_202__8_) );
INVX1 INVX1_3014 ( .gnd(gnd), .vdd(vdd), .A(data_50__9_), .Y(_6936_) );
NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_6936_), .B(_6910_), .Y(_6937_) );
NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_6912__bF_buf0), .Y(_6938_) );
AND2X2 AND2X2_1323 ( .gnd(gnd), .vdd(vdd), .A(_6938_), .B(_6937_), .Y(_202__9_) );
INVX1 INVX1_3015 ( .gnd(gnd), .vdd(vdd), .A(data_50__10_), .Y(_6939_) );
NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_6939_), .B(_6910_), .Y(_6940_) );
NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_6912__bF_buf3), .Y(_6941_) );
AND2X2 AND2X2_1324 ( .gnd(gnd), .vdd(vdd), .A(_6941_), .B(_6940_), .Y(_202__10_) );
INVX1 INVX1_3016 ( .gnd(gnd), .vdd(vdd), .A(data_50__11_), .Y(_6942_) );
NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_6942_), .B(_6910_), .Y(_6943_) );
NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_6912__bF_buf2), .Y(_6944_) );
AND2X2 AND2X2_1325 ( .gnd(gnd), .vdd(vdd), .A(_6944_), .B(_6943_), .Y(_202__11_) );
OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_6912__bF_buf1), .B(data_50__12_), .Y(_6945_) );
NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_6912__bF_buf0), .Y(_6946_) );
AND2X2 AND2X2_1326 ( .gnd(gnd), .vdd(vdd), .A(_6945_), .B(_6946_), .Y(_202__12_) );
INVX1 INVX1_3017 ( .gnd(gnd), .vdd(vdd), .A(data_50__13_), .Y(_6947_) );
NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_6947_), .B(_6910_), .Y(_6948_) );
NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf10), .B(_6912__bF_buf3), .Y(_6949_) );
AND2X2 AND2X2_1327 ( .gnd(gnd), .vdd(vdd), .A(_6949_), .B(_6948_), .Y(_202__13_) );
INVX1 INVX1_3018 ( .gnd(gnd), .vdd(vdd), .A(data_50__14_), .Y(_6950_) );
NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_6950_), .B(_6910_), .Y(_6951_) );
NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_6912__bF_buf2), .Y(_6952_) );
AND2X2 AND2X2_1328 ( .gnd(gnd), .vdd(vdd), .A(_6952_), .B(_6951_), .Y(_202__14_) );
INVX1 INVX1_3019 ( .gnd(gnd), .vdd(vdd), .A(data_50__15_), .Y(_6953_) );
NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_6953_), .B(_6910_), .Y(_6954_) );
NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_6912__bF_buf1), .Y(_6955_) );
AND2X2 AND2X2_1329 ( .gnd(gnd), .vdd(vdd), .A(_6955_), .B(_6954_), .Y(_202__15_) );
INVX1 INVX1_3020 ( .gnd(gnd), .vdd(vdd), .A(data_49__0_), .Y(_6956_) );
OAI21X1 OAI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_4722_), .C(_6906_), .Y(_6957_) );
NOR2X1 NOR2X1_736 ( .gnd(gnd), .vdd(vdd), .A(_6957_), .B(_5459__bF_buf1), .Y(_6958_) );
AND2X2 AND2X2_1330 ( .gnd(gnd), .vdd(vdd), .A(_6958_), .B(_6770_), .Y(_6959_) );
NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_6959_), .B(_3313__bF_buf62), .Y(_6960_) );
MUX2X1 MUX2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_6956_), .B(_14932__bF_buf7), .S(_6960_), .Y(_200__0_) );
INVX1 INVX1_3021 ( .gnd(gnd), .vdd(vdd), .A(data_49__1_), .Y(_6961_) );
MUX2X1 MUX2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_6961_), .B(_14894__bF_buf8), .S(_6960_), .Y(_200__1_) );
INVX1 INVX1_3022 ( .gnd(gnd), .vdd(vdd), .A(data_49__2_), .Y(_6962_) );
NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_6962_), .B(_6960_), .Y(_6963_) );
AND2X2 AND2X2_1331 ( .gnd(gnd), .vdd(vdd), .A(_3313__bF_buf61), .B(_6959_), .Y(_6964_) );
NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_6964_), .Y(_6965_) );
AND2X2 AND2X2_1332 ( .gnd(gnd), .vdd(vdd), .A(_6965_), .B(_6963_), .Y(_200__2_) );
INVX1 INVX1_3023 ( .gnd(gnd), .vdd(vdd), .A(data_49__3_), .Y(_6966_) );
MUX2X1 MUX2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_6966_), .B(_14899__bF_buf7), .S(_6960_), .Y(_200__3_) );
INVX1 INVX1_3024 ( .gnd(gnd), .vdd(vdd), .A(data_49__4_), .Y(_6967_) );
MUX2X1 MUX2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_6967_), .B(_14902__bF_buf9), .S(_6960_), .Y(_200__4_) );
OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_6964_), .B(data_49__5_), .Y(_6968_) );
NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_6964_), .Y(_6969_) );
AND2X2 AND2X2_1333 ( .gnd(gnd), .vdd(vdd), .A(_6968_), .B(_6969_), .Y(_200__5_) );
INVX1 INVX1_3025 ( .gnd(gnd), .vdd(vdd), .A(data_49__6_), .Y(_6970_) );
NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_6970_), .B(_6960_), .Y(_6971_) );
NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_6964_), .Y(_6972_) );
AND2X2 AND2X2_1334 ( .gnd(gnd), .vdd(vdd), .A(_6972_), .B(_6971_), .Y(_200__6_) );
OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_6964_), .B(data_49__7_), .Y(_6973_) );
NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_6964_), .Y(_6974_) );
AND2X2 AND2X2_1335 ( .gnd(gnd), .vdd(vdd), .A(_6973_), .B(_6974_), .Y(_200__7_) );
INVX1 INVX1_3026 ( .gnd(gnd), .vdd(vdd), .A(data_49__8_), .Y(_6975_) );
NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_6975_), .B(_6960_), .Y(_6976_) );
NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf9), .B(_6964_), .Y(_6977_) );
AND2X2 AND2X2_1336 ( .gnd(gnd), .vdd(vdd), .A(_6977_), .B(_6976_), .Y(_200__8_) );
AOI21X1 AOI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_6959_), .B(_3313__bF_buf60), .C(data_49__9_), .Y(_6978_) );
AOI21X1 AOI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_6964_), .C(_6978_), .Y(_200__9_) );
AOI21X1 AOI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_6959_), .B(_3313__bF_buf59), .C(data_49__10_), .Y(_6979_) );
AOI21X1 AOI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_6964_), .C(_6979_), .Y(_200__10_) );
INVX1 INVX1_3027 ( .gnd(gnd), .vdd(vdd), .A(data_49__11_), .Y(_6980_) );
MUX2X1 MUX2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_6980_), .B(_14918__bF_buf11), .S(_6960_), .Y(_200__11_) );
OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_6964_), .B(data_49__12_), .Y(_6981_) );
NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_6964_), .Y(_6982_) );
AND2X2 AND2X2_1337 ( .gnd(gnd), .vdd(vdd), .A(_6981_), .B(_6982_), .Y(_200__12_) );
AOI21X1 AOI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_6959_), .B(_3313__bF_buf58), .C(data_49__13_), .Y(_6983_) );
AOI21X1 AOI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_6964_), .C(_6983_), .Y(_200__13_) );
INVX1 INVX1_3028 ( .gnd(gnd), .vdd(vdd), .A(data_49__14_), .Y(_6984_) );
NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_6984_), .B(_6960_), .Y(_6985_) );
NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf6), .B(_6964_), .Y(_6986_) );
AND2X2 AND2X2_1338 ( .gnd(gnd), .vdd(vdd), .A(_6986_), .B(_6985_), .Y(_200__14_) );
INVX1 INVX1_3029 ( .gnd(gnd), .vdd(vdd), .A(data_49__15_), .Y(_6987_) );
NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_6987_), .B(_6960_), .Y(_6988_) );
NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_6964_), .Y(_6989_) );
AND2X2 AND2X2_1339 ( .gnd(gnd), .vdd(vdd), .A(_6989_), .B(_6988_), .Y(_200__15_) );
INVX1 INVX1_3030 ( .gnd(gnd), .vdd(vdd), .A(data_48__0_), .Y(_6990_) );
NAND3X1 NAND3X1_951 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .B(_14998__bF_buf0), .C(_14986_), .Y(_6991_) );
MUX2X1 MUX2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_6990_), .B(_14932__bF_buf6), .S(_6991_), .Y(_199__0_) );
INVX1 INVX1_3031 ( .gnd(gnd), .vdd(vdd), .A(data_48__1_), .Y(_6992_) );
MUX2X1 MUX2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_6992_), .B(_14894__bF_buf7), .S(_6991_), .Y(_199__1_) );
INVX1 INVX1_3032 ( .gnd(gnd), .vdd(vdd), .A(data_48__2_), .Y(_6993_) );
OAI21X1 OAI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf1), .C(_6993_), .Y(_6994_) );
OAI21X1 OAI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_2_bF_buf3), .B(_6991_), .C(_6994_), .Y(_6995_) );
INVX1 INVX1_3033 ( .gnd(gnd), .vdd(vdd), .A(_6995_), .Y(_199__2_) );
INVX1 INVX1_3034 ( .gnd(gnd), .vdd(vdd), .A(data_48__3_), .Y(_6996_) );
MUX2X1 MUX2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_6996_), .B(_14899__bF_buf6), .S(_6991_), .Y(_199__3_) );
INVX1 INVX1_3035 ( .gnd(gnd), .vdd(vdd), .A(data_48__4_), .Y(_6997_) );
OAI21X1 OAI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf0), .C(_6997_), .Y(_6998_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_6991_), .Y(_6999_) );
NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf8), .B(_6999_), .Y(_7000_) );
AND2X2 AND2X2_1340 ( .gnd(gnd), .vdd(vdd), .A(_7000_), .B(_6998_), .Y(_199__4_) );
INVX1 INVX1_3036 ( .gnd(gnd), .vdd(vdd), .A(data_48__5_), .Y(_7001_) );
OAI21X1 OAI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf15_bF_buf3), .C(_7001_), .Y(_7002_) );
OAI21X1 OAI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf0), .B(_6991_), .C(_7002_), .Y(_7003_) );
INVX1 INVX1_3037 ( .gnd(gnd), .vdd(vdd), .A(_7003_), .Y(_199__5_) );
INVX1 INVX1_3038 ( .gnd(gnd), .vdd(vdd), .A(data_48__6_), .Y(_7004_) );
MUX2X1 MUX2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_7004_), .B(_15049__bF_buf5), .S(_6991_), .Y(_199__6_) );
INVX1 INVX1_3039 ( .gnd(gnd), .vdd(vdd), .A(data_48__7_), .Y(_7005_) );
OAI21X1 OAI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf14_bF_buf3), .C(_7005_), .Y(_7006_) );
OAI21X1 OAI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf0), .B(_6991_), .C(_7006_), .Y(_7007_) );
INVX1 INVX1_3040 ( .gnd(gnd), .vdd(vdd), .A(_7007_), .Y(_199__7_) );
INVX1 INVX1_3041 ( .gnd(gnd), .vdd(vdd), .A(data_48__8_), .Y(_7008_) );
OAI21X1 OAI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf13_bF_buf3), .C(_7008_), .Y(_7009_) );
NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_6999_), .Y(_7010_) );
AND2X2 AND2X2_1341 ( .gnd(gnd), .vdd(vdd), .A(_7010_), .B(_7009_), .Y(_199__8_) );
NOR2X1 NOR2X1_737 ( .gnd(gnd), .vdd(vdd), .A(data_48__9_), .B(_6999_), .Y(_7011_) );
AOI21X1 AOI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf4), .B(_6999_), .C(_7011_), .Y(_199__9_) );
INVX1 INVX1_3042 ( .gnd(gnd), .vdd(vdd), .A(data_48__10_), .Y(_7012_) );
MUX2X1 MUX2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_7012_), .B(_15055__bF_buf10), .S(_6991_), .Y(_199__10_) );
INVX1 INVX1_3043 ( .gnd(gnd), .vdd(vdd), .A(data_48__11_), .Y(_7013_) );
OAI21X1 OAI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf12), .C(_7013_), .Y(_7014_) );
OAI21X1 OAI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf1), .B(_6991_), .C(_7014_), .Y(_7015_) );
INVX1 INVX1_3044 ( .gnd(gnd), .vdd(vdd), .A(_7015_), .Y(_199__11_) );
INVX1 INVX1_3045 ( .gnd(gnd), .vdd(vdd), .A(data_48__12_), .Y(_7016_) );
MUX2X1 MUX2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_7016_), .B(_14920__bF_buf11), .S(_6991_), .Y(_199__12_) );
INVX1 INVX1_3046 ( .gnd(gnd), .vdd(vdd), .A(data_48__13_), .Y(_7017_) );
MUX2X1 MUX2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_7017_), .B(_14924__bF_buf8), .S(_6991_), .Y(_199__13_) );
INVX1 INVX1_3047 ( .gnd(gnd), .vdd(vdd), .A(data_48__14_), .Y(_7018_) );
MUX2X1 MUX2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_7018_), .B(_15060__bF_buf5), .S(_6991_), .Y(_199__14_) );
INVX1 INVX1_3048 ( .gnd(gnd), .vdd(vdd), .A(data_48__15_), .Y(_7019_) );
OAI21X1 OAI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_14882__bF_buf11), .C(_7019_), .Y(_7020_) );
OAI21X1 OAI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf0), .B(_6991_), .C(_7020_), .Y(_7021_) );
INVX1 INVX1_3049 ( .gnd(gnd), .vdd(vdd), .A(_7021_), .Y(_199__15_) );
NOR2X1 NOR2X1_738 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_15170__bF_buf2), .Y(_7022_) );
NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_7022_), .Y(_7023_) );
INVX1 INVX1_3050 ( .gnd(gnd), .vdd(vdd), .A(data_47__0_), .Y(_7024_) );
NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf1), .B(_14946__bF_buf4), .Y(_7025_) );
OAI21X1 OAI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf10), .C(_7024_), .Y(_7026_) );
OAI21X1 OAI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf4), .B(_7023_), .C(_7026_), .Y(_7027_) );
INVX1 INVX1_3051 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .Y(_198__0_) );
INVX1 INVX1_3052 ( .gnd(gnd), .vdd(vdd), .A(data_47__1_), .Y(_7028_) );
OAI21X1 OAI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf9), .C(_7028_), .Y(_7029_) );
NOR2X1 NOR2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf8), .B(_7025_), .Y(_7030_) );
NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_7030_), .Y(_7031_) );
AND2X2 AND2X2_1342 ( .gnd(gnd), .vdd(vdd), .A(_7031_), .B(_7029_), .Y(_198__1_) );
NOR2X1 NOR2X1_740 ( .gnd(gnd), .vdd(vdd), .A(data_47__2_), .B(_7030_), .Y(_7032_) );
AOI21X1 AOI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf2), .B(_7030_), .C(_7032_), .Y(_198__2_) );
INVX1 INVX1_3053 ( .gnd(gnd), .vdd(vdd), .A(data_47__3_), .Y(_7033_) );
OAI21X1 OAI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf7), .C(_7033_), .Y(_7034_) );
NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_7030_), .Y(_7035_) );
AND2X2 AND2X2_1343 ( .gnd(gnd), .vdd(vdd), .A(_7035_), .B(_7034_), .Y(_198__3_) );
INVX1 INVX1_3054 ( .gnd(gnd), .vdd(vdd), .A(data_47__4_), .Y(_7036_) );
OAI21X1 OAI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf6), .C(_7036_), .Y(_7037_) );
OAI21X1 OAI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf3), .B(_7023_), .C(_7037_), .Y(_7038_) );
INVX1 INVX1_3055 ( .gnd(gnd), .vdd(vdd), .A(_7038_), .Y(_198__4_) );
INVX1 INVX1_3056 ( .gnd(gnd), .vdd(vdd), .A(data_47__5_), .Y(_7039_) );
OAI21X1 OAI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf5), .C(_7039_), .Y(_7040_) );
NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_7030_), .Y(_7041_) );
AND2X2 AND2X2_1344 ( .gnd(gnd), .vdd(vdd), .A(_7041_), .B(_7040_), .Y(_198__5_) );
INVX1 INVX1_3057 ( .gnd(gnd), .vdd(vdd), .A(data_47__6_), .Y(_7042_) );
OAI21X1 OAI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf4), .C(_7042_), .Y(_7043_) );
OAI21X1 OAI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf0), .B(_7023_), .C(_7043_), .Y(_7044_) );
INVX1 INVX1_3058 ( .gnd(gnd), .vdd(vdd), .A(_7044_), .Y(_198__6_) );
INVX1 INVX1_3059 ( .gnd(gnd), .vdd(vdd), .A(data_47__7_), .Y(_7045_) );
OAI21X1 OAI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf3), .C(_7045_), .Y(_7046_) );
OAI21X1 OAI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf5), .B(_7023_), .C(_7046_), .Y(_7047_) );
INVX1 INVX1_3060 ( .gnd(gnd), .vdd(vdd), .A(_7047_), .Y(_198__7_) );
INVX1 INVX1_3061 ( .gnd(gnd), .vdd(vdd), .A(data_47__8_), .Y(_7048_) );
OAI21X1 OAI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf2), .C(_7048_), .Y(_7049_) );
OAI21X1 OAI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf3), .B(_7023_), .C(_7049_), .Y(_7050_) );
INVX1 INVX1_3062 ( .gnd(gnd), .vdd(vdd), .A(_7050_), .Y(_198__8_) );
NOR2X1 NOR2X1_741 ( .gnd(gnd), .vdd(vdd), .A(data_47__9_), .B(_7030_), .Y(_7051_) );
AOI21X1 AOI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_7030_), .C(_7051_), .Y(_198__9_) );
INVX1 INVX1_3063 ( .gnd(gnd), .vdd(vdd), .A(data_47__10_), .Y(_7052_) );
OAI21X1 OAI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf1), .C(_7052_), .Y(_7053_) );
NAND3X1 NAND3X1_952 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_15055__bF_buf9), .C(_7022_), .Y(_7054_) );
AND2X2 AND2X2_1345 ( .gnd(gnd), .vdd(vdd), .A(_7053_), .B(_7054_), .Y(_198__10_) );
INVX1 INVX1_3064 ( .gnd(gnd), .vdd(vdd), .A(data_47__11_), .Y(_7055_) );
OAI21X1 OAI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf0), .C(_7055_), .Y(_7056_) );
OAI21X1 OAI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf0), .B(_7023_), .C(_7056_), .Y(_7057_) );
INVX1 INVX1_3065 ( .gnd(gnd), .vdd(vdd), .A(_7057_), .Y(_198__11_) );
INVX1 INVX1_3066 ( .gnd(gnd), .vdd(vdd), .A(data_47__12_), .Y(_7058_) );
OAI21X1 OAI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf15_bF_buf2), .C(_7058_), .Y(_7059_) );
OAI21X1 OAI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf0), .B(_7023_), .C(_7059_), .Y(_7060_) );
INVX1 INVX1_3067 ( .gnd(gnd), .vdd(vdd), .A(_7060_), .Y(_198__12_) );
INVX1 INVX1_3068 ( .gnd(gnd), .vdd(vdd), .A(data_47__13_), .Y(_7061_) );
OAI21X1 OAI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf14_bF_buf2), .C(_7061_), .Y(_7062_) );
NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf7), .B(_7030_), .Y(_7063_) );
AND2X2 AND2X2_1346 ( .gnd(gnd), .vdd(vdd), .A(_7063_), .B(_7062_), .Y(_198__13_) );
INVX1 INVX1_3069 ( .gnd(gnd), .vdd(vdd), .A(data_47__14_), .Y(_7064_) );
OAI21X1 OAI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf13_bF_buf2), .C(_7064_), .Y(_7065_) );
NAND3X1 NAND3X1_953 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf5), .B(_15060__bF_buf4), .C(_7022_), .Y(_7066_) );
AND2X2 AND2X2_1347 ( .gnd(gnd), .vdd(vdd), .A(_7065_), .B(_7066_), .Y(_198__14_) );
INVX1 INVX1_3070 ( .gnd(gnd), .vdd(vdd), .A(data_47__15_), .Y(_7067_) );
OAI21X1 OAI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_7025_), .B(_14882__bF_buf12), .C(_7067_), .Y(_7068_) );
NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf10), .B(_7030_), .Y(_7069_) );
AND2X2 AND2X2_1348 ( .gnd(gnd), .vdd(vdd), .A(_7069_), .B(_7068_), .Y(_198__15_) );
NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf3), .B(_15793__bF_buf0), .Y(_7070_) );
INVX1 INVX1_3071 ( .gnd(gnd), .vdd(vdd), .A(data_46__0_), .Y(_7071_) );
OAI21X1 OAI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15170__bF_buf1), .C(_7071_), .Y(_7072_) );
OAI21X1 OAI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf3), .B(_7070_), .C(_7072_), .Y(_7073_) );
INVX1 INVX1_3072 ( .gnd(gnd), .vdd(vdd), .A(_7073_), .Y(_197__0_) );
INVX1 INVX1_3073 ( .gnd(gnd), .vdd(vdd), .A(data_46__1_), .Y(_7074_) );
OAI21X1 OAI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15170__bF_buf0), .C(_7074_), .Y(_7075_) );
NOR2X1 NOR2X1_742 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf3), .B(_15788__bF_buf8), .Y(_7076_) );
NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_7076_), .Y(_7077_) );
AND2X2 AND2X2_1349 ( .gnd(gnd), .vdd(vdd), .A(_7077_), .B(_7075_), .Y(_197__1_) );
NOR2X1 NOR2X1_743 ( .gnd(gnd), .vdd(vdd), .A(data_46__2_), .B(_7076_), .Y(_7078_) );
AOI21X1 AOI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_7076_), .C(_7078_), .Y(_197__2_) );
NOR2X1 NOR2X1_744 ( .gnd(gnd), .vdd(vdd), .A(data_46__3_), .B(_7076_), .Y(_7079_) );
NOR2X1 NOR2X1_745 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf4), .B(_7070_), .Y(_7080_) );
NOR2X1 NOR2X1_746 ( .gnd(gnd), .vdd(vdd), .A(_7080_), .B(_7079_), .Y(_197__3_) );
INVX1 INVX1_3074 ( .gnd(gnd), .vdd(vdd), .A(data_46__4_), .Y(_7081_) );
OAI21X1 OAI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15170__bF_buf2), .C(_7081_), .Y(_7082_) );
OAI21X1 OAI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf2), .B(_7070_), .C(_7082_), .Y(_7083_) );
INVX1 INVX1_3075 ( .gnd(gnd), .vdd(vdd), .A(_7083_), .Y(_197__4_) );
INVX1 INVX1_3076 ( .gnd(gnd), .vdd(vdd), .A(data_46__5_), .Y(_7084_) );
OAI21X1 OAI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15170__bF_buf1), .C(_7084_), .Y(_7085_) );
NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_7076_), .Y(_7086_) );
AND2X2 AND2X2_1350 ( .gnd(gnd), .vdd(vdd), .A(_7086_), .B(_7085_), .Y(_197__5_) );
INVX1 INVX1_3077 ( .gnd(gnd), .vdd(vdd), .A(data_46__6_), .Y(_7087_) );
OAI21X1 OAI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15170__bF_buf0), .C(_7087_), .Y(_7088_) );
NAND3X1 NAND3X1_954 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf4), .B(_14946__bF_buf2), .C(_15793__bF_buf5), .Y(_7089_) );
AND2X2 AND2X2_1351 ( .gnd(gnd), .vdd(vdd), .A(_7088_), .B(_7089_), .Y(_197__6_) );
INVX1 INVX1_3078 ( .gnd(gnd), .vdd(vdd), .A(data_46__7_), .Y(_7090_) );
OAI21X1 OAI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15170__bF_buf3), .C(_7090_), .Y(_7091_) );
OAI21X1 OAI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf4), .B(_7070_), .C(_7091_), .Y(_7092_) );
INVX1 INVX1_3079 ( .gnd(gnd), .vdd(vdd), .A(_7092_), .Y(_197__7_) );
INVX1 INVX1_3080 ( .gnd(gnd), .vdd(vdd), .A(data_46__8_), .Y(_7093_) );
OAI21X1 OAI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15170__bF_buf2), .C(_7093_), .Y(_7094_) );
NAND3X1 NAND3X1_955 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_14946__bF_buf1), .C(_15793__bF_buf4), .Y(_7095_) );
AND2X2 AND2X2_1352 ( .gnd(gnd), .vdd(vdd), .A(_7094_), .B(_7095_), .Y(_197__8_) );
NOR2X1 NOR2X1_747 ( .gnd(gnd), .vdd(vdd), .A(data_46__9_), .B(_7076_), .Y(_7096_) );
AOI21X1 AOI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_7076_), .C(_7096_), .Y(_197__9_) );
INVX1 INVX1_3081 ( .gnd(gnd), .vdd(vdd), .A(data_46__10_), .Y(_7097_) );
OAI21X1 OAI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15170__bF_buf1), .C(_7097_), .Y(_7098_) );
NAND3X1 NAND3X1_956 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_14946__bF_buf0), .C(_15793__bF_buf3), .Y(_7099_) );
AND2X2 AND2X2_1353 ( .gnd(gnd), .vdd(vdd), .A(_7098_), .B(_7099_), .Y(_197__10_) );
INVX1 INVX1_3082 ( .gnd(gnd), .vdd(vdd), .A(data_46__11_), .Y(_7100_) );
OAI21X1 OAI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15170__bF_buf0), .C(_7100_), .Y(_7101_) );
NAND3X1 NAND3X1_957 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_14946__bF_buf4), .C(_15793__bF_buf2), .Y(_7102_) );
AND2X2 AND2X2_1354 ( .gnd(gnd), .vdd(vdd), .A(_7101_), .B(_7102_), .Y(_197__11_) );
INVX1 INVX1_3083 ( .gnd(gnd), .vdd(vdd), .A(data_46__12_), .Y(_7103_) );
OAI21X1 OAI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15170__bF_buf3), .C(_7103_), .Y(_7104_) );
NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf10), .B(_7076_), .Y(_7105_) );
AND2X2 AND2X2_1355 ( .gnd(gnd), .vdd(vdd), .A(_7105_), .B(_7104_), .Y(_197__12_) );
INVX1 INVX1_3084 ( .gnd(gnd), .vdd(vdd), .A(data_46__13_), .Y(_7106_) );
OAI21X1 OAI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15170__bF_buf2), .C(_7106_), .Y(_7107_) );
OAI21X1 OAI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf3), .B(_7070_), .C(_7107_), .Y(_7108_) );
INVX1 INVX1_3085 ( .gnd(gnd), .vdd(vdd), .A(_7108_), .Y(_197__13_) );
INVX1 INVX1_3086 ( .gnd(gnd), .vdd(vdd), .A(data_46__14_), .Y(_7109_) );
OAI21X1 OAI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15170__bF_buf1), .C(_7109_), .Y(_7110_) );
OAI21X1 OAI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf0), .B(_7070_), .C(_7110_), .Y(_7111_) );
INVX1 INVX1_3087 ( .gnd(gnd), .vdd(vdd), .A(_7111_), .Y(_197__14_) );
NOR2X1 NOR2X1_748 ( .gnd(gnd), .vdd(vdd), .A(data_46__15_), .B(_7076_), .Y(_7112_) );
NOR2X1 NOR2X1_749 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf5), .B(_7070_), .Y(_7113_) );
NOR2X1 NOR2X1_750 ( .gnd(gnd), .vdd(vdd), .A(_7113_), .B(_7112_), .Y(_197__15_) );
INVX1 INVX1_3088 ( .gnd(gnd), .vdd(vdd), .A(data_45__0_), .Y(_7114_) );
NOR2X1 NOR2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf0), .B(_3942_), .Y(_7115_) );
AOI21X1 AOI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(_3313__bF_buf57), .C(_7115_), .Y(_7116_) );
AOI21X1 AOI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf3), .B(_3983_), .C(_3317_), .Y(_7117_) );
NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_7117_), .B(_7116_), .Y(_7118_) );
NOR2X1 NOR2X1_752 ( .gnd(gnd), .vdd(vdd), .A(_3353__bF_buf3), .B(_3393__bF_buf52), .Y(_7119_) );
OAI21X1 OAI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_15078_), .B(_14957_), .C(_14946__bF_buf2), .Y(_7120_) );
NAND3X1 NAND3X1_958 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_7025_), .C(_7120_), .Y(_7121_) );
NOR2X1 NOR2X1_753 ( .gnd(gnd), .vdd(vdd), .A(_7121_), .B(_3386_), .Y(_7122_) );
NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_7122_), .B(_7119_), .Y(_7123_) );
OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf3), .B(_7118__bF_buf9), .Y(_7124_) );
NOR3X1 NOR3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf8), .B(IDATA_PROG_data_0_bF_buf2), .C(_7123__bF_buf2), .Y(_7125_) );
AOI21X1 AOI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_7114_), .B(_7124_), .C(_7125_), .Y(_196__0_) );
INVX1 INVX1_3089 ( .gnd(gnd), .vdd(vdd), .A(data_45__1_), .Y(_7126_) );
NOR3X1 NOR3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf7), .B(IDATA_PROG_data_1_bF_buf3), .C(_7123__bF_buf1), .Y(_7127_) );
AOI21X1 AOI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_7126_), .B(_7124_), .C(_7127_), .Y(_196__1_) );
INVX1 INVX1_3090 ( .gnd(gnd), .vdd(vdd), .A(data_45__2_), .Y(_7128_) );
OAI21X1 OAI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf0), .B(_7118__bF_buf6), .C(_7128_), .Y(_7129_) );
OAI21X1 OAI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_2_bF_buf2), .C(_7129_), .Y(_7130_) );
INVX1 INVX1_3091 ( .gnd(gnd), .vdd(vdd), .A(_7130_), .Y(_196__2_) );
INVX1 INVX1_3092 ( .gnd(gnd), .vdd(vdd), .A(data_45__3_), .Y(_7131_) );
NOR3X1 NOR3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf5), .B(IDATA_PROG_data_3_bF_buf3), .C(_7123__bF_buf3), .Y(_7132_) );
AOI21X1 AOI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_7131_), .B(_7124_), .C(_7132_), .Y(_196__3_) );
INVX1 INVX1_3093 ( .gnd(gnd), .vdd(vdd), .A(data_45__4_), .Y(_7133_) );
NOR3X1 NOR3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf4), .B(IDATA_PROG_data_4_bF_buf1), .C(_7123__bF_buf2), .Y(_7134_) );
AOI21X1 AOI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_7133_), .B(_7124_), .C(_7134_), .Y(_196__4_) );
INVX1 INVX1_3094 ( .gnd(gnd), .vdd(vdd), .A(data_45__5_), .Y(_7135_) );
NOR3X1 NOR3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf3), .B(IDATA_PROG_data_5_bF_buf4), .C(_7123__bF_buf1), .Y(_7136_) );
AOI21X1 AOI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_7135_), .B(_7124_), .C(_7136_), .Y(_196__5_) );
INVX1 INVX1_3095 ( .gnd(gnd), .vdd(vdd), .A(data_45__6_), .Y(_7137_) );
OAI21X1 OAI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf0), .B(_7118__bF_buf2), .C(_7137_), .Y(_7138_) );
OAI21X1 OAI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_6_bF_buf4), .C(_7138_), .Y(_7139_) );
INVX1 INVX1_3096 ( .gnd(gnd), .vdd(vdd), .A(_7139_), .Y(_196__6_) );
INVX1 INVX1_3097 ( .gnd(gnd), .vdd(vdd), .A(data_45__7_), .Y(_7140_) );
NOR3X1 NOR3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf1), .B(IDATA_PROG_data_7_bF_buf3), .C(_7123__bF_buf3), .Y(_7141_) );
AOI21X1 AOI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_7140_), .B(_7124_), .C(_7141_), .Y(_196__7_) );
INVX1 INVX1_3098 ( .gnd(gnd), .vdd(vdd), .A(data_45__8_), .Y(_7142_) );
OAI21X1 OAI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf2), .B(_7118__bF_buf0), .C(_7142_), .Y(_7143_) );
OAI21X1 OAI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_8_bF_buf2), .C(_7143_), .Y(_7144_) );
INVX1 INVX1_3099 ( .gnd(gnd), .vdd(vdd), .A(_7144_), .Y(_196__8_) );
INVX1 INVX1_3100 ( .gnd(gnd), .vdd(vdd), .A(data_45__9_), .Y(_7145_) );
OAI21X1 OAI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf1), .B(_7118__bF_buf9), .C(_7145_), .Y(_7146_) );
OAI21X1 OAI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_9_bF_buf1), .C(_7146_), .Y(_7147_) );
INVX1 INVX1_3101 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .Y(_196__9_) );
INVX1 INVX1_3102 ( .gnd(gnd), .vdd(vdd), .A(data_45__10_), .Y(_7148_) );
OAI21X1 OAI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf0), .B(_7118__bF_buf8), .C(_7148_), .Y(_7149_) );
OAI21X1 OAI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_10_bF_buf1), .C(_7149_), .Y(_7150_) );
INVX1 INVX1_3103 ( .gnd(gnd), .vdd(vdd), .A(_7150_), .Y(_196__10_) );
INVX1 INVX1_3104 ( .gnd(gnd), .vdd(vdd), .A(data_45__11_), .Y(_7151_) );
NOR3X1 NOR3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf7), .B(IDATA_PROG_data_11_bF_buf4), .C(_7123__bF_buf3), .Y(_7152_) );
AOI21X1 AOI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_7151_), .B(_7124_), .C(_7152_), .Y(_196__11_) );
INVX1 INVX1_3105 ( .gnd(gnd), .vdd(vdd), .A(data_45__12_), .Y(_7153_) );
NOR3X1 NOR3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf6), .B(IDATA_PROG_data_12_bF_buf4), .C(_7123__bF_buf2), .Y(_7154_) );
AOI21X1 AOI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_7153_), .B(_7124_), .C(_7154_), .Y(_196__12_) );
INVX1 INVX1_3106 ( .gnd(gnd), .vdd(vdd), .A(data_45__13_), .Y(_7155_) );
OAI21X1 OAI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf1), .B(_7118__bF_buf5), .C(_7155_), .Y(_7156_) );
OAI21X1 OAI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_13_bF_buf2), .C(_7156_), .Y(_7157_) );
INVX1 INVX1_3107 ( .gnd(gnd), .vdd(vdd), .A(_7157_), .Y(_196__13_) );
INVX1 INVX1_3108 ( .gnd(gnd), .vdd(vdd), .A(data_45__14_), .Y(_7158_) );
OAI21X1 OAI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf0), .B(_7118__bF_buf4), .C(_7158_), .Y(_7159_) );
OAI21X1 OAI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_14_bF_buf4), .C(_7159_), .Y(_7160_) );
INVX1 INVX1_3109 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .Y(_196__14_) );
INVX1 INVX1_3110 ( .gnd(gnd), .vdd(vdd), .A(data_45__15_), .Y(_7161_) );
OAI21X1 OAI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_7123__bF_buf3), .B(_7118__bF_buf3), .C(_7161_), .Y(_7162_) );
OAI21X1 OAI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_7124_), .B(IDATA_PROG_data_15_bF_buf4), .C(_7162_), .Y(_7163_) );
INVX1 INVX1_3111 ( .gnd(gnd), .vdd(vdd), .A(_7163_), .Y(_196__15_) );
INVX1 INVX1_3112 ( .gnd(gnd), .vdd(vdd), .A(data_44__0_), .Y(_7164_) );
OAI21X1 OAI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_14957_), .B(_14961_), .C(_14946__bF_buf1), .Y(_7165_) );
NOR2X1 NOR2X1_754 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf11), .B(_3386_), .Y(_7166_) );
NAND3X1 NAND3X1_959 ( .gnd(gnd), .vdd(vdd), .A(_7165_), .B(_7166_), .C(_7119_), .Y(_7167_) );
OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf3), .B(_7118__bF_buf2), .Y(_7168_) );
NOR3X1 NOR3X1_156 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf1), .B(_7118__bF_buf1), .C(_7167__bF_buf2), .Y(_7169_) );
AOI21X1 AOI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_7164_), .B(_7168_), .C(_7169_), .Y(_195__0_) );
INVX1 INVX1_3113 ( .gnd(gnd), .vdd(vdd), .A(data_44__1_), .Y(_7170_) );
NOR3X1 NOR3X1_157 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf2), .B(_7118__bF_buf0), .C(_7167__bF_buf1), .Y(_7171_) );
AOI21X1 AOI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_7170_), .B(_7168_), .C(_7171_), .Y(_195__1_) );
INVX1 INVX1_3114 ( .gnd(gnd), .vdd(vdd), .A(data_44__2_), .Y(_7172_) );
OAI21X1 OAI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf0), .B(_7118__bF_buf9), .C(_7172_), .Y(_7173_) );
OAI21X1 OAI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_2_bF_buf1), .C(_7173_), .Y(_7174_) );
INVX1 INVX1_3115 ( .gnd(gnd), .vdd(vdd), .A(_7174_), .Y(_195__2_) );
INVX1 INVX1_3116 ( .gnd(gnd), .vdd(vdd), .A(data_44__3_), .Y(_7175_) );
NOR3X1 NOR3X1_158 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf2), .B(_7118__bF_buf8), .C(_7167__bF_buf3), .Y(_7176_) );
AOI21X1 AOI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_7175_), .B(_7168_), .C(_7176_), .Y(_195__3_) );
INVX1 INVX1_3117 ( .gnd(gnd), .vdd(vdd), .A(data_44__4_), .Y(_7177_) );
NOR3X1 NOR3X1_159 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf0), .B(_7118__bF_buf7), .C(_7167__bF_buf2), .Y(_7178_) );
AOI21X1 AOI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_7177_), .B(_7168_), .C(_7178_), .Y(_195__4_) );
INVX1 INVX1_3118 ( .gnd(gnd), .vdd(vdd), .A(data_44__5_), .Y(_7179_) );
NOR3X1 NOR3X1_160 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf3), .B(_7118__bF_buf6), .C(_7167__bF_buf1), .Y(_7180_) );
AOI21X1 AOI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_7179_), .B(_7168_), .C(_7180_), .Y(_195__5_) );
INVX1 INVX1_3119 ( .gnd(gnd), .vdd(vdd), .A(data_44__6_), .Y(_7181_) );
OAI21X1 OAI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf0), .B(_7118__bF_buf5), .C(_7181_), .Y(_7182_) );
OAI21X1 OAI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_6_bF_buf3), .C(_7182_), .Y(_7183_) );
INVX1 INVX1_3120 ( .gnd(gnd), .vdd(vdd), .A(_7183_), .Y(_195__6_) );
INVX1 INVX1_3121 ( .gnd(gnd), .vdd(vdd), .A(data_44__7_), .Y(_7184_) );
NOR3X1 NOR3X1_161 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf2), .B(_7118__bF_buf4), .C(_7167__bF_buf3), .Y(_7185_) );
AOI21X1 AOI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_7184_), .B(_7168_), .C(_7185_), .Y(_195__7_) );
INVX1 INVX1_3122 ( .gnd(gnd), .vdd(vdd), .A(data_44__8_), .Y(_7186_) );
OAI21X1 OAI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf2), .B(_7118__bF_buf3), .C(_7186_), .Y(_7187_) );
OAI21X1 OAI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_8_bF_buf1), .C(_7187_), .Y(_7188_) );
INVX1 INVX1_3123 ( .gnd(gnd), .vdd(vdd), .A(_7188_), .Y(_195__8_) );
INVX1 INVX1_3124 ( .gnd(gnd), .vdd(vdd), .A(data_44__9_), .Y(_7189_) );
OAI21X1 OAI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf1), .B(_7118__bF_buf2), .C(_7189_), .Y(_7190_) );
OAI21X1 OAI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_9_bF_buf0), .C(_7190_), .Y(_7191_) );
INVX1 INVX1_3125 ( .gnd(gnd), .vdd(vdd), .A(_7191_), .Y(_195__9_) );
INVX1 INVX1_3126 ( .gnd(gnd), .vdd(vdd), .A(data_44__10_), .Y(_7192_) );
OAI21X1 OAI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf0), .B(_7118__bF_buf1), .C(_7192_), .Y(_7193_) );
OAI21X1 OAI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_10_bF_buf0), .C(_7193_), .Y(_7194_) );
INVX1 INVX1_3127 ( .gnd(gnd), .vdd(vdd), .A(_7194_), .Y(_195__10_) );
INVX1 INVX1_3128 ( .gnd(gnd), .vdd(vdd), .A(data_44__11_), .Y(_7195_) );
NOR3X1 NOR3X1_162 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf3), .B(_7118__bF_buf0), .C(_7167__bF_buf3), .Y(_7196_) );
AOI21X1 AOI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_7195_), .B(_7168_), .C(_7196_), .Y(_195__11_) );
INVX1 INVX1_3129 ( .gnd(gnd), .vdd(vdd), .A(data_44__12_), .Y(_7197_) );
NOR3X1 NOR3X1_163 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf3), .B(_7118__bF_buf9), .C(_7167__bF_buf2), .Y(_7198_) );
AOI21X1 AOI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_7197_), .B(_7168_), .C(_7198_), .Y(_195__12_) );
INVX1 INVX1_3130 ( .gnd(gnd), .vdd(vdd), .A(data_44__13_), .Y(_7199_) );
OAI21X1 OAI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf1), .B(_7118__bF_buf8), .C(_7199_), .Y(_7200_) );
OAI21X1 OAI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_13_bF_buf1), .C(_7200_), .Y(_7201_) );
INVX1 INVX1_3131 ( .gnd(gnd), .vdd(vdd), .A(_7201_), .Y(_195__13_) );
INVX1 INVX1_3132 ( .gnd(gnd), .vdd(vdd), .A(data_44__14_), .Y(_7202_) );
OAI21X1 OAI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf0), .B(_7118__bF_buf7), .C(_7202_), .Y(_7203_) );
OAI21X1 OAI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_14_bF_buf3), .C(_7203_), .Y(_7204_) );
INVX1 INVX1_3133 ( .gnd(gnd), .vdd(vdd), .A(_7204_), .Y(_195__14_) );
INVX1 INVX1_3134 ( .gnd(gnd), .vdd(vdd), .A(data_44__15_), .Y(_7205_) );
OAI21X1 OAI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_7167__bF_buf3), .B(_7118__bF_buf6), .C(_7205_), .Y(_7206_) );
OAI21X1 OAI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_7168_), .B(IDATA_PROG_data_15_bF_buf3), .C(_7206_), .Y(_7207_) );
INVX1 INVX1_3135 ( .gnd(gnd), .vdd(vdd), .A(_7207_), .Y(_195__15_) );
INVX1 INVX1_3136 ( .gnd(gnd), .vdd(vdd), .A(data_43__0_), .Y(_7208_) );
OAI21X1 OAI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_14945_), .B(_14943_), .C(IDATA_PROG_write_bF_buf3), .Y(_7209_) );
NOR2X1 NOR2X1_755 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf10), .B(_14963__bF_buf3), .Y(_7210_) );
OAI21X1 OAI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_14982_), .B(_14989_), .C(_7210_), .Y(_7211_) );
OAI21X1 OAI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_7211_), .C(_7209_), .Y(_7212_) );
NAND3X1 NAND3X1_960 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .B(_7212_), .C(_7119_), .Y(_7213_) );
OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf3), .B(_7118__bF_buf5), .Y(_7214_) );
NOR3X1 NOR3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf4), .B(IDATA_PROG_data_0_bF_buf0), .C(_7213__bF_buf2), .Y(_7215_) );
AOI21X1 AOI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_7208_), .B(_7214_), .C(_7215_), .Y(_194__0_) );
INVX1 INVX1_3137 ( .gnd(gnd), .vdd(vdd), .A(data_43__1_), .Y(_7216_) );
NOR3X1 NOR3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf3), .B(IDATA_PROG_data_1_bF_buf1), .C(_7213__bF_buf1), .Y(_7217_) );
AOI21X1 AOI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_7216_), .B(_7214_), .C(_7217_), .Y(_194__1_) );
INVX1 INVX1_3138 ( .gnd(gnd), .vdd(vdd), .A(data_43__2_), .Y(_7218_) );
OAI21X1 OAI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf0), .B(_7118__bF_buf2), .C(_7218_), .Y(_7219_) );
OAI21X1 OAI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_2_bF_buf0), .C(_7219_), .Y(_7220_) );
INVX1 INVX1_3139 ( .gnd(gnd), .vdd(vdd), .A(_7220_), .Y(_194__2_) );
INVX1 INVX1_3140 ( .gnd(gnd), .vdd(vdd), .A(data_43__3_), .Y(_7221_) );
NOR3X1 NOR3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf1), .B(IDATA_PROG_data_3_bF_buf1), .C(_7213__bF_buf3), .Y(_7222_) );
AOI21X1 AOI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_7221_), .B(_7214_), .C(_7222_), .Y(_194__3_) );
INVX1 INVX1_3141 ( .gnd(gnd), .vdd(vdd), .A(data_43__4_), .Y(_7223_) );
NOR3X1 NOR3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf0), .B(IDATA_PROG_data_4_bF_buf4), .C(_7213__bF_buf2), .Y(_7224_) );
AOI21X1 AOI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_7223_), .B(_7214_), .C(_7224_), .Y(_194__4_) );
INVX1 INVX1_3142 ( .gnd(gnd), .vdd(vdd), .A(data_43__5_), .Y(_7225_) );
NOR3X1 NOR3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf9), .B(IDATA_PROG_data_5_bF_buf2), .C(_7213__bF_buf1), .Y(_7226_) );
AOI21X1 AOI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_7225_), .B(_7214_), .C(_7226_), .Y(_194__5_) );
INVX1 INVX1_3143 ( .gnd(gnd), .vdd(vdd), .A(data_43__6_), .Y(_7227_) );
OAI21X1 OAI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf0), .B(_7118__bF_buf8), .C(_7227_), .Y(_7228_) );
OAI21X1 OAI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_6_bF_buf2), .C(_7228_), .Y(_7229_) );
INVX1 INVX1_3144 ( .gnd(gnd), .vdd(vdd), .A(_7229_), .Y(_194__6_) );
INVX1 INVX1_3145 ( .gnd(gnd), .vdd(vdd), .A(data_43__7_), .Y(_7230_) );
NOR3X1 NOR3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf7), .B(IDATA_PROG_data_7_bF_buf1), .C(_7213__bF_buf3), .Y(_7231_) );
AOI21X1 AOI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_7230_), .B(_7214_), .C(_7231_), .Y(_194__7_) );
INVX1 INVX1_3146 ( .gnd(gnd), .vdd(vdd), .A(data_43__8_), .Y(_7232_) );
OAI21X1 OAI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf2), .B(_7118__bF_buf6), .C(_7232_), .Y(_7233_) );
OAI21X1 OAI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_8_bF_buf0), .C(_7233_), .Y(_7234_) );
INVX1 INVX1_3147 ( .gnd(gnd), .vdd(vdd), .A(_7234_), .Y(_194__8_) );
INVX1 INVX1_3148 ( .gnd(gnd), .vdd(vdd), .A(data_43__9_), .Y(_7235_) );
OAI21X1 OAI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf1), .B(_7118__bF_buf5), .C(_7235_), .Y(_7236_) );
OAI21X1 OAI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_9_bF_buf4), .C(_7236_), .Y(_7237_) );
INVX1 INVX1_3149 ( .gnd(gnd), .vdd(vdd), .A(_7237_), .Y(_194__9_) );
INVX1 INVX1_3150 ( .gnd(gnd), .vdd(vdd), .A(data_43__10_), .Y(_7238_) );
OAI21X1 OAI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf0), .B(_7118__bF_buf4), .C(_7238_), .Y(_7239_) );
OAI21X1 OAI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_10_bF_buf4), .C(_7239_), .Y(_7240_) );
INVX1 INVX1_3151 ( .gnd(gnd), .vdd(vdd), .A(_7240_), .Y(_194__10_) );
INVX1 INVX1_3152 ( .gnd(gnd), .vdd(vdd), .A(data_43__11_), .Y(_7241_) );
NOR3X1 NOR3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf3), .B(IDATA_PROG_data_11_bF_buf2), .C(_7213__bF_buf3), .Y(_7242_) );
AOI21X1 AOI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_7241_), .B(_7214_), .C(_7242_), .Y(_194__11_) );
INVX1 INVX1_3153 ( .gnd(gnd), .vdd(vdd), .A(data_43__12_), .Y(_7243_) );
NOR3X1 NOR3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf2), .B(IDATA_PROG_data_12_bF_buf2), .C(_7213__bF_buf2), .Y(_7244_) );
AOI21X1 AOI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_7243_), .B(_7214_), .C(_7244_), .Y(_194__12_) );
INVX1 INVX1_3154 ( .gnd(gnd), .vdd(vdd), .A(data_43__13_), .Y(_7245_) );
OAI21X1 OAI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf1), .B(_7118__bF_buf1), .C(_7245_), .Y(_7246_) );
OAI21X1 OAI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_13_bF_buf0), .C(_7246_), .Y(_7247_) );
INVX1 INVX1_3155 ( .gnd(gnd), .vdd(vdd), .A(_7247_), .Y(_194__13_) );
INVX1 INVX1_3156 ( .gnd(gnd), .vdd(vdd), .A(data_43__14_), .Y(_7248_) );
OAI21X1 OAI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf0), .B(_7118__bF_buf0), .C(_7248_), .Y(_7249_) );
OAI21X1 OAI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_14_bF_buf2), .C(_7249_), .Y(_7250_) );
INVX1 INVX1_3157 ( .gnd(gnd), .vdd(vdd), .A(_7250_), .Y(_194__14_) );
INVX1 INVX1_3158 ( .gnd(gnd), .vdd(vdd), .A(data_43__15_), .Y(_7251_) );
OAI21X1 OAI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_7213__bF_buf3), .B(_7118__bF_buf9), .C(_7251_), .Y(_7252_) );
OAI21X1 OAI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_7214_), .B(IDATA_PROG_data_15_bF_buf2), .C(_7252_), .Y(_7253_) );
INVX1 INVX1_3159 ( .gnd(gnd), .vdd(vdd), .A(_7253_), .Y(_194__15_) );
INVX1 INVX1_3160 ( .gnd(gnd), .vdd(vdd), .A(data_42__0_), .Y(_7254_) );
NOR2X1 NOR2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_14989_), .B(_15170__bF_buf3), .Y(_7255_) );
INVX1 INVX1_3161 ( .gnd(gnd), .vdd(vdd), .A(_7209_), .Y(_7256_) );
OAI21X1 OAI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_7256_), .C(_15069_), .Y(_7257_) );
AOI21X1 AOI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_14949_), .B(_7255_), .C(_7257_), .Y(_7258_) );
NAND3X1 NAND3X1_961 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .B(_7258_), .C(_7119_), .Y(_7259_) );
OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf3), .B(_7118__bF_buf8), .Y(_7260_) );
NOR3X1 NOR3X1_172 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf4), .B(_7118__bF_buf7), .C(_7259__bF_buf2), .Y(_7261_) );
AOI21X1 AOI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_7254_), .B(_7260_), .C(_7261_), .Y(_193__0_) );
INVX1 INVX1_3162 ( .gnd(gnd), .vdd(vdd), .A(data_42__1_), .Y(_7262_) );
NOR3X1 NOR3X1_173 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf0), .B(_7118__bF_buf6), .C(_7259__bF_buf1), .Y(_7263_) );
AOI21X1 AOI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_7262_), .B(_7260_), .C(_7263_), .Y(_193__1_) );
INVX1 INVX1_3163 ( .gnd(gnd), .vdd(vdd), .A(data_42__2_), .Y(_7264_) );
OAI21X1 OAI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf0), .B(_7118__bF_buf5), .C(_7264_), .Y(_7265_) );
OAI21X1 OAI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_2_bF_buf3), .C(_7265_), .Y(_7266_) );
INVX1 INVX1_3164 ( .gnd(gnd), .vdd(vdd), .A(_7266_), .Y(_193__2_) );
INVX1 INVX1_3165 ( .gnd(gnd), .vdd(vdd), .A(data_42__3_), .Y(_7267_) );
NOR3X1 NOR3X1_174 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf0), .B(_7118__bF_buf4), .C(_7259__bF_buf3), .Y(_7268_) );
AOI21X1 AOI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_7267_), .B(_7260_), .C(_7268_), .Y(_193__3_) );
INVX1 INVX1_3166 ( .gnd(gnd), .vdd(vdd), .A(data_42__4_), .Y(_7269_) );
NOR3X1 NOR3X1_175 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf3), .B(_7118__bF_buf3), .C(_7259__bF_buf2), .Y(_7270_) );
AOI21X1 AOI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_7269_), .B(_7260_), .C(_7270_), .Y(_193__4_) );
INVX1 INVX1_3167 ( .gnd(gnd), .vdd(vdd), .A(data_42__5_), .Y(_7271_) );
NOR3X1 NOR3X1_176 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf1), .B(_7118__bF_buf2), .C(_7259__bF_buf1), .Y(_7272_) );
AOI21X1 AOI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_7271_), .B(_7260_), .C(_7272_), .Y(_193__5_) );
INVX1 INVX1_3168 ( .gnd(gnd), .vdd(vdd), .A(data_42__6_), .Y(_7273_) );
OAI21X1 OAI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf0), .B(_7118__bF_buf1), .C(_7273_), .Y(_7274_) );
OAI21X1 OAI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_6_bF_buf1), .C(_7274_), .Y(_7275_) );
INVX1 INVX1_3169 ( .gnd(gnd), .vdd(vdd), .A(_7275_), .Y(_193__6_) );
INVX1 INVX1_3170 ( .gnd(gnd), .vdd(vdd), .A(data_42__7_), .Y(_7276_) );
NOR3X1 NOR3X1_177 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf0), .B(_7118__bF_buf0), .C(_7259__bF_buf3), .Y(_7277_) );
AOI21X1 AOI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_7276_), .B(_7260_), .C(_7277_), .Y(_193__7_) );
INVX1 INVX1_3171 ( .gnd(gnd), .vdd(vdd), .A(data_42__8_), .Y(_7278_) );
OAI21X1 OAI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf2), .B(_7118__bF_buf9), .C(_7278_), .Y(_7279_) );
OAI21X1 OAI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_8_bF_buf4), .C(_7279_), .Y(_7280_) );
INVX1 INVX1_3172 ( .gnd(gnd), .vdd(vdd), .A(_7280_), .Y(_193__8_) );
INVX1 INVX1_3173 ( .gnd(gnd), .vdd(vdd), .A(data_42__9_), .Y(_7281_) );
OAI21X1 OAI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf1), .B(_7118__bF_buf8), .C(_7281_), .Y(_7282_) );
OAI21X1 OAI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_9_bF_buf3), .C(_7282_), .Y(_7283_) );
INVX1 INVX1_3174 ( .gnd(gnd), .vdd(vdd), .A(_7283_), .Y(_193__9_) );
INVX1 INVX1_3175 ( .gnd(gnd), .vdd(vdd), .A(data_42__10_), .Y(_7284_) );
OAI21X1 OAI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf0), .B(_7118__bF_buf7), .C(_7284_), .Y(_7285_) );
OAI21X1 OAI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_10_bF_buf3), .C(_7285_), .Y(_7286_) );
INVX1 INVX1_3176 ( .gnd(gnd), .vdd(vdd), .A(_7286_), .Y(_193__10_) );
INVX1 INVX1_3177 ( .gnd(gnd), .vdd(vdd), .A(data_42__11_), .Y(_7287_) );
NOR3X1 NOR3X1_178 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf1), .B(_7118__bF_buf6), .C(_7259__bF_buf3), .Y(_7288_) );
AOI21X1 AOI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_7287_), .B(_7260_), .C(_7288_), .Y(_193__11_) );
INVX1 INVX1_3178 ( .gnd(gnd), .vdd(vdd), .A(data_42__12_), .Y(_7289_) );
NOR3X1 NOR3X1_179 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf1), .B(_7118__bF_buf5), .C(_7259__bF_buf2), .Y(_7290_) );
AOI21X1 AOI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_7289_), .B(_7260_), .C(_7290_), .Y(_193__12_) );
INVX1 INVX1_3179 ( .gnd(gnd), .vdd(vdd), .A(data_42__13_), .Y(_7291_) );
OAI21X1 OAI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf1), .B(_7118__bF_buf4), .C(_7291_), .Y(_7292_) );
OAI21X1 OAI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_13_bF_buf4), .C(_7292_), .Y(_7293_) );
INVX1 INVX1_3180 ( .gnd(gnd), .vdd(vdd), .A(_7293_), .Y(_193__13_) );
INVX1 INVX1_3181 ( .gnd(gnd), .vdd(vdd), .A(data_42__14_), .Y(_7294_) );
OAI21X1 OAI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf0), .B(_7118__bF_buf3), .C(_7294_), .Y(_7295_) );
OAI21X1 OAI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_14_bF_buf1), .C(_7295_), .Y(_7296_) );
INVX1 INVX1_3182 ( .gnd(gnd), .vdd(vdd), .A(_7296_), .Y(_193__14_) );
INVX1 INVX1_3183 ( .gnd(gnd), .vdd(vdd), .A(data_42__15_), .Y(_7297_) );
OAI21X1 OAI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_7259__bF_buf3), .B(_7118__bF_buf2), .C(_7297_), .Y(_7298_) );
OAI21X1 OAI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_7260_), .B(IDATA_PROG_data_15_bF_buf1), .C(_7298_), .Y(_7299_) );
INVX1 INVX1_3184 ( .gnd(gnd), .vdd(vdd), .A(_7299_), .Y(_193__15_) );
INVX1 INVX1_3185 ( .gnd(gnd), .vdd(vdd), .A(data_41__0_), .Y(_7300_) );
AOI21X1 AOI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf0), .B(_15285_), .C(_7257_), .Y(_7301_) );
NAND3X1 NAND3X1_962 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .B(_7301_), .C(_7119_), .Y(_7302_) );
OR2X2 OR2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf3), .B(_7118__bF_buf1), .Y(_7303_) );
NOR3X1 NOR3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf0), .B(IDATA_PROG_data_0_bF_buf3), .C(_7302__bF_buf2), .Y(_7304_) );
AOI21X1 AOI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_7300_), .B(_7303_), .C(_7304_), .Y(_192__0_) );
INVX1 INVX1_3186 ( .gnd(gnd), .vdd(vdd), .A(data_41__1_), .Y(_7305_) );
NOR3X1 NOR3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf9), .B(IDATA_PROG_data_1_bF_buf4), .C(_7302__bF_buf1), .Y(_7306_) );
AOI21X1 AOI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_7305_), .B(_7303_), .C(_7306_), .Y(_192__1_) );
INVX1 INVX1_3187 ( .gnd(gnd), .vdd(vdd), .A(data_41__2_), .Y(_7307_) );
OAI21X1 OAI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf0), .B(_7118__bF_buf8), .C(_7307_), .Y(_7308_) );
OAI21X1 OAI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_2_bF_buf2), .C(_7308_), .Y(_7309_) );
INVX1 INVX1_3188 ( .gnd(gnd), .vdd(vdd), .A(_7309_), .Y(_192__2_) );
INVX1 INVX1_3189 ( .gnd(gnd), .vdd(vdd), .A(data_41__3_), .Y(_7310_) );
NOR3X1 NOR3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf7), .B(IDATA_PROG_data_3_bF_buf4), .C(_7302__bF_buf3), .Y(_7311_) );
AOI21X1 AOI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_7310_), .B(_7303_), .C(_7311_), .Y(_192__3_) );
INVX1 INVX1_3190 ( .gnd(gnd), .vdd(vdd), .A(data_41__4_), .Y(_7312_) );
NOR3X1 NOR3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf6), .B(IDATA_PROG_data_4_bF_buf2), .C(_7302__bF_buf2), .Y(_7313_) );
AOI21X1 AOI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_7312_), .B(_7303_), .C(_7313_), .Y(_192__4_) );
INVX1 INVX1_3191 ( .gnd(gnd), .vdd(vdd), .A(data_41__5_), .Y(_7314_) );
NOR3X1 NOR3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf5), .B(IDATA_PROG_data_5_bF_buf0), .C(_7302__bF_buf1), .Y(_7315_) );
AOI21X1 AOI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_7314_), .B(_7303_), .C(_7315_), .Y(_192__5_) );
INVX1 INVX1_3192 ( .gnd(gnd), .vdd(vdd), .A(data_41__6_), .Y(_7316_) );
OAI21X1 OAI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf0), .B(_7118__bF_buf4), .C(_7316_), .Y(_7317_) );
OAI21X1 OAI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_6_bF_buf0), .C(_7317_), .Y(_7318_) );
INVX1 INVX1_3193 ( .gnd(gnd), .vdd(vdd), .A(_7318_), .Y(_192__6_) );
INVX1 INVX1_3194 ( .gnd(gnd), .vdd(vdd), .A(data_41__7_), .Y(_7319_) );
NOR3X1 NOR3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf3), .B(IDATA_PROG_data_7_bF_buf5), .C(_7302__bF_buf3), .Y(_7320_) );
AOI21X1 AOI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_7319_), .B(_7303_), .C(_7320_), .Y(_192__7_) );
INVX1 INVX1_3195 ( .gnd(gnd), .vdd(vdd), .A(data_41__8_), .Y(_7321_) );
OAI21X1 OAI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf2), .B(_7118__bF_buf2), .C(_7321_), .Y(_7322_) );
OAI21X1 OAI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_8_bF_buf3), .C(_7322_), .Y(_7323_) );
INVX1 INVX1_3196 ( .gnd(gnd), .vdd(vdd), .A(_7323_), .Y(_192__8_) );
INVX1 INVX1_3197 ( .gnd(gnd), .vdd(vdd), .A(data_41__9_), .Y(_7324_) );
OAI21X1 OAI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf1), .B(_7118__bF_buf1), .C(_7324_), .Y(_7325_) );
OAI21X1 OAI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_9_bF_buf2), .C(_7325_), .Y(_7326_) );
INVX1 INVX1_3198 ( .gnd(gnd), .vdd(vdd), .A(_7326_), .Y(_192__9_) );
INVX1 INVX1_3199 ( .gnd(gnd), .vdd(vdd), .A(data_41__10_), .Y(_7327_) );
OAI21X1 OAI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf0), .B(_7118__bF_buf0), .C(_7327_), .Y(_7328_) );
OAI21X1 OAI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_10_bF_buf2), .C(_7328_), .Y(_7329_) );
INVX1 INVX1_3200 ( .gnd(gnd), .vdd(vdd), .A(_7329_), .Y(_192__10_) );
INVX1 INVX1_3201 ( .gnd(gnd), .vdd(vdd), .A(data_41__11_), .Y(_7330_) );
NOR3X1 NOR3X1_186 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf9), .B(IDATA_PROG_data_11_bF_buf0), .C(_7302__bF_buf3), .Y(_7331_) );
AOI21X1 AOI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_7330_), .B(_7303_), .C(_7331_), .Y(_192__11_) );
INVX1 INVX1_3202 ( .gnd(gnd), .vdd(vdd), .A(data_41__12_), .Y(_7332_) );
NOR3X1 NOR3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf8), .B(IDATA_PROG_data_12_bF_buf0), .C(_7302__bF_buf2), .Y(_7333_) );
AOI21X1 AOI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_7332_), .B(_7303_), .C(_7333_), .Y(_192__12_) );
INVX1 INVX1_3203 ( .gnd(gnd), .vdd(vdd), .A(data_41__13_), .Y(_7334_) );
OAI21X1 OAI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf1), .B(_7118__bF_buf7), .C(_7334_), .Y(_7335_) );
OAI21X1 OAI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_13_bF_buf3), .C(_7335_), .Y(_7336_) );
INVX1 INVX1_3204 ( .gnd(gnd), .vdd(vdd), .A(_7336_), .Y(_192__13_) );
INVX1 INVX1_3205 ( .gnd(gnd), .vdd(vdd), .A(data_41__14_), .Y(_7337_) );
OAI21X1 OAI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf0), .B(_7118__bF_buf6), .C(_7337_), .Y(_7338_) );
OAI21X1 OAI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_14_bF_buf0), .C(_7338_), .Y(_7339_) );
INVX1 INVX1_3206 ( .gnd(gnd), .vdd(vdd), .A(_7339_), .Y(_192__14_) );
INVX1 INVX1_3207 ( .gnd(gnd), .vdd(vdd), .A(data_41__15_), .Y(_7340_) );
OAI21X1 OAI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_7302__bF_buf3), .B(_7118__bF_buf5), .C(_7340_), .Y(_7341_) );
OAI21X1 OAI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_7303_), .B(IDATA_PROG_data_15_bF_buf0), .C(_7341_), .Y(_7342_) );
INVX1 INVX1_3208 ( .gnd(gnd), .vdd(vdd), .A(_7342_), .Y(_192__15_) );
INVX1 INVX1_3209 ( .gnd(gnd), .vdd(vdd), .A(data_40__0_), .Y(_7343_) );
NOR2X1 NOR2X1_757 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_3386_), .Y(_7344_) );
NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_7344_), .B(_7119_), .Y(_7345_) );
OR2X2 OR2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf3), .B(_7118__bF_buf4), .Y(_7346_) );
NOR3X1 NOR3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf3), .B(IDATA_PROG_data_0_bF_buf2), .C(_7345__bF_buf2), .Y(_7347_) );
AOI21X1 AOI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_7343_), .B(_7346_), .C(_7347_), .Y(_191__0_) );
INVX1 INVX1_3210 ( .gnd(gnd), .vdd(vdd), .A(data_40__1_), .Y(_7348_) );
NOR3X1 NOR3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf2), .B(IDATA_PROG_data_1_bF_buf3), .C(_7345__bF_buf1), .Y(_7349_) );
AOI21X1 AOI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_7348_), .B(_7346_), .C(_7349_), .Y(_191__1_) );
INVX1 INVX1_3211 ( .gnd(gnd), .vdd(vdd), .A(data_40__2_), .Y(_7350_) );
OAI21X1 OAI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf0), .B(_7118__bF_buf1), .C(_7350_), .Y(_7351_) );
OAI21X1 OAI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_2_bF_buf1), .C(_7351_), .Y(_7352_) );
INVX1 INVX1_3212 ( .gnd(gnd), .vdd(vdd), .A(_7352_), .Y(_191__2_) );
INVX1 INVX1_3213 ( .gnd(gnd), .vdd(vdd), .A(data_40__3_), .Y(_7353_) );
NOR3X1 NOR3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf0), .B(IDATA_PROG_data_3_bF_buf3), .C(_7345__bF_buf3), .Y(_7354_) );
AOI21X1 AOI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_7353_), .B(_7346_), .C(_7354_), .Y(_191__3_) );
INVX1 INVX1_3214 ( .gnd(gnd), .vdd(vdd), .A(data_40__4_), .Y(_7355_) );
NOR3X1 NOR3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf9), .B(IDATA_PROG_data_4_bF_buf1), .C(_7345__bF_buf2), .Y(_7356_) );
AOI21X1 AOI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_7355_), .B(_7346_), .C(_7356_), .Y(_191__4_) );
INVX1 INVX1_3215 ( .gnd(gnd), .vdd(vdd), .A(data_40__5_), .Y(_7357_) );
NOR3X1 NOR3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf8), .B(IDATA_PROG_data_5_bF_buf4), .C(_7345__bF_buf1), .Y(_7358_) );
AOI21X1 AOI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_7357_), .B(_7346_), .C(_7358_), .Y(_191__5_) );
INVX1 INVX1_3216 ( .gnd(gnd), .vdd(vdd), .A(data_40__6_), .Y(_7359_) );
OAI21X1 OAI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf0), .B(_7118__bF_buf7), .C(_7359_), .Y(_7360_) );
OAI21X1 OAI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_6_bF_buf4), .C(_7360_), .Y(_7361_) );
INVX1 INVX1_3217 ( .gnd(gnd), .vdd(vdd), .A(_7361_), .Y(_191__6_) );
INVX1 INVX1_3218 ( .gnd(gnd), .vdd(vdd), .A(data_40__7_), .Y(_7362_) );
NOR3X1 NOR3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf6), .B(IDATA_PROG_data_7_bF_buf4), .C(_7345__bF_buf3), .Y(_7363_) );
AOI21X1 AOI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_7362_), .B(_7346_), .C(_7363_), .Y(_191__7_) );
INVX1 INVX1_3219 ( .gnd(gnd), .vdd(vdd), .A(data_40__8_), .Y(_7364_) );
OAI21X1 OAI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf2), .B(_7118__bF_buf5), .C(_7364_), .Y(_7365_) );
OAI21X1 OAI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_8_bF_buf2), .C(_7365_), .Y(_7366_) );
INVX1 INVX1_3220 ( .gnd(gnd), .vdd(vdd), .A(_7366_), .Y(_191__8_) );
INVX1 INVX1_3221 ( .gnd(gnd), .vdd(vdd), .A(data_40__9_), .Y(_7367_) );
OAI21X1 OAI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf1), .B(_7118__bF_buf4), .C(_7367_), .Y(_7368_) );
OAI21X1 OAI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_9_bF_buf1), .C(_7368_), .Y(_7369_) );
INVX1 INVX1_3222 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .Y(_191__9_) );
INVX1 INVX1_3223 ( .gnd(gnd), .vdd(vdd), .A(data_40__10_), .Y(_7370_) );
OAI21X1 OAI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf0), .B(_7118__bF_buf3), .C(_7370_), .Y(_7371_) );
OAI21X1 OAI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_10_bF_buf1), .C(_7371_), .Y(_7372_) );
INVX1 INVX1_3224 ( .gnd(gnd), .vdd(vdd), .A(_7372_), .Y(_191__10_) );
INVX1 INVX1_3225 ( .gnd(gnd), .vdd(vdd), .A(data_40__11_), .Y(_7373_) );
NOR3X1 NOR3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf2), .B(IDATA_PROG_data_11_bF_buf4), .C(_7345__bF_buf3), .Y(_7374_) );
AOI21X1 AOI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_7373_), .B(_7346_), .C(_7374_), .Y(_191__11_) );
INVX1 INVX1_3226 ( .gnd(gnd), .vdd(vdd), .A(data_40__12_), .Y(_7375_) );
NOR3X1 NOR3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_7118__bF_buf1), .B(IDATA_PROG_data_12_bF_buf4), .C(_7345__bF_buf2), .Y(_7376_) );
AOI21X1 AOI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_7375_), .B(_7346_), .C(_7376_), .Y(_191__12_) );
INVX1 INVX1_3227 ( .gnd(gnd), .vdd(vdd), .A(data_40__13_), .Y(_7377_) );
OAI21X1 OAI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf1), .B(_7118__bF_buf0), .C(_7377_), .Y(_7378_) );
OAI21X1 OAI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_13_bF_buf2), .C(_7378_), .Y(_7379_) );
INVX1 INVX1_3228 ( .gnd(gnd), .vdd(vdd), .A(_7379_), .Y(_191__13_) );
INVX1 INVX1_3229 ( .gnd(gnd), .vdd(vdd), .A(data_40__14_), .Y(_7380_) );
OAI21X1 OAI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf0), .B(_7118__bF_buf9), .C(_7380_), .Y(_7381_) );
OAI21X1 OAI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_14_bF_buf4), .C(_7381_), .Y(_7382_) );
INVX1 INVX1_3230 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .Y(_191__14_) );
INVX1 INVX1_3231 ( .gnd(gnd), .vdd(vdd), .A(data_40__15_), .Y(_7383_) );
OAI21X1 OAI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_7345__bF_buf3), .B(_7118__bF_buf8), .C(_7383_), .Y(_7384_) );
OAI21X1 OAI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_7346_), .B(IDATA_PROG_data_15_bF_buf5), .C(_7384_), .Y(_7385_) );
INVX1 INVX1_3232 ( .gnd(gnd), .vdd(vdd), .A(_7385_), .Y(_191__15_) );
INVX1 INVX1_3233 ( .gnd(gnd), .vdd(vdd), .A(data_39__0_), .Y(_7386_) );
NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf4), .B(_16156_), .Y(_7387_) );
OAI21X1 OAI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_3400_), .C(_7387_), .Y(_7388_) );
OR2X2 OR2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_3317_), .B(_15072_), .Y(_7389_) );
AOI21X1 AOI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_14946__bF_buf3), .B(_15363_), .C(_7389_), .Y(_7390_) );
NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf2), .B(_7390_), .Y(_7391_) );
NOR2X1 NOR2X1_758 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .B(_7391_), .Y(_7392_) );
NAND3X1 NAND3X1_963 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf2), .B(_7392_), .C(_3313__bF_buf56), .Y(_7393_) );
OAI21X1 OAI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7386_), .Y(_7394_) );
OR2X2 OR2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_7391_), .B(_3386_), .Y(_7395_) );
NOR3X1 NOR3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf50), .B(_3353__bF_buf2), .C(_7395_), .Y(_7396_) );
NAND3X1 NAND3X1_964 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf5), .B(_7116_), .C(_7396_), .Y(_7397_) );
AND2X2 AND2X2_1356 ( .gnd(gnd), .vdd(vdd), .A(_7397_), .B(_7394_), .Y(_189__0_) );
INVX1 INVX1_3234 ( .gnd(gnd), .vdd(vdd), .A(data_39__1_), .Y(_7398_) );
OAI21X1 OAI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7398_), .Y(_7399_) );
NAND3X1 NAND3X1_965 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_7116_), .C(_7396_), .Y(_7400_) );
AND2X2 AND2X2_1357 ( .gnd(gnd), .vdd(vdd), .A(_7400_), .B(_7399_), .Y(_189__1_) );
NOR2X1 NOR2X1_759 ( .gnd(gnd), .vdd(vdd), .A(_7393_), .B(_7388_), .Y(_7401_) );
NOR2X1 NOR2X1_760 ( .gnd(gnd), .vdd(vdd), .A(data_39__2_), .B(_7401_), .Y(_7402_) );
AOI21X1 AOI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_7401_), .C(_7402_), .Y(_189__2_) );
INVX1 INVX1_3235 ( .gnd(gnd), .vdd(vdd), .A(data_39__3_), .Y(_7403_) );
OAI21X1 OAI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7403_), .Y(_7404_) );
NAND3X1 NAND3X1_966 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_7116_), .C(_7396_), .Y(_7405_) );
AND2X2 AND2X2_1358 ( .gnd(gnd), .vdd(vdd), .A(_7405_), .B(_7404_), .Y(_189__3_) );
INVX1 INVX1_3236 ( .gnd(gnd), .vdd(vdd), .A(data_39__4_), .Y(_7406_) );
OAI21X1 OAI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7406_), .Y(_7407_) );
NAND3X1 NAND3X1_967 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_7116_), .C(_7396_), .Y(_7408_) );
AND2X2 AND2X2_1359 ( .gnd(gnd), .vdd(vdd), .A(_7408_), .B(_7407_), .Y(_189__4_) );
INVX1 INVX1_3237 ( .gnd(gnd), .vdd(vdd), .A(data_39__5_), .Y(_7409_) );
OAI21X1 OAI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7409_), .Y(_7410_) );
NAND3X1 NAND3X1_968 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_7116_), .C(_7396_), .Y(_7411_) );
AND2X2 AND2X2_1360 ( .gnd(gnd), .vdd(vdd), .A(_7411_), .B(_7410_), .Y(_189__5_) );
NOR2X1 NOR2X1_761 ( .gnd(gnd), .vdd(vdd), .A(data_39__6_), .B(_7401_), .Y(_7412_) );
AOI21X1 AOI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf3), .B(_7401_), .C(_7412_), .Y(_189__6_) );
INVX1 INVX1_3238 ( .gnd(gnd), .vdd(vdd), .A(data_39__7_), .Y(_7413_) );
OAI21X1 OAI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7413_), .Y(_7414_) );
NAND3X1 NAND3X1_969 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf10), .B(_7116_), .C(_7396_), .Y(_7415_) );
AND2X2 AND2X2_1361 ( .gnd(gnd), .vdd(vdd), .A(_7415_), .B(_7414_), .Y(_189__7_) );
NOR2X1 NOR2X1_762 ( .gnd(gnd), .vdd(vdd), .A(data_39__8_), .B(_7401_), .Y(_7416_) );
AOI21X1 AOI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf6), .B(_7401_), .C(_7416_), .Y(_189__8_) );
NOR2X1 NOR2X1_763 ( .gnd(gnd), .vdd(vdd), .A(data_39__9_), .B(_7401_), .Y(_7417_) );
AOI21X1 AOI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf1), .B(_7401_), .C(_7417_), .Y(_189__9_) );
NOR2X1 NOR2X1_764 ( .gnd(gnd), .vdd(vdd), .A(data_39__10_), .B(_7401_), .Y(_7418_) );
AOI21X1 AOI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_7401_), .C(_7418_), .Y(_189__10_) );
INVX1 INVX1_3239 ( .gnd(gnd), .vdd(vdd), .A(data_39__11_), .Y(_7419_) );
OAI21X1 OAI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7419_), .Y(_7420_) );
NAND3X1 NAND3X1_970 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_7116_), .C(_7396_), .Y(_7421_) );
AND2X2 AND2X2_1362 ( .gnd(gnd), .vdd(vdd), .A(_7421_), .B(_7420_), .Y(_189__11_) );
INVX1 INVX1_3240 ( .gnd(gnd), .vdd(vdd), .A(data_39__12_), .Y(_7422_) );
OAI21X1 OAI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_7388_), .B(_7393_), .C(_7422_), .Y(_7423_) );
NAND3X1 NAND3X1_971 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_7116_), .C(_7396_), .Y(_7424_) );
AND2X2 AND2X2_1363 ( .gnd(gnd), .vdd(vdd), .A(_7424_), .B(_7423_), .Y(_189__12_) );
NOR2X1 NOR2X1_765 ( .gnd(gnd), .vdd(vdd), .A(data_39__13_), .B(_7401_), .Y(_7425_) );
AOI21X1 AOI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf6), .B(_7401_), .C(_7425_), .Y(_189__13_) );
NOR2X1 NOR2X1_766 ( .gnd(gnd), .vdd(vdd), .A(data_39__14_), .B(_7401_), .Y(_7426_) );
AOI21X1 AOI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_7401_), .C(_7426_), .Y(_189__14_) );
NOR2X1 NOR2X1_767 ( .gnd(gnd), .vdd(vdd), .A(data_39__15_), .B(_7401_), .Y(_7427_) );
AOI21X1 AOI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf9), .B(_7401_), .C(_7427_), .Y(_189__15_) );
OAI21X1 OAI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_7256_), .C(_3318_), .Y(_7428_) );
NOR2X1 NOR2X1_768 ( .gnd(gnd), .vdd(vdd), .A(_7428_), .B(_3386_), .Y(_7429_) );
NAND3X1 NAND3X1_972 ( .gnd(gnd), .vdd(vdd), .A(_3395__bF_buf1), .B(_7429_), .C(_3313__bF_buf55), .Y(_7430_) );
NOR2X1 NOR2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_7430_), .B(_7388_), .Y(_7431_) );
NOR2X1 NOR2X1_770 ( .gnd(gnd), .vdd(vdd), .A(data_38__0_), .B(_7431__bF_buf4), .Y(_7432_) );
AOI21X1 AOI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_7431__bF_buf3), .C(_7432_), .Y(_188__0_) );
NOR2X1 NOR2X1_771 ( .gnd(gnd), .vdd(vdd), .A(data_38__1_), .B(_7431__bF_buf2), .Y(_7433_) );
AOI21X1 AOI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_7431__bF_buf1), .C(_7433_), .Y(_188__1_) );
NOR2X1 NOR2X1_772 ( .gnd(gnd), .vdd(vdd), .A(data_38__2_), .B(_7431__bF_buf0), .Y(_7434_) );
AOI21X1 AOI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf14), .B(_7431__bF_buf4), .C(_7434_), .Y(_188__2_) );
NOR2X1 NOR2X1_773 ( .gnd(gnd), .vdd(vdd), .A(data_38__3_), .B(_7431__bF_buf3), .Y(_7435_) );
AOI21X1 AOI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_7431__bF_buf2), .C(_7435_), .Y(_188__3_) );
NOR2X1 NOR2X1_774 ( .gnd(gnd), .vdd(vdd), .A(data_38__4_), .B(_7431__bF_buf1), .Y(_7436_) );
AOI21X1 AOI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_7431__bF_buf0), .C(_7436_), .Y(_188__4_) );
NOR2X1 NOR2X1_775 ( .gnd(gnd), .vdd(vdd), .A(data_38__5_), .B(_7431__bF_buf4), .Y(_7437_) );
AOI21X1 AOI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf8), .B(_7431__bF_buf3), .C(_7437_), .Y(_188__5_) );
NOR2X1 NOR2X1_776 ( .gnd(gnd), .vdd(vdd), .A(data_38__6_), .B(_7431__bF_buf2), .Y(_7438_) );
AOI21X1 AOI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_7431__bF_buf1), .C(_7438_), .Y(_188__6_) );
NOR2X1 NOR2X1_777 ( .gnd(gnd), .vdd(vdd), .A(data_38__7_), .B(_7431__bF_buf0), .Y(_7439_) );
AOI21X1 AOI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_7431__bF_buf4), .C(_7439_), .Y(_188__7_) );
NOR2X1 NOR2X1_778 ( .gnd(gnd), .vdd(vdd), .A(data_38__8_), .B(_7431__bF_buf3), .Y(_7440_) );
AOI21X1 AOI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf5), .B(_7431__bF_buf2), .C(_7440_), .Y(_188__8_) );
NOR2X1 NOR2X1_779 ( .gnd(gnd), .vdd(vdd), .A(data_38__9_), .B(_7431__bF_buf1), .Y(_7441_) );
AOI21X1 AOI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_7431__bF_buf0), .C(_7441_), .Y(_188__9_) );
NOR2X1 NOR2X1_780 ( .gnd(gnd), .vdd(vdd), .A(data_38__10_), .B(_7431__bF_buf4), .Y(_7442_) );
AOI21X1 AOI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf6), .B(_7431__bF_buf3), .C(_7442_), .Y(_188__10_) );
NOR2X1 NOR2X1_781 ( .gnd(gnd), .vdd(vdd), .A(data_38__11_), .B(_7431__bF_buf2), .Y(_7443_) );
AOI21X1 AOI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_7431__bF_buf1), .C(_7443_), .Y(_188__11_) );
NOR2X1 NOR2X1_782 ( .gnd(gnd), .vdd(vdd), .A(data_38__12_), .B(_7431__bF_buf0), .Y(_7444_) );
AOI21X1 AOI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_7431__bF_buf4), .C(_7444_), .Y(_188__12_) );
NOR2X1 NOR2X1_783 ( .gnd(gnd), .vdd(vdd), .A(data_38__13_), .B(_7431__bF_buf3), .Y(_7445_) );
AOI21X1 AOI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_7431__bF_buf2), .C(_7445_), .Y(_188__13_) );
NOR2X1 NOR2X1_784 ( .gnd(gnd), .vdd(vdd), .A(data_38__14_), .B(_7431__bF_buf1), .Y(_7446_) );
AOI21X1 AOI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_7431__bF_buf0), .C(_7446_), .Y(_188__14_) );
NOR2X1 NOR2X1_785 ( .gnd(gnd), .vdd(vdd), .A(data_38__15_), .B(_7431__bF_buf4), .Y(_7447_) );
AOI21X1 AOI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_7431__bF_buf3), .C(_7447_), .Y(_188__15_) );
NOR2X1 NOR2X1_786 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf9), .B(_7387_), .Y(_7448_) );
NOR2X1 NOR2X1_787 ( .gnd(gnd), .vdd(vdd), .A(data_37__0_), .B(_7448__bF_buf3), .Y(_7449_) );
AOI21X1 AOI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_7448__bF_buf2), .C(_7449_), .Y(_187__0_) );
INVX1 INVX1_3241 ( .gnd(gnd), .vdd(vdd), .A(data_37__1_), .Y(_7450_) );
OAI21X1 OAI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_14882__bF_buf8), .C(_7450_), .Y(_7451_) );
NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_7448__bF_buf1), .Y(_7452_) );
AND2X2 AND2X2_1364 ( .gnd(gnd), .vdd(vdd), .A(_7452_), .B(_7451_), .Y(_187__1_) );
NOR2X1 NOR2X1_788 ( .gnd(gnd), .vdd(vdd), .A(data_37__2_), .B(_7448__bF_buf0), .Y(_7453_) );
AOI21X1 AOI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf13), .B(_7448__bF_buf3), .C(_7453_), .Y(_187__2_) );
NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_7115_), .Y(_7454_) );
INVX1 INVX1_3242 ( .gnd(gnd), .vdd(vdd), .A(data_37__3_), .Y(_7455_) );
OAI21X1 OAI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_14882__bF_buf7), .C(_7455_), .Y(_7456_) );
OAI21X1 OAI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_7454_), .B(IDATA_PROG_data_3_bF_buf2), .C(_7456_), .Y(_7457_) );
INVX1 INVX1_3243 ( .gnd(gnd), .vdd(vdd), .A(_7457_), .Y(_187__3_) );
INVX1 INVX1_3244 ( .gnd(gnd), .vdd(vdd), .A(data_37__4_), .Y(_7458_) );
OAI21X1 OAI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_14882__bF_buf6), .C(_7458_), .Y(_7459_) );
OAI21X1 OAI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_7454_), .B(IDATA_PROG_data_4_bF_buf0), .C(_7459_), .Y(_7460_) );
INVX1 INVX1_3245 ( .gnd(gnd), .vdd(vdd), .A(_7460_), .Y(_187__4_) );
INVX1 INVX1_3246 ( .gnd(gnd), .vdd(vdd), .A(data_37__5_), .Y(_7461_) );
OAI21X1 OAI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_14882__bF_buf5), .C(_7461_), .Y(_7462_) );
OAI21X1 OAI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_7454_), .B(IDATA_PROG_data_5_bF_buf3), .C(_7462_), .Y(_7463_) );
INVX1 INVX1_3247 ( .gnd(gnd), .vdd(vdd), .A(_7463_), .Y(_187__5_) );
NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_7448__bF_buf2), .Y(_7464_) );
OAI21X1 OAI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(data_37__6_), .B(_7448__bF_buf1), .C(_7464_), .Y(_7465_) );
INVX1 INVX1_3248 ( .gnd(gnd), .vdd(vdd), .A(_7465_), .Y(_187__6_) );
INVX1 INVX1_3249 ( .gnd(gnd), .vdd(vdd), .A(data_37__7_), .Y(_7466_) );
OAI21X1 OAI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_7387_), .B(_14882__bF_buf4), .C(_7466_), .Y(_7467_) );
OAI21X1 OAI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_7454_), .B(IDATA_PROG_data_7_bF_buf3), .C(_7467_), .Y(_7468_) );
INVX1 INVX1_3250 ( .gnd(gnd), .vdd(vdd), .A(_7468_), .Y(_187__7_) );
NOR2X1 NOR2X1_789 ( .gnd(gnd), .vdd(vdd), .A(data_37__8_), .B(_7448__bF_buf0), .Y(_7469_) );
NOR2X1 NOR2X1_790 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf1), .B(_7454_), .Y(_7470_) );
NOR2X1 NOR2X1_791 ( .gnd(gnd), .vdd(vdd), .A(_7469_), .B(_7470_), .Y(_187__8_) );
NOR2X1 NOR2X1_792 ( .gnd(gnd), .vdd(vdd), .A(data_37__9_), .B(_7448__bF_buf3), .Y(_7471_) );
AOI21X1 AOI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf14), .B(_7448__bF_buf2), .C(_7471_), .Y(_187__9_) );
NOR2X1 NOR2X1_793 ( .gnd(gnd), .vdd(vdd), .A(data_37__10_), .B(_7448__bF_buf1), .Y(_7472_) );
NOR2X1 NOR2X1_794 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf0), .B(_7454_), .Y(_7473_) );
NOR2X1 NOR2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_7472_), .B(_7473_), .Y(_187__10_) );
NOR2X1 NOR2X1_796 ( .gnd(gnd), .vdd(vdd), .A(data_37__11_), .B(_7448__bF_buf0), .Y(_7474_) );
NOR2X1 NOR2X1_797 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf3), .B(_7454_), .Y(_7475_) );
NOR2X1 NOR2X1_798 ( .gnd(gnd), .vdd(vdd), .A(_7474_), .B(_7475_), .Y(_187__11_) );
NOR2X1 NOR2X1_799 ( .gnd(gnd), .vdd(vdd), .A(data_37__12_), .B(_7448__bF_buf3), .Y(_7476_) );
NOR2X1 NOR2X1_800 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf3), .B(_7454_), .Y(_7477_) );
NOR2X1 NOR2X1_801 ( .gnd(gnd), .vdd(vdd), .A(_7476_), .B(_7477_), .Y(_187__12_) );
NOR2X1 NOR2X1_802 ( .gnd(gnd), .vdd(vdd), .A(data_37__13_), .B(_7448__bF_buf2), .Y(_7478_) );
NOR2X1 NOR2X1_803 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf1), .B(_7454_), .Y(_7479_) );
NOR2X1 NOR2X1_804 ( .gnd(gnd), .vdd(vdd), .A(_7478_), .B(_7479_), .Y(_187__13_) );
NOR2X1 NOR2X1_805 ( .gnd(gnd), .vdd(vdd), .A(data_37__14_), .B(_7448__bF_buf1), .Y(_7480_) );
AOI21X1 AOI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_7448__bF_buf0), .C(_7480_), .Y(_187__14_) );
NOR2X1 NOR2X1_806 ( .gnd(gnd), .vdd(vdd), .A(data_37__15_), .B(_7448__bF_buf3), .Y(_7481_) );
NOR2X1 NOR2X1_807 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf4), .B(_7454_), .Y(_7482_) );
NOR2X1 NOR2X1_808 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .B(_7482_), .Y(_187__15_) );
INVX1 INVX1_3251 ( .gnd(gnd), .vdd(vdd), .A(data_36__0_), .Y(_7483_) );
NAND3X1 NAND3X1_973 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf0), .B(_14946__bF_buf2), .C(_16157_), .Y(_7484_) );
MUX2X1 MUX2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_7483_), .B(_14932__bF_buf2), .S(_7484_), .Y(_186__0_) );
INVX1 INVX1_3252 ( .gnd(gnd), .vdd(vdd), .A(data_36__1_), .Y(_7485_) );
MUX2X1 MUX2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_7485_), .B(_14894__bF_buf1), .S(_7484_), .Y(_186__1_) );
INVX1 INVX1_3253 ( .gnd(gnd), .vdd(vdd), .A(data_36__2_), .Y(_7486_) );
MUX2X1 MUX2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_7486_), .B(_14897__bF_buf12), .S(_7484_), .Y(_186__2_) );
INVX1 INVX1_3254 ( .gnd(gnd), .vdd(vdd), .A(data_36__3_), .Y(_7487_) );
MUX2X1 MUX2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_7487_), .B(_14899__bF_buf2), .S(_7484_), .Y(_186__3_) );
INVX1 INVX1_3255 ( .gnd(gnd), .vdd(vdd), .A(data_36__4_), .Y(_7488_) );
MUX2X1 MUX2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_7488_), .B(_14902__bF_buf5), .S(_7484_), .Y(_186__4_) );
INVX1 INVX1_3256 ( .gnd(gnd), .vdd(vdd), .A(data_36__5_), .Y(_7489_) );
MUX2X1 MUX2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_7489_), .B(_14903__bF_buf7), .S(_7484_), .Y(_186__5_) );
INVX1 INVX1_3257 ( .gnd(gnd), .vdd(vdd), .A(data_36__6_), .Y(_7490_) );
OAI21X1 OAI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_14882__bF_buf3), .C(_7490_), .Y(_7491_) );
OAI21X1 OAI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf3), .B(_7484_), .C(_7491_), .Y(_7492_) );
INVX1 INVX1_3258 ( .gnd(gnd), .vdd(vdd), .A(_7492_), .Y(_186__6_) );
INVX1 INVX1_3259 ( .gnd(gnd), .vdd(vdd), .A(data_36__7_), .Y(_7493_) );
MUX2X1 MUX2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_7493_), .B(_14908__bF_buf8), .S(_7484_), .Y(_186__7_) );
INVX1 INVX1_3260 ( .gnd(gnd), .vdd(vdd), .A(data_36__8_), .Y(_7494_) );
OAI21X1 OAI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_14882__bF_buf2), .C(_7494_), .Y(_7495_) );
OAI21X1 OAI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf0), .B(_7484_), .C(_7495_), .Y(_7496_) );
INVX1 INVX1_3261 ( .gnd(gnd), .vdd(vdd), .A(_7496_), .Y(_186__8_) );
INVX1 INVX1_3262 ( .gnd(gnd), .vdd(vdd), .A(data_36__9_), .Y(_7497_) );
MUX2X1 MUX2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_7497_), .B(_14913__bF_buf13), .S(_7484_), .Y(_186__9_) );
INVX1 INVX1_3263 ( .gnd(gnd), .vdd(vdd), .A(data_36__10_), .Y(_7498_) );
MUX2X1 MUX2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_7498_), .B(_15055__bF_buf5), .S(_7484_), .Y(_186__10_) );
INVX1 INVX1_3264 ( .gnd(gnd), .vdd(vdd), .A(data_36__11_), .Y(_7499_) );
MUX2X1 MUX2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_7499_), .B(_14918__bF_buf7), .S(_7484_), .Y(_186__11_) );
INVX1 INVX1_3265 ( .gnd(gnd), .vdd(vdd), .A(data_36__12_), .Y(_7500_) );
MUX2X1 MUX2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_7500_), .B(_14920__bF_buf7), .S(_7484_), .Y(_186__12_) );
INVX1 INVX1_3266 ( .gnd(gnd), .vdd(vdd), .A(data_36__13_), .Y(_7501_) );
MUX2X1 MUX2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_7501_), .B(_14924__bF_buf4), .S(_7484_), .Y(_186__13_) );
INVX1 INVX1_3267 ( .gnd(gnd), .vdd(vdd), .A(data_36__14_), .Y(_7502_) );
MUX2X1 MUX2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_7502_), .B(_15060__bF_buf0), .S(_7484_), .Y(_186__14_) );
INVX1 INVX1_3268 ( .gnd(gnd), .vdd(vdd), .A(data_36__15_), .Y(_7503_) );
OAI21X1 OAI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_14882__bF_buf1), .C(_7503_), .Y(_7504_) );
OAI21X1 OAI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf3), .B(_7484_), .C(_7504_), .Y(_7505_) );
INVX1 INVX1_3269 ( .gnd(gnd), .vdd(vdd), .A(_7505_), .Y(_186__15_) );
INVX1 INVX1_3270 ( .gnd(gnd), .vdd(vdd), .A(data_35__0_), .Y(_7506_) );
NOR2X1 NOR2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_15580_), .B(_15572_), .Y(_7507_) );
NOR2X1 NOR2X1_810 ( .gnd(gnd), .vdd(vdd), .A(_14998__bF_buf3), .B(_6483_), .Y(_7508_) );
OAI21X1 OAI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_14942__bF_buf0), .B(_15175__bF_buf1), .C(_7508_), .Y(_7509_) );
INVX1 INVX1_3271 ( .gnd(gnd), .vdd(vdd), .A(_7509_), .Y(_7510_) );
OAI21X1 OAI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf2), .B(_7507_), .C(_7510_), .Y(_7511_) );
NOR2X1 NOR2X1_811 ( .gnd(gnd), .vdd(vdd), .A(_7511_), .B(_5459__bF_buf0), .Y(_7512_) );
NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_3313__bF_buf54), .Y(_7513_) );
MUX2X1 MUX2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_7506_), .B(_14932__bF_buf1), .S(_7513_), .Y(_185__0_) );
INVX1 INVX1_3272 ( .gnd(gnd), .vdd(vdd), .A(data_35__1_), .Y(_7514_) );
MUX2X1 MUX2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_7514_), .B(_14894__bF_buf0), .S(_7513_), .Y(_185__1_) );
INVX1 INVX1_3273 ( .gnd(gnd), .vdd(vdd), .A(data_35__2_), .Y(_7515_) );
MUX2X1 MUX2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_7515_), .B(_14897__bF_buf11), .S(_7513_), .Y(_185__2_) );
INVX1 INVX1_3274 ( .gnd(gnd), .vdd(vdd), .A(data_35__3_), .Y(_7516_) );
MUX2X1 MUX2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_7516_), .B(_14899__bF_buf1), .S(_7513_), .Y(_185__3_) );
INVX1 INVX1_3275 ( .gnd(gnd), .vdd(vdd), .A(data_35__4_), .Y(_7517_) );
MUX2X1 MUX2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_7517_), .B(_14902__bF_buf4), .S(_7513_), .Y(_185__4_) );
INVX1 INVX1_3276 ( .gnd(gnd), .vdd(vdd), .A(data_35__5_), .Y(_7518_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .Y(_7519_) );
OAI21X1 OAI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_7519_), .C(_7518_), .Y(_7520_) );
NAND3X1 NAND3X1_974 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_7512_), .C(_3313__bF_buf53), .Y(_7521_) );
AND2X2 AND2X2_1365 ( .gnd(gnd), .vdd(vdd), .A(_7520_), .B(_7521_), .Y(_185__5_) );
INVX1 INVX1_3277 ( .gnd(gnd), .vdd(vdd), .A(data_35__6_), .Y(_7522_) );
MUX2X1 MUX2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_7522_), .B(_15049__bF_buf0), .S(_7513_), .Y(_185__6_) );
INVX1 INVX1_3278 ( .gnd(gnd), .vdd(vdd), .A(data_35__7_), .Y(_7523_) );
OAI21X1 OAI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_7519_), .C(_7523_), .Y(_7524_) );
NAND3X1 NAND3X1_975 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_7512_), .C(_3313__bF_buf52), .Y(_7525_) );
AND2X2 AND2X2_1366 ( .gnd(gnd), .vdd(vdd), .A(_7524_), .B(_7525_), .Y(_185__7_) );
INVX1 INVX1_3279 ( .gnd(gnd), .vdd(vdd), .A(data_35__8_), .Y(_7526_) );
MUX2X1 MUX2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_7526_), .B(_15052__bF_buf4), .S(_7513_), .Y(_185__8_) );
NOR2X1 NOR2X1_812 ( .gnd(gnd), .vdd(vdd), .A(_7519_), .B(_3393__bF_buf47), .Y(_7527_) );
AOI21X1 AOI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_3313__bF_buf51), .C(data_35__9_), .Y(_7528_) );
AOI21X1 AOI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_7527_), .C(_7528_), .Y(_185__9_) );
AOI21X1 AOI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_3313__bF_buf50), .C(data_35__10_), .Y(_7529_) );
AOI21X1 AOI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_7527_), .C(_7529_), .Y(_185__10_) );
INVX1 INVX1_3280 ( .gnd(gnd), .vdd(vdd), .A(data_35__11_), .Y(_7530_) );
MUX2X1 MUX2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_7530_), .B(_14918__bF_buf6), .S(_7513_), .Y(_185__11_) );
INVX1 INVX1_3281 ( .gnd(gnd), .vdd(vdd), .A(data_35__12_), .Y(_7531_) );
OAI21X1 OAI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_7519_), .C(_7531_), .Y(_7532_) );
NAND3X1 NAND3X1_976 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_7512_), .C(_3313__bF_buf49), .Y(_7533_) );
AND2X2 AND2X2_1367 ( .gnd(gnd), .vdd(vdd), .A(_7532_), .B(_7533_), .Y(_185__12_) );
AOI21X1 AOI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_7512_), .B(_3313__bF_buf48), .C(data_35__13_), .Y(_7534_) );
AOI21X1 AOI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_7527_), .C(_7534_), .Y(_185__13_) );
INVX1 INVX1_3282 ( .gnd(gnd), .vdd(vdd), .A(data_35__14_), .Y(_7535_) );
MUX2X1 MUX2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_7535_), .B(_15060__bF_buf14), .S(_7513_), .Y(_185__14_) );
INVX1 INVX1_3283 ( .gnd(gnd), .vdd(vdd), .A(data_35__15_), .Y(_7536_) );
MUX2X1 MUX2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_7536_), .B(_15062__bF_buf7), .S(_7513_), .Y(_185__15_) );
INVX1 INVX1_3284 ( .gnd(gnd), .vdd(vdd), .A(data_34__0_), .Y(_7537_) );
NOR2X1 NOR2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf1), .B(_15572_), .Y(_7538_) );
NOR2X1 NOR2X1_814 ( .gnd(gnd), .vdd(vdd), .A(_7509_), .B(_5459__bF_buf3), .Y(_7539_) );
OAI21X1 OAI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf1), .B(_7538_), .C(_7539_), .Y(_7540_) );
OAI21X1 OAI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_7540_), .C(_7537_), .Y(_7541_) );
INVX4 INVX4_35 ( .gnd(gnd), .vdd(vdd), .A(_7540_), .Y(_7542_) );
NAND3X1 NAND3X1_977 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_7542_), .C(_3313__bF_buf47), .Y(_7543_) );
AND2X2 AND2X2_1368 ( .gnd(gnd), .vdd(vdd), .A(_7541_), .B(_7543_), .Y(_184__0_) );
INVX1 INVX1_3285 ( .gnd(gnd), .vdd(vdd), .A(data_34__1_), .Y(_7544_) );
OAI21X1 OAI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_7540_), .C(_7544_), .Y(_7545_) );
NAND3X1 NAND3X1_978 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_7542_), .C(_3313__bF_buf46), .Y(_7546_) );
AND2X2 AND2X2_1369 ( .gnd(gnd), .vdd(vdd), .A(_7545_), .B(_7546_), .Y(_184__1_) );
INVX1 INVX1_3286 ( .gnd(gnd), .vdd(vdd), .A(data_34__2_), .Y(_7547_) );
NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_7542_), .B(_3313__bF_buf45), .Y(_7548_) );
MUX2X1 MUX2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_7547_), .B(_14897__bF_buf10), .S(_7548_), .Y(_184__2_) );
INVX1 INVX1_3287 ( .gnd(gnd), .vdd(vdd), .A(data_34__3_), .Y(_7549_) );
OAI21X1 OAI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_7540_), .C(_7549_), .Y(_7550_) );
NAND3X1 NAND3X1_979 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_7542_), .C(_3313__bF_buf44), .Y(_7551_) );
AND2X2 AND2X2_1370 ( .gnd(gnd), .vdd(vdd), .A(_7550_), .B(_7551_), .Y(_184__3_) );
INVX1 INVX1_3288 ( .gnd(gnd), .vdd(vdd), .A(data_34__4_), .Y(_7552_) );
OAI21X1 OAI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_7540_), .C(_7552_), .Y(_7553_) );
NAND3X1 NAND3X1_980 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_7542_), .C(_3313__bF_buf43), .Y(_7554_) );
AND2X2 AND2X2_1371 ( .gnd(gnd), .vdd(vdd), .A(_7553_), .B(_7554_), .Y(_184__4_) );
INVX1 INVX1_3289 ( .gnd(gnd), .vdd(vdd), .A(data_34__5_), .Y(_7555_) );
OAI21X1 OAI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_7540_), .C(_7555_), .Y(_7556_) );
NAND3X1 NAND3X1_981 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_7542_), .C(_3313__bF_buf42), .Y(_7557_) );
AND2X2 AND2X2_1372 ( .gnd(gnd), .vdd(vdd), .A(_7556_), .B(_7557_), .Y(_184__5_) );
INVX1 INVX1_3290 ( .gnd(gnd), .vdd(vdd), .A(data_34__6_), .Y(_7558_) );
MUX2X1 MUX2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_7558_), .B(_15049__bF_buf14), .S(_7548_), .Y(_184__6_) );
INVX1 INVX1_3291 ( .gnd(gnd), .vdd(vdd), .A(data_34__7_), .Y(_7559_) );
OAI21X1 OAI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_7540_), .C(_7559_), .Y(_7560_) );
NAND3X1 NAND3X1_982 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_7542_), .C(_3313__bF_buf41), .Y(_7561_) );
AND2X2 AND2X2_1373 ( .gnd(gnd), .vdd(vdd), .A(_7560_), .B(_7561_), .Y(_184__7_) );
INVX1 INVX1_3292 ( .gnd(gnd), .vdd(vdd), .A(data_34__8_), .Y(_7562_) );
MUX2X1 MUX2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_7562_), .B(_15052__bF_buf3), .S(_7548_), .Y(_184__8_) );
INVX1 INVX1_3293 ( .gnd(gnd), .vdd(vdd), .A(data_34__9_), .Y(_7563_) );
MUX2X1 MUX2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_7563_), .B(_14913__bF_buf11), .S(_7548_), .Y(_184__9_) );
INVX1 INVX1_3294 ( .gnd(gnd), .vdd(vdd), .A(data_34__10_), .Y(_7564_) );
MUX2X1 MUX2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_7564_), .B(_15055__bF_buf3), .S(_7548_), .Y(_184__10_) );
INVX1 INVX1_3295 ( .gnd(gnd), .vdd(vdd), .A(data_34__11_), .Y(_7565_) );
OAI21X1 OAI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_7540_), .C(_7565_), .Y(_7566_) );
NAND3X1 NAND3X1_983 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_7542_), .C(_3313__bF_buf40), .Y(_7567_) );
AND2X2 AND2X2_1374 ( .gnd(gnd), .vdd(vdd), .A(_7566_), .B(_7567_), .Y(_184__11_) );
INVX1 INVX1_3296 ( .gnd(gnd), .vdd(vdd), .A(data_34__12_), .Y(_7568_) );
OAI21X1 OAI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_7540_), .C(_7568_), .Y(_7569_) );
NAND3X1 NAND3X1_984 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_7542_), .C(_3313__bF_buf39), .Y(_7570_) );
AND2X2 AND2X2_1375 ( .gnd(gnd), .vdd(vdd), .A(_7569_), .B(_7570_), .Y(_184__12_) );
INVX1 INVX1_3297 ( .gnd(gnd), .vdd(vdd), .A(data_34__13_), .Y(_7571_) );
MUX2X1 MUX2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_7571_), .B(_14924__bF_buf2), .S(_7548_), .Y(_184__13_) );
INVX1 INVX1_3298 ( .gnd(gnd), .vdd(vdd), .A(data_34__14_), .Y(_7572_) );
MUX2X1 MUX2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_7572_), .B(_15060__bF_buf13), .S(_7548_), .Y(_184__14_) );
INVX1 INVX1_3299 ( .gnd(gnd), .vdd(vdd), .A(data_34__15_), .Y(_7573_) );
MUX2X1 MUX2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_7573_), .B(_15062__bF_buf6), .S(_7548_), .Y(_184__15_) );
INVX1 INVX1_3300 ( .gnd(gnd), .vdd(vdd), .A(data_33__0_), .Y(_7574_) );
NOR2X1 NOR2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_14978__bF_buf0), .B(_15684_), .Y(_7575_) );
OAI21X1 OAI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_15170__bF_buf0), .B(_7575_), .C(_7539_), .Y(_7576_) );
OAI21X1 OAI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_7576_), .C(_7574_), .Y(_7577_) );
INVX4 INVX4_36 ( .gnd(gnd), .vdd(vdd), .A(_7576_), .Y(_7578_) );
NAND3X1 NAND3X1_985 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf14), .B(_7578_), .C(_3313__bF_buf38), .Y(_7579_) );
AND2X2 AND2X2_1376 ( .gnd(gnd), .vdd(vdd), .A(_7577_), .B(_7579_), .Y(_183__0_) );
INVX1 INVX1_3301 ( .gnd(gnd), .vdd(vdd), .A(data_33__1_), .Y(_7580_) );
OAI21X1 OAI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_7576_), .C(_7580_), .Y(_7581_) );
NAND3X1 NAND3X1_986 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf13), .B(_7578_), .C(_3313__bF_buf37), .Y(_7582_) );
AND2X2 AND2X2_1377 ( .gnd(gnd), .vdd(vdd), .A(_7581_), .B(_7582_), .Y(_183__1_) );
INVX1 INVX1_3302 ( .gnd(gnd), .vdd(vdd), .A(data_33__2_), .Y(_7583_) );
NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_7578_), .B(_3313__bF_buf36), .Y(_7584_) );
MUX2X1 MUX2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_7583_), .B(_14897__bF_buf9), .S(_7584_), .Y(_183__2_) );
INVX1 INVX1_3303 ( .gnd(gnd), .vdd(vdd), .A(data_33__3_), .Y(_7585_) );
OAI21X1 OAI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_7576_), .C(_7585_), .Y(_7586_) );
NAND3X1 NAND3X1_987 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_7578_), .C(_3313__bF_buf35), .Y(_7587_) );
AND2X2 AND2X2_1378 ( .gnd(gnd), .vdd(vdd), .A(_7586_), .B(_7587_), .Y(_183__3_) );
INVX1 INVX1_3304 ( .gnd(gnd), .vdd(vdd), .A(data_33__4_), .Y(_7588_) );
OAI21X1 OAI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf34), .B(_7576_), .C(_7588_), .Y(_7589_) );
NAND3X1 NAND3X1_988 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf2), .B(_7578_), .C(_3313__bF_buf34), .Y(_7590_) );
AND2X2 AND2X2_1379 ( .gnd(gnd), .vdd(vdd), .A(_7589_), .B(_7590_), .Y(_183__4_) );
INVX1 INVX1_3305 ( .gnd(gnd), .vdd(vdd), .A(data_33__5_), .Y(_7591_) );
OAI21X1 OAI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf33), .B(_7576_), .C(_7591_), .Y(_7592_) );
NAND3X1 NAND3X1_989 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_7578_), .C(_3313__bF_buf33), .Y(_7593_) );
AND2X2 AND2X2_1380 ( .gnd(gnd), .vdd(vdd), .A(_7592_), .B(_7593_), .Y(_183__5_) );
INVX1 INVX1_3306 ( .gnd(gnd), .vdd(vdd), .A(data_33__6_), .Y(_7594_) );
MUX2X1 MUX2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_7594_), .B(_15049__bF_buf13), .S(_7584_), .Y(_183__6_) );
INVX1 INVX1_3307 ( .gnd(gnd), .vdd(vdd), .A(data_33__7_), .Y(_7595_) );
OAI21X1 OAI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf32), .B(_7576_), .C(_7595_), .Y(_7596_) );
NAND3X1 NAND3X1_990 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_7578_), .C(_3313__bF_buf32), .Y(_7597_) );
AND2X2 AND2X2_1381 ( .gnd(gnd), .vdd(vdd), .A(_7596_), .B(_7597_), .Y(_183__7_) );
INVX1 INVX1_3308 ( .gnd(gnd), .vdd(vdd), .A(data_33__8_), .Y(_7598_) );
MUX2X1 MUX2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_7598_), .B(_15052__bF_buf2), .S(_7584_), .Y(_183__8_) );
INVX1 INVX1_3309 ( .gnd(gnd), .vdd(vdd), .A(data_33__9_), .Y(_7599_) );
MUX2X1 MUX2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_7599_), .B(_14913__bF_buf10), .S(_7584_), .Y(_183__9_) );
INVX1 INVX1_3310 ( .gnd(gnd), .vdd(vdd), .A(data_33__10_), .Y(_7600_) );
MUX2X1 MUX2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_7600_), .B(_15055__bF_buf2), .S(_7584_), .Y(_183__10_) );
INVX1 INVX1_3311 ( .gnd(gnd), .vdd(vdd), .A(data_33__11_), .Y(_7601_) );
OAI21X1 OAI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf31), .B(_7576_), .C(_7601_), .Y(_7602_) );
NAND3X1 NAND3X1_991 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_7578_), .C(_3313__bF_buf31), .Y(_7603_) );
AND2X2 AND2X2_1382 ( .gnd(gnd), .vdd(vdd), .A(_7602_), .B(_7603_), .Y(_183__11_) );
INVX1 INVX1_3312 ( .gnd(gnd), .vdd(vdd), .A(data_33__12_), .Y(_7604_) );
OAI21X1 OAI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf30), .B(_7576_), .C(_7604_), .Y(_7605_) );
NAND3X1 NAND3X1_992 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_7578_), .C(_3313__bF_buf30), .Y(_7606_) );
AND2X2 AND2X2_1383 ( .gnd(gnd), .vdd(vdd), .A(_7605_), .B(_7606_), .Y(_183__12_) );
INVX1 INVX1_3313 ( .gnd(gnd), .vdd(vdd), .A(data_33__13_), .Y(_7607_) );
MUX2X1 MUX2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_7607_), .B(_14924__bF_buf1), .S(_7584_), .Y(_183__13_) );
INVX1 INVX1_3314 ( .gnd(gnd), .vdd(vdd), .A(data_33__14_), .Y(_7608_) );
MUX2X1 MUX2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_7608_), .B(_15060__bF_buf12), .S(_7584_), .Y(_183__14_) );
INVX1 INVX1_3315 ( .gnd(gnd), .vdd(vdd), .A(data_33__15_), .Y(_7609_) );
MUX2X1 MUX2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_7609_), .B(_15062__bF_buf5), .S(_7584_), .Y(_183__15_) );
NAND3X1 NAND3X1_993 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf8), .B(_14986_), .C(_14946__bF_buf1), .Y(_7610_) );
INVX1 INVX1_3316 ( .gnd(gnd), .vdd(vdd), .A(data_32__0_), .Y(_7611_) );
NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_14986_), .B(_14946__bF_buf0), .Y(_7612_) );
OAI21X1 OAI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf0), .C(_7611_), .Y(_7613_) );
OAI21X1 OAI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf1), .B(_7610_), .C(_7613_), .Y(_7614_) );
INVX1 INVX1_3317 ( .gnd(gnd), .vdd(vdd), .A(_7614_), .Y(_182__0_) );
INVX1 INVX1_3318 ( .gnd(gnd), .vdd(vdd), .A(data_32__1_), .Y(_7615_) );
OAI21X1 OAI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf15_bF_buf1), .C(_7615_), .Y(_7616_) );
OAI21X1 OAI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf2), .B(_7610_), .C(_7616_), .Y(_7617_) );
INVX1 INVX1_3319 ( .gnd(gnd), .vdd(vdd), .A(_7617_), .Y(_182__1_) );
INVX1 INVX1_3320 ( .gnd(gnd), .vdd(vdd), .A(data_32__2_), .Y(_7618_) );
MUX2X1 MUX2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_7618_), .B(_14897__bF_buf8), .S(_7610_), .Y(_182__2_) );
INVX1 INVX1_3321 ( .gnd(gnd), .vdd(vdd), .A(data_32__3_), .Y(_7619_) );
OAI21X1 OAI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf14_bF_buf1), .C(_7619_), .Y(_7620_) );
OAI21X1 OAI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_3_bF_buf1), .B(_7610_), .C(_7620_), .Y(_7621_) );
INVX1 INVX1_3322 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .Y(_182__3_) );
INVX1 INVX1_3323 ( .gnd(gnd), .vdd(vdd), .A(data_32__4_), .Y(_7622_) );
OAI21X1 OAI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf13_bF_buf1), .C(_7622_), .Y(_7623_) );
OAI21X1 OAI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf4), .B(_7610_), .C(_7623_), .Y(_7624_) );
INVX1 INVX1_3324 ( .gnd(gnd), .vdd(vdd), .A(_7624_), .Y(_182__4_) );
INVX1 INVX1_3325 ( .gnd(gnd), .vdd(vdd), .A(data_32__5_), .Y(_7625_) );
MUX2X1 MUX2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_7625_), .B(_14903__bF_buf3), .S(_7610_), .Y(_182__5_) );
INVX1 INVX1_3326 ( .gnd(gnd), .vdd(vdd), .A(data_32__6_), .Y(_7626_) );
OAI21X1 OAI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf12), .C(_7626_), .Y(_7627_) );
OAI21X1 OAI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf2), .B(_7610_), .C(_7627_), .Y(_7628_) );
INVX1 INVX1_3327 ( .gnd(gnd), .vdd(vdd), .A(_7628_), .Y(_182__6_) );
INVX1 INVX1_3328 ( .gnd(gnd), .vdd(vdd), .A(data_32__7_), .Y(_7629_) );
OAI21X1 OAI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf11), .C(_7629_), .Y(_7630_) );
OAI21X1 OAI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf2), .B(_7610_), .C(_7630_), .Y(_7631_) );
INVX1 INVX1_3329 ( .gnd(gnd), .vdd(vdd), .A(_7631_), .Y(_182__7_) );
INVX1 INVX1_3330 ( .gnd(gnd), .vdd(vdd), .A(data_32__8_), .Y(_7632_) );
OAI21X1 OAI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf10), .C(_7632_), .Y(_7633_) );
OAI21X1 OAI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf4), .B(_7610_), .C(_7633_), .Y(_7634_) );
INVX1 INVX1_3331 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .Y(_182__8_) );
INVX1 INVX1_3332 ( .gnd(gnd), .vdd(vdd), .A(data_32__9_), .Y(_7635_) );
OAI21X1 OAI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf9), .C(_7635_), .Y(_7636_) );
OAI21X1 OAI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf0), .B(_7610_), .C(_7636_), .Y(_7637_) );
INVX1 INVX1_3333 ( .gnd(gnd), .vdd(vdd), .A(_7637_), .Y(_182__9_) );
INVX1 INVX1_3334 ( .gnd(gnd), .vdd(vdd), .A(data_32__10_), .Y(_7638_) );
OAI21X1 OAI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf8), .C(_7638_), .Y(_7639_) );
OAI21X1 OAI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf4), .B(_7610_), .C(_7639_), .Y(_7640_) );
INVX1 INVX1_3335 ( .gnd(gnd), .vdd(vdd), .A(_7640_), .Y(_182__10_) );
INVX1 INVX1_3336 ( .gnd(gnd), .vdd(vdd), .A(data_32__11_), .Y(_7641_) );
OAI21X1 OAI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf7), .C(_7641_), .Y(_7642_) );
OAI21X1 OAI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf2), .B(_7610_), .C(_7642_), .Y(_7643_) );
INVX1 INVX1_3337 ( .gnd(gnd), .vdd(vdd), .A(_7643_), .Y(_182__11_) );
INVX1 INVX1_3338 ( .gnd(gnd), .vdd(vdd), .A(data_32__12_), .Y(_7644_) );
OAI21X1 OAI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf6), .C(_7644_), .Y(_7645_) );
OAI21X1 OAI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf2), .B(_7610_), .C(_7645_), .Y(_7646_) );
INVX1 INVX1_3339 ( .gnd(gnd), .vdd(vdd), .A(_7646_), .Y(_182__12_) );
INVX1 INVX1_3340 ( .gnd(gnd), .vdd(vdd), .A(data_32__13_), .Y(_7647_) );
OAI21X1 OAI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf5), .C(_7647_), .Y(_7648_) );
OAI21X1 OAI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf0), .B(_7610_), .C(_7648_), .Y(_7649_) );
INVX1 INVX1_3341 ( .gnd(gnd), .vdd(vdd), .A(_7649_), .Y(_182__13_) );
MUX2X1 MUX2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(data_32__14_), .B(IDATA_PROG_data_14_bF_buf3), .S(_7610_), .Y(_7650_) );
INVX1 INVX1_3342 ( .gnd(gnd), .vdd(vdd), .A(_7650_), .Y(_182__14_) );
INVX1 INVX1_3343 ( .gnd(gnd), .vdd(vdd), .A(data_32__15_), .Y(_7651_) );
OAI21X1 OAI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_7612_), .B(_14882__bF_buf4), .C(_7651_), .Y(_7652_) );
OAI21X1 OAI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf2), .B(_7610_), .C(_7652_), .Y(_7653_) );
INVX1 INVX1_3344 ( .gnd(gnd), .vdd(vdd), .A(_7653_), .Y(_182__15_) );
NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf0), .B(_14984__bF_buf0), .Y(_7654_) );
NOR2X1 NOR2X1_816 ( .gnd(gnd), .vdd(vdd), .A(_14882__bF_buf3), .B(_7654_), .Y(_7655_) );
NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf13), .B(_7655__bF_buf3), .Y(_7656_) );
OAI21X1 OAI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(data_31__0_), .B(_7655__bF_buf2), .C(_7656_), .Y(_7657_) );
INVX1 INVX1_3345 ( .gnd(gnd), .vdd(vdd), .A(_7657_), .Y(_181__0_) );
INVX1 INVX1_3346 ( .gnd(gnd), .vdd(vdd), .A(data_31__1_), .Y(_7658_) );
OAI21X1 OAI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf2), .C(_7658_), .Y(_7659_) );
NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_7655__bF_buf1), .Y(_7660_) );
AND2X2 AND2X2_1384 ( .gnd(gnd), .vdd(vdd), .A(_7660_), .B(_7659_), .Y(_181__1_) );
NOR2X1 NOR2X1_817 ( .gnd(gnd), .vdd(vdd), .A(_15177_), .B(_15175__bF_buf0), .Y(_7661_) );
NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf7), .B(_7661_), .Y(_7662_) );
INVX1 INVX1_3347 ( .gnd(gnd), .vdd(vdd), .A(data_31__2_), .Y(_7663_) );
OAI21X1 OAI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf1), .C(_7663_), .Y(_7664_) );
OAI21X1 OAI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(IDATA_PROG_data_2_bF_buf0), .C(_7664_), .Y(_7665_) );
INVX1 INVX1_3348 ( .gnd(gnd), .vdd(vdd), .A(_7665_), .Y(_181__2_) );
NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_7655__bF_buf0), .Y(_7666_) );
OAI21X1 OAI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(data_31__3_), .B(_7655__bF_buf3), .C(_7666_), .Y(_7667_) );
INVX1 INVX1_3349 ( .gnd(gnd), .vdd(vdd), .A(_7667_), .Y(_181__3_) );
INVX1 INVX1_3350 ( .gnd(gnd), .vdd(vdd), .A(data_31__4_), .Y(_7668_) );
OAI21X1 OAI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf0), .C(_7668_), .Y(_7669_) );
OAI21X1 OAI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(IDATA_PROG_data_4_bF_buf3), .C(_7669_), .Y(_7670_) );
INVX1 INVX1_3351 ( .gnd(gnd), .vdd(vdd), .A(_7670_), .Y(_181__4_) );
INVX1 INVX1_3352 ( .gnd(gnd), .vdd(vdd), .A(data_31__5_), .Y(_7671_) );
OAI21X1 OAI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf15_bF_buf0), .C(_7671_), .Y(_7672_) );
NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_7655__bF_buf2), .Y(_7673_) );
AND2X2 AND2X2_1385 ( .gnd(gnd), .vdd(vdd), .A(_7673_), .B(_7672_), .Y(_181__5_) );
NOR2X1 NOR2X1_818 ( .gnd(gnd), .vdd(vdd), .A(data_31__6_), .B(_7655__bF_buf1), .Y(_7674_) );
AOI21X1 AOI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf12), .B(_7655__bF_buf0), .C(_7674_), .Y(_181__6_) );
NOR2X1 NOR2X1_819 ( .gnd(gnd), .vdd(vdd), .A(data_31__7_), .B(_7655__bF_buf3), .Y(_7675_) );
AOI21X1 AOI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_7655__bF_buf2), .C(_7675_), .Y(_181__7_) );
INVX1 INVX1_3353 ( .gnd(gnd), .vdd(vdd), .A(data_31__8_), .Y(_7676_) );
OAI21X1 OAI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf14_bF_buf0), .C(_7676_), .Y(_7677_) );
NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_7655__bF_buf1), .Y(_7678_) );
AND2X2 AND2X2_1386 ( .gnd(gnd), .vdd(vdd), .A(_7678_), .B(_7677_), .Y(_181__8_) );
NOR2X1 NOR2X1_820 ( .gnd(gnd), .vdd(vdd), .A(data_31__9_), .B(_7655__bF_buf0), .Y(_7679_) );
AOI21X1 AOI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_7655__bF_buf3), .C(_7679_), .Y(_181__9_) );
INVX1 INVX1_3354 ( .gnd(gnd), .vdd(vdd), .A(data_31__10_), .Y(_7680_) );
OAI21X1 OAI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf13_bF_buf0), .C(_7680_), .Y(_7681_) );
NAND3X1 NAND3X1_994 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf6), .B(_15055__bF_buf1), .C(_7661_), .Y(_7682_) );
AND2X2 AND2X2_1387 ( .gnd(gnd), .vdd(vdd), .A(_7682_), .B(_7681_), .Y(_181__10_) );
INVX1 INVX1_3355 ( .gnd(gnd), .vdd(vdd), .A(data_31__11_), .Y(_7683_) );
OAI21X1 OAI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf12), .C(_7683_), .Y(_7684_) );
NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_7655__bF_buf2), .Y(_7685_) );
AND2X2 AND2X2_1388 ( .gnd(gnd), .vdd(vdd), .A(_7685_), .B(_7684_), .Y(_181__11_) );
NOR2X1 NOR2X1_821 ( .gnd(gnd), .vdd(vdd), .A(data_31__12_), .B(_7655__bF_buf1), .Y(_7686_) );
AOI21X1 AOI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_7655__bF_buf0), .C(_7686_), .Y(_181__12_) );
INVX1 INVX1_3356 ( .gnd(gnd), .vdd(vdd), .A(data_31__13_), .Y(_7687_) );
OAI21X1 OAI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_7654_), .B(_14882__bF_buf11), .C(_7687_), .Y(_7688_) );
OAI21X1 OAI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(IDATA_PROG_data_13_bF_buf4), .C(_7688_), .Y(_7689_) );
INVX1 INVX1_3357 ( .gnd(gnd), .vdd(vdd), .A(_7689_), .Y(_181__13_) );
OR2X2 OR2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_7655__bF_buf3), .B(data_31__14_), .Y(_7690_) );
OAI21X1 OAI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_7662_), .B(IDATA_PROG_data_14_bF_buf2), .C(_7690_), .Y(_7691_) );
INVX1 INVX1_3358 ( .gnd(gnd), .vdd(vdd), .A(_7691_), .Y(_181__14_) );
NOR2X1 NOR2X1_822 ( .gnd(gnd), .vdd(vdd), .A(data_31__15_), .B(_7655__bF_buf2), .Y(_7692_) );
AOI21X1 AOI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_7655__bF_buf1), .C(_7692_), .Y(_181__15_) );
NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf4), .B(_15793__bF_buf1), .Y(_7693_) );
INVX1 INVX1_3359 ( .gnd(gnd), .vdd(vdd), .A(data_30__0_), .Y(_7694_) );
OAI21X1 OAI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15175__bF_buf4), .C(_7694_), .Y(_7695_) );
OAI21X1 OAI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf0), .B(_7693_), .C(_7695_), .Y(_7696_) );
INVX1 INVX1_3360 ( .gnd(gnd), .vdd(vdd), .A(_7696_), .Y(_180__0_) );
INVX1 INVX1_3361 ( .gnd(gnd), .vdd(vdd), .A(data_30__1_), .Y(_7697_) );
OAI21X1 OAI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15175__bF_buf3), .C(_7697_), .Y(_7698_) );
NOR2X1 NOR2X1_823 ( .gnd(gnd), .vdd(vdd), .A(_15175__bF_buf2), .B(_15788__bF_buf5), .Y(_7699_) );
NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_7699_), .Y(_7700_) );
AND2X2 AND2X2_1389 ( .gnd(gnd), .vdd(vdd), .A(_7700_), .B(_7698_), .Y(_180__1_) );
NOR2X1 NOR2X1_824 ( .gnd(gnd), .vdd(vdd), .A(data_30__2_), .B(_7699_), .Y(_7701_) );
AOI21X1 AOI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_7699_), .C(_7701_), .Y(_180__2_) );
INVX1 INVX1_3362 ( .gnd(gnd), .vdd(vdd), .A(data_30__3_), .Y(_7702_) );
OAI21X1 OAI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15175__bF_buf1), .C(_7702_), .Y(_7703_) );
NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf12), .B(_7699_), .Y(_7704_) );
AND2X2 AND2X2_1390 ( .gnd(gnd), .vdd(vdd), .A(_7704_), .B(_7703_), .Y(_180__3_) );
INVX1 INVX1_3363 ( .gnd(gnd), .vdd(vdd), .A(data_30__4_), .Y(_7705_) );
OAI21X1 OAI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15175__bF_buf0), .C(_7705_), .Y(_7706_) );
OAI21X1 OAI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf2), .B(_7693_), .C(_7706_), .Y(_7707_) );
INVX1 INVX1_3364 ( .gnd(gnd), .vdd(vdd), .A(_7707_), .Y(_180__4_) );
INVX1 INVX1_3365 ( .gnd(gnd), .vdd(vdd), .A(data_30__5_), .Y(_7708_) );
OAI21X1 OAI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15175__bF_buf4), .C(_7708_), .Y(_7709_) );
NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_7699_), .Y(_7710_) );
AND2X2 AND2X2_1391 ( .gnd(gnd), .vdd(vdd), .A(_7710_), .B(_7709_), .Y(_180__5_) );
INVX1 INVX1_3366 ( .gnd(gnd), .vdd(vdd), .A(data_30__6_), .Y(_7711_) );
OAI21X1 OAI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15175__bF_buf3), .C(_7711_), .Y(_7712_) );
NAND3X1 NAND3X1_995 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_14984__bF_buf3), .C(_15793__bF_buf0), .Y(_7713_) );
AND2X2 AND2X2_1392 ( .gnd(gnd), .vdd(vdd), .A(_7712_), .B(_7713_), .Y(_180__6_) );
INVX1 INVX1_3367 ( .gnd(gnd), .vdd(vdd), .A(data_30__7_), .Y(_7714_) );
OAI21X1 OAI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15175__bF_buf2), .C(_7714_), .Y(_7715_) );
NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf3), .B(_7699_), .Y(_7716_) );
AND2X2 AND2X2_1393 ( .gnd(gnd), .vdd(vdd), .A(_7716_), .B(_7715_), .Y(_180__7_) );
INVX1 INVX1_3368 ( .gnd(gnd), .vdd(vdd), .A(data_30__8_), .Y(_7717_) );
OAI21X1 OAI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15175__bF_buf1), .C(_7717_), .Y(_7718_) );
NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_7699_), .Y(_7719_) );
AND2X2 AND2X2_1394 ( .gnd(gnd), .vdd(vdd), .A(_7719_), .B(_7718_), .Y(_180__8_) );
INVX1 INVX1_3369 ( .gnd(gnd), .vdd(vdd), .A(data_30__9_), .Y(_7720_) );
OAI21X1 OAI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15175__bF_buf0), .C(_7720_), .Y(_7721_) );
NAND3X1 NAND3X1_996 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_14984__bF_buf2), .C(_15793__bF_buf5), .Y(_7722_) );
AND2X2 AND2X2_1395 ( .gnd(gnd), .vdd(vdd), .A(_7721_), .B(_7722_), .Y(_180__9_) );
INVX1 INVX1_3370 ( .gnd(gnd), .vdd(vdd), .A(data_30__10_), .Y(_7723_) );
OAI21X1 OAI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15175__bF_buf4), .C(_7723_), .Y(_7724_) );
OAI21X1 OAI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf3), .B(_7693_), .C(_7724_), .Y(_7725_) );
INVX1 INVX1_3371 ( .gnd(gnd), .vdd(vdd), .A(_7725_), .Y(_180__10_) );
INVX1 INVX1_3372 ( .gnd(gnd), .vdd(vdd), .A(data_30__11_), .Y(_7726_) );
OAI21X1 OAI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15175__bF_buf3), .C(_7726_), .Y(_7727_) );
NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_7699_), .Y(_7728_) );
AND2X2 AND2X2_1396 ( .gnd(gnd), .vdd(vdd), .A(_7728_), .B(_7727_), .Y(_180__11_) );
INVX1 INVX1_3373 ( .gnd(gnd), .vdd(vdd), .A(data_30__12_), .Y(_7729_) );
OAI21X1 OAI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15175__bF_buf2), .C(_7729_), .Y(_7730_) );
OAI21X1 OAI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf1), .B(_7693_), .C(_7730_), .Y(_7731_) );
INVX1 INVX1_3374 ( .gnd(gnd), .vdd(vdd), .A(_7731_), .Y(_180__12_) );
INVX1 INVX1_3375 ( .gnd(gnd), .vdd(vdd), .A(data_30__13_), .Y(_7732_) );
OAI21X1 OAI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15175__bF_buf1), .C(_7732_), .Y(_7733_) );
NAND3X1 NAND3X1_997 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_14984__bF_buf1), .C(_15793__bF_buf4), .Y(_7734_) );
AND2X2 AND2X2_1397 ( .gnd(gnd), .vdd(vdd), .A(_7733_), .B(_7734_), .Y(_180__13_) );
AOI21X1 AOI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf0), .B(_15793__bF_buf3), .C(data_30__14_), .Y(_7735_) );
NOR2X1 NOR2X1_825 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf1), .B(_7693_), .Y(_7736_) );
NOR2X1 NOR2X1_826 ( .gnd(gnd), .vdd(vdd), .A(_7735_), .B(_7736_), .Y(_180__14_) );
INVX1 INVX1_3376 ( .gnd(gnd), .vdd(vdd), .A(data_30__15_), .Y(_7737_) );
OAI21X1 OAI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15175__bF_buf0), .C(_7737_), .Y(_7738_) );
NAND3X1 NAND3X1_998 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf3), .B(_14984__bF_buf4), .C(_15793__bF_buf2), .Y(_7739_) );
AND2X2 AND2X2_1398 ( .gnd(gnd), .vdd(vdd), .A(_7738_), .B(_7739_), .Y(_180__15_) );
INVX1 INVX1_3377 ( .gnd(gnd), .vdd(vdd), .A(data_29__0_), .Y(_7740_) );
OAI21X1 OAI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_addr_3_bF_buf2), .B(IDATA_PROG_addr[2]), .C(_14984__bF_buf3), .Y(_7741_) );
OAI21X1 OAI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_7741_), .B(_14963__bF_buf2), .C(_7508_), .Y(_7742_) );
INVX1 INVX1_3378 ( .gnd(gnd), .vdd(vdd), .A(_7742_), .Y(_7743_) );
AOI21X1 AOI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf2), .B(_15078_), .C(_15178_), .Y(_7744_) );
NAND3X1 NAND3X1_999 ( .gnd(gnd), .vdd(vdd), .A(_14979_), .B(_7744_), .C(_7743_), .Y(_7745_) );
NOR2X1 NOR2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_7745_), .B(_5459__bF_buf2), .Y(_7746_) );
NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .B(_3313__bF_buf29), .Y(_7747_) );
MUX2X1 MUX2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_7740_), .B(_14932__bF_buf12), .S(_7747_), .Y(_178__0_) );
INVX1 INVX1_3379 ( .gnd(gnd), .vdd(vdd), .A(data_29__1_), .Y(_7748_) );
MUX2X1 MUX2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_7748_), .B(_14894__bF_buf10), .S(_7747_), .Y(_178__1_) );
INVX1 INVX1_3380 ( .gnd(gnd), .vdd(vdd), .A(data_29__2_), .Y(_7749_) );
MUX2X1 MUX2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_7749_), .B(_14897__bF_buf6), .S(_7747_), .Y(_178__2_) );
INVX1 INVX1_3381 ( .gnd(gnd), .vdd(vdd), .A(data_29__3_), .Y(_7750_) );
MUX2X1 MUX2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_7750_), .B(_14899__bF_buf11), .S(_7747_), .Y(_178__3_) );
INVX1 INVX1_3382 ( .gnd(gnd), .vdd(vdd), .A(data_29__4_), .Y(_7751_) );
MUX2X1 MUX2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_7751_), .B(_14902__bF_buf1), .S(_7747_), .Y(_178__4_) );
INVX1 INVX1_3383 ( .gnd(gnd), .vdd(vdd), .A(data_29__5_), .Y(_7752_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(_7746_), .Y(_7753_) );
OAI21X1 OAI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf29), .B(_7753_), .C(_7752_), .Y(_7754_) );
NAND3X1 NAND3X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_7746_), .C(_3313__bF_buf28), .Y(_7755_) );
AND2X2 AND2X2_1399 ( .gnd(gnd), .vdd(vdd), .A(_7754_), .B(_7755_), .Y(_178__5_) );
INVX1 INVX1_3384 ( .gnd(gnd), .vdd(vdd), .A(data_29__6_), .Y(_7756_) );
MUX2X1 MUX2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_7756_), .B(_15049__bF_buf10), .S(_7747_), .Y(_178__6_) );
INVX1 INVX1_3385 ( .gnd(gnd), .vdd(vdd), .A(data_29__7_), .Y(_7757_) );
OAI21X1 OAI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf28), .B(_7753_), .C(_7757_), .Y(_7758_) );
NAND3X1 NAND3X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf2), .B(_7746_), .C(_3313__bF_buf27), .Y(_7759_) );
AND2X2 AND2X2_1400 ( .gnd(gnd), .vdd(vdd), .A(_7758_), .B(_7759_), .Y(_178__7_) );
INVX1 INVX1_3386 ( .gnd(gnd), .vdd(vdd), .A(data_29__8_), .Y(_7760_) );
MUX2X1 MUX2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_7760_), .B(_15052__bF_buf13), .S(_7747_), .Y(_178__8_) );
INVX1 INVX1_3387 ( .gnd(gnd), .vdd(vdd), .A(data_29__9_), .Y(_7761_) );
MUX2X1 MUX2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_7761_), .B(_14913__bF_buf7), .S(_7747_), .Y(_178__9_) );
INVX1 INVX1_3388 ( .gnd(gnd), .vdd(vdd), .A(data_29__10_), .Y(_7762_) );
MUX2X1 MUX2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_7762_), .B(_15055__bF_buf0), .S(_7747_), .Y(_178__10_) );
INVX1 INVX1_3389 ( .gnd(gnd), .vdd(vdd), .A(data_29__11_), .Y(_7763_) );
MUX2X1 MUX2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_7763_), .B(_14918__bF_buf1), .S(_7747_), .Y(_178__11_) );
INVX1 INVX1_3390 ( .gnd(gnd), .vdd(vdd), .A(data_29__12_), .Y(_7764_) );
OAI21X1 OAI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf27), .B(_7753_), .C(_7764_), .Y(_7765_) );
NAND3X1 NAND3X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_7746_), .C(_3313__bF_buf26), .Y(_7766_) );
AND2X2 AND2X2_1401 ( .gnd(gnd), .vdd(vdd), .A(_7765_), .B(_7766_), .Y(_178__12_) );
INVX1 INVX1_3391 ( .gnd(gnd), .vdd(vdd), .A(data_29__13_), .Y(_7767_) );
MUX2X1 MUX2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_7767_), .B(_14924__bF_buf13), .S(_7747_), .Y(_178__13_) );
INVX1 INVX1_3392 ( .gnd(gnd), .vdd(vdd), .A(data_29__14_), .Y(_7768_) );
MUX2X1 MUX2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_7768_), .B(_15060__bF_buf11), .S(_7747_), .Y(_178__14_) );
INVX1 INVX1_3393 ( .gnd(gnd), .vdd(vdd), .A(data_29__15_), .Y(_7769_) );
MUX2X1 MUX2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_7769_), .B(_15062__bF_buf2), .S(_7747_), .Y(_178__15_) );
INVX1 INVX1_3394 ( .gnd(gnd), .vdd(vdd), .A(data_28__0_), .Y(_7770_) );
NOR2X1 NOR2X1_828 ( .gnd(gnd), .vdd(vdd), .A(_14988_), .B(_5459__bF_buf1), .Y(_7771_) );
NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_7743_), .B(_7771_), .Y(_7772_) );
OAI21X1 OAI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf26), .B(_7772_), .C(_7770_), .Y(_7773_) );
INVX8 INVX8_32 ( .gnd(gnd), .vdd(vdd), .A(_7772_), .Y(_7774_) );
NAND3X1 NAND3X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_7774_), .C(_3313__bF_buf25), .Y(_7775_) );
AND2X2 AND2X2_1402 ( .gnd(gnd), .vdd(vdd), .A(_7773_), .B(_7775_), .Y(_177__0_) );
INVX1 INVX1_3395 ( .gnd(gnd), .vdd(vdd), .A(data_28__1_), .Y(_7776_) );
OAI21X1 OAI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf25), .B(_7772_), .C(_7776_), .Y(_7777_) );
NAND3X1 NAND3X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_7774_), .C(_3313__bF_buf24), .Y(_7778_) );
AND2X2 AND2X2_1403 ( .gnd(gnd), .vdd(vdd), .A(_7777_), .B(_7778_), .Y(_177__1_) );
NOR2X1 NOR2X1_829 ( .gnd(gnd), .vdd(vdd), .A(_7772_), .B(_3393__bF_buf24), .Y(_7779_) );
AOI21X1 AOI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf23), .C(data_28__2_), .Y(_7780_) );
AOI21X1 AOI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf5), .B(_7779_), .C(_7780_), .Y(_177__2_) );
INVX1 INVX1_3396 ( .gnd(gnd), .vdd(vdd), .A(data_28__3_), .Y(_7781_) );
OAI21X1 OAI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf23), .B(_7772_), .C(_7781_), .Y(_7782_) );
NAND3X1 NAND3X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf10), .B(_7774_), .C(_3313__bF_buf22), .Y(_7783_) );
AND2X2 AND2X2_1404 ( .gnd(gnd), .vdd(vdd), .A(_7782_), .B(_7783_), .Y(_177__3_) );
INVX1 INVX1_3397 ( .gnd(gnd), .vdd(vdd), .A(data_28__4_), .Y(_7784_) );
OAI21X1 OAI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf22), .B(_7772_), .C(_7784_), .Y(_7785_) );
NAND3X1 NAND3X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_7774_), .C(_3313__bF_buf21), .Y(_7786_) );
AND2X2 AND2X2_1405 ( .gnd(gnd), .vdd(vdd), .A(_7785_), .B(_7786_), .Y(_177__4_) );
AOI21X1 AOI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf20), .C(data_28__5_), .Y(_7787_) );
AOI21X1 AOI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf13), .B(_7779_), .C(_7787_), .Y(_177__5_) );
AOI21X1 AOI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf19), .C(data_28__6_), .Y(_7788_) );
AOI21X1 AOI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_7779_), .C(_7788_), .Y(_177__6_) );
AOI21X1 AOI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf18), .C(data_28__7_), .Y(_7789_) );
AOI21X1 AOI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_7779_), .C(_7789_), .Y(_177__7_) );
AOI21X1 AOI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf17), .C(data_28__8_), .Y(_7790_) );
AOI21X1 AOI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf12), .B(_7779_), .C(_7790_), .Y(_177__8_) );
INVX1 INVX1_3398 ( .gnd(gnd), .vdd(vdd), .A(data_28__9_), .Y(_7791_) );
NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf16), .Y(_7792_) );
MUX2X1 MUX2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_7791_), .B(_14913__bF_buf6), .S(_7792_), .Y(_177__9_) );
INVX1 INVX1_3399 ( .gnd(gnd), .vdd(vdd), .A(data_28__10_), .Y(_7793_) );
MUX2X1 MUX2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_7793_), .B(_15055__bF_buf13), .S(_7792_), .Y(_177__10_) );
INVX1 INVX1_3400 ( .gnd(gnd), .vdd(vdd), .A(data_28__11_), .Y(_7794_) );
OAI21X1 OAI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf21), .B(_7772_), .C(_7794_), .Y(_7795_) );
NAND3X1 NAND3X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf0), .B(_7774_), .C(_3313__bF_buf15), .Y(_7796_) );
AND2X2 AND2X2_1406 ( .gnd(gnd), .vdd(vdd), .A(_7795_), .B(_7796_), .Y(_177__11_) );
AOI21X1 AOI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf14), .C(data_28__12_), .Y(_7797_) );
AOI21X1 AOI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf1), .B(_7779_), .C(_7797_), .Y(_177__12_) );
INVX1 INVX1_3401 ( .gnd(gnd), .vdd(vdd), .A(data_28__13_), .Y(_7798_) );
MUX2X1 MUX2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_7798_), .B(_14924__bF_buf12), .S(_7792_), .Y(_177__13_) );
AOI21X1 AOI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf13), .C(data_28__14_), .Y(_7799_) );
AOI21X1 AOI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_7779_), .C(_7799_), .Y(_177__14_) );
AOI21X1 AOI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_7774_), .B(_3313__bF_buf12), .C(data_28__15_), .Y(_7800_) );
AOI21X1 AOI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_7779_), .C(_7800_), .Y(_177__15_) );
INVX1 INVX1_3402 ( .gnd(gnd), .vdd(vdd), .A(data_27__0_), .Y(_7801_) );
INVX1 INVX1_3403 ( .gnd(gnd), .vdd(vdd), .A(_7771_), .Y(_7802_) );
INVX1 INVX1_3404 ( .gnd(gnd), .vdd(vdd), .A(_7508_), .Y(_7803_) );
AOI21X1 AOI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf1), .B(_15161_), .C(_7803_), .Y(_7804_) );
OAI21X1 OAI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_15175__bF_buf4), .C(_7804_), .Y(_7805_) );
OR2X2 OR2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_7802_), .B(_7805_), .Y(_7806_) );
OAI21X1 OAI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf20), .C(_7801_), .Y(_7807_) );
NOR2X1 NOR2X1_830 ( .gnd(gnd), .vdd(vdd), .A(_7805_), .B(_7802_), .Y(_7808_) );
NAND3X1 NAND3X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf10), .B(_7808_), .C(_3313__bF_buf11), .Y(_7809_) );
AND2X2 AND2X2_1407 ( .gnd(gnd), .vdd(vdd), .A(_7807_), .B(_7809_), .Y(_176__0_) );
INVX1 INVX1_3405 ( .gnd(gnd), .vdd(vdd), .A(data_27__1_), .Y(_7810_) );
OAI21X1 OAI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf19), .C(_7810_), .Y(_7811_) );
NAND3X1 NAND3X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf8), .B(_7808_), .C(_3313__bF_buf10), .Y(_7812_) );
AND2X2 AND2X2_1408 ( .gnd(gnd), .vdd(vdd), .A(_7811_), .B(_7812_), .Y(_176__1_) );
INVX1 INVX1_3406 ( .gnd(gnd), .vdd(vdd), .A(data_27__2_), .Y(_7813_) );
NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_7808_), .B(_3313__bF_buf9), .Y(_7814_) );
MUX2X1 MUX2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_7813_), .B(_14897__bF_buf4), .S(_7814_), .Y(_176__2_) );
INVX1 INVX1_3407 ( .gnd(gnd), .vdd(vdd), .A(data_27__3_), .Y(_7815_) );
OAI21X1 OAI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf18), .C(_7815_), .Y(_7816_) );
NAND3X1 NAND3X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_7808_), .C(_3313__bF_buf8), .Y(_7817_) );
AND2X2 AND2X2_1409 ( .gnd(gnd), .vdd(vdd), .A(_7816_), .B(_7817_), .Y(_176__3_) );
INVX1 INVX1_3408 ( .gnd(gnd), .vdd(vdd), .A(data_27__4_), .Y(_7818_) );
OAI21X1 OAI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf17), .C(_7818_), .Y(_7819_) );
NAND3X1 NAND3X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf13), .B(_7808_), .C(_3313__bF_buf7), .Y(_7820_) );
AND2X2 AND2X2_1410 ( .gnd(gnd), .vdd(vdd), .A(_7819_), .B(_7820_), .Y(_176__4_) );
INVX1 INVX1_3409 ( .gnd(gnd), .vdd(vdd), .A(data_27__5_), .Y(_7821_) );
OAI21X1 OAI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf16), .C(_7821_), .Y(_7822_) );
NAND3X1 NAND3X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_7808_), .C(_3313__bF_buf6), .Y(_7823_) );
AND2X2 AND2X2_1411 ( .gnd(gnd), .vdd(vdd), .A(_7822_), .B(_7823_), .Y(_176__5_) );
INVX1 INVX1_3410 ( .gnd(gnd), .vdd(vdd), .A(data_27__6_), .Y(_7824_) );
MUX2X1 MUX2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_7824_), .B(_15049__bF_buf8), .S(_7814_), .Y(_176__6_) );
INVX1 INVX1_3411 ( .gnd(gnd), .vdd(vdd), .A(data_27__7_), .Y(_7825_) );
OAI21X1 OAI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf15), .C(_7825_), .Y(_7826_) );
NAND3X1 NAND3X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf0), .B(_7808_), .C(_3313__bF_buf5), .Y(_7827_) );
AND2X2 AND2X2_1412 ( .gnd(gnd), .vdd(vdd), .A(_7826_), .B(_7827_), .Y(_176__7_) );
INVX1 INVX1_3412 ( .gnd(gnd), .vdd(vdd), .A(data_27__8_), .Y(_7828_) );
MUX2X1 MUX2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_7828_), .B(_15052__bF_buf11), .S(_7814_), .Y(_176__8_) );
INVX1 INVX1_3413 ( .gnd(gnd), .vdd(vdd), .A(data_27__9_), .Y(_7829_) );
MUX2X1 MUX2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_7829_), .B(_14913__bF_buf5), .S(_7814_), .Y(_176__9_) );
INVX1 INVX1_3414 ( .gnd(gnd), .vdd(vdd), .A(data_27__10_), .Y(_7830_) );
MUX2X1 MUX2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_7830_), .B(_15055__bF_buf12), .S(_7814_), .Y(_176__10_) );
INVX1 INVX1_3415 ( .gnd(gnd), .vdd(vdd), .A(data_27__11_), .Y(_7831_) );
OAI21X1 OAI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf14), .C(_7831_), .Y(_7832_) );
NAND3X1 NAND3X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_7808_), .C(_3313__bF_buf4), .Y(_7833_) );
AND2X2 AND2X2_1413 ( .gnd(gnd), .vdd(vdd), .A(_7832_), .B(_7833_), .Y(_176__11_) );
INVX1 INVX1_3416 ( .gnd(gnd), .vdd(vdd), .A(data_27__12_), .Y(_7834_) );
OAI21X1 OAI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_7806_), .B(_3393__bF_buf13), .C(_7834_), .Y(_7835_) );
NAND3X1 NAND3X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_7808_), .C(_3313__bF_buf3), .Y(_7836_) );
AND2X2 AND2X2_1414 ( .gnd(gnd), .vdd(vdd), .A(_7835_), .B(_7836_), .Y(_176__12_) );
INVX1 INVX1_3417 ( .gnd(gnd), .vdd(vdd), .A(data_27__13_), .Y(_7837_) );
MUX2X1 MUX2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_7837_), .B(_14924__bF_buf11), .S(_7814_), .Y(_176__13_) );
INVX1 INVX1_3418 ( .gnd(gnd), .vdd(vdd), .A(data_27__14_), .Y(_7838_) );
MUX2X1 MUX2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_7838_), .B(_15060__bF_buf9), .S(_7814_), .Y(_176__14_) );
INVX1 INVX1_3419 ( .gnd(gnd), .vdd(vdd), .A(data_27__15_), .Y(_7839_) );
MUX2X1 MUX2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_7839_), .B(_15062__bF_buf0), .S(_7814_), .Y(_176__15_) );
INVX1 INVX1_3420 ( .gnd(gnd), .vdd(vdd), .A(data_26__0_), .Y(_7840_) );
OAI21X1 OAI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_14964_), .B(_15175__bF_buf3), .C(_7508_), .Y(_7841_) );
INVX1 INVX1_3421 ( .gnd(gnd), .vdd(vdd), .A(_7841_), .Y(_7842_) );
OAI21X1 OAI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_14952__bF_buf3), .C(_14984__bF_buf0), .Y(_7843_) );
NAND3X1 NAND3X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_7842_), .B(_7843_), .C(_7771_), .Y(_7844_) );
OAI21X1 OAI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf12), .B(_7844_), .C(_7840_), .Y(_7845_) );
INVX4 INVX4_37 ( .gnd(gnd), .vdd(vdd), .A(_7844_), .Y(_7846_) );
NAND3X1 NAND3X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf9), .B(_7846_), .C(_3313__bF_buf2), .Y(_7847_) );
AND2X2 AND2X2_1415 ( .gnd(gnd), .vdd(vdd), .A(_7845_), .B(_7847_), .Y(_175__0_) );
INVX1 INVX1_3422 ( .gnd(gnd), .vdd(vdd), .A(data_26__1_), .Y(_7848_) );
OAI21X1 OAI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf11), .B(_7844_), .C(_7848_), .Y(_7849_) );
NAND3X1 NAND3X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf7), .B(_7846_), .C(_3313__bF_buf1), .Y(_7850_) );
AND2X2 AND2X2_1416 ( .gnd(gnd), .vdd(vdd), .A(_7849_), .B(_7850_), .Y(_175__1_) );
INVX1 INVX1_3423 ( .gnd(gnd), .vdd(vdd), .A(data_26__2_), .Y(_7851_) );
NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_7846_), .B(_3313__bF_buf0), .Y(_7852_) );
MUX2X1 MUX2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_7851_), .B(_14897__bF_buf3), .S(_7852_), .Y(_175__2_) );
INVX1 INVX1_3424 ( .gnd(gnd), .vdd(vdd), .A(data_26__3_), .Y(_7853_) );
OAI21X1 OAI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf10), .B(_7844_), .C(_7853_), .Y(_7854_) );
NAND3X1 NAND3X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf8), .B(_7846_), .C(_3313__bF_buf91), .Y(_7855_) );
AND2X2 AND2X2_1417 ( .gnd(gnd), .vdd(vdd), .A(_7854_), .B(_7855_), .Y(_175__3_) );
INVX1 INVX1_3425 ( .gnd(gnd), .vdd(vdd), .A(data_26__4_), .Y(_7856_) );
OAI21X1 OAI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf9), .B(_7844_), .C(_7856_), .Y(_7857_) );
NAND3X1 NAND3X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf12), .B(_7846_), .C(_3313__bF_buf90), .Y(_7858_) );
AND2X2 AND2X2_1418 ( .gnd(gnd), .vdd(vdd), .A(_7857_), .B(_7858_), .Y(_175__4_) );
INVX1 INVX1_3426 ( .gnd(gnd), .vdd(vdd), .A(data_26__5_), .Y(_7859_) );
OAI21X1 OAI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf8), .B(_7844_), .C(_7859_), .Y(_7860_) );
NAND3X1 NAND3X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf11), .B(_7846_), .C(_3313__bF_buf89), .Y(_7861_) );
AND2X2 AND2X2_1419 ( .gnd(gnd), .vdd(vdd), .A(_7860_), .B(_7861_), .Y(_175__5_) );
INVX1 INVX1_3427 ( .gnd(gnd), .vdd(vdd), .A(data_26__6_), .Y(_7862_) );
MUX2X1 MUX2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_7862_), .B(_15049__bF_buf7), .S(_7852_), .Y(_175__6_) );
INVX1 INVX1_3428 ( .gnd(gnd), .vdd(vdd), .A(data_26__7_), .Y(_7863_) );
OAI21X1 OAI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf7), .B(_7844_), .C(_7863_), .Y(_7864_) );
NAND3X1 NAND3X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf13), .B(_7846_), .C(_3313__bF_buf88), .Y(_7865_) );
AND2X2 AND2X2_1420 ( .gnd(gnd), .vdd(vdd), .A(_7864_), .B(_7865_), .Y(_175__7_) );
INVX1 INVX1_3429 ( .gnd(gnd), .vdd(vdd), .A(data_26__8_), .Y(_7866_) );
MUX2X1 MUX2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_7866_), .B(_15052__bF_buf10), .S(_7852_), .Y(_175__8_) );
INVX1 INVX1_3430 ( .gnd(gnd), .vdd(vdd), .A(data_26__9_), .Y(_7867_) );
MUX2X1 MUX2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_7867_), .B(_14913__bF_buf4), .S(_7852_), .Y(_175__9_) );
INVX1 INVX1_3431 ( .gnd(gnd), .vdd(vdd), .A(data_26__10_), .Y(_7868_) );
MUX2X1 MUX2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_7868_), .B(_15055__bF_buf11), .S(_7852_), .Y(_175__10_) );
INVX1 INVX1_3432 ( .gnd(gnd), .vdd(vdd), .A(data_26__11_), .Y(_7869_) );
OAI21X1 OAI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf6), .B(_7844_), .C(_7869_), .Y(_7870_) );
NAND3X1 NAND3X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf12), .B(_7846_), .C(_3313__bF_buf87), .Y(_7871_) );
AND2X2 AND2X2_1421 ( .gnd(gnd), .vdd(vdd), .A(_7870_), .B(_7871_), .Y(_175__11_) );
INVX1 INVX1_3433 ( .gnd(gnd), .vdd(vdd), .A(data_26__12_), .Y(_7872_) );
OAI21X1 OAI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf5), .B(_7844_), .C(_7872_), .Y(_7873_) );
NAND3X1 NAND3X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf13), .B(_7846_), .C(_3313__bF_buf86), .Y(_7874_) );
AND2X2 AND2X2_1422 ( .gnd(gnd), .vdd(vdd), .A(_7873_), .B(_7874_), .Y(_175__12_) );
INVX1 INVX1_3434 ( .gnd(gnd), .vdd(vdd), .A(data_26__13_), .Y(_7875_) );
MUX2X1 MUX2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_7875_), .B(_14924__bF_buf10), .S(_7852_), .Y(_175__13_) );
INVX1 INVX1_3435 ( .gnd(gnd), .vdd(vdd), .A(data_26__14_), .Y(_7876_) );
MUX2X1 MUX2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_7876_), .B(_15060__bF_buf8), .S(_7852_), .Y(_175__14_) );
INVX1 INVX1_3436 ( .gnd(gnd), .vdd(vdd), .A(data_26__15_), .Y(_7877_) );
MUX2X1 MUX2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_7877_), .B(_15062__bF_buf13), .S(_7852_), .Y(_175__15_) );
INVX1 INVX1_3437 ( .gnd(gnd), .vdd(vdd), .A(data_25__0_), .Y(_7878_) );
OAI21X1 OAI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_15285_), .B(_14952__bF_buf2), .C(_14984__bF_buf4), .Y(_7879_) );
NAND3X1 NAND3X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_7842_), .B(_7879_), .C(_7771_), .Y(_7880_) );
OAI21X1 OAI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf4), .B(_7880_), .C(_7878_), .Y(_7881_) );
INVX4 INVX4_38 ( .gnd(gnd), .vdd(vdd), .A(_7880_), .Y(_7882_) );
NAND3X1 NAND3X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_7882_), .C(_3313__bF_buf85), .Y(_7883_) );
AND2X2 AND2X2_1423 ( .gnd(gnd), .vdd(vdd), .A(_7881_), .B(_7883_), .Y(_174__0_) );
INVX1 INVX1_3438 ( .gnd(gnd), .vdd(vdd), .A(data_25__1_), .Y(_7884_) );
OAI21X1 OAI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf3), .B(_7880_), .C(_7884_), .Y(_7885_) );
NAND3X1 NAND3X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_7882_), .C(_3313__bF_buf84), .Y(_7886_) );
AND2X2 AND2X2_1424 ( .gnd(gnd), .vdd(vdd), .A(_7885_), .B(_7886_), .Y(_174__1_) );
INVX1 INVX1_3439 ( .gnd(gnd), .vdd(vdd), .A(data_25__2_), .Y(_7887_) );
NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_7882_), .B(_3313__bF_buf83), .Y(_7888_) );
MUX2X1 MUX2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_7887_), .B(_14897__bF_buf2), .S(_7888_), .Y(_174__2_) );
INVX1 INVX1_3440 ( .gnd(gnd), .vdd(vdd), .A(data_25__3_), .Y(_7889_) );
OAI21X1 OAI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf2), .B(_7880_), .C(_7889_), .Y(_7890_) );
NAND3X1 NAND3X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf7), .B(_7882_), .C(_3313__bF_buf82), .Y(_7891_) );
AND2X2 AND2X2_1425 ( .gnd(gnd), .vdd(vdd), .A(_7890_), .B(_7891_), .Y(_174__3_) );
INVX1 INVX1_3441 ( .gnd(gnd), .vdd(vdd), .A(data_25__4_), .Y(_7892_) );
OAI21X1 OAI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf1), .B(_7880_), .C(_7892_), .Y(_7893_) );
NAND3X1 NAND3X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_7882_), .C(_3313__bF_buf81), .Y(_7894_) );
AND2X2 AND2X2_1426 ( .gnd(gnd), .vdd(vdd), .A(_7893_), .B(_7894_), .Y(_174__4_) );
INVX1 INVX1_3442 ( .gnd(gnd), .vdd(vdd), .A(data_25__5_), .Y(_7895_) );
OAI21X1 OAI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf0), .B(_7880_), .C(_7895_), .Y(_7896_) );
NAND3X1 NAND3X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf10), .B(_7882_), .C(_3313__bF_buf80), .Y(_7897_) );
AND2X2 AND2X2_1427 ( .gnd(gnd), .vdd(vdd), .A(_7896_), .B(_7897_), .Y(_174__5_) );
INVX1 INVX1_3443 ( .gnd(gnd), .vdd(vdd), .A(data_25__6_), .Y(_7898_) );
MUX2X1 MUX2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_7898_), .B(_15049__bF_buf6), .S(_7888_), .Y(_174__6_) );
INVX1 INVX1_3444 ( .gnd(gnd), .vdd(vdd), .A(data_25__7_), .Y(_7899_) );
OAI21X1 OAI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf69), .B(_7880_), .C(_7899_), .Y(_7900_) );
NAND3X1 NAND3X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_7882_), .C(_3313__bF_buf79), .Y(_7901_) );
AND2X2 AND2X2_1428 ( .gnd(gnd), .vdd(vdd), .A(_7900_), .B(_7901_), .Y(_174__7_) );
INVX1 INVX1_3445 ( .gnd(gnd), .vdd(vdd), .A(data_25__8_), .Y(_7902_) );
MUX2X1 MUX2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_7902_), .B(_15052__bF_buf9), .S(_7888_), .Y(_174__8_) );
INVX1 INVX1_3446 ( .gnd(gnd), .vdd(vdd), .A(data_25__9_), .Y(_7903_) );
MUX2X1 MUX2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_7903_), .B(_14913__bF_buf3), .S(_7888_), .Y(_174__9_) );
INVX1 INVX1_3447 ( .gnd(gnd), .vdd(vdd), .A(data_25__10_), .Y(_7904_) );
MUX2X1 MUX2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7904_), .B(_15055__bF_buf10), .S(_7888_), .Y(_174__10_) );
INVX1 INVX1_3448 ( .gnd(gnd), .vdd(vdd), .A(data_25__11_), .Y(_7905_) );
OAI21X1 OAI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf68), .B(_7880_), .C(_7905_), .Y(_7906_) );
NAND3X1 NAND3X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf11), .B(_7882_), .C(_3313__bF_buf78), .Y(_7907_) );
AND2X2 AND2X2_1429 ( .gnd(gnd), .vdd(vdd), .A(_7906_), .B(_7907_), .Y(_174__11_) );
INVX1 INVX1_3449 ( .gnd(gnd), .vdd(vdd), .A(data_25__12_), .Y(_7908_) );
OAI21X1 OAI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf67), .B(_7880_), .C(_7908_), .Y(_7909_) );
NAND3X1 NAND3X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf12), .B(_7882_), .C(_3313__bF_buf77), .Y(_7910_) );
AND2X2 AND2X2_1430 ( .gnd(gnd), .vdd(vdd), .A(_7909_), .B(_7910_), .Y(_174__12_) );
INVX1 INVX1_3450 ( .gnd(gnd), .vdd(vdd), .A(data_25__13_), .Y(_7911_) );
MUX2X1 MUX2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_7911_), .B(_14924__bF_buf9), .S(_7888_), .Y(_174__13_) );
INVX1 INVX1_3451 ( .gnd(gnd), .vdd(vdd), .A(data_25__14_), .Y(_7912_) );
MUX2X1 MUX2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_7912_), .B(_15060__bF_buf7), .S(_7888_), .Y(_174__14_) );
INVX1 INVX1_3452 ( .gnd(gnd), .vdd(vdd), .A(data_25__15_), .Y(_7913_) );
MUX2X1 MUX2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_7913_), .B(_15062__bF_buf12), .S(_7888_), .Y(_174__15_) );
INVX1 INVX1_3453 ( .gnd(gnd), .vdd(vdd), .A(data_24__0_), .Y(_7914_) );
OAI21X1 OAI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_14977__bF_buf0), .B(_15175__bF_buf2), .C(_7508_), .Y(_7915_) );
NAND3X1 NAND3X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_15179_), .B(_14992_), .C(_14973_), .Y(_7916_) );
NOR2X1 NOR2X1_831 ( .gnd(gnd), .vdd(vdd), .A(_7915_), .B(_7916_), .Y(_7917_) );
INVX4 INVX4_39 ( .gnd(gnd), .vdd(vdd), .A(_7917_), .Y(_7918_) );
OAI21X1 OAI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf66), .B(_7918_), .C(_7914_), .Y(_7919_) );
NAND3X1 NAND3X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_7917_), .C(_3313__bF_buf76), .Y(_7920_) );
AND2X2 AND2X2_1431 ( .gnd(gnd), .vdd(vdd), .A(_7919_), .B(_7920_), .Y(_167__0_) );
INVX1 INVX1_3454 ( .gnd(gnd), .vdd(vdd), .A(data_24__1_), .Y(_7921_) );
OAI21X1 OAI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf65), .B(_7918_), .C(_7921_), .Y(_7922_) );
NAND3X1 NAND3X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf5), .B(_7917_), .C(_3313__bF_buf75), .Y(_7923_) );
AND2X2 AND2X2_1432 ( .gnd(gnd), .vdd(vdd), .A(_7922_), .B(_7923_), .Y(_167__1_) );
INVX1 INVX1_3455 ( .gnd(gnd), .vdd(vdd), .A(data_24__2_), .Y(_7924_) );
NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_7917_), .B(_3313__bF_buf74), .Y(_7925_) );
MUX2X1 MUX2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_7924_), .B(_14897__bF_buf1), .S(_7925_), .Y(_167__2_) );
INVX1 INVX1_3456 ( .gnd(gnd), .vdd(vdd), .A(data_24__3_), .Y(_7926_) );
OAI21X1 OAI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf64), .B(_7918_), .C(_7926_), .Y(_7927_) );
NAND3X1 NAND3X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_7917_), .C(_3313__bF_buf73), .Y(_7928_) );
AND2X2 AND2X2_1433 ( .gnd(gnd), .vdd(vdd), .A(_7927_), .B(_7928_), .Y(_167__3_) );
INVX1 INVX1_3457 ( .gnd(gnd), .vdd(vdd), .A(data_24__4_), .Y(_7929_) );
OAI21X1 OAI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf63), .B(_7918_), .C(_7929_), .Y(_7930_) );
NAND3X1 NAND3X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf10), .B(_7917_), .C(_3313__bF_buf72), .Y(_7931_) );
AND2X2 AND2X2_1434 ( .gnd(gnd), .vdd(vdd), .A(_7930_), .B(_7931_), .Y(_167__4_) );
INVX1 INVX1_3458 ( .gnd(gnd), .vdd(vdd), .A(data_24__5_), .Y(_7932_) );
OAI21X1 OAI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf62), .B(_7918_), .C(_7932_), .Y(_7933_) );
NAND3X1 NAND3X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_7917_), .C(_3313__bF_buf71), .Y(_7934_) );
AND2X2 AND2X2_1435 ( .gnd(gnd), .vdd(vdd), .A(_7933_), .B(_7934_), .Y(_167__5_) );
INVX1 INVX1_3459 ( .gnd(gnd), .vdd(vdd), .A(data_24__6_), .Y(_7935_) );
MUX2X1 MUX2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_7935_), .B(_15049__bF_buf5), .S(_7925_), .Y(_167__6_) );
INVX1 INVX1_3460 ( .gnd(gnd), .vdd(vdd), .A(data_24__7_), .Y(_7936_) );
OAI21X1 OAI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf61), .B(_7918_), .C(_7936_), .Y(_7937_) );
NAND3X1 NAND3X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf11), .B(_7917_), .C(_3313__bF_buf70), .Y(_7938_) );
AND2X2 AND2X2_1436 ( .gnd(gnd), .vdd(vdd), .A(_7937_), .B(_7938_), .Y(_167__7_) );
INVX1 INVX1_3461 ( .gnd(gnd), .vdd(vdd), .A(data_24__8_), .Y(_7939_) );
MUX2X1 MUX2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_7939_), .B(_15052__bF_buf8), .S(_7925_), .Y(_167__8_) );
INVX1 INVX1_3462 ( .gnd(gnd), .vdd(vdd), .A(data_24__9_), .Y(_7940_) );
MUX2X1 MUX2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_7940_), .B(_14913__bF_buf2), .S(_7925_), .Y(_167__9_) );
INVX1 INVX1_3463 ( .gnd(gnd), .vdd(vdd), .A(data_24__10_), .Y(_7941_) );
MUX2X1 MUX2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_7941_), .B(_15055__bF_buf9), .S(_7925_), .Y(_167__10_) );
INVX1 INVX1_3464 ( .gnd(gnd), .vdd(vdd), .A(data_24__11_), .Y(_7942_) );
OAI21X1 OAI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf60), .B(_7918_), .C(_7942_), .Y(_7943_) );
NAND3X1 NAND3X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_7917_), .C(_3313__bF_buf69), .Y(_7944_) );
AND2X2 AND2X2_1437 ( .gnd(gnd), .vdd(vdd), .A(_7943_), .B(_7944_), .Y(_167__11_) );
INVX1 INVX1_3465 ( .gnd(gnd), .vdd(vdd), .A(data_24__12_), .Y(_7945_) );
OAI21X1 OAI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf59), .B(_7918_), .C(_7945_), .Y(_7946_) );
NAND3X1 NAND3X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_7917_), .C(_3313__bF_buf68), .Y(_7947_) );
AND2X2 AND2X2_1438 ( .gnd(gnd), .vdd(vdd), .A(_7946_), .B(_7947_), .Y(_167__12_) );
INVX1 INVX1_3466 ( .gnd(gnd), .vdd(vdd), .A(data_24__13_), .Y(_7948_) );
MUX2X1 MUX2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_7948_), .B(_14924__bF_buf8), .S(_7925_), .Y(_167__13_) );
INVX1 INVX1_3467 ( .gnd(gnd), .vdd(vdd), .A(data_24__14_), .Y(_7949_) );
MUX2X1 MUX2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_7949_), .B(_15060__bF_buf6), .S(_7925_), .Y(_167__14_) );
INVX1 INVX1_3468 ( .gnd(gnd), .vdd(vdd), .A(data_24__15_), .Y(_7950_) );
MUX2X1 MUX2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_7950_), .B(_15062__bF_buf11), .S(_7925_), .Y(_167__15_) );
INVX1 INVX1_3469 ( .gnd(gnd), .vdd(vdd), .A(data_23__0_), .Y(_7951_) );
OAI21X1 OAI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_15175__bF_buf1), .B(_15360_), .C(_7508_), .Y(_7952_) );
AOI21X1 AOI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf3), .B(_15364_), .C(_7952_), .Y(_7953_) );
NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_7953_), .B(_7771_), .Y(_7954_) );
OAI21X1 OAI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf58), .B(_7954_), .C(_7951_), .Y(_7955_) );
INVX4 INVX4_40 ( .gnd(gnd), .vdd(vdd), .A(_7954_), .Y(_7956_) );
NAND3X1 NAND3X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf6), .B(_7956_), .C(_3313__bF_buf67), .Y(_7957_) );
AND2X2 AND2X2_1439 ( .gnd(gnd), .vdd(vdd), .A(_7955_), .B(_7957_), .Y(_156__0_) );
INVX1 INVX1_3470 ( .gnd(gnd), .vdd(vdd), .A(data_23__1_), .Y(_7958_) );
OAI21X1 OAI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf57), .B(_7954_), .C(_7958_), .Y(_7959_) );
NAND3X1 NAND3X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf4), .B(_7956_), .C(_3313__bF_buf66), .Y(_7960_) );
AND2X2 AND2X2_1440 ( .gnd(gnd), .vdd(vdd), .A(_7959_), .B(_7960_), .Y(_156__1_) );
INVX1 INVX1_3471 ( .gnd(gnd), .vdd(vdd), .A(data_23__2_), .Y(_7961_) );
NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_7956_), .B(_3313__bF_buf65), .Y(_7962_) );
MUX2X1 MUX2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_7961_), .B(_14897__bF_buf0), .S(_7962_), .Y(_156__2_) );
INVX1 INVX1_3472 ( .gnd(gnd), .vdd(vdd), .A(data_23__3_), .Y(_7963_) );
OAI21X1 OAI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf56), .B(_7954_), .C(_7963_), .Y(_7964_) );
NAND3X1 NAND3X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf5), .B(_7956_), .C(_3313__bF_buf64), .Y(_7965_) );
AND2X2 AND2X2_1441 ( .gnd(gnd), .vdd(vdd), .A(_7964_), .B(_7965_), .Y(_156__3_) );
INVX1 INVX1_3473 ( .gnd(gnd), .vdd(vdd), .A(data_23__4_), .Y(_7966_) );
OAI21X1 OAI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf55), .B(_7954_), .C(_7966_), .Y(_7967_) );
NAND3X1 NAND3X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf9), .B(_7956_), .C(_3313__bF_buf63), .Y(_7968_) );
AND2X2 AND2X2_1442 ( .gnd(gnd), .vdd(vdd), .A(_7967_), .B(_7968_), .Y(_156__4_) );
INVX1 INVX1_3474 ( .gnd(gnd), .vdd(vdd), .A(data_23__5_), .Y(_7969_) );
MUX2X1 MUX2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_7969_), .B(_14903__bF_buf8), .S(_7962_), .Y(_156__5_) );
INVX1 INVX1_3475 ( .gnd(gnd), .vdd(vdd), .A(data_23__6_), .Y(_7970_) );
MUX2X1 MUX2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_7970_), .B(_15049__bF_buf4), .S(_7962_), .Y(_156__6_) );
INVX1 INVX1_3476 ( .gnd(gnd), .vdd(vdd), .A(data_23__7_), .Y(_7971_) );
MUX2X1 MUX2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_7971_), .B(_14908__bF_buf10), .S(_7962_), .Y(_156__7_) );
INVX1 INVX1_3477 ( .gnd(gnd), .vdd(vdd), .A(data_23__8_), .Y(_7972_) );
MUX2X1 MUX2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_7972_), .B(_15052__bF_buf7), .S(_7962_), .Y(_156__8_) );
INVX1 INVX1_3478 ( .gnd(gnd), .vdd(vdd), .A(data_23__9_), .Y(_7973_) );
MUX2X1 MUX2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_7973_), .B(_14913__bF_buf1), .S(_7962_), .Y(_156__9_) );
INVX1 INVX1_3479 ( .gnd(gnd), .vdd(vdd), .A(data_23__10_), .Y(_7974_) );
MUX2X1 MUX2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_7974_), .B(_15055__bF_buf8), .S(_7962_), .Y(_156__10_) );
INVX1 INVX1_3480 ( .gnd(gnd), .vdd(vdd), .A(data_23__11_), .Y(_7975_) );
OAI21X1 OAI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf54), .B(_7954_), .C(_7975_), .Y(_7976_) );
NAND3X1 NAND3X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf9), .B(_7956_), .C(_3313__bF_buf62), .Y(_7977_) );
AND2X2 AND2X2_1443 ( .gnd(gnd), .vdd(vdd), .A(_7976_), .B(_7977_), .Y(_156__11_) );
INVX1 INVX1_3481 ( .gnd(gnd), .vdd(vdd), .A(data_23__12_), .Y(_7978_) );
MUX2X1 MUX2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_7978_), .B(_14920__bF_buf10), .S(_7962_), .Y(_156__12_) );
INVX1 INVX1_3482 ( .gnd(gnd), .vdd(vdd), .A(data_23__13_), .Y(_7979_) );
MUX2X1 MUX2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_7979_), .B(_14924__bF_buf7), .S(_7962_), .Y(_156__13_) );
INVX1 INVX1_3483 ( .gnd(gnd), .vdd(vdd), .A(data_23__14_), .Y(_7980_) );
MUX2X1 MUX2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_7980_), .B(_15060__bF_buf5), .S(_7962_), .Y(_156__14_) );
INVX1 INVX1_3484 ( .gnd(gnd), .vdd(vdd), .A(data_23__15_), .Y(_7981_) );
MUX2X1 MUX2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_7981_), .B(_15062__bF_buf10), .S(_7962_), .Y(_156__15_) );
INVX1 INVX1_3485 ( .gnd(gnd), .vdd(vdd), .A(data_22__0_), .Y(_7982_) );
OAI21X1 OAI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_14958_), .B(_15175__bF_buf0), .C(_7508_), .Y(_7983_) );
AOI21X1 AOI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf2), .B(_888_), .C(_7983_), .Y(_7984_) );
INVX1 INVX1_3486 ( .gnd(gnd), .vdd(vdd), .A(_7984_), .Y(_7985_) );
NOR2X1 NOR2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_7985_), .B(_7916_), .Y(_7986_) );
NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .B(_3313__bF_buf61), .Y(_7987_) );
MUX2X1 MUX2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_7982_), .B(_14932__bF_buf5), .S(_7987_), .Y(_145__0_) );
INVX1 INVX1_3487 ( .gnd(gnd), .vdd(vdd), .A(data_22__1_), .Y(_7988_) );
MUX2X1 MUX2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_7988_), .B(_14894__bF_buf3), .S(_7987_), .Y(_145__1_) );
INVX1 INVX1_3488 ( .gnd(gnd), .vdd(vdd), .A(data_22__2_), .Y(_7989_) );
MUX2X1 MUX2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_7989_), .B(_14897__bF_buf14), .S(_7987_), .Y(_145__2_) );
INVX1 INVX1_3489 ( .gnd(gnd), .vdd(vdd), .A(data_22__3_), .Y(_7990_) );
INVX4 INVX4_41 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .Y(_7991_) );
OAI21X1 OAI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf53), .B(_7991_), .C(_7990_), .Y(_7992_) );
NAND3X1 NAND3X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf4), .B(_7986_), .C(_3313__bF_buf60), .Y(_7993_) );
AND2X2 AND2X2_1444 ( .gnd(gnd), .vdd(vdd), .A(_7992_), .B(_7993_), .Y(_145__3_) );
INVX1 INVX1_3490 ( .gnd(gnd), .vdd(vdd), .A(data_22__4_), .Y(_7994_) );
MUX2X1 MUX2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_7994_), .B(_14902__bF_buf8), .S(_7987_), .Y(_145__4_) );
INVX1 INVX1_3491 ( .gnd(gnd), .vdd(vdd), .A(data_22__5_), .Y(_7995_) );
OAI21X1 OAI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf52), .B(_7991_), .C(_7995_), .Y(_7996_) );
NAND3X1 NAND3X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf7), .B(_7986_), .C(_3313__bF_buf59), .Y(_7997_) );
AND2X2 AND2X2_1445 ( .gnd(gnd), .vdd(vdd), .A(_7996_), .B(_7997_), .Y(_145__5_) );
INVX1 INVX1_3492 ( .gnd(gnd), .vdd(vdd), .A(data_22__6_), .Y(_7998_) );
MUX2X1 MUX2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_7998_), .B(_15049__bF_buf3), .S(_7987_), .Y(_145__6_) );
INVX1 INVX1_3493 ( .gnd(gnd), .vdd(vdd), .A(data_22__7_), .Y(_7999_) );
OAI21X1 OAI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf51), .B(_7991_), .C(_7999_), .Y(_8000_) );
NAND3X1 NAND3X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf9), .B(_7986_), .C(_3313__bF_buf58), .Y(_8001_) );
AND2X2 AND2X2_1446 ( .gnd(gnd), .vdd(vdd), .A(_8000_), .B(_8001_), .Y(_145__7_) );
INVX1 INVX1_3494 ( .gnd(gnd), .vdd(vdd), .A(data_22__8_), .Y(_8002_) );
MUX2X1 MUX2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_8002_), .B(_15052__bF_buf6), .S(_7987_), .Y(_145__8_) );
NOR2X1 NOR2X1_833 ( .gnd(gnd), .vdd(vdd), .A(_7991_), .B(_3393__bF_buf50), .Y(_8003_) );
AOI21X1 AOI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .B(_3313__bF_buf57), .C(data_22__9_), .Y(_8004_) );
AOI21X1 AOI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf0), .B(_8003_), .C(_8004_), .Y(_145__9_) );
AOI21X1 AOI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_7986_), .B(_3313__bF_buf56), .C(data_22__10_), .Y(_8005_) );
AOI21X1 AOI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf7), .B(_8003_), .C(_8005_), .Y(_145__10_) );
INVX1 INVX1_3495 ( .gnd(gnd), .vdd(vdd), .A(data_22__11_), .Y(_8006_) );
OAI21X1 OAI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf49), .B(_7991_), .C(_8006_), .Y(_8007_) );
NAND3X1 NAND3X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf8), .B(_7986_), .C(_3313__bF_buf55), .Y(_8008_) );
AND2X2 AND2X2_1447 ( .gnd(gnd), .vdd(vdd), .A(_8007_), .B(_8008_), .Y(_145__11_) );
INVX1 INVX1_3496 ( .gnd(gnd), .vdd(vdd), .A(data_22__12_), .Y(_8009_) );
OAI21X1 OAI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf48), .B(_7991_), .C(_8009_), .Y(_8010_) );
NAND3X1 NAND3X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf9), .B(_7986_), .C(_3313__bF_buf54), .Y(_8011_) );
AND2X2 AND2X2_1448 ( .gnd(gnd), .vdd(vdd), .A(_8010_), .B(_8011_), .Y(_145__12_) );
INVX1 INVX1_3497 ( .gnd(gnd), .vdd(vdd), .A(data_22__13_), .Y(_8012_) );
MUX2X1 MUX2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_8012_), .B(_14924__bF_buf6), .S(_7987_), .Y(_145__13_) );
INVX1 INVX1_3498 ( .gnd(gnd), .vdd(vdd), .A(data_22__14_), .Y(_8013_) );
MUX2X1 MUX2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_8013_), .B(_15060__bF_buf4), .S(_7987_), .Y(_145__14_) );
INVX1 INVX1_3499 ( .gnd(gnd), .vdd(vdd), .A(data_22__15_), .Y(_8014_) );
MUX2X1 MUX2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_8014_), .B(_15062__bF_buf9), .S(_7987_), .Y(_145__15_) );
INVX1 INVX1_3500 ( .gnd(gnd), .vdd(vdd), .A(data_21__0_), .Y(_8015_) );
AOI21X1 AOI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_14984__bF_buf1), .B(_911_), .C(_7983_), .Y(_8016_) );
NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_15179_), .B(_8016_), .Y(_8017_) );
NOR2X1 NOR2X1_834 ( .gnd(gnd), .vdd(vdd), .A(_8017_), .B(_5459__bF_buf0), .Y(_8018_) );
INVX4 INVX4_42 ( .gnd(gnd), .vdd(vdd), .A(_8018_), .Y(_8019_) );
OAI21X1 OAI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf47), .B(_8019_), .C(_8015_), .Y(_8020_) );
NAND3X1 NAND3X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_8018_), .C(_3313__bF_buf53), .Y(_8021_) );
AND2X2 AND2X2_1449 ( .gnd(gnd), .vdd(vdd), .A(_8020_), .B(_8021_), .Y(_134__0_) );
INVX1 INVX1_3501 ( .gnd(gnd), .vdd(vdd), .A(data_21__1_), .Y(_8022_) );
OAI21X1 OAI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf46), .B(_8019_), .C(_8022_), .Y(_8023_) );
NAND3X1 NAND3X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_8018_), .C(_3313__bF_buf52), .Y(_8024_) );
AND2X2 AND2X2_1450 ( .gnd(gnd), .vdd(vdd), .A(_8023_), .B(_8024_), .Y(_134__1_) );
INVX1 INVX1_3502 ( .gnd(gnd), .vdd(vdd), .A(data_21__2_), .Y(_8025_) );
NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_8018_), .B(_3313__bF_buf51), .Y(_8026_) );
MUX2X1 MUX2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_8025_), .B(_14897__bF_buf13), .S(_8026_), .Y(_134__2_) );
INVX1 INVX1_3503 ( .gnd(gnd), .vdd(vdd), .A(data_21__3_), .Y(_8027_) );
OAI21X1 OAI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf45), .B(_8019_), .C(_8027_), .Y(_8028_) );
NAND3X1 NAND3X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf3), .B(_8018_), .C(_3313__bF_buf50), .Y(_8029_) );
AND2X2 AND2X2_1451 ( .gnd(gnd), .vdd(vdd), .A(_8028_), .B(_8029_), .Y(_134__3_) );
INVX1 INVX1_3504 ( .gnd(gnd), .vdd(vdd), .A(data_21__4_), .Y(_8030_) );
OAI21X1 OAI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf44), .B(_8019_), .C(_8030_), .Y(_8031_) );
NAND3X1 NAND3X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_8018_), .C(_3313__bF_buf49), .Y(_8032_) );
AND2X2 AND2X2_1452 ( .gnd(gnd), .vdd(vdd), .A(_8031_), .B(_8032_), .Y(_134__4_) );
INVX1 INVX1_3505 ( .gnd(gnd), .vdd(vdd), .A(data_21__5_), .Y(_8033_) );
OAI21X1 OAI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf43), .B(_8019_), .C(_8033_), .Y(_8034_) );
NAND3X1 NAND3X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf6), .B(_8018_), .C(_3313__bF_buf48), .Y(_8035_) );
AND2X2 AND2X2_1453 ( .gnd(gnd), .vdd(vdd), .A(_8034_), .B(_8035_), .Y(_134__5_) );
INVX1 INVX1_3506 ( .gnd(gnd), .vdd(vdd), .A(data_21__6_), .Y(_8036_) );
MUX2X1 MUX2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_8036_), .B(_15049__bF_buf2), .S(_8026_), .Y(_134__6_) );
INVX1 INVX1_3507 ( .gnd(gnd), .vdd(vdd), .A(data_21__7_), .Y(_8037_) );
OAI21X1 OAI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf42), .B(_8019_), .C(_8037_), .Y(_8038_) );
NAND3X1 NAND3X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_8018_), .C(_3313__bF_buf47), .Y(_8039_) );
AND2X2 AND2X2_1454 ( .gnd(gnd), .vdd(vdd), .A(_8038_), .B(_8039_), .Y(_134__7_) );
INVX1 INVX1_3508 ( .gnd(gnd), .vdd(vdd), .A(data_21__8_), .Y(_8040_) );
MUX2X1 MUX2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_8040_), .B(_15052__bF_buf5), .S(_8026_), .Y(_134__8_) );
INVX1 INVX1_3509 ( .gnd(gnd), .vdd(vdd), .A(data_21__9_), .Y(_8041_) );
MUX2X1 MUX2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_8041_), .B(_14913__bF_buf14), .S(_8026_), .Y(_134__9_) );
INVX1 INVX1_3510 ( .gnd(gnd), .vdd(vdd), .A(data_21__10_), .Y(_8042_) );
MUX2X1 MUX2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_8042_), .B(_15055__bF_buf6), .S(_8026_), .Y(_134__10_) );
INVX1 INVX1_3511 ( .gnd(gnd), .vdd(vdd), .A(data_21__11_), .Y(_8043_) );
OAI21X1 OAI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf41), .B(_8019_), .C(_8043_), .Y(_8044_) );
NAND3X1 NAND3X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf7), .B(_8018_), .C(_3313__bF_buf46), .Y(_8045_) );
AND2X2 AND2X2_1455 ( .gnd(gnd), .vdd(vdd), .A(_8044_), .B(_8045_), .Y(_134__11_) );
INVX1 INVX1_3512 ( .gnd(gnd), .vdd(vdd), .A(data_21__12_), .Y(_8046_) );
OAI21X1 OAI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf40), .B(_8019_), .C(_8046_), .Y(_8047_) );
NAND3X1 NAND3X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf8), .B(_8018_), .C(_3313__bF_buf45), .Y(_8048_) );
AND2X2 AND2X2_1456 ( .gnd(gnd), .vdd(vdd), .A(_8047_), .B(_8048_), .Y(_134__12_) );
INVX1 INVX1_3513 ( .gnd(gnd), .vdd(vdd), .A(data_21__13_), .Y(_8049_) );
MUX2X1 MUX2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_8049_), .B(_14924__bF_buf5), .S(_8026_), .Y(_134__13_) );
INVX1 INVX1_3514 ( .gnd(gnd), .vdd(vdd), .A(data_21__14_), .Y(_8050_) );
MUX2X1 MUX2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_8050_), .B(_15060__bF_buf3), .S(_8026_), .Y(_134__14_) );
INVX1 INVX1_3515 ( .gnd(gnd), .vdd(vdd), .A(data_21__15_), .Y(_8051_) );
MUX2X1 MUX2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_8051_), .B(_15062__bF_buf8), .S(_8026_), .Y(_134__15_) );
INVX1 INVX1_3516 ( .gnd(gnd), .vdd(vdd), .A(data_20__0_), .Y(_8052_) );
INVX4 INVX4_43 ( .gnd(gnd), .vdd(vdd), .A(_15739_), .Y(_8053_) );
OAI21X1 OAI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf39), .B(_8053_), .C(_8052_), .Y(_8054_) );
NAND3X1 NAND3X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_15739_), .C(_3313__bF_buf44), .Y(_8055_) );
AND2X2 AND2X2_1457 ( .gnd(gnd), .vdd(vdd), .A(_8054_), .B(_8055_), .Y(_123__0_) );
INVX1 INVX1_3517 ( .gnd(gnd), .vdd(vdd), .A(data_20__1_), .Y(_8056_) );
OAI21X1 OAI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf38), .B(_8053_), .C(_8056_), .Y(_8057_) );
NAND3X1 NAND3X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_15739_), .C(_3313__bF_buf43), .Y(_8058_) );
AND2X2 AND2X2_1458 ( .gnd(gnd), .vdd(vdd), .A(_8057_), .B(_8058_), .Y(_123__1_) );
INVX1 INVX1_3518 ( .gnd(gnd), .vdd(vdd), .A(data_20__2_), .Y(_8059_) );
NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_15739_), .B(_3313__bF_buf42), .Y(_8060_) );
MUX2X1 MUX2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_8059_), .B(_14897__bF_buf12), .S(_8060_), .Y(_123__2_) );
INVX1 INVX1_3519 ( .gnd(gnd), .vdd(vdd), .A(data_20__3_), .Y(_8061_) );
MUX2X1 MUX2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8061_), .B(_14899__bF_buf2), .S(_8060_), .Y(_123__3_) );
INVX1 INVX1_3520 ( .gnd(gnd), .vdd(vdd), .A(data_20__4_), .Y(_8062_) );
OAI21X1 OAI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf37), .B(_8053_), .C(_8062_), .Y(_8063_) );
NAND3X1 NAND3X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_15739_), .C(_3313__bF_buf41), .Y(_8064_) );
AND2X2 AND2X2_1459 ( .gnd(gnd), .vdd(vdd), .A(_8063_), .B(_8064_), .Y(_123__4_) );
INVX1 INVX1_3521 ( .gnd(gnd), .vdd(vdd), .A(data_20__5_), .Y(_8065_) );
OAI21X1 OAI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf36), .B(_8053_), .C(_8065_), .Y(_8066_) );
NAND3X1 NAND3X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_15739_), .C(_3313__bF_buf40), .Y(_8067_) );
AND2X2 AND2X2_1460 ( .gnd(gnd), .vdd(vdd), .A(_8066_), .B(_8067_), .Y(_123__5_) );
INVX1 INVX1_3522 ( .gnd(gnd), .vdd(vdd), .A(data_20__6_), .Y(_8068_) );
MUX2X1 MUX2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_8068_), .B(_15049__bF_buf1), .S(_8060_), .Y(_123__6_) );
INVX1 INVX1_3523 ( .gnd(gnd), .vdd(vdd), .A(data_20__7_), .Y(_8069_) );
OAI21X1 OAI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf35), .B(_8053_), .C(_8069_), .Y(_8070_) );
NAND3X1 NAND3X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_15739_), .C(_3313__bF_buf39), .Y(_8071_) );
AND2X2 AND2X2_1461 ( .gnd(gnd), .vdd(vdd), .A(_8070_), .B(_8071_), .Y(_123__7_) );
INVX1 INVX1_3524 ( .gnd(gnd), .vdd(vdd), .A(data_20__8_), .Y(_8072_) );
MUX2X1 MUX2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_8072_), .B(_15052__bF_buf4), .S(_8060_), .Y(_123__8_) );
INVX1 INVX1_3525 ( .gnd(gnd), .vdd(vdd), .A(data_20__9_), .Y(_8073_) );
MUX2X1 MUX2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_8073_), .B(_14913__bF_buf13), .S(_8060_), .Y(_123__9_) );
INVX1 INVX1_3526 ( .gnd(gnd), .vdd(vdd), .A(data_20__10_), .Y(_8074_) );
MUX2X1 MUX2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_8074_), .B(_15055__bF_buf5), .S(_8060_), .Y(_123__10_) );
INVX1 INVX1_3527 ( .gnd(gnd), .vdd(vdd), .A(data_20__11_), .Y(_8075_) );
MUX2X1 MUX2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_8075_), .B(_14918__bF_buf6), .S(_8060_), .Y(_123__11_) );
INVX1 INVX1_3528 ( .gnd(gnd), .vdd(vdd), .A(data_20__12_), .Y(_8076_) );
OAI21X1 OAI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_3393__bF_buf34), .B(_8053_), .C(_8076_), .Y(_8077_) );
NAND3X1 NAND3X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_15739_), .C(_3313__bF_buf38), .Y(_8078_) );
AND2X2 AND2X2_1462 ( .gnd(gnd), .vdd(vdd), .A(_8077_), .B(_8078_), .Y(_123__12_) );
NOR2X1 NOR2X1_835 ( .gnd(gnd), .vdd(vdd), .A(_8053_), .B(_3393__bF_buf33), .Y(_8079_) );
AOI21X1 AOI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_15739_), .B(_3313__bF_buf37), .C(data_20__13_), .Y(_8080_) );
AOI21X1 AOI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_8079_), .C(_8080_), .Y(_123__13_) );
INVX1 INVX1_3529 ( .gnd(gnd), .vdd(vdd), .A(data_20__14_), .Y(_8081_) );
MUX2X1 MUX2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_8081_), .B(_15060__bF_buf2), .S(_8060_), .Y(_123__14_) );
INVX1 INVX1_3530 ( .gnd(gnd), .vdd(vdd), .A(data_20__15_), .Y(_8082_) );
MUX2X1 MUX2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_8082_), .B(_15062__bF_buf7), .S(_8060_), .Y(_123__15_) );
INVX1 INVX1_3531 ( .gnd(gnd), .vdd(vdd), .A(data_19__0_), .Y(_8083_) );
INVX4 INVX4_44 ( .gnd(gnd), .vdd(vdd), .A(_3309_), .Y(_8084_) );
OAI21X1 OAI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_15034_), .B(_15031__bF_buf1), .C(IDATA_PROG_write_bF_buf5), .Y(_8085_) );
AOI21X1 AOI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_14963__bF_buf1), .B(_15011__bF_buf0), .C(_8085_), .Y(_8086_) );
OAI21X1 OAI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_7507_), .B(_15175__bF_buf4), .C(_8086_), .Y(_8087_) );
NOR3X1 NOR3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8087_), .C(_15074__bF_buf0), .Y(_8088_) );
NAND3X1 NAND3X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_8088_), .C(_3391__bF_buf5), .Y(_8089_) );
MUX2X1 MUX2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_8083_), .B(_14932__bF_buf2), .S(_8089_), .Y(_111__0_) );
INVX1 INVX1_3532 ( .gnd(gnd), .vdd(vdd), .A(data_19__1_), .Y(_8090_) );
MUX2X1 MUX2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_8090_), .B(_14894__bF_buf0), .S(_8089_), .Y(_111__1_) );
INVX1 INVX1_3533 ( .gnd(gnd), .vdd(vdd), .A(data_19__2_), .Y(_8091_) );
MUX2X1 MUX2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_8091_), .B(_14897__bF_buf11), .S(_8089_), .Y(_111__2_) );
INVX1 INVX1_3534 ( .gnd(gnd), .vdd(vdd), .A(data_19__3_), .Y(_8092_) );
MUX2X1 MUX2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_8092_), .B(_14899__bF_buf1), .S(_8089_), .Y(_111__3_) );
INVX1 INVX1_3535 ( .gnd(gnd), .vdd(vdd), .A(data_19__4_), .Y(_8093_) );
MUX2X1 MUX2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_8093_), .B(_14902__bF_buf5), .S(_8089_), .Y(_111__4_) );
INVX1 INVX1_3536 ( .gnd(gnd), .vdd(vdd), .A(data_19__5_), .Y(_8094_) );
MUX2X1 MUX2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_8094_), .B(_14903__bF_buf4), .S(_8089_), .Y(_111__5_) );
INVX1 INVX1_3537 ( .gnd(gnd), .vdd(vdd), .A(data_19__6_), .Y(_8095_) );
MUX2X1 MUX2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_8095_), .B(_15049__bF_buf0), .S(_8089_), .Y(_111__6_) );
INVX1 INVX1_3538 ( .gnd(gnd), .vdd(vdd), .A(data_19__7_), .Y(_8096_) );
MUX2X1 MUX2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_8096_), .B(_14908__bF_buf6), .S(_8089_), .Y(_111__7_) );
INVX1 INVX1_3539 ( .gnd(gnd), .vdd(vdd), .A(data_19__8_), .Y(_8097_) );
MUX2X1 MUX2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_8097_), .B(_15052__bF_buf3), .S(_8089_), .Y(_111__8_) );
INVX1 INVX1_3540 ( .gnd(gnd), .vdd(vdd), .A(data_19__9_), .Y(_8098_) );
MUX2X1 MUX2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_8098_), .B(_14913__bF_buf12), .S(_8089_), .Y(_111__9_) );
INVX1 INVX1_3541 ( .gnd(gnd), .vdd(vdd), .A(data_19__10_), .Y(_8099_) );
MUX2X1 MUX2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_8099_), .B(_15055__bF_buf4), .S(_8089_), .Y(_111__10_) );
INVX1 INVX1_3542 ( .gnd(gnd), .vdd(vdd), .A(data_19__11_), .Y(_8100_) );
MUX2X1 MUX2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_8100_), .B(_14918__bF_buf5), .S(_8089_), .Y(_111__11_) );
INVX1 INVX1_3543 ( .gnd(gnd), .vdd(vdd), .A(data_19__12_), .Y(_8101_) );
MUX2X1 MUX2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_8101_), .B(_14920__bF_buf6), .S(_8089_), .Y(_111__12_) );
INVX1 INVX1_3544 ( .gnd(gnd), .vdd(vdd), .A(data_19__13_), .Y(_8102_) );
MUX2X1 MUX2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_8102_), .B(_14924__bF_buf3), .S(_8089_), .Y(_111__13_) );
INVX1 INVX1_3545 ( .gnd(gnd), .vdd(vdd), .A(data_19__14_), .Y(_8103_) );
MUX2X1 MUX2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_8103_), .B(_15060__bF_buf1), .S(_8089_), .Y(_111__14_) );
INVX1 INVX1_3546 ( .gnd(gnd), .vdd(vdd), .A(data_19__15_), .Y(_8104_) );
MUX2X1 MUX2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_8104_), .B(_15062__bF_buf6), .S(_8089_), .Y(_111__15_) );
INVX1 INVX1_3547 ( .gnd(gnd), .vdd(vdd), .A(data_18__0_), .Y(_8105_) );
OAI21X1 OAI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_7538_), .B(_15175__bF_buf3), .C(_8086_), .Y(_8106_) );
NOR3X1 NOR3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8106_), .C(_15074__bF_buf12), .Y(_8107_) );
NAND3X1 NAND3X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_8107_), .C(_3391__bF_buf4), .Y(_8108_) );
MUX2X1 MUX2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_8105_), .B(_14932__bF_buf1), .S(_8108_), .Y(_100__0_) );
INVX1 INVX1_3548 ( .gnd(gnd), .vdd(vdd), .A(data_18__1_), .Y(_8109_) );
MUX2X1 MUX2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_8109_), .B(_14894__bF_buf14), .S(_8108_), .Y(_100__1_) );
INVX1 INVX1_3549 ( .gnd(gnd), .vdd(vdd), .A(data_18__2_), .Y(_8110_) );
MUX2X1 MUX2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_8110_), .B(_14897__bF_buf10), .S(_8108_), .Y(_100__2_) );
INVX1 INVX1_3550 ( .gnd(gnd), .vdd(vdd), .A(data_18__3_), .Y(_8111_) );
MUX2X1 MUX2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_8111_), .B(_14899__bF_buf0), .S(_8108_), .Y(_100__3_) );
INVX1 INVX1_3551 ( .gnd(gnd), .vdd(vdd), .A(data_18__4_), .Y(_8112_) );
MUX2X1 MUX2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_8112_), .B(_14902__bF_buf4), .S(_8108_), .Y(_100__4_) );
INVX1 INVX1_3552 ( .gnd(gnd), .vdd(vdd), .A(data_18__5_), .Y(_8113_) );
MUX2X1 MUX2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_8113_), .B(_14903__bF_buf3), .S(_8108_), .Y(_100__5_) );
INVX1 INVX1_3553 ( .gnd(gnd), .vdd(vdd), .A(data_18__6_), .Y(_8114_) );
MUX2X1 MUX2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_8114_), .B(_15049__bF_buf14), .S(_8108_), .Y(_100__6_) );
INVX1 INVX1_3554 ( .gnd(gnd), .vdd(vdd), .A(data_18__7_), .Y(_8115_) );
MUX2X1 MUX2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_8115_), .B(_14908__bF_buf5), .S(_8108_), .Y(_100__7_) );
INVX1 INVX1_3555 ( .gnd(gnd), .vdd(vdd), .A(data_18__8_), .Y(_8116_) );
MUX2X1 MUX2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_8116_), .B(_15052__bF_buf2), .S(_8108_), .Y(_100__8_) );
INVX1 INVX1_3556 ( .gnd(gnd), .vdd(vdd), .A(data_18__9_), .Y(_8117_) );
MUX2X1 MUX2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_8117_), .B(_14913__bF_buf11), .S(_8108_), .Y(_100__9_) );
INVX1 INVX1_3557 ( .gnd(gnd), .vdd(vdd), .A(data_18__10_), .Y(_8118_) );
MUX2X1 MUX2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_8118_), .B(_15055__bF_buf3), .S(_8108_), .Y(_100__10_) );
INVX1 INVX1_3558 ( .gnd(gnd), .vdd(vdd), .A(data_18__11_), .Y(_8119_) );
MUX2X1 MUX2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_8119_), .B(_14918__bF_buf4), .S(_8108_), .Y(_100__11_) );
INVX1 INVX1_3559 ( .gnd(gnd), .vdd(vdd), .A(data_18__12_), .Y(_8120_) );
MUX2X1 MUX2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_8120_), .B(_14920__bF_buf5), .S(_8108_), .Y(_100__12_) );
INVX1 INVX1_3560 ( .gnd(gnd), .vdd(vdd), .A(data_18__13_), .Y(_8121_) );
MUX2X1 MUX2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_8121_), .B(_14924__bF_buf2), .S(_8108_), .Y(_100__13_) );
INVX1 INVX1_3561 ( .gnd(gnd), .vdd(vdd), .A(data_18__14_), .Y(_8122_) );
MUX2X1 MUX2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_8122_), .B(_15060__bF_buf0), .S(_8108_), .Y(_100__14_) );
INVX1 INVX1_3562 ( .gnd(gnd), .vdd(vdd), .A(data_18__15_), .Y(_8123_) );
MUX2X1 MUX2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_8123_), .B(_15062__bF_buf5), .S(_8108_), .Y(_100__15_) );
INVX1 INVX1_3563 ( .gnd(gnd), .vdd(vdd), .A(data_17__0_), .Y(_8124_) );
NOR2X1 NOR2X1_836 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_3306__bF_buf5), .Y(_8125_) );
NAND3X1 NAND3X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_15001_), .B(_3309_), .C(_14973_), .Y(_8126_) );
OAI21X1 OAI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_15175__bF_buf2), .B(_7575_), .C(_8086_), .Y(_8127_) );
NOR2X1 NOR2X1_837 ( .gnd(gnd), .vdd(vdd), .A(_8127_), .B(_8126_), .Y(_8128_) );
NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_8128_), .B(_8125__bF_buf5), .Y(_8129_) );
MUX2X1 MUX2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_8124_), .B(_14932__bF_buf0), .S(_8129_), .Y(_89__0_) );
INVX1 INVX1_3564 ( .gnd(gnd), .vdd(vdd), .A(data_17__1_), .Y(_8130_) );
MUX2X1 MUX2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_8130_), .B(_14894__bF_buf13), .S(_8129_), .Y(_89__1_) );
INVX1 INVX1_3565 ( .gnd(gnd), .vdd(vdd), .A(data_17__2_), .Y(_8131_) );
MUX2X1 MUX2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_8131_), .B(_14897__bF_buf9), .S(_8129_), .Y(_89__2_) );
INVX1 INVX1_3566 ( .gnd(gnd), .vdd(vdd), .A(data_17__3_), .Y(_8132_) );
MUX2X1 MUX2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_8132_), .B(_14899__bF_buf14), .S(_8129_), .Y(_89__3_) );
INVX1 INVX1_3567 ( .gnd(gnd), .vdd(vdd), .A(data_17__4_), .Y(_8133_) );
MUX2X1 MUX2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_8133_), .B(_14902__bF_buf3), .S(_8129_), .Y(_89__4_) );
INVX1 INVX1_3568 ( .gnd(gnd), .vdd(vdd), .A(data_17__5_), .Y(_8134_) );
MUX2X1 MUX2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_8134_), .B(_14903__bF_buf2), .S(_8129_), .Y(_89__5_) );
INVX1 INVX1_3569 ( .gnd(gnd), .vdd(vdd), .A(data_17__6_), .Y(_8135_) );
MUX2X1 MUX2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_8135_), .B(_15049__bF_buf13), .S(_8129_), .Y(_89__6_) );
INVX1 INVX1_3570 ( .gnd(gnd), .vdd(vdd), .A(data_17__7_), .Y(_8136_) );
MUX2X1 MUX2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_8136_), .B(_14908__bF_buf4), .S(_8129_), .Y(_89__7_) );
INVX1 INVX1_3571 ( .gnd(gnd), .vdd(vdd), .A(data_17__8_), .Y(_8137_) );
MUX2X1 MUX2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_8137_), .B(_15052__bF_buf1), .S(_8129_), .Y(_89__8_) );
INVX1 INVX1_3572 ( .gnd(gnd), .vdd(vdd), .A(data_17__9_), .Y(_8138_) );
MUX2X1 MUX2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_8138_), .B(_14913__bF_buf10), .S(_8129_), .Y(_89__9_) );
INVX1 INVX1_3573 ( .gnd(gnd), .vdd(vdd), .A(data_17__10_), .Y(_8139_) );
MUX2X1 MUX2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_8139_), .B(_15055__bF_buf2), .S(_8129_), .Y(_89__10_) );
INVX1 INVX1_3574 ( .gnd(gnd), .vdd(vdd), .A(data_17__11_), .Y(_8140_) );
MUX2X1 MUX2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_8140_), .B(_14918__bF_buf3), .S(_8129_), .Y(_89__11_) );
INVX1 INVX1_3575 ( .gnd(gnd), .vdd(vdd), .A(data_17__12_), .Y(_8141_) );
MUX2X1 MUX2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_8141_), .B(_14920__bF_buf4), .S(_8129_), .Y(_89__12_) );
INVX1 INVX1_3576 ( .gnd(gnd), .vdd(vdd), .A(data_17__13_), .Y(_8142_) );
MUX2X1 MUX2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_8142_), .B(_14924__bF_buf1), .S(_8129_), .Y(_89__13_) );
INVX1 INVX1_3577 ( .gnd(gnd), .vdd(vdd), .A(data_17__14_), .Y(_8143_) );
MUX2X1 MUX2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_8143_), .B(_15060__bF_buf14), .S(_8129_), .Y(_89__14_) );
INVX1 INVX1_3578 ( .gnd(gnd), .vdd(vdd), .A(data_17__15_), .Y(_8144_) );
MUX2X1 MUX2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_8144_), .B(_15062__bF_buf4), .S(_8129_), .Y(_89__15_) );
NAND3X1 NAND3X1_1070 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf4), .B(_14986_), .C(_14984__bF_buf0), .Y(_8145_) );
INVX1 INVX1_3579 ( .gnd(gnd), .vdd(vdd), .A(data_16__0_), .Y(_8146_) );
NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_8146_), .B(_8145__bF_buf3), .Y(_8147_) );
OAI21X1 OAI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_0_bF_buf4), .B(_8145__bF_buf2), .C(_8147_), .Y(_8148_) );
INVX1 INVX1_3580 ( .gnd(gnd), .vdd(vdd), .A(_8148_), .Y(_78__0_) );
INVX4 INVX4_45 ( .gnd(gnd), .vdd(vdd), .A(_8145__bF_buf1), .Y(_8149_) );
OR2X2 OR2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_8149_), .B(data_16__1_), .Y(_8150_) );
OAI21X1 OAI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf1), .B(_8145__bF_buf0), .C(_8150_), .Y(_8151_) );
INVX1 INVX1_3581 ( .gnd(gnd), .vdd(vdd), .A(_8151_), .Y(_78__1_) );
NOR2X1 NOR2X1_838 ( .gnd(gnd), .vdd(vdd), .A(data_16__2_), .B(_8149_), .Y(_8152_) );
AOI21X1 AOI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_8149_), .C(_8152_), .Y(_78__2_) );
NOR2X1 NOR2X1_839 ( .gnd(gnd), .vdd(vdd), .A(data_16__3_), .B(_8149_), .Y(_8153_) );
AOI21X1 AOI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_8149_), .C(_8153_), .Y(_78__3_) );
OR2X2 OR2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_8149_), .B(data_16__4_), .Y(_8154_) );
OAI21X1 OAI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf1), .B(_8145__bF_buf3), .C(_8154_), .Y(_8155_) );
INVX1 INVX1_3582 ( .gnd(gnd), .vdd(vdd), .A(_8155_), .Y(_78__4_) );
INVX1 INVX1_3583 ( .gnd(gnd), .vdd(vdd), .A(data_16__5_), .Y(_8156_) );
NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_8156_), .B(_8145__bF_buf2), .Y(_8157_) );
OAI21X1 OAI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf2), .B(_8145__bF_buf1), .C(_8157_), .Y(_8158_) );
INVX1 INVX1_3584 ( .gnd(gnd), .vdd(vdd), .A(_8158_), .Y(_78__5_) );
INVX1 INVX1_3585 ( .gnd(gnd), .vdd(vdd), .A(data_16__6_), .Y(_8159_) );
NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_8159_), .B(_8145__bF_buf0), .Y(_8160_) );
OAI21X1 OAI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf1), .B(_8145__bF_buf3), .C(_8160_), .Y(_8161_) );
INVX1 INVX1_3586 ( .gnd(gnd), .vdd(vdd), .A(_8161_), .Y(_78__6_) );
INVX1 INVX1_3587 ( .gnd(gnd), .vdd(vdd), .A(data_16__7_), .Y(_8162_) );
NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_8162_), .B(_8145__bF_buf2), .Y(_8163_) );
OAI21X1 OAI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf1), .B(_8145__bF_buf1), .C(_8163_), .Y(_8164_) );
INVX1 INVX1_3588 ( .gnd(gnd), .vdd(vdd), .A(_8164_), .Y(_78__7_) );
INVX1 INVX1_3589 ( .gnd(gnd), .vdd(vdd), .A(data_16__8_), .Y(_8165_) );
NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_8165_), .B(_8145__bF_buf0), .Y(_8166_) );
OAI21X1 OAI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf3), .B(_8145__bF_buf3), .C(_8166_), .Y(_8167_) );
INVX1 INVX1_3590 ( .gnd(gnd), .vdd(vdd), .A(_8167_), .Y(_78__8_) );
INVX1 INVX1_3591 ( .gnd(gnd), .vdd(vdd), .A(data_16__9_), .Y(_8168_) );
NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_8168_), .B(_8145__bF_buf2), .Y(_8169_) );
OAI21X1 OAI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf4), .B(_8145__bF_buf1), .C(_8169_), .Y(_8170_) );
INVX1 INVX1_3592 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .Y(_78__9_) );
INVX1 INVX1_3593 ( .gnd(gnd), .vdd(vdd), .A(data_16__10_), .Y(_8171_) );
NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_8171_), .B(_8145__bF_buf0), .Y(_8172_) );
OAI21X1 OAI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf2), .B(_8145__bF_buf3), .C(_8172_), .Y(_8173_) );
INVX1 INVX1_3594 ( .gnd(gnd), .vdd(vdd), .A(_8173_), .Y(_78__10_) );
INVX1 INVX1_3595 ( .gnd(gnd), .vdd(vdd), .A(data_16__11_), .Y(_8174_) );
NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_8174_), .B(_8145__bF_buf2), .Y(_8175_) );
OAI21X1 OAI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_11_bF_buf1), .B(_8145__bF_buf1), .C(_8175_), .Y(_8176_) );
INVX1 INVX1_3596 ( .gnd(gnd), .vdd(vdd), .A(_8176_), .Y(_78__11_) );
OR2X2 OR2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_8149_), .B(data_16__12_), .Y(_8177_) );
OAI21X1 OAI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_12_bF_buf0), .B(_8145__bF_buf0), .C(_8177_), .Y(_8178_) );
INVX1 INVX1_3597 ( .gnd(gnd), .vdd(vdd), .A(_8178_), .Y(_78__12_) );
NOR2X1 NOR2X1_840 ( .gnd(gnd), .vdd(vdd), .A(data_16__13_), .B(_8149_), .Y(_8179_) );
NOR2X1 NOR2X1_841 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf3), .B(_8145__bF_buf3), .Y(_8180_) );
NOR2X1 NOR2X1_842 ( .gnd(gnd), .vdd(vdd), .A(_8180_), .B(_8179_), .Y(_78__13_) );
NOR2X1 NOR2X1_843 ( .gnd(gnd), .vdd(vdd), .A(data_16__14_), .B(_8149_), .Y(_8181_) );
NOR2X1 NOR2X1_844 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf0), .B(_8145__bF_buf2), .Y(_8182_) );
NOR2X1 NOR2X1_845 ( .gnd(gnd), .vdd(vdd), .A(_8182_), .B(_8181_), .Y(_78__14_) );
INVX1 INVX1_3598 ( .gnd(gnd), .vdd(vdd), .A(data_16__15_), .Y(_8183_) );
NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_8183_), .B(_8145__bF_buf1), .Y(_8184_) );
OAI21X1 OAI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf1), .B(_8145__bF_buf0), .C(_8184_), .Y(_8185_) );
INVX1 INVX1_3599 ( .gnd(gnd), .vdd(vdd), .A(_8185_), .Y(_78__15_) );
INVX1 INVX1_3600 ( .gnd(gnd), .vdd(vdd), .A(data_15__0_), .Y(_8186_) );
NAND3X1 NAND3X1_1071 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf3), .B(_14888__bF_buf3), .C(_15011__bF_buf3), .Y(_8187_) );
MUX2X1 MUX2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_8186_), .B(_14932__bF_buf14), .S(_8187_), .Y(_67__0_) );
INVX4 INVX4_46 ( .gnd(gnd), .vdd(vdd), .A(_8187_), .Y(_8188_) );
NOR2X1 NOR2X1_846 ( .gnd(gnd), .vdd(vdd), .A(data_15__1_), .B(_8188_), .Y(_8189_) );
AOI21X1 AOI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf12), .B(_8188_), .C(_8189_), .Y(_67__1_) );
INVX1 INVX1_3601 ( .gnd(gnd), .vdd(vdd), .A(data_15__2_), .Y(_8190_) );
NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_14888__bF_buf2), .B(_15011__bF_buf2), .Y(_8191_) );
OAI21X1 OAI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_14882__bF_buf10), .C(_8190_), .Y(_8192_) );
NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf7), .B(_8188_), .Y(_8193_) );
AND2X2 AND2X2_1463 ( .gnd(gnd), .vdd(vdd), .A(_8193_), .B(_8192_), .Y(_67__2_) );
INVX1 INVX1_3602 ( .gnd(gnd), .vdd(vdd), .A(data_15__3_), .Y(_8194_) );
MUX2X1 MUX2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_8194_), .B(_14899__bF_buf12), .S(_8187_), .Y(_67__3_) );
INVX1 INVX1_3603 ( .gnd(gnd), .vdd(vdd), .A(data_15__4_), .Y(_8195_) );
MUX2X1 MUX2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_8195_), .B(_14902__bF_buf2), .S(_8187_), .Y(_67__4_) );
INVX1 INVX1_3604 ( .gnd(gnd), .vdd(vdd), .A(data_15__5_), .Y(_8196_) );
MUX2X1 MUX2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_8196_), .B(_14903__bF_buf1), .S(_8187_), .Y(_67__5_) );
INVX1 INVX1_3605 ( .gnd(gnd), .vdd(vdd), .A(data_15__6_), .Y(_8197_) );
MUX2X1 MUX2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_8197_), .B(_15049__bF_buf12), .S(_8187_), .Y(_67__6_) );
INVX1 INVX1_3606 ( .gnd(gnd), .vdd(vdd), .A(data_15__7_), .Y(_8198_) );
MUX2X1 MUX2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_8198_), .B(_14908__bF_buf3), .S(_8187_), .Y(_67__7_) );
INVX1 INVX1_3607 ( .gnd(gnd), .vdd(vdd), .A(data_15__8_), .Y(_8199_) );
OAI21X1 OAI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_14882__bF_buf9), .C(_8199_), .Y(_8200_) );
NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_8188_), .Y(_8201_) );
AND2X2 AND2X2_1464 ( .gnd(gnd), .vdd(vdd), .A(_8201_), .B(_8200_), .Y(_67__8_) );
NOR2X1 NOR2X1_847 ( .gnd(gnd), .vdd(vdd), .A(data_15__9_), .B(_8188_), .Y(_8202_) );
AOI21X1 AOI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf9), .B(_8188_), .C(_8202_), .Y(_67__9_) );
INVX1 INVX1_3608 ( .gnd(gnd), .vdd(vdd), .A(data_15__10_), .Y(_8203_) );
OAI21X1 OAI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_14882__bF_buf8), .C(_8203_), .Y(_8204_) );
NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_8188_), .Y(_8205_) );
AND2X2 AND2X2_1465 ( .gnd(gnd), .vdd(vdd), .A(_8205_), .B(_8204_), .Y(_67__10_) );
INVX1 INVX1_3609 ( .gnd(gnd), .vdd(vdd), .A(data_15__11_), .Y(_8206_) );
MUX2X1 MUX2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_8206_), .B(_14918__bF_buf2), .S(_8187_), .Y(_67__11_) );
INVX1 INVX1_3610 ( .gnd(gnd), .vdd(vdd), .A(data_15__12_), .Y(_8207_) );
OAI21X1 OAI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_14882__bF_buf7), .C(_8207_), .Y(_8208_) );
NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_8188_), .Y(_8209_) );
AND2X2 AND2X2_1466 ( .gnd(gnd), .vdd(vdd), .A(_8209_), .B(_8208_), .Y(_67__12_) );
INVX1 INVX1_3611 ( .gnd(gnd), .vdd(vdd), .A(data_15__13_), .Y(_8210_) );
OAI21X1 OAI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_8191_), .B(_14882__bF_buf6), .C(_8210_), .Y(_8211_) );
NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf0), .B(_8188_), .Y(_8212_) );
AND2X2 AND2X2_1467 ( .gnd(gnd), .vdd(vdd), .A(_8212_), .B(_8211_), .Y(_67__13_) );
INVX1 INVX1_3612 ( .gnd(gnd), .vdd(vdd), .A(data_15__14_), .Y(_8213_) );
MUX2X1 MUX2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_8213_), .B(_15060__bF_buf13), .S(_8187_), .Y(_67__14_) );
INVX1 INVX1_3613 ( .gnd(gnd), .vdd(vdd), .A(data_15__15_), .Y(_8214_) );
MUX2X1 MUX2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_8214_), .B(_15062__bF_buf3), .S(_8187_), .Y(_67__15_) );
INVX1 INVX1_3614 ( .gnd(gnd), .vdd(vdd), .A(data_14__0_), .Y(_8215_) );
NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_15011__bF_buf1), .B(_15793__bF_buf1), .Y(_8216_) );
MUX2X1 MUX2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_8215_), .B(_14932__bF_buf13), .S(_8216_), .Y(_56__0_) );
INVX1 INVX1_3615 ( .gnd(gnd), .vdd(vdd), .A(data_14__1_), .Y(_8217_) );
OAI21X1 OAI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15031__bF_buf0), .C(_8217_), .Y(_8218_) );
NAND3X1 NAND3X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf11), .B(_15011__bF_buf0), .C(_15793__bF_buf0), .Y(_8219_) );
AND2X2 AND2X2_1468 ( .gnd(gnd), .vdd(vdd), .A(_8218_), .B(_8219_), .Y(_56__1_) );
NOR2X1 NOR2X1_848 ( .gnd(gnd), .vdd(vdd), .A(_15031__bF_buf3), .B(_15788__bF_buf1), .Y(_8220_) );
NOR2X1 NOR2X1_849 ( .gnd(gnd), .vdd(vdd), .A(data_14__2_), .B(_8220_), .Y(_8221_) );
AOI21X1 AOI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf6), .B(_8220_), .C(_8221_), .Y(_56__2_) );
NOR2X1 NOR2X1_850 ( .gnd(gnd), .vdd(vdd), .A(data_14__3_), .B(_8220_), .Y(_8222_) );
AOI21X1 AOI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf11), .B(_8220_), .C(_8222_), .Y(_56__3_) );
INVX1 INVX1_3616 ( .gnd(gnd), .vdd(vdd), .A(data_14__4_), .Y(_8223_) );
OAI21X1 OAI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15031__bF_buf2), .C(_8223_), .Y(_8224_) );
OAI21X1 OAI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_4_bF_buf0), .B(_8216_), .C(_8224_), .Y(_8225_) );
INVX1 INVX1_3617 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .Y(_56__4_) );
INVX1 INVX1_3618 ( .gnd(gnd), .vdd(vdd), .A(data_14__5_), .Y(_8226_) );
OAI21X1 OAI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf9), .B(_15031__bF_buf1), .C(_8226_), .Y(_8227_) );
NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf0), .B(_8220_), .Y(_8228_) );
AND2X2 AND2X2_1469 ( .gnd(gnd), .vdd(vdd), .A(_8228_), .B(_8227_), .Y(_56__5_) );
INVX1 INVX1_3619 ( .gnd(gnd), .vdd(vdd), .A(data_14__6_), .Y(_8229_) );
OAI21X1 OAI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf8), .B(_15031__bF_buf0), .C(_8229_), .Y(_8230_) );
NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf11), .B(_8220_), .Y(_8231_) );
AND2X2 AND2X2_1470 ( .gnd(gnd), .vdd(vdd), .A(_8231_), .B(_8230_), .Y(_56__6_) );
INVX1 INVX1_3620 ( .gnd(gnd), .vdd(vdd), .A(data_14__7_), .Y(_8232_) );
OAI21X1 OAI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf7), .B(_15031__bF_buf3), .C(_8232_), .Y(_8233_) );
OAI21X1 OAI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_7_bF_buf0), .B(_8216_), .C(_8233_), .Y(_8234_) );
INVX1 INVX1_3621 ( .gnd(gnd), .vdd(vdd), .A(_8234_), .Y(_56__7_) );
INVX1 INVX1_3622 ( .gnd(gnd), .vdd(vdd), .A(data_14__8_), .Y(_8235_) );
OAI21X1 OAI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf6), .B(_15031__bF_buf2), .C(_8235_), .Y(_8236_) );
NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf13), .B(_8220_), .Y(_8237_) );
AND2X2 AND2X2_1471 ( .gnd(gnd), .vdd(vdd), .A(_8237_), .B(_8236_), .Y(_56__8_) );
NOR2X1 NOR2X1_851 ( .gnd(gnd), .vdd(vdd), .A(data_14__9_), .B(_8220_), .Y(_8238_) );
AOI21X1 AOI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf8), .B(_8220_), .C(_8238_), .Y(_56__9_) );
INVX1 INVX1_3623 ( .gnd(gnd), .vdd(vdd), .A(data_14__10_), .Y(_8239_) );
OAI21X1 OAI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf5), .B(_15031__bF_buf1), .C(_8239_), .Y(_8240_) );
NAND3X1 NAND3X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf0), .B(_15011__bF_buf3), .C(_15793__bF_buf5), .Y(_8241_) );
AND2X2 AND2X2_1472 ( .gnd(gnd), .vdd(vdd), .A(_8240_), .B(_8241_), .Y(_56__10_) );
INVX1 INVX1_3624 ( .gnd(gnd), .vdd(vdd), .A(data_14__11_), .Y(_8242_) );
OAI21X1 OAI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf4), .B(_15031__bF_buf0), .C(_8242_), .Y(_8243_) );
NAND3X1 NAND3X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf1), .B(_15011__bF_buf2), .C(_15793__bF_buf4), .Y(_8244_) );
AND2X2 AND2X2_1473 ( .gnd(gnd), .vdd(vdd), .A(_8243_), .B(_8244_), .Y(_56__11_) );
INVX1 INVX1_3625 ( .gnd(gnd), .vdd(vdd), .A(data_14__12_), .Y(_8245_) );
OAI21X1 OAI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf3), .B(_15031__bF_buf3), .C(_8245_), .Y(_8246_) );
NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf2), .B(_8220_), .Y(_8247_) );
AND2X2 AND2X2_1474 ( .gnd(gnd), .vdd(vdd), .A(_8247_), .B(_8246_), .Y(_56__12_) );
INVX1 INVX1_3626 ( .gnd(gnd), .vdd(vdd), .A(data_14__13_), .Y(_8248_) );
OAI21X1 OAI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf2), .B(_15031__bF_buf2), .C(_8248_), .Y(_8249_) );
OAI21X1 OAI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_13_bF_buf2), .B(_8216_), .C(_8249_), .Y(_8250_) );
INVX1 INVX1_3627 ( .gnd(gnd), .vdd(vdd), .A(_8250_), .Y(_56__13_) );
INVX1 INVX1_3628 ( .gnd(gnd), .vdd(vdd), .A(data_14__14_), .Y(_8251_) );
OAI21X1 OAI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf1), .B(_15031__bF_buf1), .C(_8251_), .Y(_8252_) );
OAI21X1 OAI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf4), .B(_8216_), .C(_8252_), .Y(_8253_) );
INVX1 INVX1_3629 ( .gnd(gnd), .vdd(vdd), .A(_8253_), .Y(_56__14_) );
INVX1 INVX1_3630 ( .gnd(gnd), .vdd(vdd), .A(data_14__15_), .Y(_8254_) );
OAI21X1 OAI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_15788__bF_buf0), .B(_15031__bF_buf0), .C(_8254_), .Y(_8255_) );
OAI21X1 OAI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf0), .B(_8216_), .C(_8255_), .Y(_8256_) );
INVX1 INVX1_3631 ( .gnd(gnd), .vdd(vdd), .A(_8256_), .Y(_56__15_) );
INVX1 INVX1_3632 ( .gnd(gnd), .vdd(vdd), .A(data_13__0_), .Y(_8257_) );
OAI21X1 OAI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_15835_), .B(_15031__bF_buf3), .C(_15013_), .Y(_8258_) );
INVX1 INVX1_3633 ( .gnd(gnd), .vdd(vdd), .A(_8085_), .Y(_8259_) );
OAI21X1 OAI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_15175__bF_buf1), .C(_8259_), .Y(_8260_) );
OR2X2 OR2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_8260_), .B(_8258_), .Y(_8261_) );
NOR3X1 NOR3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8261_), .C(_15074__bF_buf11), .Y(_8262_) );
NAND3X1 NAND3X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_8262_), .C(_3391__bF_buf3), .Y(_8263_) );
MUX2X1 MUX2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_8257_), .B(_14932__bF_buf12), .S(_8263_), .Y(_45__0_) );
INVX1 INVX1_3634 ( .gnd(gnd), .vdd(vdd), .A(data_13__1_), .Y(_8264_) );
MUX2X1 MUX2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_8264_), .B(_14894__bF_buf10), .S(_8263_), .Y(_45__1_) );
INVX1 INVX1_3635 ( .gnd(gnd), .vdd(vdd), .A(data_13__2_), .Y(_8265_) );
MUX2X1 MUX2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_8265_), .B(_14897__bF_buf5), .S(_8263_), .Y(_45__2_) );
INVX1 INVX1_3636 ( .gnd(gnd), .vdd(vdd), .A(data_13__3_), .Y(_8266_) );
MUX2X1 MUX2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_8266_), .B(_14899__bF_buf10), .S(_8263_), .Y(_45__3_) );
INVX1 INVX1_3637 ( .gnd(gnd), .vdd(vdd), .A(data_13__4_), .Y(_8267_) );
MUX2X1 MUX2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_8267_), .B(_14902__bF_buf1), .S(_8263_), .Y(_45__4_) );
INVX1 INVX1_3638 ( .gnd(gnd), .vdd(vdd), .A(data_13__5_), .Y(_8268_) );
MUX2X1 MUX2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_8268_), .B(_14903__bF_buf13), .S(_8263_), .Y(_45__5_) );
INVX1 INVX1_3639 ( .gnd(gnd), .vdd(vdd), .A(data_13__6_), .Y(_8269_) );
MUX2X1 MUX2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_8269_), .B(_15049__bF_buf10), .S(_8263_), .Y(_45__6_) );
INVX1 INVX1_3640 ( .gnd(gnd), .vdd(vdd), .A(data_13__7_), .Y(_8270_) );
MUX2X1 MUX2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_8270_), .B(_14908__bF_buf2), .S(_8263_), .Y(_45__7_) );
INVX1 INVX1_3641 ( .gnd(gnd), .vdd(vdd), .A(data_13__8_), .Y(_8271_) );
MUX2X1 MUX2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_8271_), .B(_15052__bF_buf12), .S(_8263_), .Y(_45__8_) );
INVX1 INVX1_3642 ( .gnd(gnd), .vdd(vdd), .A(data_13__9_), .Y(_8272_) );
MUX2X1 MUX2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_8272_), .B(_14913__bF_buf7), .S(_8263_), .Y(_45__9_) );
INVX1 INVX1_3643 ( .gnd(gnd), .vdd(vdd), .A(data_13__10_), .Y(_8273_) );
MUX2X1 MUX2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_8273_), .B(_15055__bF_buf13), .S(_8263_), .Y(_45__10_) );
INVX1 INVX1_3644 ( .gnd(gnd), .vdd(vdd), .A(data_13__11_), .Y(_8274_) );
MUX2X1 MUX2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_8274_), .B(_14918__bF_buf0), .S(_8263_), .Y(_45__11_) );
INVX1 INVX1_3645 ( .gnd(gnd), .vdd(vdd), .A(data_13__12_), .Y(_8275_) );
MUX2X1 MUX2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_8275_), .B(_14920__bF_buf1), .S(_8263_), .Y(_45__12_) );
INVX1 INVX1_3646 ( .gnd(gnd), .vdd(vdd), .A(data_13__13_), .Y(_8276_) );
MUX2X1 MUX2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_8276_), .B(_14924__bF_buf13), .S(_8263_), .Y(_45__13_) );
INVX1 INVX1_3647 ( .gnd(gnd), .vdd(vdd), .A(data_13__14_), .Y(_8277_) );
MUX2X1 MUX2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_8277_), .B(_15060__bF_buf12), .S(_8263_), .Y(_45__14_) );
INVX1 INVX1_3648 ( .gnd(gnd), .vdd(vdd), .A(data_13__15_), .Y(_8278_) );
MUX2X1 MUX2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_8278_), .B(_15062__bF_buf2), .S(_8263_), .Y(_45__15_) );
NOR3X1 NOR3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .B(_8085_), .C(_8126_), .Y(_8279_) );
AND2X2 AND2X2_1475 ( .gnd(gnd), .vdd(vdd), .A(_8125__bF_buf4), .B(_8279__bF_buf3), .Y(_8280_) );
AOI21X1 AOI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf2), .B(_8125__bF_buf3), .C(data_12__0_), .Y(_8281_) );
AOI21X1 AOI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf11), .B(_8280_), .C(_8281_), .Y(_34__0_) );
AOI21X1 AOI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf1), .B(_8125__bF_buf2), .C(data_12__1_), .Y(_8282_) );
AOI21X1 AOI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf9), .B(_8280_), .C(_8282_), .Y(_34__1_) );
AOI21X1 AOI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf0), .B(_8125__bF_buf1), .C(data_12__2_), .Y(_8283_) );
AOI21X1 AOI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf4), .B(_8280_), .C(_8283_), .Y(_34__2_) );
AOI21X1 AOI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf3), .B(_8125__bF_buf0), .C(data_12__3_), .Y(_8284_) );
AOI21X1 AOI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf9), .B(_8280_), .C(_8284_), .Y(_34__3_) );
AOI21X1 AOI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf2), .B(_8125__bF_buf5), .C(data_12__4_), .Y(_8285_) );
AOI21X1 AOI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf0), .B(_8280_), .C(_8285_), .Y(_34__4_) );
AOI21X1 AOI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf1), .B(_8125__bF_buf4), .C(data_12__5_), .Y(_8286_) );
AOI21X1 AOI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf12), .B(_8280_), .C(_8286_), .Y(_34__5_) );
AOI21X1 AOI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf0), .B(_8125__bF_buf3), .C(data_12__6_), .Y(_8287_) );
AOI21X1 AOI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf9), .B(_8280_), .C(_8287_), .Y(_34__6_) );
AOI21X1 AOI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf3), .B(_8125__bF_buf2), .C(data_12__7_), .Y(_8288_) );
AOI21X1 AOI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf1), .B(_8280_), .C(_8288_), .Y(_34__7_) );
AOI21X1 AOI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf2), .B(_8125__bF_buf1), .C(data_12__8_), .Y(_8289_) );
AOI21X1 AOI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf11), .B(_8280_), .C(_8289_), .Y(_34__8_) );
AOI21X1 AOI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf1), .B(_8125__bF_buf0), .C(data_12__9_), .Y(_8290_) );
AOI21X1 AOI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf6), .B(_8280_), .C(_8290_), .Y(_34__9_) );
AOI21X1 AOI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf0), .B(_8125__bF_buf5), .C(data_12__10_), .Y(_8291_) );
AOI21X1 AOI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf12), .B(_8280_), .C(_8291_), .Y(_34__10_) );
AOI21X1 AOI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf3), .B(_8125__bF_buf4), .C(data_12__11_), .Y(_8292_) );
AOI21X1 AOI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf13), .B(_8280_), .C(_8292_), .Y(_34__11_) );
AOI21X1 AOI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf2), .B(_8125__bF_buf3), .C(data_12__12_), .Y(_8293_) );
AOI21X1 AOI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf0), .B(_8280_), .C(_8293_), .Y(_34__12_) );
AOI21X1 AOI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf1), .B(_8125__bF_buf2), .C(data_12__13_), .Y(_8294_) );
AOI21X1 AOI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf12), .B(_8280_), .C(_8294_), .Y(_34__13_) );
AOI21X1 AOI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf0), .B(_8125__bF_buf1), .C(data_12__14_), .Y(_8295_) );
AOI21X1 AOI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf11), .B(_8280_), .C(_8295_), .Y(_34__14_) );
AOI21X1 AOI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_8279__bF_buf3), .B(_8125__bF_buf0), .C(data_12__15_), .Y(_8296_) );
AOI21X1 AOI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf1), .B(_8280_), .C(_8296_), .Y(_34__15_) );
INVX1 INVX1_3649 ( .gnd(gnd), .vdd(vdd), .A(data_11__0_), .Y(_8297_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .Y(_8298_) );
OAI21X1 OAI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_15031__bF_buf2), .B(_14977__bF_buf3), .C(IDATA_PROG_write_bF_buf2), .Y(_8299_) );
INVX1 INVX1_3650 ( .gnd(gnd), .vdd(vdd), .A(_8299_), .Y(_8300_) );
OAI21X1 OAI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_15160_), .B(_15031__bF_buf1), .C(_8300_), .Y(_8301_) );
AOI21X1 AOI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_15011__bF_buf1), .B(_15163_), .C(_8301_), .Y(_8302_) );
NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_8298_), .B(_8302_), .Y(_8303_) );
NOR2X1 NOR2X1_852 ( .gnd(gnd), .vdd(vdd), .A(_8303_), .B(_8126_), .Y(_8304_) );
NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_8304_), .B(_8125__bF_buf5), .Y(_8305_) );
MUX2X1 MUX2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_8297_), .B(_14932__bF_buf10), .S(_8305_), .Y(_23__0_) );
INVX1 INVX1_3651 ( .gnd(gnd), .vdd(vdd), .A(data_11__1_), .Y(_8306_) );
MUX2X1 MUX2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_8306_), .B(_14894__bF_buf8), .S(_8305_), .Y(_23__1_) );
INVX1 INVX1_3652 ( .gnd(gnd), .vdd(vdd), .A(data_11__2_), .Y(_8307_) );
NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_8307_), .B(_8305_), .Y(_8308_) );
AND2X2 AND2X2_1476 ( .gnd(gnd), .vdd(vdd), .A(_8125__bF_buf4), .B(_8304_), .Y(_8309_) );
NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf3), .B(_8309_), .Y(_8310_) );
AND2X2 AND2X2_1477 ( .gnd(gnd), .vdd(vdd), .A(_8310_), .B(_8308_), .Y(_23__2_) );
INVX1 INVX1_3653 ( .gnd(gnd), .vdd(vdd), .A(data_11__3_), .Y(_8311_) );
MUX2X1 MUX2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_8311_), .B(_14899__bF_buf8), .S(_8305_), .Y(_23__3_) );
INVX1 INVX1_3654 ( .gnd(gnd), .vdd(vdd), .A(data_11__4_), .Y(_8312_) );
MUX2X1 MUX2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_8312_), .B(_14902__bF_buf13), .S(_8305_), .Y(_23__4_) );
INVX1 INVX1_3655 ( .gnd(gnd), .vdd(vdd), .A(data_11__5_), .Y(_8313_) );
MUX2X1 MUX2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_8313_), .B(_14903__bF_buf11), .S(_8305_), .Y(_23__5_) );
INVX1 INVX1_3656 ( .gnd(gnd), .vdd(vdd), .A(data_11__6_), .Y(_8314_) );
NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_8314_), .B(_8305_), .Y(_8315_) );
NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf8), .B(_8309_), .Y(_8316_) );
AND2X2 AND2X2_1478 ( .gnd(gnd), .vdd(vdd), .A(_8316_), .B(_8315_), .Y(_23__6_) );
INVX1 INVX1_3657 ( .gnd(gnd), .vdd(vdd), .A(data_11__7_), .Y(_8317_) );
MUX2X1 MUX2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_8317_), .B(_14908__bF_buf0), .S(_8305_), .Y(_23__7_) );
INVX1 INVX1_3658 ( .gnd(gnd), .vdd(vdd), .A(data_11__8_), .Y(_8318_) );
NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_8318_), .B(_8305_), .Y(_8319_) );
NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf10), .B(_8309_), .Y(_8320_) );
AND2X2 AND2X2_1479 ( .gnd(gnd), .vdd(vdd), .A(_8320_), .B(_8319_), .Y(_23__8_) );
INVX1 INVX1_3659 ( .gnd(gnd), .vdd(vdd), .A(data_11__9_), .Y(_8321_) );
NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_8321_), .B(_8305_), .Y(_8322_) );
NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf5), .B(_8309_), .Y(_8323_) );
AND2X2 AND2X2_1480 ( .gnd(gnd), .vdd(vdd), .A(_8323_), .B(_8322_), .Y(_23__9_) );
INVX1 INVX1_3660 ( .gnd(gnd), .vdd(vdd), .A(data_11__10_), .Y(_8324_) );
NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_8324_), .B(_8305_), .Y(_8325_) );
NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf11), .B(_8309_), .Y(_8326_) );
AND2X2 AND2X2_1481 ( .gnd(gnd), .vdd(vdd), .A(_8326_), .B(_8325_), .Y(_23__10_) );
INVX1 INVX1_3661 ( .gnd(gnd), .vdd(vdd), .A(data_11__11_), .Y(_8327_) );
MUX2X1 MUX2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_8327_), .B(_14918__bF_buf12), .S(_8305_), .Y(_23__11_) );
INVX1 INVX1_3662 ( .gnd(gnd), .vdd(vdd), .A(data_11__12_), .Y(_8328_) );
MUX2X1 MUX2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_8328_), .B(_14920__bF_buf13), .S(_8305_), .Y(_23__12_) );
INVX1 INVX1_3663 ( .gnd(gnd), .vdd(vdd), .A(data_11__13_), .Y(_8329_) );
NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_8329_), .B(_8305_), .Y(_8330_) );
NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf11), .B(_8309_), .Y(_8331_) );
AND2X2 AND2X2_1482 ( .gnd(gnd), .vdd(vdd), .A(_8331_), .B(_8330_), .Y(_23__13_) );
INVX1 INVX1_3664 ( .gnd(gnd), .vdd(vdd), .A(data_11__14_), .Y(_8332_) );
NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_8332_), .B(_8305_), .Y(_8333_) );
NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf10), .B(_8309_), .Y(_8334_) );
AND2X2 AND2X2_1483 ( .gnd(gnd), .vdd(vdd), .A(_8334_), .B(_8333_), .Y(_23__14_) );
INVX1 INVX1_3665 ( .gnd(gnd), .vdd(vdd), .A(data_11__15_), .Y(_8335_) );
NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_8335_), .B(_8305_), .Y(_8336_) );
NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf0), .B(_8309_), .Y(_8337_) );
AND2X2 AND2X2_1484 ( .gnd(gnd), .vdd(vdd), .A(_8337_), .B(_8336_), .Y(_23__15_) );
INVX1 INVX1_3666 ( .gnd(gnd), .vdd(vdd), .A(data_10__0_), .Y(_8338_) );
AOI21X1 AOI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_14991_), .B(_15011__bF_buf0), .C(_8299_), .Y(_8339_) );
AOI21X1 AOI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_15161_), .B(_15011__bF_buf3), .C(_15014_), .Y(_8340_) );
NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_8339_), .B(_8340_), .Y(_8341_) );
NOR2X1 NOR2X1_853 ( .gnd(gnd), .vdd(vdd), .A(_8341_), .B(_8126_), .Y(_8342_) );
NAND3X1 NAND3X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_3391__bF_buf2), .B(_3307_), .C(_8342_), .Y(_8343_) );
MUX2X1 MUX2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_8338_), .B(_14932__bF_buf9), .S(_8343_), .Y(_12__0_) );
INVX1 INVX1_3667 ( .gnd(gnd), .vdd(vdd), .A(data_10__1_), .Y(_8344_) );
MUX2X1 MUX2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_8344_), .B(_14894__bF_buf7), .S(_8343_), .Y(_12__1_) );
INVX1 INVX1_3668 ( .gnd(gnd), .vdd(vdd), .A(data_10__2_), .Y(_8345_) );
MUX2X1 MUX2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_8345_), .B(_14897__bF_buf2), .S(_8343_), .Y(_12__2_) );
INVX1 INVX1_3669 ( .gnd(gnd), .vdd(vdd), .A(data_10__3_), .Y(_8346_) );
MUX2X1 MUX2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_8346_), .B(_14899__bF_buf7), .S(_8343_), .Y(_12__3_) );
INVX1 INVX1_3670 ( .gnd(gnd), .vdd(vdd), .A(data_10__4_), .Y(_8347_) );
MUX2X1 MUX2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_8347_), .B(_14902__bF_buf12), .S(_8343_), .Y(_12__4_) );
INVX1 INVX1_3671 ( .gnd(gnd), .vdd(vdd), .A(data_10__5_), .Y(_8348_) );
MUX2X1 MUX2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_8348_), .B(_14903__bF_buf10), .S(_8343_), .Y(_12__5_) );
INVX1 INVX1_3672 ( .gnd(gnd), .vdd(vdd), .A(data_10__6_), .Y(_8349_) );
MUX2X1 MUX2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_8349_), .B(_15049__bF_buf7), .S(_8343_), .Y(_12__6_) );
INVX1 INVX1_3673 ( .gnd(gnd), .vdd(vdd), .A(data_10__7_), .Y(_8350_) );
MUX2X1 MUX2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_8350_), .B(_14908__bF_buf13), .S(_8343_), .Y(_12__7_) );
INVX1 INVX1_3674 ( .gnd(gnd), .vdd(vdd), .A(data_10__8_), .Y(_8351_) );
MUX2X1 MUX2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_8351_), .B(_15052__bF_buf9), .S(_8343_), .Y(_12__8_) );
INVX1 INVX1_3675 ( .gnd(gnd), .vdd(vdd), .A(data_10__9_), .Y(_8352_) );
MUX2X1 MUX2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_8352_), .B(_14913__bF_buf4), .S(_8343_), .Y(_12__9_) );
INVX1 INVX1_3676 ( .gnd(gnd), .vdd(vdd), .A(data_10__10_), .Y(_8353_) );
MUX2X1 MUX2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_8353_), .B(_15055__bF_buf10), .S(_8343_), .Y(_12__10_) );
INVX1 INVX1_3677 ( .gnd(gnd), .vdd(vdd), .A(data_10__11_), .Y(_8354_) );
MUX2X1 MUX2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_8354_), .B(_14918__bF_buf11), .S(_8343_), .Y(_12__11_) );
INVX1 INVX1_3678 ( .gnd(gnd), .vdd(vdd), .A(data_10__12_), .Y(_8355_) );
MUX2X1 MUX2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_8355_), .B(_14920__bF_buf12), .S(_8343_), .Y(_12__12_) );
INVX1 INVX1_3679 ( .gnd(gnd), .vdd(vdd), .A(data_10__13_), .Y(_8356_) );
MUX2X1 MUX2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_8356_), .B(_14924__bF_buf10), .S(_8343_), .Y(_12__13_) );
INVX1 INVX1_3680 ( .gnd(gnd), .vdd(vdd), .A(data_10__14_), .Y(_8357_) );
MUX2X1 MUX2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_8357_), .B(_15060__bF_buf9), .S(_8343_), .Y(_12__14_) );
INVX1 INVX1_3681 ( .gnd(gnd), .vdd(vdd), .A(data_10__15_), .Y(_8358_) );
MUX2X1 MUX2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_8358_), .B(_15062__bF_buf13), .S(_8343_), .Y(_12__15_) );
INVX1 INVX1_3682 ( .gnd(gnd), .vdd(vdd), .A(data_9__0_), .Y(_8359_) );
NOR2X1 NOR2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_15074__bF_buf10), .Y(_8360_) );
INVX1 INVX1_3683 ( .gnd(gnd), .vdd(vdd), .A(_15285_), .Y(_8361_) );
OAI21X1 OAI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_8361_), .B(_15031__bF_buf0), .C(_8339_), .Y(_8362_) );
INVX1 INVX1_3684 ( .gnd(gnd), .vdd(vdd), .A(_8362_), .Y(_8363_) );
NAND3X1 NAND3X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_8298_), .B(_8363_), .C(_8360_), .Y(_8364_) );
OAI21X1 OAI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf4), .B(_8364__bF_buf3), .C(_8359_), .Y(_8365_) );
NOR2X1 NOR2X1_855 ( .gnd(gnd), .vdd(vdd), .A(_8364__bF_buf2), .B(_3989__bF_buf3), .Y(_8366_) );
NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf8), .B(_8366_), .Y(_8367_) );
AND2X2 AND2X2_1485 ( .gnd(gnd), .vdd(vdd), .A(_8367_), .B(_8365_), .Y(_256__0_) );
INVX1 INVX1_3685 ( .gnd(gnd), .vdd(vdd), .A(data_9__1_), .Y(_8368_) );
OAI21X1 OAI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf2), .B(_8364__bF_buf1), .C(_8368_), .Y(_8369_) );
NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf6), .B(_8366_), .Y(_8370_) );
AND2X2 AND2X2_1486 ( .gnd(gnd), .vdd(vdd), .A(_8370_), .B(_8369_), .Y(_256__1_) );
INVX1 INVX1_3686 ( .gnd(gnd), .vdd(vdd), .A(data_9__2_), .Y(_8371_) );
OAI21X1 OAI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf1), .B(_8364__bF_buf0), .C(_8371_), .Y(_8372_) );
NOR3X1 NOR3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_15014_), .B(_8362_), .C(_8126_), .Y(_8373_) );
NAND3X1 NAND3X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf1), .B(_8373_), .C(_8125__bF_buf3), .Y(_8374_) );
AND2X2 AND2X2_1487 ( .gnd(gnd), .vdd(vdd), .A(_8372_), .B(_8374_), .Y(_256__2_) );
INVX1 INVX1_3687 ( .gnd(gnd), .vdd(vdd), .A(data_9__3_), .Y(_8375_) );
OAI21X1 OAI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf0), .B(_8364__bF_buf3), .C(_8375_), .Y(_8376_) );
NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf6), .B(_8366_), .Y(_8377_) );
AND2X2 AND2X2_1488 ( .gnd(gnd), .vdd(vdd), .A(_8377_), .B(_8376_), .Y(_256__3_) );
INVX1 INVX1_3688 ( .gnd(gnd), .vdd(vdd), .A(data_9__4_), .Y(_8378_) );
OAI21X1 OAI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf4), .B(_8364__bF_buf2), .C(_8378_), .Y(_8379_) );
NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf11), .B(_8366_), .Y(_8380_) );
AND2X2 AND2X2_1489 ( .gnd(gnd), .vdd(vdd), .A(_8380_), .B(_8379_), .Y(_256__4_) );
INVX1 INVX1_3689 ( .gnd(gnd), .vdd(vdd), .A(data_9__5_), .Y(_8381_) );
OAI21X1 OAI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf3), .B(_8364__bF_buf1), .C(_8381_), .Y(_8382_) );
NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf9), .B(_8366_), .Y(_8383_) );
AND2X2 AND2X2_1490 ( .gnd(gnd), .vdd(vdd), .A(_8383_), .B(_8382_), .Y(_256__5_) );
INVX1 INVX1_3690 ( .gnd(gnd), .vdd(vdd), .A(data_9__6_), .Y(_8384_) );
OAI21X1 OAI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf2), .B(_8364__bF_buf0), .C(_8384_), .Y(_8385_) );
NAND3X1 NAND3X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf6), .B(_8373_), .C(_8125__bF_buf2), .Y(_8386_) );
AND2X2 AND2X2_1491 ( .gnd(gnd), .vdd(vdd), .A(_8385_), .B(_8386_), .Y(_256__6_) );
INVX1 INVX1_3691 ( .gnd(gnd), .vdd(vdd), .A(data_9__7_), .Y(_8387_) );
OAI21X1 OAI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf1), .B(_8364__bF_buf3), .C(_8387_), .Y(_8388_) );
NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf12), .B(_8366_), .Y(_8389_) );
AND2X2 AND2X2_1492 ( .gnd(gnd), .vdd(vdd), .A(_8389_), .B(_8388_), .Y(_256__7_) );
INVX1 INVX1_3692 ( .gnd(gnd), .vdd(vdd), .A(data_9__8_), .Y(_8390_) );
OAI21X1 OAI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf0), .B(_8364__bF_buf2), .C(_8390_), .Y(_8391_) );
NAND3X1 NAND3X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf8), .B(_8373_), .C(_8125__bF_buf1), .Y(_8392_) );
AND2X2 AND2X2_1493 ( .gnd(gnd), .vdd(vdd), .A(_8391_), .B(_8392_), .Y(_256__8_) );
INVX1 INVX1_3693 ( .gnd(gnd), .vdd(vdd), .A(data_9__9_), .Y(_8393_) );
OAI21X1 OAI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf4), .B(_8364__bF_buf1), .C(_8393_), .Y(_8394_) );
NAND3X1 NAND3X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf3), .B(_8373_), .C(_8125__bF_buf0), .Y(_8395_) );
AND2X2 AND2X2_1494 ( .gnd(gnd), .vdd(vdd), .A(_8394_), .B(_8395_), .Y(_256__9_) );
INVX1 INVX1_3694 ( .gnd(gnd), .vdd(vdd), .A(data_9__10_), .Y(_8396_) );
OAI21X1 OAI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf3), .B(_8364__bF_buf0), .C(_8396_), .Y(_8397_) );
NAND3X1 NAND3X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf9), .B(_8373_), .C(_8125__bF_buf5), .Y(_8398_) );
AND2X2 AND2X2_1495 ( .gnd(gnd), .vdd(vdd), .A(_8397_), .B(_8398_), .Y(_256__10_) );
INVX1 INVX1_3695 ( .gnd(gnd), .vdd(vdd), .A(data_9__11_), .Y(_8399_) );
OAI21X1 OAI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf2), .B(_8364__bF_buf3), .C(_8399_), .Y(_8400_) );
NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf10), .B(_8366_), .Y(_8401_) );
AND2X2 AND2X2_1496 ( .gnd(gnd), .vdd(vdd), .A(_8401_), .B(_8400_), .Y(_256__11_) );
INVX1 INVX1_3696 ( .gnd(gnd), .vdd(vdd), .A(data_9__12_), .Y(_8402_) );
OAI21X1 OAI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf1), .B(_8364__bF_buf2), .C(_8402_), .Y(_8403_) );
NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf11), .B(_8366_), .Y(_8404_) );
AND2X2 AND2X2_1497 ( .gnd(gnd), .vdd(vdd), .A(_8404_), .B(_8403_), .Y(_256__12_) );
INVX1 INVX1_3697 ( .gnd(gnd), .vdd(vdd), .A(data_9__13_), .Y(_8405_) );
OAI21X1 OAI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf0), .B(_8364__bF_buf1), .C(_8405_), .Y(_8406_) );
NAND3X1 NAND3X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf9), .B(_8373_), .C(_8125__bF_buf4), .Y(_8407_) );
AND2X2 AND2X2_1498 ( .gnd(gnd), .vdd(vdd), .A(_8406_), .B(_8407_), .Y(_256__13_) );
INVX1 INVX1_3698 ( .gnd(gnd), .vdd(vdd), .A(data_9__14_), .Y(_8408_) );
OAI21X1 OAI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf4), .B(_8364__bF_buf0), .C(_8408_), .Y(_8409_) );
NAND3X1 NAND3X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf8), .B(_8373_), .C(_8125__bF_buf3), .Y(_8410_) );
AND2X2 AND2X2_1499 ( .gnd(gnd), .vdd(vdd), .A(_8409_), .B(_8410_), .Y(_256__14_) );
INVX1 INVX1_3699 ( .gnd(gnd), .vdd(vdd), .A(data_9__15_), .Y(_8411_) );
OAI21X1 OAI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf3), .B(_8364__bF_buf3), .C(_8411_), .Y(_8412_) );
NAND3X1 NAND3X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf12), .B(_8373_), .C(_8125__bF_buf2), .Y(_8413_) );
AND2X2 AND2X2_1500 ( .gnd(gnd), .vdd(vdd), .A(_8412_), .B(_8413_), .Y(_256__15_) );
NAND3X1 NAND3X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_15015_), .B(_8300_), .C(_8298_), .Y(_8414_) );
OR2X2 OR2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_8126_), .B(_8414_), .Y(_8415_) );
NOR2X1 NOR2X1_856 ( .gnd(gnd), .vdd(vdd), .A(_8415_), .B(_3989__bF_buf2), .Y(_8416_) );
NOR2X1 NOR2X1_857 ( .gnd(gnd), .vdd(vdd), .A(_8414_), .B(_8126_), .Y(_8417_) );
AOI21X1 AOI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .B(_8125__bF_buf1), .C(data_8__0_), .Y(_8418_) );
AOI21X1 AOI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf7), .B(_8416_), .C(_8418_), .Y(_245__0_) );
INVX1 INVX1_3700 ( .gnd(gnd), .vdd(vdd), .A(data_8__1_), .Y(_8419_) );
NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_8417_), .B(_8125__bF_buf0), .Y(_8420_) );
MUX2X1 MUX2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_8419_), .B(_14894__bF_buf5), .S(_8420_), .Y(_245__1_) );
INVX1 INVX1_3701 ( .gnd(gnd), .vdd(vdd), .A(data_8__2_), .Y(_8421_) );
OAI21X1 OAI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf1), .B(_8415_), .C(_8421_), .Y(_8422_) );
NAND3X1 NAND3X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf0), .B(_8417_), .C(_8125__bF_buf5), .Y(_8423_) );
AND2X2 AND2X2_1501 ( .gnd(gnd), .vdd(vdd), .A(_8422_), .B(_8423_), .Y(_245__2_) );
INVX1 INVX1_3702 ( .gnd(gnd), .vdd(vdd), .A(data_8__3_), .Y(_8424_) );
MUX2X1 MUX2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_8424_), .B(_14899__bF_buf5), .S(_8420_), .Y(_245__3_) );
INVX1 INVX1_3703 ( .gnd(gnd), .vdd(vdd), .A(data_8__4_), .Y(_8425_) );
MUX2X1 MUX2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_8425_), .B(_14902__bF_buf10), .S(_8420_), .Y(_245__4_) );
INVX1 INVX1_3704 ( .gnd(gnd), .vdd(vdd), .A(data_8__5_), .Y(_8426_) );
MUX2X1 MUX2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_8426_), .B(_14903__bF_buf8), .S(_8420_), .Y(_245__5_) );
INVX1 INVX1_3705 ( .gnd(gnd), .vdd(vdd), .A(data_8__6_), .Y(_8427_) );
OAI21X1 OAI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf0), .B(_8415_), .C(_8427_), .Y(_8428_) );
NAND3X1 NAND3X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf5), .B(_8417_), .C(_8125__bF_buf4), .Y(_8429_) );
AND2X2 AND2X2_1502 ( .gnd(gnd), .vdd(vdd), .A(_8428_), .B(_8429_), .Y(_245__6_) );
INVX1 INVX1_3706 ( .gnd(gnd), .vdd(vdd), .A(data_8__7_), .Y(_8430_) );
MUX2X1 MUX2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_8430_), .B(_14908__bF_buf11), .S(_8420_), .Y(_245__7_) );
INVX1 INVX1_3707 ( .gnd(gnd), .vdd(vdd), .A(data_8__8_), .Y(_8431_) );
OAI21X1 OAI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf4), .B(_8415_), .C(_8431_), .Y(_8432_) );
NAND3X1 NAND3X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf7), .B(_8417_), .C(_8125__bF_buf3), .Y(_8433_) );
AND2X2 AND2X2_1503 ( .gnd(gnd), .vdd(vdd), .A(_8432_), .B(_8433_), .Y(_245__8_) );
INVX1 INVX1_3708 ( .gnd(gnd), .vdd(vdd), .A(data_8__9_), .Y(_8434_) );
OAI21X1 OAI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf3), .B(_8415_), .C(_8434_), .Y(_8435_) );
NAND3X1 NAND3X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf2), .B(_8417_), .C(_8125__bF_buf2), .Y(_8436_) );
AND2X2 AND2X2_1504 ( .gnd(gnd), .vdd(vdd), .A(_8435_), .B(_8436_), .Y(_245__9_) );
INVX1 INVX1_3709 ( .gnd(gnd), .vdd(vdd), .A(data_8__10_), .Y(_8437_) );
OAI21X1 OAI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf2), .B(_8415_), .C(_8437_), .Y(_8438_) );
NAND3X1 NAND3X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf8), .B(_8417_), .C(_8125__bF_buf1), .Y(_8439_) );
AND2X2 AND2X2_1505 ( .gnd(gnd), .vdd(vdd), .A(_8438_), .B(_8439_), .Y(_245__10_) );
INVX1 INVX1_3710 ( .gnd(gnd), .vdd(vdd), .A(data_8__11_), .Y(_8440_) );
MUX2X1 MUX2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_8440_), .B(_14918__bF_buf9), .S(_8420_), .Y(_245__11_) );
INVX1 INVX1_3711 ( .gnd(gnd), .vdd(vdd), .A(data_8__12_), .Y(_8441_) );
MUX2X1 MUX2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_8441_), .B(_14920__bF_buf10), .S(_8420_), .Y(_245__12_) );
INVX1 INVX1_3712 ( .gnd(gnd), .vdd(vdd), .A(data_8__13_), .Y(_8442_) );
OAI21X1 OAI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf1), .B(_8415_), .C(_8442_), .Y(_8443_) );
NAND3X1 NAND3X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf8), .B(_8417_), .C(_8125__bF_buf0), .Y(_8444_) );
AND2X2 AND2X2_1506 ( .gnd(gnd), .vdd(vdd), .A(_8443_), .B(_8444_), .Y(_245__13_) );
INVX1 INVX1_3713 ( .gnd(gnd), .vdd(vdd), .A(data_8__14_), .Y(_8445_) );
OAI21X1 OAI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf0), .B(_8415_), .C(_8445_), .Y(_8446_) );
NAND3X1 NAND3X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf7), .B(_8417_), .C(_8125__bF_buf5), .Y(_8447_) );
AND2X2 AND2X2_1507 ( .gnd(gnd), .vdd(vdd), .A(_8446_), .B(_8447_), .Y(_245__14_) );
INVX1 INVX1_3714 ( .gnd(gnd), .vdd(vdd), .A(data_8__15_), .Y(_8448_) );
OAI21X1 OAI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_3989__bF_buf4), .B(_8415_), .C(_8448_), .Y(_8449_) );
NAND3X1 NAND3X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf11), .B(_8417_), .C(_8125__bF_buf4), .Y(_8450_) );
AND2X2 AND2X2_1508 ( .gnd(gnd), .vdd(vdd), .A(_8449_), .B(_8450_), .Y(_245__15_) );
INVX1 INVX1_3715 ( .gnd(gnd), .vdd(vdd), .A(data_7__0_), .Y(_8451_) );
AOI21X1 AOI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_15011__bF_buf2), .B(_15363_), .C(_15014_), .Y(_8452_) );
AOI21X1 AOI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_15011__bF_buf1), .B(_1989_), .C(_14882__bF_buf5), .Y(_8453_) );
NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_8453_), .B(_8452_), .Y(_8454_) );
NOR3X1 NOR3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8454_), .C(_15074__bF_buf9), .Y(_8455_) );
NAND3X1 NAND3X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .B(_8455_), .C(_3391__bF_buf1), .Y(_8456_) );
MUX2X1 MUX2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_8451_), .B(_14932__bF_buf6), .S(_8456_), .Y(_234__0_) );
INVX1 INVX1_3716 ( .gnd(gnd), .vdd(vdd), .A(data_7__1_), .Y(_8457_) );
MUX2X1 MUX2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_8457_), .B(_14894__bF_buf4), .S(_8456_), .Y(_234__1_) );
INVX1 INVX1_3717 ( .gnd(gnd), .vdd(vdd), .A(data_7__2_), .Y(_8458_) );
MUX2X1 MUX2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_8458_), .B(_14897__bF_buf14), .S(_8456_), .Y(_234__2_) );
INVX1 INVX1_3718 ( .gnd(gnd), .vdd(vdd), .A(data_7__3_), .Y(_8459_) );
MUX2X1 MUX2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_8459_), .B(_14899__bF_buf4), .S(_8456_), .Y(_234__3_) );
INVX1 INVX1_3719 ( .gnd(gnd), .vdd(vdd), .A(data_7__4_), .Y(_8460_) );
MUX2X1 MUX2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_8460_), .B(_14902__bF_buf9), .S(_8456_), .Y(_234__4_) );
INVX1 INVX1_3720 ( .gnd(gnd), .vdd(vdd), .A(data_7__5_), .Y(_8461_) );
MUX2X1 MUX2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_8461_), .B(_14903__bF_buf7), .S(_8456_), .Y(_234__5_) );
INVX1 INVX1_3721 ( .gnd(gnd), .vdd(vdd), .A(data_7__6_), .Y(_8462_) );
MUX2X1 MUX2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_8462_), .B(_15049__bF_buf4), .S(_8456_), .Y(_234__6_) );
INVX1 INVX1_3722 ( .gnd(gnd), .vdd(vdd), .A(data_7__7_), .Y(_8463_) );
MUX2X1 MUX2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_8463_), .B(_14908__bF_buf10), .S(_8456_), .Y(_234__7_) );
INVX1 INVX1_3723 ( .gnd(gnd), .vdd(vdd), .A(data_7__8_), .Y(_8464_) );
MUX2X1 MUX2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_8464_), .B(_15052__bF_buf6), .S(_8456_), .Y(_234__8_) );
INVX1 INVX1_3724 ( .gnd(gnd), .vdd(vdd), .A(data_7__9_), .Y(_8465_) );
MUX2X1 MUX2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_8465_), .B(_14913__bF_buf1), .S(_8456_), .Y(_234__9_) );
INVX1 INVX1_3725 ( .gnd(gnd), .vdd(vdd), .A(data_7__10_), .Y(_8466_) );
MUX2X1 MUX2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_8466_), .B(_15055__bF_buf7), .S(_8456_), .Y(_234__10_) );
INVX1 INVX1_3726 ( .gnd(gnd), .vdd(vdd), .A(data_7__11_), .Y(_8467_) );
MUX2X1 MUX2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_8467_), .B(_14918__bF_buf8), .S(_8456_), .Y(_234__11_) );
INVX1 INVX1_3727 ( .gnd(gnd), .vdd(vdd), .A(data_7__12_), .Y(_8468_) );
MUX2X1 MUX2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_8468_), .B(_14920__bF_buf9), .S(_8456_), .Y(_234__12_) );
INVX1 INVX1_3728 ( .gnd(gnd), .vdd(vdd), .A(data_7__13_), .Y(_8469_) );
MUX2X1 MUX2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_8469_), .B(_14924__bF_buf7), .S(_8456_), .Y(_234__13_) );
INVX1 INVX1_3729 ( .gnd(gnd), .vdd(vdd), .A(data_7__14_), .Y(_8470_) );
MUX2X1 MUX2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_8470_), .B(_15060__bF_buf6), .S(_8456_), .Y(_234__14_) );
INVX1 INVX1_3730 ( .gnd(gnd), .vdd(vdd), .A(data_7__15_), .Y(_8471_) );
MUX2X1 MUX2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_8471_), .B(_15062__bF_buf10), .S(_8456_), .Y(_234__15_) );
INVX1 INVX1_3731 ( .gnd(gnd), .vdd(vdd), .A(data_6__0_), .Y(_8472_) );
AOI21X1 AOI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_14996_), .B(_15011__bF_buf0), .C(_15014_), .Y(_8473_) );
NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_8453_), .B(_8473_), .Y(_8474_) );
NOR2X1 NOR2X1_858 ( .gnd(gnd), .vdd(vdd), .A(_8474_), .B(_8126_), .Y(_8475_) );
NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_8475_), .B(_8125__bF_buf3), .Y(_8476_) );
MUX2X1 MUX2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8472_), .B(_14932__bF_buf5), .S(_8476__bF_buf3), .Y(_223__0_) );
INVX1 INVX1_3732 ( .gnd(gnd), .vdd(vdd), .A(data_6__1_), .Y(_8477_) );
NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_8477_), .B(_8476__bF_buf2), .Y(_8478_) );
OR2X2 OR2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_8476__bF_buf1), .B(IDATA_PROG_data_1_bF_buf0), .Y(_8479_) );
AND2X2 AND2X2_1509 ( .gnd(gnd), .vdd(vdd), .A(_8479_), .B(_8478_), .Y(_223__1_) );
INVX1 INVX1_3733 ( .gnd(gnd), .vdd(vdd), .A(data_6__2_), .Y(_8480_) );
MUX2X1 MUX2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_8480_), .B(_14897__bF_buf13), .S(_8476__bF_buf0), .Y(_223__2_) );
INVX1 INVX1_3734 ( .gnd(gnd), .vdd(vdd), .A(data_6__3_), .Y(_8481_) );
MUX2X1 MUX2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_8481_), .B(_14899__bF_buf3), .S(_8476__bF_buf3), .Y(_223__3_) );
INVX1 INVX1_3735 ( .gnd(gnd), .vdd(vdd), .A(data_6__4_), .Y(_8482_) );
MUX2X1 MUX2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_8482_), .B(_14902__bF_buf8), .S(_8476__bF_buf2), .Y(_223__4_) );
INVX1 INVX1_3736 ( .gnd(gnd), .vdd(vdd), .A(data_6__5_), .Y(_8483_) );
MUX2X1 MUX2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_8483_), .B(_14903__bF_buf6), .S(_8476__bF_buf1), .Y(_223__5_) );
INVX1 INVX1_3737 ( .gnd(gnd), .vdd(vdd), .A(data_6__6_), .Y(_8484_) );
MUX2X1 MUX2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_8484_), .B(_15049__bF_buf3), .S(_8476__bF_buf0), .Y(_223__6_) );
INVX1 INVX1_3738 ( .gnd(gnd), .vdd(vdd), .A(data_6__7_), .Y(_8485_) );
MUX2X1 MUX2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_8485_), .B(_14908__bF_buf9), .S(_8476__bF_buf3), .Y(_223__7_) );
INVX1 INVX1_3739 ( .gnd(gnd), .vdd(vdd), .A(data_6__8_), .Y(_8486_) );
MUX2X1 MUX2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_8486_), .B(_15052__bF_buf5), .S(_8476__bF_buf2), .Y(_223__8_) );
INVX1 INVX1_3740 ( .gnd(gnd), .vdd(vdd), .A(data_6__9_), .Y(_8487_) );
MUX2X1 MUX2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_8487_), .B(_14913__bF_buf0), .S(_8476__bF_buf1), .Y(_223__9_) );
INVX1 INVX1_3741 ( .gnd(gnd), .vdd(vdd), .A(data_6__10_), .Y(_8488_) );
MUX2X1 MUX2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_8488_), .B(_15055__bF_buf6), .S(_8476__bF_buf0), .Y(_223__10_) );
INVX1 INVX1_3742 ( .gnd(gnd), .vdd(vdd), .A(data_6__11_), .Y(_8489_) );
MUX2X1 MUX2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_8489_), .B(_14918__bF_buf7), .S(_8476__bF_buf3), .Y(_223__11_) );
INVX1 INVX1_3743 ( .gnd(gnd), .vdd(vdd), .A(data_6__12_), .Y(_8490_) );
MUX2X1 MUX2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_8490_), .B(_14920__bF_buf8), .S(_8476__bF_buf2), .Y(_223__12_) );
INVX1 INVX1_3744 ( .gnd(gnd), .vdd(vdd), .A(data_6__13_), .Y(_8491_) );
MUX2X1 MUX2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_8491_), .B(_14924__bF_buf6), .S(_8476__bF_buf1), .Y(_223__13_) );
INVX1 INVX1_3745 ( .gnd(gnd), .vdd(vdd), .A(data_6__14_), .Y(_8492_) );
MUX2X1 MUX2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_8492_), .B(_15060__bF_buf5), .S(_8476__bF_buf0), .Y(_223__14_) );
INVX1 INVX1_3746 ( .gnd(gnd), .vdd(vdd), .A(data_6__15_), .Y(_8493_) );
MUX2X1 MUX2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_8493_), .B(_15062__bF_buf9), .S(_8476__bF_buf3), .Y(_223__15_) );
INVX1 INVX1_3747 ( .gnd(gnd), .vdd(vdd), .A(data_5__0_), .Y(_8494_) );
INVX1 INVX1_3748 ( .gnd(gnd), .vdd(vdd), .A(_15015_), .Y(_8495_) );
OAI21X1 OAI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_14947_), .B(_14882__bF_buf4), .C(_8299_), .Y(_8496_) );
NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_8496_), .B(_8473_), .Y(_8497_) );
NOR3X1 NOR3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_8495_), .B(_8497_), .C(_8126_), .Y(_8498_) );
AND2X2 AND2X2_1510 ( .gnd(gnd), .vdd(vdd), .A(_8125__bF_buf2), .B(_8498_), .Y(_8499_) );
MUX2X1 MUX2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf4), .B(_8494_), .S(_8499_), .Y(_212__0_) );
INVX1 INVX1_3749 ( .gnd(gnd), .vdd(vdd), .A(data_5__1_), .Y(_8500_) );
MUX2X1 MUX2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf3), .B(_8500_), .S(_8499_), .Y(_212__1_) );
AOI21X1 AOI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf1), .C(data_5__2_), .Y(_8501_) );
AOI21X1 AOI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf12), .B(_8499_), .C(_8501_), .Y(_212__2_) );
INVX1 INVX1_3750 ( .gnd(gnd), .vdd(vdd), .A(data_5__3_), .Y(_8502_) );
MUX2X1 MUX2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf2), .B(_8502_), .S(_8499_), .Y(_212__3_) );
INVX1 INVX1_3751 ( .gnd(gnd), .vdd(vdd), .A(data_5__4_), .Y(_8503_) );
MUX2X1 MUX2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf7), .B(_8503_), .S(_8499_), .Y(_212__4_) );
INVX1 INVX1_3752 ( .gnd(gnd), .vdd(vdd), .A(data_5__5_), .Y(_8504_) );
MUX2X1 MUX2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf5), .B(_8504_), .S(_8499_), .Y(_212__5_) );
AOI21X1 AOI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf0), .C(data_5__6_), .Y(_8505_) );
AOI21X1 AOI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf2), .B(_8499_), .C(_8505_), .Y(_212__6_) );
INVX1 INVX1_3753 ( .gnd(gnd), .vdd(vdd), .A(data_5__7_), .Y(_8506_) );
MUX2X1 MUX2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf8), .B(_8506_), .S(_8499_), .Y(_212__7_) );
AOI21X1 AOI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf5), .C(data_5__8_), .Y(_8507_) );
AOI21X1 AOI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf4), .B(_8499_), .C(_8507_), .Y(_212__8_) );
AOI21X1 AOI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf4), .C(data_5__9_), .Y(_8508_) );
AOI21X1 AOI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf14), .B(_8499_), .C(_8508_), .Y(_212__9_) );
AOI21X1 AOI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf3), .C(data_5__10_), .Y(_8509_) );
AOI21X1 AOI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf5), .B(_8499_), .C(_8509_), .Y(_212__10_) );
INVX1 INVX1_3754 ( .gnd(gnd), .vdd(vdd), .A(data_5__11_), .Y(_8510_) );
MUX2X1 MUX2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf6), .B(_8510_), .S(_8499_), .Y(_212__11_) );
INVX1 INVX1_3755 ( .gnd(gnd), .vdd(vdd), .A(data_5__12_), .Y(_8511_) );
MUX2X1 MUX2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf7), .B(_8511_), .S(_8499_), .Y(_212__12_) );
AOI21X1 AOI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf2), .C(data_5__13_), .Y(_8512_) );
AOI21X1 AOI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf5), .B(_8499_), .C(_8512_), .Y(_212__13_) );
AOI21X1 AOI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf1), .C(data_5__14_), .Y(_8513_) );
AOI21X1 AOI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf4), .B(_8499_), .C(_8513_), .Y(_212__14_) );
AOI21X1 AOI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_8498_), .B(_8125__bF_buf0), .C(data_5__15_), .Y(_8514_) );
AOI21X1 AOI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf8), .B(_8499_), .C(_8514_), .Y(_212__15_) );
INVX1 INVX1_3756 ( .gnd(gnd), .vdd(vdd), .A(data_4__0_), .Y(_8515_) );
NAND3X1 NAND3X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_15507_), .B(_15514_), .C(_15183__bF_buf3), .Y(_8516_) );
NOR3X1 NOR3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_3306__bF_buf4), .B(_3308_), .C(_8516_), .Y(_8517_) );
MUX2X1 MUX2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf3), .B(_8515_), .S(_8517_), .Y(_201__0_) );
INVX1 INVX1_3757 ( .gnd(gnd), .vdd(vdd), .A(data_4__1_), .Y(_8518_) );
MUX2X1 MUX2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf2), .B(_8518_), .S(_8517_), .Y(_201__1_) );
INVX1 INVX1_3758 ( .gnd(gnd), .vdd(vdd), .A(data_4__2_), .Y(_8519_) );
MUX2X1 MUX2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf11), .B(_8519_), .S(_8517_), .Y(_201__2_) );
INVX1 INVX1_3759 ( .gnd(gnd), .vdd(vdd), .A(data_4__3_), .Y(_8520_) );
MUX2X1 MUX2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf1), .B(_8520_), .S(_8517_), .Y(_201__3_) );
INVX1 INVX1_3760 ( .gnd(gnd), .vdd(vdd), .A(data_4__4_), .Y(_8521_) );
MUX2X1 MUX2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf6), .B(_8521_), .S(_8517_), .Y(_201__4_) );
INVX1 INVX1_3761 ( .gnd(gnd), .vdd(vdd), .A(data_4__5_), .Y(_8522_) );
MUX2X1 MUX2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf4), .B(_8522_), .S(_8517_), .Y(_201__5_) );
INVX1 INVX1_3762 ( .gnd(gnd), .vdd(vdd), .A(data_4__6_), .Y(_8523_) );
MUX2X1 MUX2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf1), .B(_8523_), .S(_8517_), .Y(_201__6_) );
INVX1 INVX1_3763 ( .gnd(gnd), .vdd(vdd), .A(data_4__7_), .Y(_8524_) );
MUX2X1 MUX2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf7), .B(_8524_), .S(_8517_), .Y(_201__7_) );
INVX1 INVX1_3764 ( .gnd(gnd), .vdd(vdd), .A(data_4__8_), .Y(_8525_) );
MUX2X1 MUX2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf3), .B(_8525_), .S(_8517_), .Y(_201__8_) );
INVX1 INVX1_3765 ( .gnd(gnd), .vdd(vdd), .A(data_4__9_), .Y(_8526_) );
MUX2X1 MUX2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf13), .B(_8526_), .S(_8517_), .Y(_201__9_) );
INVX1 INVX1_3766 ( .gnd(gnd), .vdd(vdd), .A(data_4__10_), .Y(_8527_) );
MUX2X1 MUX2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf4), .B(_8527_), .S(_8517_), .Y(_201__10_) );
INVX1 INVX1_3767 ( .gnd(gnd), .vdd(vdd), .A(data_4__11_), .Y(_8528_) );
MUX2X1 MUX2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf5), .B(_8528_), .S(_8517_), .Y(_201__11_) );
INVX1 INVX1_3768 ( .gnd(gnd), .vdd(vdd), .A(data_4__12_), .Y(_8529_) );
MUX2X1 MUX2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf6), .B(_8529_), .S(_8517_), .Y(_201__12_) );
INVX1 INVX1_3769 ( .gnd(gnd), .vdd(vdd), .A(data_4__13_), .Y(_8530_) );
MUX2X1 MUX2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf4), .B(_8530_), .S(_8517_), .Y(_201__13_) );
INVX1 INVX1_3770 ( .gnd(gnd), .vdd(vdd), .A(data_4__14_), .Y(_8531_) );
MUX2X1 MUX2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf3), .B(_8531_), .S(_8517_), .Y(_201__14_) );
INVX1 INVX1_3771 ( .gnd(gnd), .vdd(vdd), .A(data_4__15_), .Y(_8532_) );
MUX2X1 MUX2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf7), .B(_8532_), .S(_8517_), .Y(_201__15_) );
INVX1 INVX1_3772 ( .gnd(gnd), .vdd(vdd), .A(data_3__0_), .Y(_8533_) );
INVX1 INVX1_3773 ( .gnd(gnd), .vdd(vdd), .A(_15123_), .Y(_8534_) );
OAI21X1 OAI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_15572_), .B(_15580_), .C(_15011__bF_buf3), .Y(_8535_) );
NAND3X1 NAND3X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_8534_), .B(_8535_), .C(_15507_), .Y(_8536_) );
INVX1 INVX1_3774 ( .gnd(gnd), .vdd(vdd), .A(_8536_), .Y(_8537_) );
NAND3X1 NAND3X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_3309_), .B(_15183__bF_buf2), .C(_8537_), .Y(_8538_) );
OAI21X1 OAI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf3), .C(_8533_), .Y(_8539_) );
NOR3X1 NOR3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_8084_), .B(_8536_), .C(_15074__bF_buf8), .Y(_8540_) );
NAND3X1 NAND3X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf2), .B(_8540_), .C(_3391__bF_buf0), .Y(_8541_) );
AND2X2 AND2X2_1511 ( .gnd(gnd), .vdd(vdd), .A(_8539_), .B(_8541_), .Y(_190__0_) );
INVX1 INVX1_3775 ( .gnd(gnd), .vdd(vdd), .A(data_3__1_), .Y(_8542_) );
OAI21X1 OAI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf2), .C(_8542_), .Y(_8543_) );
NAND3X1 NAND3X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf1), .B(_8540_), .C(_3391__bF_buf6), .Y(_8544_) );
AND2X2 AND2X2_1512 ( .gnd(gnd), .vdd(vdd), .A(_8543_), .B(_8544_), .Y(_190__1_) );
INVX1 INVX1_3776 ( .gnd(gnd), .vdd(vdd), .A(data_3__2_), .Y(_8545_) );
OAI21X1 OAI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf1), .C(_8545_), .Y(_8546_) );
NAND3X1 NAND3X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf10), .B(_8540_), .C(_3391__bF_buf5), .Y(_8547_) );
AND2X2 AND2X2_1513 ( .gnd(gnd), .vdd(vdd), .A(_8546_), .B(_8547_), .Y(_190__2_) );
INVX1 INVX1_3777 ( .gnd(gnd), .vdd(vdd), .A(data_3__3_), .Y(_8548_) );
OAI21X1 OAI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf0), .C(_8548_), .Y(_8549_) );
NAND3X1 NAND3X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf0), .B(_8540_), .C(_3391__bF_buf4), .Y(_8550_) );
AND2X2 AND2X2_1514 ( .gnd(gnd), .vdd(vdd), .A(_8549_), .B(_8550_), .Y(_190__3_) );
INVX1 INVX1_3778 ( .gnd(gnd), .vdd(vdd), .A(data_3__4_), .Y(_8551_) );
OAI21X1 OAI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf6), .C(_8551_), .Y(_8552_) );
NAND3X1 NAND3X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf5), .B(_8540_), .C(_3391__bF_buf3), .Y(_8553_) );
AND2X2 AND2X2_1515 ( .gnd(gnd), .vdd(vdd), .A(_8552_), .B(_8553_), .Y(_190__4_) );
INVX1 INVX1_3779 ( .gnd(gnd), .vdd(vdd), .A(data_3__5_), .Y(_8554_) );
OAI21X1 OAI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf5), .C(_8554_), .Y(_8555_) );
NAND3X1 NAND3X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf3), .B(_8540_), .C(_3391__bF_buf2), .Y(_8556_) );
AND2X2 AND2X2_1516 ( .gnd(gnd), .vdd(vdd), .A(_8555_), .B(_8556_), .Y(_190__5_) );
INVX1 INVX1_3780 ( .gnd(gnd), .vdd(vdd), .A(data_3__6_), .Y(_8557_) );
OAI21X1 OAI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf4), .C(_8557_), .Y(_8558_) );
NAND3X1 NAND3X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf0), .B(_8540_), .C(_3391__bF_buf1), .Y(_8559_) );
AND2X2 AND2X2_1517 ( .gnd(gnd), .vdd(vdd), .A(_8558_), .B(_8559_), .Y(_190__6_) );
INVX1 INVX1_3781 ( .gnd(gnd), .vdd(vdd), .A(data_3__7_), .Y(_8560_) );
OAI21X1 OAI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf3), .C(_8560_), .Y(_8561_) );
NAND3X1 NAND3X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf6), .B(_8540_), .C(_3391__bF_buf0), .Y(_8562_) );
AND2X2 AND2X2_1518 ( .gnd(gnd), .vdd(vdd), .A(_8561_), .B(_8562_), .Y(_190__7_) );
INVX1 INVX1_3782 ( .gnd(gnd), .vdd(vdd), .A(data_3__8_), .Y(_8563_) );
OAI21X1 OAI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf2), .C(_8563_), .Y(_8564_) );
NAND3X1 NAND3X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf2), .B(_8540_), .C(_3391__bF_buf6), .Y(_8565_) );
AND2X2 AND2X2_1519 ( .gnd(gnd), .vdd(vdd), .A(_8564_), .B(_8565_), .Y(_190__8_) );
INVX1 INVX1_3783 ( .gnd(gnd), .vdd(vdd), .A(data_3__9_), .Y(_8566_) );
OAI21X1 OAI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf1), .C(_8566_), .Y(_8567_) );
NAND3X1 NAND3X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf12), .B(_8540_), .C(_3391__bF_buf5), .Y(_8568_) );
AND2X2 AND2X2_1520 ( .gnd(gnd), .vdd(vdd), .A(_8567_), .B(_8568_), .Y(_190__9_) );
INVX1 INVX1_3784 ( .gnd(gnd), .vdd(vdd), .A(data_3__10_), .Y(_8569_) );
OAI21X1 OAI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf0), .C(_8569_), .Y(_8570_) );
NAND3X1 NAND3X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf3), .B(_8540_), .C(_3391__bF_buf4), .Y(_8571_) );
AND2X2 AND2X2_1521 ( .gnd(gnd), .vdd(vdd), .A(_8570_), .B(_8571_), .Y(_190__10_) );
INVX1 INVX1_3785 ( .gnd(gnd), .vdd(vdd), .A(data_3__11_), .Y(_8572_) );
OAI21X1 OAI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf6), .C(_8572_), .Y(_8573_) );
NAND3X1 NAND3X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf4), .B(_8540_), .C(_3391__bF_buf3), .Y(_8574_) );
AND2X2 AND2X2_1522 ( .gnd(gnd), .vdd(vdd), .A(_8573_), .B(_8574_), .Y(_190__11_) );
INVX1 INVX1_3786 ( .gnd(gnd), .vdd(vdd), .A(data_3__12_), .Y(_8575_) );
OAI21X1 OAI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf5), .C(_8575_), .Y(_8576_) );
NAND3X1 NAND3X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf5), .B(_8540_), .C(_3391__bF_buf2), .Y(_8577_) );
AND2X2 AND2X2_1523 ( .gnd(gnd), .vdd(vdd), .A(_8576_), .B(_8577_), .Y(_190__12_) );
INVX1 INVX1_3787 ( .gnd(gnd), .vdd(vdd), .A(data_3__13_), .Y(_8578_) );
OAI21X1 OAI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf4), .C(_8578_), .Y(_8579_) );
NAND3X1 NAND3X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf3), .B(_8540_), .C(_3391__bF_buf1), .Y(_8580_) );
AND2X2 AND2X2_1524 ( .gnd(gnd), .vdd(vdd), .A(_8579_), .B(_8580_), .Y(_190__13_) );
INVX1 INVX1_3788 ( .gnd(gnd), .vdd(vdd), .A(data_3__14_), .Y(_8581_) );
OAI21X1 OAI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf3), .C(_8581_), .Y(_8582_) );
NAND3X1 NAND3X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf2), .B(_8540_), .C(_3391__bF_buf0), .Y(_8583_) );
AND2X2 AND2X2_1525 ( .gnd(gnd), .vdd(vdd), .A(_8582_), .B(_8583_), .Y(_190__14_) );
INVX1 INVX1_3789 ( .gnd(gnd), .vdd(vdd), .A(data_3__15_), .Y(_8584_) );
OAI21X1 OAI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_8538_), .B(_3306__bF_buf2), .C(_8584_), .Y(_8585_) );
NAND3X1 NAND3X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf6), .B(_8540_), .C(_3391__bF_buf6), .Y(_8586_) );
AND2X2 AND2X2_1526 ( .gnd(gnd), .vdd(vdd), .A(_8585_), .B(_8586_), .Y(_190__15_) );
INVX1 INVX1_3790 ( .gnd(gnd), .vdd(vdd), .A(data_2__0_), .Y(_8587_) );
INVX1 INVX1_3791 ( .gnd(gnd), .vdd(vdd), .A(_7538_), .Y(_8588_) );
AOI21X1 AOI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_15011__bF_buf2), .B(_8588_), .C(_15123_), .Y(_8589_) );
AND2X2 AND2X2_1527 ( .gnd(gnd), .vdd(vdd), .A(_8589_), .B(_15018_), .Y(_8590_) );
NAND3X1 NAND3X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_15120__bF_buf1), .B(_8590_), .C(_15183__bF_buf1), .Y(_8591_) );
OAI21X1 OAI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf1), .C(_8587_), .Y(_8592_) );
NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_15018_), .B(_8589_), .Y(_8593_) );
NOR3X1 NOR3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_8593_), .B(_15028_), .C(_15074__bF_buf7), .Y(_8594_) );
NAND3X1 NAND3X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf1), .B(_8594_), .C(_3391__bF_buf5), .Y(_8595_) );
AND2X2 AND2X2_1528 ( .gnd(gnd), .vdd(vdd), .A(_8595_), .B(_8592_), .Y(_179__0_) );
INVX1 INVX1_3792 ( .gnd(gnd), .vdd(vdd), .A(data_2__1_), .Y(_8596_) );
OAI21X1 OAI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf0), .C(_8596_), .Y(_8597_) );
NAND3X1 NAND3X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf0), .B(_8594_), .C(_3391__bF_buf4), .Y(_8598_) );
AND2X2 AND2X2_1529 ( .gnd(gnd), .vdd(vdd), .A(_8598_), .B(_8597_), .Y(_179__1_) );
INVX1 INVX1_3793 ( .gnd(gnd), .vdd(vdd), .A(data_2__2_), .Y(_8599_) );
OAI21X1 OAI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf6), .C(_8599_), .Y(_8600_) );
NAND3X1 NAND3X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf9), .B(_8594_), .C(_3391__bF_buf3), .Y(_8601_) );
AND2X2 AND2X2_1530 ( .gnd(gnd), .vdd(vdd), .A(_8601_), .B(_8600_), .Y(_179__2_) );
INVX1 INVX1_3794 ( .gnd(gnd), .vdd(vdd), .A(data_2__3_), .Y(_8602_) );
OAI21X1 OAI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf5), .C(_8602_), .Y(_8603_) );
NAND3X1 NAND3X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf14), .B(_8594_), .C(_3391__bF_buf2), .Y(_8604_) );
AND2X2 AND2X2_1531 ( .gnd(gnd), .vdd(vdd), .A(_8604_), .B(_8603_), .Y(_179__3_) );
INVX1 INVX1_3795 ( .gnd(gnd), .vdd(vdd), .A(data_2__4_), .Y(_8605_) );
OAI21X1 OAI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf4), .C(_8605_), .Y(_8606_) );
NAND3X1 NAND3X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf4), .B(_8594_), .C(_3391__bF_buf1), .Y(_8607_) );
AND2X2 AND2X2_1532 ( .gnd(gnd), .vdd(vdd), .A(_8607_), .B(_8606_), .Y(_179__4_) );
INVX1 INVX1_3796 ( .gnd(gnd), .vdd(vdd), .A(data_2__5_), .Y(_8608_) );
OAI21X1 OAI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf3), .C(_8608_), .Y(_8609_) );
NAND3X1 NAND3X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf2), .B(_8594_), .C(_3391__bF_buf0), .Y(_8610_) );
AND2X2 AND2X2_1533 ( .gnd(gnd), .vdd(vdd), .A(_8610_), .B(_8609_), .Y(_179__5_) );
INVX1 INVX1_3797 ( .gnd(gnd), .vdd(vdd), .A(data_2__6_), .Y(_8611_) );
OAI21X1 OAI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf2), .C(_8611_), .Y(_8612_) );
NAND3X1 NAND3X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf14), .B(_8594_), .C(_3391__bF_buf6), .Y(_8613_) );
AND2X2 AND2X2_1534 ( .gnd(gnd), .vdd(vdd), .A(_8613_), .B(_8612_), .Y(_179__6_) );
INVX1 INVX1_3798 ( .gnd(gnd), .vdd(vdd), .A(data_2__7_), .Y(_8614_) );
OAI21X1 OAI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf1), .C(_8614_), .Y(_8615_) );
NAND3X1 NAND3X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf5), .B(_8594_), .C(_3391__bF_buf5), .Y(_8616_) );
AND2X2 AND2X2_1535 ( .gnd(gnd), .vdd(vdd), .A(_8616_), .B(_8615_), .Y(_179__7_) );
INVX1 INVX1_3799 ( .gnd(gnd), .vdd(vdd), .A(data_2__8_), .Y(_8617_) );
OAI21X1 OAI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf0), .C(_8617_), .Y(_8618_) );
NAND3X1 NAND3X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf1), .B(_8594_), .C(_3391__bF_buf4), .Y(_8619_) );
AND2X2 AND2X2_1536 ( .gnd(gnd), .vdd(vdd), .A(_8619_), .B(_8618_), .Y(_179__8_) );
INVX1 INVX1_3800 ( .gnd(gnd), .vdd(vdd), .A(data_2__9_), .Y(_8620_) );
OAI21X1 OAI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf6), .C(_8620_), .Y(_8621_) );
NAND3X1 NAND3X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf11), .B(_8594_), .C(_3391__bF_buf3), .Y(_8622_) );
AND2X2 AND2X2_1537 ( .gnd(gnd), .vdd(vdd), .A(_8622_), .B(_8621_), .Y(_179__9_) );
INVX1 INVX1_3801 ( .gnd(gnd), .vdd(vdd), .A(data_2__10_), .Y(_8623_) );
OAI21X1 OAI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf5), .C(_8623_), .Y(_8624_) );
NAND3X1 NAND3X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf2), .B(_8594_), .C(_3391__bF_buf2), .Y(_8625_) );
AND2X2 AND2X2_1538 ( .gnd(gnd), .vdd(vdd), .A(_8625_), .B(_8624_), .Y(_179__10_) );
INVX1 INVX1_3802 ( .gnd(gnd), .vdd(vdd), .A(data_2__11_), .Y(_8626_) );
OAI21X1 OAI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf4), .C(_8626_), .Y(_8627_) );
NAND3X1 NAND3X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf3), .B(_8594_), .C(_3391__bF_buf1), .Y(_8628_) );
AND2X2 AND2X2_1539 ( .gnd(gnd), .vdd(vdd), .A(_8628_), .B(_8627_), .Y(_179__11_) );
INVX1 INVX1_3803 ( .gnd(gnd), .vdd(vdd), .A(data_2__12_), .Y(_8629_) );
OAI21X1 OAI21X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf3), .C(_8629_), .Y(_8630_) );
NAND3X1 NAND3X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf4), .B(_8594_), .C(_3391__bF_buf0), .Y(_8631_) );
AND2X2 AND2X2_1540 ( .gnd(gnd), .vdd(vdd), .A(_8631_), .B(_8630_), .Y(_179__12_) );
INVX1 INVX1_3804 ( .gnd(gnd), .vdd(vdd), .A(data_2__13_), .Y(_8632_) );
OAI21X1 OAI21X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf2), .C(_8632_), .Y(_8633_) );
NAND3X1 NAND3X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf2), .B(_8594_), .C(_3391__bF_buf6), .Y(_8634_) );
AND2X2 AND2X2_1541 ( .gnd(gnd), .vdd(vdd), .A(_8634_), .B(_8633_), .Y(_179__13_) );
INVX1 INVX1_3805 ( .gnd(gnd), .vdd(vdd), .A(data_2__14_), .Y(_8635_) );
OAI21X1 OAI21X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf1), .C(_8635_), .Y(_8636_) );
NAND3X1 NAND3X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf1), .B(_8594_), .C(_3391__bF_buf5), .Y(_8637_) );
AND2X2 AND2X2_1542 ( .gnd(gnd), .vdd(vdd), .A(_8637_), .B(_8636_), .Y(_179__14_) );
INVX1 INVX1_3806 ( .gnd(gnd), .vdd(vdd), .A(data_2__15_), .Y(_8638_) );
OAI21X1 OAI21X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_8591_), .B(_3306__bF_buf0), .C(_8638_), .Y(_8639_) );
NAND3X1 NAND3X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf5), .B(_8594_), .C(_3391__bF_buf4), .Y(_8640_) );
AND2X2 AND2X2_1543 ( .gnd(gnd), .vdd(vdd), .A(_8640_), .B(_8639_), .Y(_179__15_) );
INVX1 INVX1_3807 ( .gnd(gnd), .vdd(vdd), .A(data_1__0_), .Y(_8641_) );
INVX1 INVX1_3808 ( .gnd(gnd), .vdd(vdd), .A(_7575_), .Y(_8642_) );
AOI21X1 AOI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_15011__bF_buf1), .B(_8642_), .C(_15123_), .Y(_8643_) );
NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_8643_), .B(_15018_), .Y(_8644_) );
INVX1 INVX1_3809 ( .gnd(gnd), .vdd(vdd), .A(_8644_), .Y(_8645_) );
NAND3X1 NAND3X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_15183__bF_buf0), .B(_15120__bF_buf0), .C(_8645_), .Y(_8646_) );
OAI21X1 OAI21X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf6), .C(_8641_), .Y(_8647_) );
NOR3X1 NOR3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_15028_), .B(_8644_), .C(_15074__bF_buf6), .Y(_8648_) );
NAND3X1 NAND3X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_14932__bF_buf0), .B(_8648_), .C(_3391__bF_buf3), .Y(_8649_) );
AND2X2 AND2X2_1544 ( .gnd(gnd), .vdd(vdd), .A(_8647_), .B(_8649_), .Y(_112__0_) );
INVX1 INVX1_3810 ( .gnd(gnd), .vdd(vdd), .A(data_1__1_), .Y(_8650_) );
OAI21X1 OAI21X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf5), .C(_8650_), .Y(_8651_) );
NAND3X1 NAND3X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_14894__bF_buf14), .B(_8648_), .C(_3391__bF_buf2), .Y(_8652_) );
AND2X2 AND2X2_1545 ( .gnd(gnd), .vdd(vdd), .A(_8651_), .B(_8652_), .Y(_112__1_) );
INVX1 INVX1_3811 ( .gnd(gnd), .vdd(vdd), .A(data_1__2_), .Y(_8653_) );
OAI21X1 OAI21X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf4), .C(_8653_), .Y(_8654_) );
NAND3X1 NAND3X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_14897__bF_buf8), .B(_8648_), .C(_3391__bF_buf1), .Y(_8655_) );
AND2X2 AND2X2_1546 ( .gnd(gnd), .vdd(vdd), .A(_8654_), .B(_8655_), .Y(_112__2_) );
INVX1 INVX1_3812 ( .gnd(gnd), .vdd(vdd), .A(data_1__3_), .Y(_8656_) );
OAI21X1 OAI21X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf3), .C(_8656_), .Y(_8657_) );
NAND3X1 NAND3X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_14899__bF_buf13), .B(_8648_), .C(_3391__bF_buf0), .Y(_8658_) );
AND2X2 AND2X2_1547 ( .gnd(gnd), .vdd(vdd), .A(_8657_), .B(_8658_), .Y(_112__3_) );
INVX1 INVX1_3813 ( .gnd(gnd), .vdd(vdd), .A(data_1__4_), .Y(_8659_) );
OAI21X1 OAI21X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf2), .C(_8659_), .Y(_8660_) );
NAND3X1 NAND3X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_14902__bF_buf3), .B(_8648_), .C(_3391__bF_buf6), .Y(_8661_) );
AND2X2 AND2X2_1548 ( .gnd(gnd), .vdd(vdd), .A(_8660_), .B(_8661_), .Y(_112__4_) );
INVX1 INVX1_3814 ( .gnd(gnd), .vdd(vdd), .A(data_1__5_), .Y(_8662_) );
OAI21X1 OAI21X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf1), .C(_8662_), .Y(_8663_) );
NAND3X1 NAND3X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_14903__bF_buf1), .B(_8648_), .C(_3391__bF_buf5), .Y(_8664_) );
AND2X2 AND2X2_1549 ( .gnd(gnd), .vdd(vdd), .A(_8663_), .B(_8664_), .Y(_112__5_) );
INVX1 INVX1_3815 ( .gnd(gnd), .vdd(vdd), .A(data_1__6_), .Y(_8665_) );
OAI21X1 OAI21X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf0), .C(_8665_), .Y(_8666_) );
NAND3X1 NAND3X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_15049__bF_buf13), .B(_8648_), .C(_3391__bF_buf4), .Y(_8667_) );
AND2X2 AND2X2_1550 ( .gnd(gnd), .vdd(vdd), .A(_8666_), .B(_8667_), .Y(_112__6_) );
INVX1 INVX1_3816 ( .gnd(gnd), .vdd(vdd), .A(data_1__7_), .Y(_8668_) );
OAI21X1 OAI21X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf6), .C(_8668_), .Y(_8669_) );
NAND3X1 NAND3X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_14908__bF_buf4), .B(_8648_), .C(_3391__bF_buf3), .Y(_8670_) );
AND2X2 AND2X2_1551 ( .gnd(gnd), .vdd(vdd), .A(_8669_), .B(_8670_), .Y(_112__7_) );
INVX1 INVX1_3817 ( .gnd(gnd), .vdd(vdd), .A(data_1__8_), .Y(_8671_) );
OAI21X1 OAI21X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf5), .C(_8671_), .Y(_8672_) );
NAND3X1 NAND3X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_15052__bF_buf0), .B(_8648_), .C(_3391__bF_buf2), .Y(_8673_) );
AND2X2 AND2X2_1552 ( .gnd(gnd), .vdd(vdd), .A(_8672_), .B(_8673_), .Y(_112__8_) );
INVX1 INVX1_3818 ( .gnd(gnd), .vdd(vdd), .A(data_1__9_), .Y(_8674_) );
OAI21X1 OAI21X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf4), .C(_8674_), .Y(_8675_) );
NAND3X1 NAND3X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_14913__bF_buf10), .B(_8648_), .C(_3391__bF_buf1), .Y(_8676_) );
AND2X2 AND2X2_1553 ( .gnd(gnd), .vdd(vdd), .A(_8675_), .B(_8676_), .Y(_112__9_) );
INVX1 INVX1_3819 ( .gnd(gnd), .vdd(vdd), .A(data_1__10_), .Y(_8677_) );
OAI21X1 OAI21X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf3), .C(_8677_), .Y(_8678_) );
NAND3X1 NAND3X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_15055__bF_buf1), .B(_8648_), .C(_3391__bF_buf0), .Y(_8679_) );
AND2X2 AND2X2_1554 ( .gnd(gnd), .vdd(vdd), .A(_8678_), .B(_8679_), .Y(_112__10_) );
INVX1 INVX1_3820 ( .gnd(gnd), .vdd(vdd), .A(data_1__11_), .Y(_8680_) );
OAI21X1 OAI21X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf2), .C(_8680_), .Y(_8681_) );
NAND3X1 NAND3X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_14918__bF_buf2), .B(_8648_), .C(_3391__bF_buf6), .Y(_8682_) );
AND2X2 AND2X2_1555 ( .gnd(gnd), .vdd(vdd), .A(_8681_), .B(_8682_), .Y(_112__11_) );
INVX1 INVX1_3821 ( .gnd(gnd), .vdd(vdd), .A(data_1__12_), .Y(_8683_) );
OAI21X1 OAI21X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf1), .C(_8683_), .Y(_8684_) );
NAND3X1 NAND3X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_14920__bF_buf3), .B(_8648_), .C(_3391__bF_buf5), .Y(_8685_) );
AND2X2 AND2X2_1556 ( .gnd(gnd), .vdd(vdd), .A(_8684_), .B(_8685_), .Y(_112__12_) );
INVX1 INVX1_3822 ( .gnd(gnd), .vdd(vdd), .A(data_1__13_), .Y(_8686_) );
OAI21X1 OAI21X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf0), .C(_8686_), .Y(_8687_) );
NAND3X1 NAND3X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_14924__bF_buf1), .B(_8648_), .C(_3391__bF_buf4), .Y(_8688_) );
AND2X2 AND2X2_1557 ( .gnd(gnd), .vdd(vdd), .A(_8687_), .B(_8688_), .Y(_112__13_) );
INVX1 INVX1_3823 ( .gnd(gnd), .vdd(vdd), .A(data_1__14_), .Y(_8689_) );
OAI21X1 OAI21X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf6), .C(_8689_), .Y(_8690_) );
NAND3X1 NAND3X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_15060__bF_buf0), .B(_8648_), .C(_3391__bF_buf3), .Y(_8691_) );
AND2X2 AND2X2_1558 ( .gnd(gnd), .vdd(vdd), .A(_8690_), .B(_8691_), .Y(_112__14_) );
INVX1 INVX1_3824 ( .gnd(gnd), .vdd(vdd), .A(data_1__15_), .Y(_8692_) );
OAI21X1 OAI21X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_8646_), .B(_3306__bF_buf5), .C(_8692_), .Y(_8693_) );
NAND3X1 NAND3X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_15062__bF_buf4), .B(_8648_), .C(_3391__bF_buf2), .Y(_8694_) );
AND2X2 AND2X2_1559 ( .gnd(gnd), .vdd(vdd), .A(_8693_), .B(_8694_), .Y(_112__15_) );
INVX1 INVX1_3825 ( .gnd(gnd), .vdd(vdd), .A(data_0__0_), .Y(_8695_) );
NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_write_bF_buf1), .B(_15032_), .Y(_8696_) );
MUX2X1 MUX2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_8695_), .B(_14932__bF_buf14), .S(_8696_), .Y(_1__0_) );
INVX1 INVX1_3826 ( .gnd(gnd), .vdd(vdd), .A(data_0__1_), .Y(_8697_) );
OAI21X1 OAI21X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf3), .C(_8697_), .Y(_8698_) );
OAI21X1 OAI21X1_2367 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_1_bF_buf4), .B(_8696_), .C(_8698_), .Y(_8699_) );
INVX1 INVX1_3827 ( .gnd(gnd), .vdd(vdd), .A(_8699_), .Y(_1__1_) );
INVX1 INVX1_3828 ( .gnd(gnd), .vdd(vdd), .A(data_0__2_), .Y(_8700_) );
MUX2X1 MUX2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_8700_), .B(_14897__bF_buf7), .S(_8696_), .Y(_1__2_) );
INVX1 INVX1_3829 ( .gnd(gnd), .vdd(vdd), .A(data_0__3_), .Y(_8701_) );
MUX2X1 MUX2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_8701_), .B(_14899__bF_buf12), .S(_8696_), .Y(_1__3_) );
INVX1 INVX1_3830 ( .gnd(gnd), .vdd(vdd), .A(data_0__4_), .Y(_8702_) );
MUX2X1 MUX2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_8702_), .B(_14902__bF_buf2), .S(_8696_), .Y(_1__4_) );
INVX1 INVX1_3831 ( .gnd(gnd), .vdd(vdd), .A(data_0__5_), .Y(_8703_) );
MUX2X1 MUX2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_8703_), .B(_14903__bF_buf0), .S(_8696_), .Y(_1__5_) );
INVX1 INVX1_3832 ( .gnd(gnd), .vdd(vdd), .A(data_0__6_), .Y(_8704_) );
OAI21X1 OAI21X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf2), .C(_8704_), .Y(_8705_) );
OAI21X1 OAI21X1_2369 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_6_bF_buf0), .B(_8696_), .C(_8705_), .Y(_8706_) );
INVX1 INVX1_3833 ( .gnd(gnd), .vdd(vdd), .A(_8706_), .Y(_1__6_) );
INVX1 INVX1_3834 ( .gnd(gnd), .vdd(vdd), .A(data_0__7_), .Y(_8707_) );
MUX2X1 MUX2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_8707_), .B(_14908__bF_buf3), .S(_8696_), .Y(_1__7_) );
INVX1 INVX1_3835 ( .gnd(gnd), .vdd(vdd), .A(data_0__8_), .Y(_8708_) );
OAI21X1 OAI21X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf1), .C(_8708_), .Y(_8709_) );
OAI21X1 OAI21X1_2371 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_8_bF_buf2), .B(_8696_), .C(_8709_), .Y(_8710_) );
INVX1 INVX1_3836 ( .gnd(gnd), .vdd(vdd), .A(_8710_), .Y(_1__8_) );
INVX1 INVX1_3837 ( .gnd(gnd), .vdd(vdd), .A(data_0__9_), .Y(_8711_) );
OAI21X1 OAI21X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf0), .C(_8711_), .Y(_8712_) );
OAI21X1 OAI21X1_2373 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_9_bF_buf3), .B(_8696_), .C(_8712_), .Y(_8713_) );
INVX1 INVX1_3838 ( .gnd(gnd), .vdd(vdd), .A(_8713_), .Y(_1__9_) );
INVX1 INVX1_3839 ( .gnd(gnd), .vdd(vdd), .A(data_0__10_), .Y(_8714_) );
OAI21X1 OAI21X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf15_bF_buf3), .C(_8714_), .Y(_8715_) );
OAI21X1 OAI21X1_2375 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_10_bF_buf1), .B(_8696_), .C(_8715_), .Y(_8716_) );
INVX1 INVX1_3840 ( .gnd(gnd), .vdd(vdd), .A(_8716_), .Y(_1__10_) );
INVX1 INVX1_3841 ( .gnd(gnd), .vdd(vdd), .A(data_0__11_), .Y(_8717_) );
MUX2X1 MUX2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_8717_), .B(_14918__bF_buf1), .S(_8696_), .Y(_1__11_) );
INVX1 INVX1_3842 ( .gnd(gnd), .vdd(vdd), .A(data_0__12_), .Y(_8718_) );
MUX2X1 MUX2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_8718_), .B(_14920__bF_buf2), .S(_8696_), .Y(_1__12_) );
INVX1 INVX1_3843 ( .gnd(gnd), .vdd(vdd), .A(data_0__13_), .Y(_8719_) );
MUX2X1 MUX2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_8719_), .B(_14924__bF_buf0), .S(_8696_), .Y(_1__13_) );
INVX1 INVX1_3844 ( .gnd(gnd), .vdd(vdd), .A(data_0__14_), .Y(_8720_) );
OAI21X1 OAI21X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf14_bF_buf3), .C(_8720_), .Y(_8721_) );
OAI21X1 OAI21X1_2377 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_14_bF_buf3), .B(_8696_), .C(_8721_), .Y(_8722_) );
INVX1 INVX1_3845 ( .gnd(gnd), .vdd(vdd), .A(_8722_), .Y(_1__14_) );
INVX1 INVX1_3846 ( .gnd(gnd), .vdd(vdd), .A(data_0__15_), .Y(_8723_) );
OAI21X1 OAI21X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_15033_), .B(_14882__bF_buf13_bF_buf3), .C(_8723_), .Y(_8724_) );
OAI21X1 OAI21X1_2379 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_15_bF_buf5), .B(_8696_), .C(_8724_), .Y(_8725_) );
INVX1 INVX1_3847 ( .gnd(gnd), .vdd(vdd), .A(_8725_), .Y(_1__15_) );
NOR2X1 NOR2X1_859 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[1]), .B(IDATA_CORE_addr[0]), .Y(_8726_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(_8726_), .Y(_8727_) );
NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[2]), .B(IDATA_CORE_addr[3]), .Y(_8728_) );
NOR2X1 NOR2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_8728_), .B(_8727_), .Y(_8729_) );
INVX8 INVX8_33 ( .gnd(gnd), .vdd(vdd), .A(_8729_), .Y(_8730_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[4]), .Y(_8731_) );
NOR2X1 NOR2X1_861 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[5]), .B(_8731_), .Y(_8732_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[7]), .Y(_8733_) );
NOR2X1 NOR2X1_862 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[6]), .B(_8733_), .Y(_8734_) );
NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_8732_), .B(_8734_), .Y(_8735_) );
NOR2X1 NOR2X1_863 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8730_), .Y(_8736_) );
NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__0_), .Y(_8737_) );
INVX1 INVX1_3848 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[2]), .Y(_8738_) );
NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[3]), .B(_8738_), .Y(_8739_) );
NOR2X1 NOR2X1_864 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_8727_), .Y(_8740_) );
INVX8 INVX8_34 ( .gnd(gnd), .vdd(vdd), .A(_8740_), .Y(_8741_) );
NOR2X1 NOR2X1_865 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8741_), .Y(_8742_) );
NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__0_), .Y(_8743_) );
NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_8737_), .B(_8743_), .Y(_8744_) );
NOR2X1 NOR2X1_866 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[3]), .B(_8738_), .Y(_8745_) );
INVX1 INVX1_3849 ( .gnd(gnd), .vdd(vdd), .A(_8745_), .Y(_8746_) );
NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[1]), .B(IDATA_CORE_addr[0]), .Y(_8747_) );
NOR2X1 NOR2X1_867 ( .gnd(gnd), .vdd(vdd), .A(_8747_), .B(_8746_), .Y(_8748_) );
INVX8 INVX8_35 ( .gnd(gnd), .vdd(vdd), .A(_8748_), .Y(_8749_) );
NOR2X1 NOR2X1_868 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8749_), .Y(_8750_) );
NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__0_), .Y(_8751_) );
INVX1 INVX1_3850 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[0]), .Y(_8752_) );
NOR2X1 NOR2X1_869 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[1]), .B(_8752_), .Y(_8753_) );
INVX1 INVX1_3851 ( .gnd(gnd), .vdd(vdd), .A(_8753_), .Y(_8754_) );
NOR2X1 NOR2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_8754_), .Y(_8755_) );
INVX8 INVX8_36 ( .gnd(gnd), .vdd(vdd), .A(_8755_), .Y(_8756_) );
NOR2X1 NOR2X1_871 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8756_), .Y(_8757_) );
NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__0_), .Y(_8758_) );
NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_8751_), .B(_8758_), .Y(_8759_) );
NOR2X1 NOR2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_8744_), .B(_8759_), .Y(_8760_) );
NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_8726_), .B(_8745_), .Y(_8761_) );
NOR2X1 NOR2X1_873 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8735_), .Y(_8762_) );
NAND3X1 NAND3X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_3258_), .B(_8762_), .C(_3256_), .Y(_8763_) );
NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_8745_), .B(_8753_), .Y(_8764_) );
NOR2X1 NOR2X1_874 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8764_), .Y(_8765_) );
NAND3X1 NAND3X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_3217_), .B(_8765_), .C(_3214_), .Y(_8766_) );
AND2X2 AND2X2_1560 ( .gnd(gnd), .vdd(vdd), .A(_8766_), .B(_8763_), .Y(_8767_) );
NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[1]), .B(_8752_), .Y(_8768_) );
NOR2X1 NOR2X1_875 ( .gnd(gnd), .vdd(vdd), .A(_8768_), .B(_8746_), .Y(_8769_) );
INVX8 INVX8_37 ( .gnd(gnd), .vdd(vdd), .A(_8769_), .Y(_8770_) );
NOR2X1 NOR2X1_876 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8770_), .Y(_8771_) );
NOR2X1 NOR2X1_877 ( .gnd(gnd), .vdd(vdd), .A(_8747_), .B(_8739_), .Y(_8772_) );
INVX8 INVX8_38 ( .gnd(gnd), .vdd(vdd), .A(_8772_), .Y(_8773_) );
NOR2X1 NOR2X1_878 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8773_), .Y(_8774_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_62__0_), .B(_8774_), .C(_57__0_), .D(_8771_), .Y(_8775_) );
NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_8767_), .B(_8775_), .Y(_8776_) );
NOR2X1 NOR2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_8728_), .B(_8754_), .Y(_8777_) );
INVX8 INVX8_39 ( .gnd(gnd), .vdd(vdd), .A(_8777_), .Y(_8778_) );
NOR2X1 NOR2X1_880 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8778_), .Y(_8779_) );
NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__0_), .Y(_8780_) );
NOR2X1 NOR2X1_881 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[2]), .B(IDATA_CORE_addr[3]), .Y(_8781_) );
NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_8781_), .B(_8753_), .Y(_8782_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[5]), .Y(_8783_) );
NOR2X1 NOR2X1_882 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[4]), .B(_8783_), .Y(_8784_) );
NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .B(_8784_), .Y(_8785_) );
NOR2X1 NOR2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf3), .B(_8785_), .Y(_8786_) );
NAND3X1 NAND3X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_2792_), .B(_8786_), .C(_2794_), .Y(_8787_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(_8781_), .Y(_8788_) );
NOR2X1 NOR2X1_884 ( .gnd(gnd), .vdd(vdd), .A(_8747_), .B(_8788_), .Y(_8789_) );
INVX8 INVX8_40 ( .gnd(gnd), .vdd(vdd), .A(_8789_), .Y(_8790_) );
NOR2X1 NOR2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8790_), .Y(_8791_) );
INVX8 INVX8_41 ( .gnd(gnd), .vdd(vdd), .A(_8791_), .Y(_8792_) );
OAI21X1 OAI21X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .B(_8792_), .C(_8787_), .Y(_8793_) );
NOR2X1 NOR2X1_886 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8785_), .Y(_8794_) );
NAND3X1 NAND3X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_8794_), .C(_2624_), .Y(_8795_) );
NOR2X1 NOR2X1_887 ( .gnd(gnd), .vdd(vdd), .A(_8768_), .B(_8788_), .Y(_8796_) );
INVX8 INVX8_42 ( .gnd(gnd), .vdd(vdd), .A(_8796_), .Y(_8797_) );
NOR2X1 NOR2X1_888 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8797_), .Y(_8798_) );
INVX8 INVX8_43 ( .gnd(gnd), .vdd(vdd), .A(_8798_), .Y(_8799_) );
OAI21X1 OAI21X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .B(_8799_), .C(_8795_), .Y(_8800_) );
NOR2X1 NOR2X1_889 ( .gnd(gnd), .vdd(vdd), .A(_8800_), .B(_8793_), .Y(_8801_) );
NOR2X1 NOR2X1_890 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8749_), .Y(_8802_) );
NOR2X1 NOR2X1_891 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8770_), .Y(_8803_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_75__0_), .B(_8802_), .C(_74__0_), .D(_8803_), .Y(_8804_) );
NOR2X1 NOR2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8773_), .Y(_8805_) );
NOR2X1 NOR2X1_893 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8778_), .Y(_8806_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_82__0_), .B(_8806_), .C(_80__0_), .D(_8805_), .Y(_8807_) );
NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_8804_), .B(_8807_), .Y(_8808_) );
INVX1 INVX1_3852 ( .gnd(gnd), .vdd(vdd), .A(_84__0_), .Y(_8809_) );
INVX1 INVX1_3853 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .Y(_8810_) );
NOR2X1 NOR2X1_894 ( .gnd(gnd), .vdd(vdd), .A(_8728_), .B(_8747_), .Y(_8811_) );
NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8810_), .Y(_8812_) );
NOR2X1 NOR2X1_895 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_8809_), .Y(_8813_) );
NOR2X1 NOR2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_8727_), .B(_8788_), .Y(_8814_) );
NOR2X1 NOR2X1_897 ( .gnd(gnd), .vdd(vdd), .A(_8731_), .B(_8783_), .Y(_8815_) );
NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .B(_8815_), .Y(_8816_) );
INVX1 INVX1_3854 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .Y(_8817_) );
NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_8817_), .Y(_8818_) );
NOR2X1 NOR2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2282_), .Y(_8819_) );
OR2X2 OR2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_8739_), .B(_8768_), .Y(_8820_) );
NOR2X1 NOR2X1_899 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8820__bF_buf3), .Y(_8821_) );
NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__0_), .Y(_8822_) );
NOR2X1 NOR2X1_900 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8816_), .Y(_8823_) );
NAND3X1 NAND3X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_8823_), .C(_2034_), .Y(_8824_) );
NOR2X1 NOR2X1_901 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8756_), .Y(_8825_) );
NAND3X1 NAND3X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1891_), .C(_1893_), .Y(_8826_) );
NAND3X1 NAND3X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_8826_), .B(_8824_), .C(_8822_), .Y(_8827_) );
NOR3X1 NOR3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_8813_), .B(_8827_), .C(_8819_), .Y(_8828_) );
NOR2X1 NOR2X1_902 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf2), .B(_8816_), .Y(_8829_) );
NAND3X1 NAND3X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_8829_), .C(_2231_), .Y(_8830_) );
NOR2X1 NOR2X1_903 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8790_), .Y(_8831_) );
NAND3X1 NAND3X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(_8831_), .C(_2125_), .Y(_8832_) );
NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_8830_), .B(_8832_), .Y(_8833_) );
NOR2X1 NOR2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8816_), .Y(_8834_) );
NAND3X1 NAND3X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .B(_8834_), .C(_2066_), .Y(_8835_) );
NOR2X1 NOR2X1_905 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8797_), .Y(_8836_) );
NAND3X1 NAND3X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_2175_), .B(_8836_), .C(_2177_), .Y(_8837_) );
NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_8835_), .B(_8837_), .Y(_8838_) );
NOR2X1 NOR2X1_906 ( .gnd(gnd), .vdd(vdd), .A(_8838_), .B(_8833_), .Y(_8839_) );
NOR2X1 NOR2X1_907 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8749_), .Y(_8840_) );
NOR2X1 NOR2X1_908 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8741_), .Y(_8841_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_94__0_), .B(_8841_), .C(_93__0_), .D(_8840_), .Y(_8842_) );
NOR2X1 NOR2X1_909 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8770_), .Y(_8843_) );
NAND2X1 NAND2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_8843_), .B(_92__0_), .Y(_8844_) );
NOR2X1 NOR2X1_910 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8730_), .Y(_8845_) );
NAND2X1 NAND2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_98__0_), .Y(_8846_) );
NAND3X1 NAND3X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_8844_), .B(_8846_), .C(_8842_), .Y(_8847_) );
NOR2X1 NOR2X1_911 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8778_), .Y(_8848_) );
NAND2X1 NAND2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__0_), .Y(_8849_) );
NAND2X1 NAND2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_8731_), .B(_8783_), .Y(_8850_) );
INVX1 INVX1_3855 ( .gnd(gnd), .vdd(vdd), .A(_8850_), .Y(_8851_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[6]), .Y(_8852_) );
NOR2X1 NOR2X1_912 ( .gnd(gnd), .vdd(vdd), .A(_8852_), .B(_8733_), .Y(_8853_) );
NAND2X1 NAND2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_8853_), .B(_8851_), .Y(_8854_) );
NOR2X1 NOR2X1_913 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8790_), .Y(_8855_) );
NAND3X1 NAND3X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1569_), .C(_1571_), .Y(_8856_) );
NOR2X1 NOR2X1_914 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8741_), .Y(_8857_) );
NAND3X1 NAND3X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_8857_), .C(_1358_), .Y(_8858_) );
NAND2X1 NAND2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_8858_), .B(_8856_), .Y(_8859_) );
NOR2X1 NOR2X1_915 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf1), .B(_8854_), .Y(_8860_) );
NAND3X1 NAND3X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1650_), .C(_1652_), .Y(_8861_) );
NOR2X1 NOR2X1_916 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8730_), .Y(_8862_) );
NAND3X1 NAND3X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_1232_), .B(_8862_), .C(_1230_), .Y(_8863_) );
NAND2X1 NAND2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_8861_), .B(_8863_), .Y(_8864_) );
OR2X2 OR2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_8864_), .B(_8859_), .Y(_8865_) );
NOR2X1 NOR2X1_917 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8778_), .Y(_8866_) );
INVX4 INVX4_47 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .Y(_8867_) );
NOR3X1 NOR3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_8867_), .C(_1199_), .Y(_8868_) );
NAND2X1 NAND2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_8852_), .B(_8733_), .Y(_8869_) );
INVX1 INVX1_3856 ( .gnd(gnd), .vdd(vdd), .A(_8869_), .Y(_8870_) );
NAND2X1 NAND2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_8870_), .Y(_8871_) );
NOR2X1 NOR2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8756_), .Y(_8872_) );
NOR2X1 NOR2X1_919 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8741_), .Y(_8873_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_191__0_), .B(_8873_), .C(_192__0_), .D(_8872_), .Y(_8874_) );
NOR2X1 NOR2X1_920 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8730_), .Y(_8875_) );
NOR2X1 NOR2X1_921 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf2), .B(_8871_), .Y(_8876_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_195__0_), .B(_8875_), .C(_193__0_), .D(_8876_), .Y(_8877_) );
NAND2X1 NAND2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_8874_), .B(_8877_), .Y(_8878_) );
NOR2X1 NOR2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8770_), .Y(_8879_) );
NAND2X1 NAND2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_8732_), .B(_8853_), .Y(_8880_) );
NOR2X1 NOR2X1_923 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8880_), .Y(_8881_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_188__0_), .B(_8879_), .C(_126__0_), .D(_8881_), .Y(_8882_) );
NOR2X1 NOR2X1_924 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8778_), .Y(_8883_) );
NOR2X1 NOR2X1_925 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8773_), .Y(_8884_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_196__0_), .B(_8883_), .C(_194__0_), .D(_8884_), .Y(_8885_) );
NAND2X1 NAND2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_8882_), .B(_8885_), .Y(_8886_) );
NOR3X1 NOR3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_8886_), .B(_8868_), .C(_8878_), .Y(_8887_) );
INVX1 INVX1_3857 ( .gnd(gnd), .vdd(vdd), .A(_8732_), .Y(_8888_) );
NOR2X1 NOR2X1_926 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[7]), .B(_8852_), .Y(_8889_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(_8889_), .Y(_8890_) );
NOR2X1 NOR2X1_927 ( .gnd(gnd), .vdd(vdd), .A(_8888_), .B(_8890_), .Y(_8891_) );
INVX8 INVX8_44 ( .gnd(gnd), .vdd(vdd), .A(_8891_), .Y(_8892_) );
NOR2X1 NOR2X1_928 ( .gnd(gnd), .vdd(vdd), .A(_8790_), .B(_8892_), .Y(_8893_) );
NAND3X1 NAND3X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_5812_), .B(_8893_), .C(_5810_), .Y(_8894_) );
INVX1 INVX1_3858 ( .gnd(gnd), .vdd(vdd), .A(_8815_), .Y(_8895_) );
NOR2X1 NOR2X1_929 ( .gnd(gnd), .vdd(vdd), .A(_8890_), .B(_8895_), .Y(_8896_) );
INVX8 INVX8_45 ( .gnd(gnd), .vdd(vdd), .A(_8896_), .Y(_8897_) );
NOR2X1 NOR2X1_930 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8897_), .Y(_8898_) );
NAND3X1 NAND3X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_4572_), .B(_8898_), .C(_4570_), .Y(_8899_) );
NAND2X1 NAND2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_8894_), .B(_8899_), .Y(_8900_) );
NOR2X1 NOR2X1_931 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .B(_8892_), .Y(_8901_) );
NAND3X1 NAND3X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_5509_), .B(_8901_), .C(_5507_), .Y(_8902_) );
NAND2X1 NAND2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_8732_), .B(_8870_), .Y(_8903_) );
NOR2X1 NOR2X1_932 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf1), .B(_8903_), .Y(_8904_) );
NAND3X1 NAND3X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_7847_), .B(_8904_), .C(_7845_), .Y(_8905_) );
NAND2X1 NAND2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_8902_), .B(_8905_), .Y(_8906_) );
NOR2X1 NOR2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_8900_), .B(_8906_), .Y(_8907_) );
NAND2X1 NAND2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_8734_), .B(_8851_), .Y(_8908_) );
NOR2X1 NOR2X1_934 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8790_), .Y(_8909_) );
NAND3X1 NAND3X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_4072_), .B(_8909_), .C(_4070_), .Y(_8910_) );
NOR2X1 NOR2X1_935 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8741_), .Y(_8911_) );
NAND3X1 NAND3X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3874_), .C(_3871_), .Y(_8912_) );
NAND2X1 NAND2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_8910_), .B(_8912_), .Y(_8913_) );
NOR2X1 NOR2X1_936 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8897_), .Y(_8914_) );
NAND3X1 NAND3X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .B(_8914_), .C(_4611_), .Y(_8915_) );
NOR2X1 NOR2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_8869_), .B(_8895_), .Y(_8916_) );
INVX8 INVX8_46 ( .gnd(gnd), .vdd(vdd), .A(_8916_), .Y(_8917_) );
NOR2X1 NOR2X1_938 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf0), .B(_8917_), .Y(_8918_) );
NAND3X1 NAND3X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_6634_), .B(_8918_), .C(_6632_), .Y(_8919_) );
NAND2X1 NAND2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_8915_), .B(_8919_), .Y(_8920_) );
NOR2X1 NOR2X1_939 ( .gnd(gnd), .vdd(vdd), .A(_8913_), .B(_8920_), .Y(_8921_) );
NAND2X1 NAND2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_8907_), .B(_8921_), .Y(_8922_) );
INVX1 INVX1_3859 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .Y(_8923_) );
NOR2X1 NOR2X1_940 ( .gnd(gnd), .vdd(vdd), .A(_8923_), .B(_8890_), .Y(_8924_) );
INVX8 INVX8_47 ( .gnd(gnd), .vdd(vdd), .A(_8924_), .Y(_8925_) );
NOR2X1 NOR2X1_941 ( .gnd(gnd), .vdd(vdd), .A(_8773_), .B(_8925_), .Y(_8926_) );
NAND3X1 NAND3X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_4953_), .B(_8926_), .C(_4950_), .Y(_8927_) );
NOR2X1 NOR2X1_942 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8903_), .Y(_8928_) );
NAND3X1 NAND3X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_8055_), .B(_8928_), .C(_8054_), .Y(_8929_) );
NAND2X1 NAND2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_8927_), .B(_8929_), .Y(_8930_) );
NOR2X1 NOR2X1_943 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_8897_), .Y(_8931_) );
NAND3X1 NAND3X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_4475_), .B(_8931_), .C(_4473_), .Y(_8932_) );
NOR2X1 NOR2X1_944 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8903_), .Y(_8933_) );
NAND3X1 NAND3X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_8021_), .B(_8933_), .C(_8020_), .Y(_8934_) );
NAND2X1 NAND2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_8932_), .B(_8934_), .Y(_8935_) );
NOR2X1 NOR2X1_945 ( .gnd(gnd), .vdd(vdd), .A(_8930_), .B(_8935_), .Y(_8936_) );
NOR2X1 NOR2X1_946 ( .gnd(gnd), .vdd(vdd), .A(_8770_), .B(_8925_), .Y(_8937_) );
NAND3X1 NAND3X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_8937_), .C(_5165_), .Y(_8938_) );
NOR2X1 NOR2X1_947 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8773_), .Y(_8939_) );
NAND3X1 NAND3X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_7809_), .B(_8939_), .C(_7807_), .Y(_8940_) );
NAND2X1 NAND2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_8938_), .B(_8940_), .Y(_8941_) );
NOR2X1 NOR2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_8749_), .B(_8925_), .Y(_8942_) );
NAND3X1 NAND3X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_5129_), .B(_8942_), .C(_5127_), .Y(_8943_) );
NOR2X1 NOR2X1_949 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf3), .B(_8925_), .Y(_8944_) );
NAND3X1 NAND3X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_4991_), .B(_8944_), .C(_4989_), .Y(_8945_) );
NAND2X1 NAND2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_8943_), .B(_8945_), .Y(_8946_) );
NOR2X1 NOR2X1_950 ( .gnd(gnd), .vdd(vdd), .A(_8946_), .B(_8941_), .Y(_8947_) );
NAND2X1 NAND2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_8936_), .B(_8947_), .Y(_8948_) );
NOR2X1 NOR2X1_951 ( .gnd(gnd), .vdd(vdd), .A(_8922_), .B(_8948_), .Y(_8949_) );
NOR2X1 NOR2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_8917_), .Y(_8950_) );
NAND3X1 NAND3X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_6705_), .B(_8950_), .C(_6703_), .Y(_8951_) );
NOR2X1 NOR2X1_953 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8749_), .Y(_8952_) );
NAND3X1 NAND3X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_3915_), .B(_8952_), .C(_3913_), .Y(_8953_) );
NAND2X1 NAND2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_8951_), .B(_8953_), .Y(_8954_) );
NOR2X1 NOR2X1_954 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf0), .B(_8892_), .Y(_8955_) );
NAND3X1 NAND3X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_5884_), .B(_8955_), .C(_5882_), .Y(_8956_) );
NOR2X1 NOR2X1_955 ( .gnd(gnd), .vdd(vdd), .A(_8756_), .B(_8917_), .Y(_8957_) );
NAND3X1 NAND3X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_6673_), .B(_8957_), .C(_6672_), .Y(_8958_) );
NAND2X1 NAND2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_8956_), .B(_8958_), .Y(_8959_) );
NOR2X1 NOR2X1_956 ( .gnd(gnd), .vdd(vdd), .A(_8959_), .B(_8954_), .Y(_8960_) );
NOR2X1 NOR2X1_957 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8730_), .Y(_8961_) );
NAND3X1 NAND3X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_7775_), .B(_8961_), .C(_7773_), .Y(_8962_) );
NOR2X1 NOR2X1_958 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8756_), .Y(_8963_) );
NAND3X1 NAND3X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .B(_8963_), .C(_3832_), .Y(_8964_) );
NAND2X1 NAND2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_8962_), .B(_8964_), .Y(_8965_) );
NOR2X1 NOR2X1_959 ( .gnd(gnd), .vdd(vdd), .A(_8797_), .B(_8892_), .Y(_8966_) );
NAND3X1 NAND3X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_5850_), .B(_8966_), .C(_5848_), .Y(_8967_) );
NOR2X1 NOR2X1_960 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8773_), .Y(_8968_) );
NAND3X1 NAND3X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_3756_), .B(_8968_), .C(_3752_), .Y(_8969_) );
NAND2X1 NAND2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_8967_), .B(_8969_), .Y(_8970_) );
NOR2X1 NOR2X1_961 ( .gnd(gnd), .vdd(vdd), .A(_8965_), .B(_8970_), .Y(_8971_) );
NAND2X1 NAND2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_8960_), .B(_8971_), .Y(_8972_) );
NOR2X1 NOR2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8749_), .Y(_8973_) );
NAND3X1 NAND3X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_7957_), .B(_8973_), .C(_7955_), .Y(_8974_) );
NOR2X1 NOR2X1_963 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8797_), .Y(_8975_) );
NAND3X1 NAND3X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_3460_), .B(_8975_), .C(_3457_), .Y(_8976_) );
NAND2X1 NAND2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_8974_), .B(_8976_), .Y(_8977_) );
NOR2X1 NOR2X1_964 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8908_), .Y(_8978_) );
NAND3X1 NAND3X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_4035_), .B(_8978_), .C(_4033_), .Y(_8979_) );
NOR2X1 NOR2X1_965 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8797_), .Y(_8980_) );
NAND3X1 NAND3X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_4109_), .B(_8980_), .C(_4107_), .Y(_8981_) );
NAND2X1 NAND2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_8981_), .B(_8979_), .Y(_8982_) );
NOR2X1 NOR2X1_966 ( .gnd(gnd), .vdd(vdd), .A(_8977_), .B(_8982_), .Y(_8983_) );
NOR2X1 NOR2X1_967 ( .gnd(gnd), .vdd(vdd), .A(_8797_), .B(_8925_), .Y(_8984_) );
NAND3X1 NAND3X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_5299_), .B(_8984_), .C(_5295_), .Y(_8985_) );
NOR2X1 NOR2X1_968 ( .gnd(gnd), .vdd(vdd), .A(_8790_), .B(_8925_), .Y(_8986_) );
NAND3X1 NAND3X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_5264_), .B(_8986_), .C(_5262_), .Y(_8987_) );
NAND2X1 NAND2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_8985_), .B(_8987_), .Y(_8988_) );
NOR2X1 NOR2X1_969 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .B(_8917_), .Y(_8989_) );
NAND3X1 NAND3X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_6561_), .B(_8989_), .C(_6559_), .Y(_8990_) );
NOR2X1 NOR2X1_970 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf3), .B(_8908_), .Y(_8991_) );
NAND3X1 NAND3X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_4145_), .B(_8991_), .C(_4143_), .Y(_8992_) );
NAND2X1 NAND2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_8990_), .B(_8992_), .Y(_8993_) );
NOR2X1 NOR2X1_971 ( .gnd(gnd), .vdd(vdd), .A(_8988_), .B(_8993_), .Y(_8994_) );
NAND2X1 NAND2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_8983_), .B(_8994_), .Y(_8995_) );
NOR2X1 NOR2X1_972 ( .gnd(gnd), .vdd(vdd), .A(_8972_), .B(_8995_), .Y(_8996_) );
NAND2X1 NAND2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_8949_), .B(_8996_), .Y(_8997_) );
NOR2X1 NOR2X1_973 ( .gnd(gnd), .vdd(vdd), .A(_8778_), .B(_8925_), .Y(_8998_) );
NAND3X1 NAND3X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_4884_), .B(_8998_), .C(_4882_), .Y(_8999_) );
NOR2X1 NOR2X1_974 ( .gnd(gnd), .vdd(vdd), .A(_8728_), .B(_8768_), .Y(_9000_) );
INVX8 INVX8_48 ( .gnd(gnd), .vdd(vdd), .A(_9000_), .Y(_9001_) );
NOR2X1 NOR2X1_975 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_8917_), .Y(_9002_) );
NAND3X1 NAND3X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_6491_), .B(_9002_), .C(_6490_), .Y(_9003_) );
NAND2X1 NAND2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_8999_), .B(_9003_), .Y(_9004_) );
NOR2X1 NOR2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_8770_), .B(_8892_), .Y(_9005_) );
NAND3X1 NAND3X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_5697_), .B(_9005_), .C(_5696_), .Y(_9006_) );
NOR2X1 NOR2X1_977 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_8925_), .Y(_9007_) );
NAND3X1 NAND3X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_4845_), .B(_9007_), .C(_4843_), .Y(_9008_) );
NAND2X1 NAND2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_9006_), .B(_9008_), .Y(_9009_) );
NOR2X1 NOR2X1_978 ( .gnd(gnd), .vdd(vdd), .A(_9004_), .B(_9009_), .Y(_9010_) );
NOR2X1 NOR2X1_979 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8892_), .Y(_9011_) );
NAND3X1 NAND3X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_5735_), .B(_9011_), .C(_5734_), .Y(_9012_) );
NOR2X1 NOR2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_8770_), .B(_8917_), .Y(_9013_) );
NAND3X1 NAND3X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_6777_), .B(_9013_), .C(_6776_), .Y(_9014_) );
NAND2X1 NAND2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_9012_), .B(_9014_), .Y(_9015_) );
NOR2X1 NOR2X1_981 ( .gnd(gnd), .vdd(vdd), .A(_8749_), .B(_8917_), .Y(_9016_) );
NAND3X1 NAND3X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_6738_), .B(_9016_), .C(_6737_), .Y(_9017_) );
NOR2X1 NOR2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_8790_), .B(_8917_), .Y(_9018_) );
NAND3X1 NAND3X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_6879_), .B(_9018_), .C(_6878_), .Y(_9019_) );
NAND2X1 NAND2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_9017_), .B(_9019_), .Y(_9020_) );
NOR2X1 NOR2X1_983 ( .gnd(gnd), .vdd(vdd), .A(_9020_), .B(_9015_), .Y(_9021_) );
NAND2X1 NAND2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_9010_), .B(_9021_), .Y(_9022_) );
NAND2X1 NAND2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_8889_), .B(_8851_), .Y(_9023_) );
NOR2X1 NOR2X1_984 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_9023_), .Y(_9024_) );
NAND3X1 NAND3X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_6261_), .B(_9024_), .C(_6259_), .Y(_9025_) );
NOR2X1 NOR2X1_985 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8790_), .Y(_9026_) );
NAND3X1 NAND3X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_6333_), .B(_9026_), .C(_6332_), .Y(_9027_) );
NAND2X1 NAND2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_9025_), .B(_9027_), .Y(_9028_) );
NOR2X1 NOR2X1_986 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8730_), .Y(_9029_) );
NAND3X1 NAND3X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_6038_), .B(_9029_), .C(_6037_), .Y(_9030_) );
NOR2X1 NOR2X1_987 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf2), .B(_9023_), .Y(_9031_) );
NAND3X1 NAND3X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_6096_), .B(_9031_), .C(_6095_), .Y(_9032_) );
NAND2X1 NAND2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_9030_), .B(_9032_), .Y(_9033_) );
NOR2X1 NOR2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_9028_), .B(_9033_), .Y(_9034_) );
NOR2X1 NOR2X1_989 ( .gnd(gnd), .vdd(vdd), .A(_8749_), .B(_8892_), .Y(_9035_) );
NAND3X1 NAND3X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_5656_), .B(_9035_), .C(_5654_), .Y(_9036_) );
NOR2X1 NOR2X1_990 ( .gnd(gnd), .vdd(vdd), .A(_8790_), .B(_8897_), .Y(_9037_) );
NAND3X1 NAND3X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_4652_), .B(_9037_), .C(_4650_), .Y(_9038_) );
NAND2X1 NAND2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_9038_), .B(_9036_), .Y(_9039_) );
NOR2X1 NOR2X1_991 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_9023_), .Y(_9040_) );
NAND3X1 NAND3X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_6297_), .B(_9040_), .C(_6295_), .Y(_9041_) );
NOR2X1 NOR2X1_992 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .B(_8897_), .Y(_9042_) );
NAND3X1 NAND3X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_4314_), .B(_9042_), .C(_4312_), .Y(_9043_) );
NAND2X1 NAND2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_9041_), .B(_9043_), .Y(_9044_) );
NOR2X1 NOR2X1_993 ( .gnd(gnd), .vdd(vdd), .A(_9044_), .B(_9039_), .Y(_9045_) );
NAND2X1 NAND2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_9034_), .B(_9045_), .Y(_9046_) );
NOR2X1 NOR2X1_994 ( .gnd(gnd), .vdd(vdd), .A(_9022_), .B(_9046_), .Y(_9047_) );
NOR2X1 NOR2X1_995 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8749_), .Y(_9048_) );
NAND3X1 NAND3X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_6185_), .B(_9048_), .C(_6184_), .Y(_9049_) );
NOR2X1 NOR2X1_996 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8741_), .Y(_9050_) );
NAND3X1 NAND3X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_7920_), .B(_9050_), .C(_7919_), .Y(_9051_) );
NAND2X1 NAND2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_9049_), .B(_9051_), .Y(_9052_) );
NOR2X1 NOR2X1_997 ( .gnd(gnd), .vdd(vdd), .A(_8778_), .B(_8892_), .Y(_9053_) );
NAND3X1 NAND3X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_5469_), .B(_9053_), .C(_5467_), .Y(_9054_) );
NOR2X1 NOR2X1_998 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8756_), .Y(_9055_) );
NAND3X1 NAND3X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_7883_), .B(_9055_), .C(_7881_), .Y(_9056_) );
NAND2X1 NAND2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_9054_), .B(_9056_), .Y(_9057_) );
NOR2X1 NOR2X1_999 ( .gnd(gnd), .vdd(vdd), .A(_9052_), .B(_9057_), .Y(_9058_) );
NOR2X1 NOR2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_8756_), .B(_8897_), .Y(_9059_) );
NAND3X1 NAND3X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .B(_9059_), .C(_4433_), .Y(_9060_) );
NOR2X1 NOR2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf1), .B(_8897_), .Y(_9061_) );
NAND3X1 NAND3X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_4395_), .B(_9061_), .C(_4394_), .Y(_9062_) );
NAND2X1 NAND2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_9060_), .B(_9062_), .Y(_9063_) );
NOR2X1 NOR2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8770_), .Y(_9064_) );
NAND3X1 NAND3X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_6223_), .B(_9064_), .C(_6222_), .Y(_9065_) );
NOR2X1 NOR2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_8773_), .B(_8897_), .Y(_9066_) );
NAND3X1 NAND3X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_4355_), .B(_9066_), .C(_4353_), .Y(_9067_) );
NAND2X1 NAND2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_9065_), .B(_9067_), .Y(_9068_) );
NOR2X1 NOR2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_9068_), .B(_9063_), .Y(_9069_) );
NAND2X1 NAND2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_9058_), .B(_9069_), .Y(_9070_) );
NOR2X1 NOR2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf2), .B(_8871_), .Y(_9071_) );
NAND3X1 NAND3X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_7579_), .B(_9071_), .C(_7577_), .Y(_9072_) );
NOR2X1 NOR2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8797_), .Y(_9073_) );
NAND3X1 NAND3X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_7543_), .B(_9073_), .C(_7541_), .Y(_9074_) );
NAND2X1 NAND2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_9072_), .B(_9074_), .Y(_9075_) );
NOR2X1 NOR2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8892_), .Y(_9076_) );
NAND3X1 NAND3X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_5773_), .B(_9076_), .C(_5771_), .Y(_9077_) );
NOR2X1 NOR2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf1), .B(_8735_), .Y(_9078_) );
NAND3X1 NAND3X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_3499_), .B(_9078_), .C(_3496_), .Y(_9079_) );
NAND2X1 NAND2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_9077_), .B(_9079_), .Y(_9080_) );
NOR2X1 NOR2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_9075_), .B(_9080_), .Y(_9081_) );
NOR2X1 NOR2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_8892_), .Y(_9082_) );
NAND3X1 NAND3X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_5428_), .B(_9082_), .C(_5427_), .Y(_9083_) );
NOR2X1 NOR2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf0), .B(_8908_), .Y(_9084_) );
NAND3X1 NAND3X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_9084_), .C(_3791_), .Y(_9085_) );
NAND2X1 NAND2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_9085_), .B(_9083_), .Y(_9086_) );
NOR2X1 NOR2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_8773_), .B(_8917_), .Y(_9087_) );
NAND3X1 NAND3X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_6594_), .B(_9087_), .C(_6593_), .Y(_9088_) );
NOR2X1 NOR2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_9001_), .Y(_9089_) );
NAND3X1 NAND3X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_3648_), .B(_9089_), .C(_3643_), .Y(_9090_) );
NAND2X1 NAND2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_9088_), .B(_9090_), .Y(_9091_) );
NOR2X1 NOR2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_9086_), .B(_9091_), .Y(_9092_) );
NAND2X1 NAND2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_9081_), .B(_9092_), .Y(_9093_) );
NOR2X1 NOR2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_9070_), .B(_9093_), .Y(_9094_) );
NAND2X1 NAND2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_9047_), .B(_9094_), .Y(_9095_) );
NOR2X1 NOR2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_8997_), .B(_9095_), .Y(_9096_) );
NOR2X1 NOR2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_8730_), .B(_8925_), .Y(_9097_) );
NAND2X1 NAND2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__0_), .Y(_9098_) );
NOR2X1 NOR2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8770_), .Y(_9099_) );
NAND3X1 NAND3X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(_9099_), .C(_3953_), .Y(_9100_) );
NAND2X1 NAND2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_9098_), .B(_9100_), .Y(_9101_) );
NOR2X1 NOR2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_8925_), .Y(_9102_) );
NAND3X1 NAND3X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_9102_), .C(_5077_), .Y(_9103_) );
NOR2X1 NOR2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8917_), .Y(_9104_) );
NAND3X1 NAND3X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_6844_), .B(_9104_), .C(_6843_), .Y(_9105_) );
NAND2X1 NAND2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_9105_), .B(_9103_), .Y(_9106_) );
NOR2X1 NOR2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_9101_), .B(_9106_), .Y(_9107_) );
NAND2X1 NAND2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_8784_), .B(_8853_), .Y(_9108_) );
NOR2X1 NOR2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8730_), .Y(_9109_) );
NAND3X1 NAND3X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_15901_), .B(_9109_), .C(_15903_), .Y(_9110_) );
NOR2X1 NOR2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_8850_), .B(_8869_), .Y(_9111_) );
INVX8 INVX8_49 ( .gnd(gnd), .vdd(vdd), .A(_9111_), .Y(_9112_) );
NOR2X1 NOR2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8756_), .Y(_9113_) );
NAND3X1 NAND3X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_8365_), .B(_9113_), .C(_8367_), .Y(_9114_) );
NOR2X1 NOR2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8741_), .Y(_9115_) );
NAND3X1 NAND3X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_16113_), .B(_9115_), .C(_16112_), .Y(_9116_) );
NAND3X1 NAND3X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_9110_), .B(_9114_), .C(_9116_), .Y(_9117_) );
NOR2X1 NOR2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8790_), .Y(_9118_) );
NAND3X1 NAND3X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_370_), .C(_374_), .Y(_9119_) );
NOR2X1 NOR2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8778_), .Y(_9120_) );
NAND3X1 NAND3X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_15839_), .B(_9120_), .C(_15845_), .Y(_9121_) );
AND2X2 AND2X2_1561 ( .gnd(gnd), .vdd(vdd), .A(_9121_), .B(_9119_), .Y(_9122_) );
NOR2X1 NOR2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf0), .B(_8903_), .Y(_9123_) );
NOR2X1 NOR2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_9112_), .Y(_9124_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_201__0_), .B(_9124_), .C(_89__0_), .D(_9123_), .Y(_9125_) );
NAND2X1 NAND2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_9122_), .B(_9125_), .Y(_9126_) );
NOR2X1 NOR2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf3), .B(_8897_), .Y(_9127_) );
NAND3X1 NAND3X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_4728_), .B(_9127_), .C(_4730_), .Y(_9128_) );
NOR2X1 NOR2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8908_), .Y(_9129_) );
NAND3X1 NAND3X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_3988_), .B(_9129_), .C(_3991_), .Y(_9130_) );
NAND2X1 NAND2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_9130_), .B(_9128_), .Y(_9131_) );
NOR3X1 NOR3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_9117_), .B(_9131_), .C(_9126_), .Y(_9132_) );
NOR2X1 NOR2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8790_), .Y(_9133_) );
NAND3X1 NAND3X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3389_), .C(_3402_), .Y(_9134_) );
NOR2X1 NOR2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_8756_), .B(_8925_), .Y(_9135_) );
NAND3X1 NAND3X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_5026_), .B(_9135_), .C(_5028_), .Y(_9136_) );
NOR2X1 NOR2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_8797_), .B(_8917_), .Y(_9137_) );
NAND3X1 NAND3X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_6911_), .B(_9137_), .C(_6913_), .Y(_9138_) );
NAND3X1 NAND3X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_9136_), .B(_9138_), .C(_9134_), .Y(_9139_) );
NOR2X1 NOR2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_8797_), .B(_8897_), .Y(_9140_) );
NOR2X1 NOR2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8925_), .Y(_9141_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_17__0_), .B(_9140_), .C(_2__0_), .D(_9141_), .Y(_9142_) );
NOR2X1 NOR2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8917_), .Y(_9143_) );
NAND2X1 NAND2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__0_), .Y(_9144_) );
NOR2X1 NOR2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf2), .B(_8917_), .Y(_9145_) );
NAND2X1 NAND2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_200__0_), .Y(_9146_) );
NAND3X1 NAND3X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_9144_), .B(_9146_), .C(_9142_), .Y(_9147_) );
NOR2X1 NOR2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_9139_), .B(_9147_), .Y(_9148_) );
NAND3X1 NAND3X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_9107_), .B(_9148_), .C(_9132_), .Y(_9149_) );
NOR2X1 NOR2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_8770_), .B(_8897_), .Y(_9150_) );
NOR2X1 NOR2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8790_), .Y(_9151_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_21__0_), .B(_9150_), .C(_185__0_), .D(_9151_), .Y(_9152_) );
NOR2X1 NOR2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_8741_), .B(_8892_), .Y(_9153_) );
NOR2X1 NOR2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf1), .B(_8925_), .Y(_9154_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_243__0_), .B(_9153_), .C(_253__0_), .D(_9154_), .Y(_9155_) );
NAND2X1 NAND2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_9152_), .B(_9155_), .Y(_9156_) );
NOR2X1 NOR2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8778_), .Y(_9157_) );
NOR2X1 NOR2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8730_), .Y(_9158_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .B(_9158_), .C(_231__0_), .D(_9157_), .Y(_9159_) );
NOR2X1 NOR2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_8756_), .B(_8892_), .Y(_9160_) );
NOR2X1 NOR2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .B(_8778_), .Y(_9161_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_47__0_), .B(_9161_), .C(_244__0_), .D(_9160_), .Y(_9162_) );
NAND2X1 NAND2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_9162_), .B(_9159_), .Y(_9163_) );
NOR2X1 NOR2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_9156_), .B(_9163_), .Y(_9164_) );
NOR2X1 NOR2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_8773_), .B(_8892_), .Y(_9165_) );
NAND2X1 NAND2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_247__0_), .Y(_9166_) );
NOR2X1 NOR2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_8897_), .Y(_9167_) );
NAND2X1 NAND2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_9167_), .B(_30__0_), .Y(_9168_) );
NOR2X1 NOR2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf0), .B(_9023_), .Y(_9169_) );
NOR2X1 NOR2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8756_), .Y(_9170_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_218__0_), .B(_9169_), .C(_227__0_), .D(_9170_), .Y(_9171_) );
NAND3X1 NAND3X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_9166_), .B(_9168_), .C(_9171_), .Y(_9172_) );
NOR2X1 NOR2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8778_), .Y(_9173_) );
NOR2X1 NOR2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_8778_), .B(_8917_), .Y(_9174_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_178__0_), .B(_9173_), .C(_214__0_), .D(_9174_), .Y(_9175_) );
NOR2X1 NOR2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_8778_), .B(_8897_), .Y(_9176_) );
NOR2X1 NOR2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8770_), .Y(_9177_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_145__0_), .B(_9177_), .C(_29__0_), .D(_9176_), .Y(_9178_) );
NAND2X1 NAND2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_9175_), .B(_9178_), .Y(_9179_) );
NOR2X1 NOR2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_9179_), .B(_9172_), .Y(_9180_) );
NAND2X1 NAND2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_9164_), .B(_9180_), .Y(_9181_) );
NOR2X1 NOR2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8749_), .Y(_9182_) );
NOR2X1 NOR2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8730_), .Y(_9183_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_234__0_), .B(_9182_), .C(_34__0_), .D(_9183_), .Y(_9184_) );
NOR2X1 NOR2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8778_), .Y(_9185_) );
NAND2X1 NAND2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__0_), .Y(_9186_) );
NAND2X1 NAND2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_8772_), .B(_9111_), .Y(_9187_) );
INVX8 INVX8_50 ( .gnd(gnd), .vdd(vdd), .A(_9187_), .Y(_9188_) );
NAND2X1 NAND2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__0_), .Y(_9189_) );
NAND3X1 NAND3X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_9186_), .B(_9189_), .C(_9184_), .Y(_9190_) );
NAND2X1 NAND2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_8815_), .B(_8853_), .Y(_9191_) );
NOR2X1 NOR2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8797_), .Y(_9192_) );
NAND3X1 NAND3X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_15633_), .B(_9192_), .C(_15635_), .Y(_9193_) );
NOR2X1 NOR2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8790_), .Y(_9194_) );
INVX4 INVX4_48 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .Y(_9195_) );
OAI21X1 OAI21X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_15587_), .B(_9195_), .C(_9193_), .Y(_9196_) );
NOR2X1 NOR2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8749_), .Y(_9197_) );
NAND2X1 NAND2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__0_), .Y(_9198_) );
NOR2X1 NOR2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf3), .B(_9191_), .Y(_9199_) );
NAND3X1 NAND3X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_15689_), .B(_9199_), .C(_15691_), .Y(_9200_) );
NAND2X1 NAND2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_9198_), .B(_9200_), .Y(_9201_) );
NOR2X1 NOR2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_9201_), .B(_9196_), .Y(_9202_) );
NOR2X1 NOR2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8741_), .Y(_9203_) );
NAND2X1 NAND2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__0_), .Y(_9204_) );
NOR2X1 NOR2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8756_), .Y(_9205_) );
INVX4 INVX4_49 ( .gnd(gnd), .vdd(vdd), .A(_9205_), .Y(_9206_) );
OAI21X1 OAI21X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_15290_), .B(_9206_), .C(_9204_), .Y(_9207_) );
NOR2X1 NOR2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8730_), .Y(_9208_) );
NAND2X1 NAND2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__0_), .Y(_9209_) );
INVX1 INVX1_3860 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .Y(_9210_) );
NAND2X1 NAND2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_9210_), .B(_8777_), .Y(_9211_) );
OAI21X1 OAI21X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_15088_), .B(_9211_), .C(_9209_), .Y(_9212_) );
NOR2X1 NOR2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_9207_), .B(_9212_), .Y(_9213_) );
NOR2X1 NOR2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8773_), .Y(_9214_) );
INVX8 INVX8_51 ( .gnd(gnd), .vdd(vdd), .A(_9214_), .Y(_9215_) );
NOR3X1 NOR3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_15956_), .B(_9215_), .C(_15959_), .Y(_9216_) );
NOR2X1 NOR2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8820__bF_buf3), .Y(_9217_) );
NAND3X1 NAND3X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_15236_), .B(_9217_), .C(_15238_), .Y(_9218_) );
NOR2X1 NOR2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8773_), .Y(_9219_) );
NAND3X1 NAND3X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_15185_), .B(_9219_), .C(_15169_), .Y(_9220_) );
NAND2X1 NAND2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_9220_), .B(_9218_), .Y(_9221_) );
NOR2X1 NOR2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_9191_), .Y(_9222_) );
NAND3X1 NAND3X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_15458_), .B(_9222_), .C(_15460_), .Y(_9223_) );
NOR2X1 NOR2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_8770_), .Y(_9224_) );
NAND3X1 NAND3X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_15406_), .B(_9224_), .C(_15404_), .Y(_9225_) );
NAND2X1 NAND2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_9223_), .B(_9225_), .Y(_9226_) );
NOR3X1 NOR3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_9216_), .B(_9226_), .C(_9221_), .Y(_9227_) );
NAND3X1 NAND3X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_9213_), .B(_9227_), .C(_9202_), .Y(_9228_) );
NOR2X1 NOR2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8770_), .Y(_9229_) );
NAND2X1 NAND2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__0_), .Y(_9230_) );
INVX4 INVX4_50 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .Y(_9231_) );
NOR2X1 NOR2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_9231_), .Y(_9232_) );
NOR2X1 NOR2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_9191_), .Y(_9233_) );
NAND3X1 NAND3X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_15516_), .B(_9233_), .C(_15518_), .Y(_9234_) );
NOR2X1 NOR2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8871_), .Y(_9235_) );
INVX1 INVX1_3861 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[3]), .Y(_9236_) );
OAI21X1 OAI21X1_2385 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[1]), .B(IDATA_CORE_addr[2]), .C(_9236_), .Y(_9237_) );
NAND3X1 NAND3X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf2), .B(_9237_), .C(_9187_), .Y(_9238_) );
INVX1 INVX1_3862 ( .gnd(gnd), .vdd(vdd), .A(IDATA_CORE_addr[1]), .Y(_9239_) );
OAI21X1 OAI21X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_9239_), .B(IDATA_CORE_addr[2]), .C(IDATA_CORE_addr[3]), .Y(_9240_) );
NAND3X1 NAND3X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_9111_), .B(_9240_), .C(_8820__bF_buf2), .Y(_9241_) );
NOR2X1 NOR2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_9241_), .B(_9238_), .Y(_9242_) );
NAND2X1 NAND2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_1__0_), .B(_9242_), .Y(_9243_) );
NOR2X1 NOR2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_9001_), .Y(_9244_) );
INVX4 INVX4_51 ( .gnd(gnd), .vdd(vdd), .A(_9244_), .Y(_9245_) );
OAI21X1 OAI21X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_7073_), .B(_9245_), .C(_9243_), .Y(_9246_) );
AOI21X1 AOI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_187__0_), .B(_9235_), .C(_9246_), .Y(_9247_) );
NOR2X1 NOR2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_9001_), .Y(_9248_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(_9248_), .Y(_9249_) );
NOR2X1 NOR2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_9001_), .B(_9112_), .Y(_9250_) );
NAND2X1 NAND2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_9250_), .B(_56__0_), .Y(_9251_) );
OAI21X1 OAI21X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_7696_), .B(_9249_), .C(_9251_), .Y(_9252_) );
INVX1 INVX1_3863 ( .gnd(gnd), .vdd(vdd), .A(_8908_), .Y(_9253_) );
NAND2X1 NAND2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_9253_), .Y(_9254_) );
NOR2X1 NOR2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_9001_), .Y(_9255_) );
NAND3X1 NAND3X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_1748_), .B(_9255_), .C(_1750_), .Y(_9256_) );
OAI21X1 OAI21X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_9254_), .C(_9256_), .Y(_9257_) );
NOR2X1 NOR2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_9257_), .B(_9252_), .Y(_9258_) );
NAND2X1 NAND2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8916_), .Y(_9259_) );
INVX4 INVX4_52 ( .gnd(gnd), .vdd(vdd), .A(_9259_), .Y(_9260_) );
NAND2X1 NAND2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__0_), .Y(_9261_) );
NOR2X1 NOR2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_9001_), .Y(_9262_) );
INVX4 INVX4_53 ( .gnd(gnd), .vdd(vdd), .A(_9262_), .Y(_9263_) );
OAI21X1 OAI21X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_9263_), .C(_9261_), .Y(_9264_) );
INVX4 INVX4_54 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .Y(_9265_) );
NOR2X1 NOR2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_8871_), .Y(_9266_) );
INVX4 INVX4_55 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .Y(_9267_) );
NOR2X1 NOR2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_9001_), .Y(_9268_) );
NAND3X1 NAND3X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_9268_), .C(_1153_), .Y(_9269_) );
OAI21X1 OAI21X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_7027_), .B(_9267_), .C(_9269_), .Y(_9270_) );
NOR2X1 NOR2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_9264_), .B(_9270_), .Y(_9271_) );
NAND3X1 NAND3X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_9247_), .B(_9271_), .C(_9258_), .Y(_9272_) );
NAND2X1 NAND2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8924_), .Y(_9273_) );
INVX4 INVX4_56 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .Y(_9274_) );
NOR2X1 NOR2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_9191_), .Y(_9275_) );
INVX4 INVX4_57 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .Y(_9276_) );
NOR2X1 NOR2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_9001_), .Y(_9277_) );
NAND3X1 NAND3X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_9277_), .C(_2889_), .Y(_9278_) );
OAI21X1 OAI21X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_14893_), .B(_9276_), .C(_9278_), .Y(_9279_) );
AOI21X1 AOI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_14__0_), .B(_9274_), .C(_9279_), .Y(_9280_) );
NOR2X1 NOR2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_9231_), .Y(_9281_) );
NAND2X1 NAND2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8896_), .Y(_9282_) );
INVX4 INVX4_58 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .Y(_9283_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_31__0_), .B(_9283_), .C(_217__0_), .D(_9281_), .Y(_9284_) );
AND2X2 AND2X2_1562 ( .gnd(gnd), .vdd(vdd), .A(_9280_), .B(_9284_), .Y(_9285_) );
NOR2X1 NOR2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_9112_), .Y(_9286_) );
NAND2X1 NAND2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__0_), .Y(_9287_) );
NAND2X1 NAND2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_8916_), .Y(_9288_) );
INVX4 INVX4_59 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .Y(_9289_) );
NAND2X1 NAND2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__0_), .Y(_9290_) );
NAND2X1 NAND2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_9287_), .B(_9290_), .Y(_9291_) );
NOR2X1 NOR2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_9001_), .Y(_9292_) );
NAND3X1 NAND3X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_15789_), .B(_9292_), .C(_15791_), .Y(_9293_) );
NOR2X1 NOR2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_8908_), .Y(_9294_) );
INVX4 INVX4_60 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .Y(_9295_) );
OAI21X1 OAI21X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_3582_), .B(_9295_), .C(_9293_), .Y(_9296_) );
NOR2X1 NOR2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_9291_), .B(_9296_), .Y(_9297_) );
NOR2X1 NOR2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8871_), .Y(_9298_) );
NAND2X1 NAND2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .B(_186__0_), .Y(_9299_) );
NOR2X1 NOR2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_9231_), .Y(_9300_) );
INVX8 INVX8_52 ( .gnd(gnd), .vdd(vdd), .A(_9300_), .Y(_9301_) );
OAI21X1 OAI21X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_7614_), .B(_9301_), .C(_9299_), .Y(_9302_) );
NOR2X1 NOR2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_9231_), .Y(_9303_) );
INVX8 INVX8_53 ( .gnd(gnd), .vdd(vdd), .A(_9303_), .Y(_9304_) );
INVX1 INVX1_3864 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .Y(_9305_) );
NAND2X1 NAND2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_9305_), .Y(_9306_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_8148_), .B(_9304_), .C(_3534_), .D(_9306_), .Y(_9307_) );
NOR2X1 NOR2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_9307_), .B(_9302_), .Y(_9308_) );
NAND3X1 NAND3X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_9297_), .B(_9308_), .C(_9285_), .Y(_9309_) );
NOR2X1 NOR2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_9023_), .Y(_9310_) );
NAND3X1 NAND3X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_5943_), .B(_9310_), .C(_5945_), .Y(_9311_) );
NAND2X1 NAND2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_8896_), .Y(_9312_) );
INVX8 INVX8_54 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .Y(_9313_) );
NAND3X1 NAND3X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_4761_), .B(_9313_), .C(_4764_), .Y(_9314_) );
NOR2X1 NOR2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_9001_), .Y(_9315_) );
NAND3X1 NAND3X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_2338_), .B(_9315_), .C(_2340_), .Y(_9316_) );
NAND3X1 NAND3X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_9314_), .B(_9316_), .C(_9311_), .Y(_9317_) );
INVX1 INVX1_3865 ( .gnd(gnd), .vdd(vdd), .A(_9317_), .Y(_9318_) );
NAND2X1 NAND2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_8811_), .B(_8891_), .Y(_9319_) );
INVX8 INVX8_55 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .Y(_9320_) );
NOR2X1 NOR2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_8903_), .Y(_9321_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_251__0_), .B(_9320_), .C(_181__0_), .D(_9321_), .Y(_9322_) );
NAND2X1 NAND2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_8891_), .Y(_9323_) );
INVX8 INVX8_56 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .Y(_9324_) );
NAND2X1 NAND2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_8814_), .B(_8924_), .Y(_9325_) );
INVX8 INVX8_57 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .Y(_9326_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_252__0_), .B(_9326_), .C(_235__0_), .D(_9324_), .Y(_9327_) );
NAND3X1 NAND3X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_9327_), .B(_9322_), .C(_9318_), .Y(_9328_) );
NOR3X1 NOR3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_9272_), .B(_9328_), .C(_9309_), .Y(_9329_) );
NAND2X1 NAND2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_9234_), .B(_9329_), .Y(_9330_) );
AOI21X1 AOI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_157__0_), .B(_9232_), .C(_9330_), .Y(_9331_) );
NOR2X1 NOR2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_9191_), .B(_9001_), .Y(_9332_) );
NOR2X1 NOR2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_9265_), .Y(_9333_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_155__0_), .B(_9333_), .C(_172__0_), .D(_9332_), .Y(_9334_) );
NAND3X1 NAND3X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_9334_), .B(_9230_), .C(_9331_), .Y(_9335_) );
NOR3X1 NOR3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_9335_), .B(_9190_), .C(_9228_), .Y(_9336_) );
NOR2X1 NOR2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_9108_), .Y(_9337_) );
NAND2X1 NAND2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__0_), .Y(_9338_) );
NOR2X1 NOR2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8797_), .Y(_9339_) );
NAND3X1 NAND3X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_9339_), .C(_428_), .Y(_9340_) );
NOR2X1 NOR2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf1), .B(_9112_), .Y(_9341_) );
NOR2X1 NOR2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8790_), .Y(_9342_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_111__0_), .B(_9342_), .C(_12__0_), .D(_9341_), .Y(_9343_) );
NAND3X1 NAND3X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_9343_), .B(_9338_), .C(_9340_), .Y(_9344_) );
NOR2X1 NOR2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_9112_), .Y(_9345_) );
NOR2X1 NOR2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_8903_), .B(_8797_), .Y(_9346_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_100__0_), .B(_9346_), .C(_212__0_), .D(_9345_), .Y(_9347_) );
NOR2X1 NOR2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8741_), .Y(_9348_) );
NOR2X1 NOR2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf1), .B(_9108_), .Y(_9349_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_245__0_), .B(_9348_), .C(_140__0_), .D(_9349_), .Y(_9350_) );
NAND2X1 NAND2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_9350_), .B(_9347_), .Y(_9351_) );
NOR2X1 NOR2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_9344_), .B(_9351_), .Y(_9352_) );
NOR2X1 NOR2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8797_), .Y(_9353_) );
NOR2X1 NOR2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_9001_), .Y(_9354_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_232__0_), .B(_9354_), .C(_219__0_), .D(_9353_), .Y(_9355_) );
NOR2X1 NOR2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf0), .B(_8892_), .Y(_9356_) );
NOR2X1 NOR2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8741_), .Y(_9357_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_246__0_), .B(_9356_), .C(_226__0_), .D(_9357_), .Y(_9358_) );
NAND2X1 NAND2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_9358_), .B(_9355_), .Y(_9359_) );
NOR2X1 NOR2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8770_), .Y(_9360_) );
INVX8 INVX8_58 ( .gnd(gnd), .vdd(vdd), .A(_9360_), .Y(_9361_) );
NOR2X1 NOR2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8749_), .Y(_9362_) );
NAND3X1 NAND3X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16164_), .C(_16166_), .Y(_9363_) );
OAI21X1 OAI21X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_16215_), .B(_9361_), .C(_9363_), .Y(_9364_) );
NOR2X1 NOR2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8756_), .Y(_9365_) );
NAND3X1 NAND3X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16060_), .C(_16063_), .Y(_9366_) );
NOR2X1 NOR2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_8820__bF_buf3), .Y(_9367_) );
NAND3X1 NAND3X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16006_), .C(_16008_), .Y(_9368_) );
NAND2X1 NAND2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_9366_), .B(_9368_), .Y(_9369_) );
NOR2X1 NOR2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_9369_), .B(_9364_), .Y(_9370_) );
NOR2X1 NOR2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf0), .B(_9112_), .Y(_9371_) );
NAND3X1 NAND3X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_8649_), .B(_9371_), .C(_8647_), .Y(_9372_) );
NOR2X1 NOR2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8790_), .Y(_9373_) );
NAND3X1 NAND3X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8541_), .C(_8539_), .Y(_9374_) );
NAND2X1 NAND2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_9374_), .B(_9372_), .Y(_9375_) );
NOR2X1 NOR2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_9112_), .B(_8797_), .Y(_9376_) );
NAND3X1 NAND3X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8592_), .C(_8595_), .Y(_9377_) );
NOR2X1 NOR2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_9108_), .Y(_9378_) );
NAND3X1 NAND3X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_289_), .C(_292_), .Y(_9379_) );
NAND2X1 NAND2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_9377_), .B(_9379_), .Y(_9380_) );
NOR2X1 NOR2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_9380_), .B(_9375_), .Y(_9381_) );
NOR2X1 NOR2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_8749_), .B(_8897_), .Y(_9382_) );
NOR2X1 NOR2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8925_), .Y(_9383_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_22__0_), .B(_9382_), .C(_3__0_), .D(_9383_), .Y(_9384_) );
NAND3X1 NAND3X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_9370_), .B(_9381_), .C(_9384_), .Y(_9385_) );
NOR2X1 NOR2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_9385_), .B(_9359_), .Y(_9386_) );
NAND3X1 NAND3X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_9352_), .B(_9386_), .C(_9336_), .Y(_9387_) );
NOR3X1 NOR3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_9149_), .B(_9181_), .C(_9387_), .Y(_9388_) );
NAND3X1 NAND3X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_8887_), .B(_9388_), .C(_9096_), .Y(_9389_) );
NOR2X1 NOR2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_8761_), .B(_8854_), .Y(_9390_) );
NAND2X1 NAND2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__0_), .Y(_9391_) );
NOR2X1 NOR2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8797_), .Y(_9392_) );
NAND2X1 NAND2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__0_), .Y(_9393_) );
NAND2X1 NAND2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_9391_), .B(_9393_), .Y(_9394_) );
NOR3X1 NOR3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_8865_), .B(_9394_), .C(_9389_), .Y(_9395_) );
NOR2X1 NOR2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_8773_), .Y(_9396_) );
INVX4 INVX4_61 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .Y(_9397_) );
NOR3X1 NOR3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_9397_), .C(_1841_), .Y(_9398_) );
NOR2X1 NOR2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_8820__bF_buf2), .B(_8854_), .Y(_9399_) );
NAND3X1 NAND3X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_1313_), .C(_1311_), .Y(_9400_) );
NOR2X1 NOR2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8773_), .Y(_9401_) );
NAND3X1 NAND3X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1273_), .C(_1271_), .Y(_9402_) );
NAND2X1 NAND2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_9400_), .B(_9402_), .Y(_9403_) );
NOR2X1 NOR2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8854_), .Y(_9404_) );
NAND3X1 NAND3X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1490_), .C(_1486_), .Y(_9405_) );
NOR2X1 NOR2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8770_), .Y(_9406_) );
NAND3X1 NAND3X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1440_), .C(_1438_), .Y(_9407_) );
NAND2X1 NAND2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_9405_), .B(_9407_), .Y(_9408_) );
NOR2X1 NOR2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_9408_), .B(_9403_), .Y(_9409_) );
NOR2X1 NOR2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8797_), .Y(_9410_) );
NOR2X1 NOR2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8790_), .Y(_9411_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_125__0_), .B(_9411_), .C(_124__0_), .D(_9410_), .Y(_9412_) );
NOR2X1 NOR2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_9231_), .Y(_9413_) );
NAND3X1 NAND3X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_1082_), .B(_9413_), .C(_1080_), .Y(_9414_) );
NOR2X1 NOR2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_9265_), .B(_8854_), .Y(_9415_) );
NAND2X1 NAND2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__0_), .Y(_9416_) );
NAND3X1 NAND3X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_9414_), .B(_9416_), .C(_9412_), .Y(_9417_) );
NOR2X1 NOR2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8756_), .Y(_9418_) );
INVX4 INVX4_62 ( .gnd(gnd), .vdd(vdd), .A(_9418_), .Y(_9419_) );
NOR2X1 NOR2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8820__bF_buf1), .Y(_9420_) );
INVX4 INVX4_63 ( .gnd(gnd), .vdd(vdd), .A(_9420_), .Y(_9421_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_9421_), .C(_796_), .D(_9419_), .Y(_9422_) );
NOR2X1 NOR2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8730_), .Y(_9423_) );
INVX4 INVX4_64 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .Y(_9424_) );
NOR2X1 NOR2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8773_), .Y(_9425_) );
INVX4 INVX4_65 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .Y(_9426_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_9426_), .C(_682_), .D(_9424_), .Y(_9427_) );
NOR2X1 NOR2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_9422_), .B(_9427_), .Y(_9428_) );
NOR2X1 NOR2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8778_), .Y(_9429_) );
NAND3X1 NAND3X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_640_), .C(_644_), .Y(_9430_) );
NOR2X1 NOR2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_9108_), .B(_9231_), .Y(_9431_) );
NAND3X1 NAND3X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_9431_), .C(_521_), .Y(_9432_) );
NOR2X1 NOR2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_9023_), .B(_8773_), .Y(_9433_) );
NOR2X1 NOR2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_9265_), .Y(_9434_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_138__0_), .B(_9434_), .C(_229__0_), .D(_9433_), .Y(_9435_) );
NAND3X1 NAND3X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_9430_), .B(_9432_), .C(_9435_), .Y(_9436_) );
NOR2X1 NOR2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_8871_), .B(_8749_), .Y(_9437_) );
NAND3X1 NAND3X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7394_), .C(_7397_), .Y(_9438_) );
NOR2X1 NOR2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8749_), .Y(_9439_) );
INVX4 INVX4_66 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .Y(_9440_) );
OAI21X1 OAI21X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_9440_), .C(_9438_), .Y(_9441_) );
NOR2X1 NOR2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_9441_), .B(_9436_), .Y(_9442_) );
NAND2X1 NAND2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_9442_), .B(_9428_), .Y(_9443_) );
NOR2X1 NOR2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_8782__bF_buf3), .B(_8880_), .Y(_9444_) );
NAND3X1 NAND3X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_9444_), .C(_1039_), .Y(_9445_) );
NOR2X1 NOR2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8770_), .Y(_9446_) );
NAND2X1 NAND2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__0_), .Y(_9447_) );
NOR2X1 NOR2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8880_), .Y(_9448_) );
NOR2X1 NOR2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_8880_), .B(_8741_), .Y(_9449_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_130__0_), .B(_9449_), .C(_127__0_), .D(_9448_), .Y(_9450_) );
NAND3X1 NAND3X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_9445_), .B(_9447_), .C(_9450_), .Y(_9451_) );
NOR3X1 NOR3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_9451_), .B(_9417_), .C(_9443_), .Y(_9452_) );
NOR2X1 NOR2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8749_), .Y(_9453_) );
NOR2X1 NOR2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_8756_), .Y(_9454_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_114__0_), .B(_9454_), .C(_110__0_), .D(_9453_), .Y(_9455_) );
NAND3X1 NAND3X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_9409_), .B(_9455_), .C(_9452_), .Y(_9456_) );
NOR2X1 NOR2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_8854_), .B(_9231_), .Y(_9457_) );
NAND3X1 NAND3X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_1693_), .B(_9457_), .C(_1695_), .Y(_9458_) );
NOR2X1 NOR2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_8816_), .B(_9265_), .Y(_9459_) );
NAND2X1 NAND2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__0_), .Y(_9460_) );
NAND2X1 NAND2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_9460_), .B(_9458_), .Y(_9461_) );
NOR3X1 NOR3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_9461_), .B(_9398_), .C(_9456_), .Y(_9462_) );
NAND3X1 NAND3X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_8849_), .B(_9462_), .C(_9395_), .Y(_9463_) );
NOR2X1 NOR2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_8847_), .B(_9463_), .Y(_9464_) );
NAND3X1 NAND3X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_8828_), .B(_8839_), .C(_9464_), .Y(_9465_) );
NOR2X1 NOR2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8820__bF_buf0), .Y(_9466_) );
NAND2X1 NAND2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__0_), .Y(_9467_) );
NOR2X1 NOR2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8730_), .Y(_9468_) );
NAND3X1 NAND3X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_2419_), .B(_9468_), .C(_2421_), .Y(_9469_) );
NAND2X1 NAND2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_9467_), .B(_9469_), .Y(_9470_) );
NOR3X1 NOR3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_8808_), .B(_9470_), .C(_9465_), .Y(_9471_) );
NAND3X1 NAND3X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_8780_), .B(_8801_), .C(_9471_), .Y(_9472_) );
NOR2X1 NOR2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_8820__bF_buf3), .Y(_9473_) );
NAND3X1 NAND3X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_3040_), .B(_9473_), .C(_3041_), .Y(_9474_) );
NOR2X1 NOR2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_8735_), .B(_9265_), .Y(_9475_) );
NAND2X1 NAND2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__0_), .Y(_9476_) );
NOR2X1 NOR2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_9231_), .Y(_9477_) );
NOR2X1 NOR2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8756_), .Y(_9478_) );
NAND2X1 NAND2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__0_), .Y(_9479_) );
NOR2X1 NOR2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_8764_), .B(_8785_), .Y(_9480_) );
NAND2X1 NAND2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__0_), .Y(_9481_) );
NOR2X1 NOR2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_8785_), .B(_8741_), .Y(_9482_) );
NAND2X1 NAND2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__0_), .Y(_9483_) );
NAND3X1 NAND3X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_9483_), .B(_9479_), .C(_9481_), .Y(_9484_) );
AOI21X1 AOI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_68__0_), .B(_9477_), .C(_9484_), .Y(_9485_) );
NAND3X1 NAND3X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_9474_), .B(_9485_), .C(_9476_), .Y(_9486_) );
NOR3X1 NOR3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_8776_), .B(_9486_), .C(_9472_), .Y(_9487_) );
AOI21X1 AOI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_8760_), .B(_9487_), .C(rst), .Y(_0__0_) );
NAND2X1 NAND2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__1_), .Y(_9488_) );
NAND2X1 NAND2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__1_), .Y(_9489_) );
NAND2X1 NAND2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_9488_), .B(_9489_), .Y(_9490_) );
NAND2X1 NAND2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_55__1_), .Y(_9491_) );
NAND2X1 NAND2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__1_), .Y(_9492_) );
NAND2X1 NAND2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_9492_), .B(_9491_), .Y(_9493_) );
NOR2X1 NOR2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_9493_), .B(_9490_), .Y(_9494_) );
NAND3X1 NAND3X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .B(_8750_), .C(_3146_), .Y(_9495_) );
NAND3X1 NAND3X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .B(_8757_), .C(_3092_), .Y(_9496_) );
NAND2X1 NAND2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_9495_), .B(_9496_), .Y(_9497_) );
NAND3X1 NAND3X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_3261_), .B(_8762_), .C(_3260_), .Y(_9498_) );
NAND3X1 NAND3X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_2989_), .B(_8774_), .C(_2988_), .Y(_9499_) );
NAND2X1 NAND2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_9498_), .B(_9499_), .Y(_9500_) );
OR2X2 OR2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_9497_), .B(_9500_), .Y(_9501_) );
NAND2X1 NAND2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__1_), .Y(_9502_) );
NAND3X1 NAND3X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_2796_), .B(_8786_), .C(_2797_), .Y(_9503_) );
OAI21X1 OAI21X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .B(_8792_), .C(_9503_), .Y(_9504_) );
NAND3X1 NAND3X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_2626_), .B(_8794_), .C(_2627_), .Y(_9505_) );
OAI21X1 OAI21X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_2744_), .B(_8799_), .C(_9505_), .Y(_9506_) );
NOR2X1 NOR2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_9506_), .B(_9504_), .Y(_9507_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_76__1_), .B(_9482_), .C(_77__1_), .D(_9478_), .Y(_9508_) );
NAND2X1 NAND2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__1_), .Y(_9509_) );
NAND2X1 NAND2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_82__1_), .Y(_9510_) );
NAND3X1 NAND3X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_9509_), .B(_9510_), .C(_9508_), .Y(_9511_) );
NAND2X1 NAND2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__1_), .Y(_9512_) );
NAND3X1 NAND3X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_2575_), .B(_8803_), .C(_2574_), .Y(_9513_) );
NAND2X1 NAND2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_9513_), .B(_9512_), .Y(_9514_) );
INVX1 INVX1_3866 ( .gnd(gnd), .vdd(vdd), .A(_84__1_), .Y(_9515_) );
NOR2X1 NOR2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_9515_), .Y(_9516_) );
NOR2X1 NOR2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2284_), .Y(_9517_) );
NAND2X1 NAND2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__1_), .Y(_9518_) );
NAND3X1 NAND3X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_1994_), .B(_8843_), .C(_1995_), .Y(_9519_) );
NAND3X1 NAND3X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1895_), .C(_1896_), .Y(_9520_) );
NAND3X1 NAND3X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_9520_), .B(_9519_), .C(_9518_), .Y(_9521_) );
NOR3X1 NOR3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_9516_), .B(_9521_), .C(_9517_), .Y(_9522_) );
NAND3X1 NAND3X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_2233_), .B(_8829_), .C(_2234_), .Y(_9523_) );
NAND3X1 NAND3X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(_8831_), .C(_2128_), .Y(_9524_) );
NAND2X1 NAND2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_9523_), .B(_9524_), .Y(_9525_) );
NAND3X1 NAND3X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_2068_), .B(_8834_), .C(_2069_), .Y(_9526_) );
NAND3X1 NAND3X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .B(_8836_), .C(_2180_), .Y(_9527_) );
NAND2X1 NAND2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_9526_), .B(_9527_), .Y(_9528_) );
NOR2X1 NOR2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_9528_), .B(_9525_), .Y(_9529_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_98__1_), .B(_8845_), .C(_93__1_), .D(_8840_), .Y(_9530_) );
NAND2X1 NAND2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_91__1_), .Y(_9531_) );
NAND2X1 NAND2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_94__1_), .Y(_9532_) );
NAND3X1 NAND3X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_9531_), .B(_9532_), .C(_9530_), .Y(_9533_) );
NAND2X1 NAND2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__1_), .Y(_9534_) );
NAND3X1 NAND3X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1529_), .C(_1530_), .Y(_9535_) );
NAND3X1 NAND3X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1614_), .C(_1615_), .Y(_9536_) );
NAND2X1 NAND2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_9535_), .B(_9536_), .Y(_9537_) );
NAND3X1 NAND3X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1654_), .C(_1655_), .Y(_9538_) );
NAND3X1 NAND3X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_8857_), .C(_1363_), .Y(_9539_) );
NAND2X1 NAND2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_9539_), .B(_9538_), .Y(_9540_) );
OR2X2 OR2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_9537_), .B(_9540_), .Y(_9541_) );
NOR3X1 NOR3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_8867_), .C(_1201_), .Y(_9542_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_191__1_), .B(_8873_), .C(_192__1_), .D(_8872_), .Y(_9543_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_195__1_), .B(_8875_), .C(_193__1_), .D(_8876_), .Y(_9544_) );
NAND2X1 NAND2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_9543_), .B(_9544_), .Y(_9545_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_188__1_), .B(_8879_), .C(_126__1_), .D(_8881_), .Y(_9546_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_196__1_), .B(_8883_), .C(_194__1_), .D(_8884_), .Y(_9547_) );
NAND2X1 NAND2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_9546_), .B(_9547_), .Y(_9548_) );
NOR3X1 NOR3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_9548_), .B(_9542_), .C(_9545_), .Y(_9549_) );
NAND3X1 NAND3X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_5815_), .B(_8893_), .C(_5814_), .Y(_9550_) );
NAND3X1 NAND3X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_4575_), .B(_8898_), .C(_4574_), .Y(_9551_) );
NAND2X1 NAND2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_9550_), .B(_9551_), .Y(_9552_) );
NAND3X1 NAND3X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_5512_), .B(_8901_), .C(_5511_), .Y(_9553_) );
NAND3X1 NAND3X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_7850_), .B(_8904_), .C(_7849_), .Y(_9554_) );
NAND2X1 NAND2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_9553_), .B(_9554_), .Y(_9555_) );
NOR2X1 NOR2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_9552_), .B(_9555_), .Y(_9556_) );
NAND3X1 NAND3X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_4075_), .B(_8909_), .C(_4074_), .Y(_9557_) );
NAND3X1 NAND3X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3877_), .C(_3876_), .Y(_9558_) );
NAND2X1 NAND2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_9557_), .B(_9558_), .Y(_9559_) );
NAND3X1 NAND3X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_4616_), .B(_8914_), .C(_4615_), .Y(_9560_) );
NAND3X1 NAND3X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_6637_), .B(_8918_), .C(_6636_), .Y(_9561_) );
NAND2X1 NAND2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_9560_), .B(_9561_), .Y(_9562_) );
NOR2X1 NOR2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_9559_), .B(_9562_), .Y(_9563_) );
NAND2X1 NAND2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_9556_), .B(_9563_), .Y(_9564_) );
NAND3X1 NAND3X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_4956_), .B(_8926_), .C(_4955_), .Y(_9565_) );
NAND3X1 NAND3X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_8058_), .B(_8928_), .C(_8057_), .Y(_9566_) );
NAND2X1 NAND2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_9565_), .B(_9566_), .Y(_9567_) );
NAND3X1 NAND3X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_4478_), .B(_8931_), .C(_4477_), .Y(_9568_) );
NAND3X1 NAND3X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_8024_), .B(_8933_), .C(_8023_), .Y(_9569_) );
NAND2X1 NAND2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_9568_), .B(_9569_), .Y(_9570_) );
NOR2X1 NOR2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_9567_), .B(_9570_), .Y(_9571_) );
NAND3X1 NAND3X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_5170_), .B(_8937_), .C(_5169_), .Y(_9572_) );
NAND3X1 NAND3X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_7812_), .B(_8939_), .C(_7811_), .Y(_9573_) );
NAND2X1 NAND2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_9572_), .B(_9573_), .Y(_9574_) );
NAND3X1 NAND3X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_8942_), .C(_5131_), .Y(_9575_) );
NAND3X1 NAND3X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_8944_), .C(_4993_), .Y(_9576_) );
NAND2X1 NAND2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_9575_), .B(_9576_), .Y(_9577_) );
NOR2X1 NOR2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_9577_), .B(_9574_), .Y(_9578_) );
NAND2X1 NAND2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_9571_), .B(_9578_), .Y(_9579_) );
NOR2X1 NOR2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_9564_), .B(_9579_), .Y(_9580_) );
NAND3X1 NAND3X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_6708_), .B(_8950_), .C(_6707_), .Y(_9581_) );
NAND3X1 NAND3X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_3918_), .B(_8952_), .C(_3917_), .Y(_9582_) );
NAND2X1 NAND2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_9581_), .B(_9582_), .Y(_9583_) );
NAND3X1 NAND3X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_5887_), .B(_8955_), .C(_5886_), .Y(_9584_) );
NAND3X1 NAND3X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_6676_), .B(_8957_), .C(_6675_), .Y(_9585_) );
NAND2X1 NAND2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_9584_), .B(_9585_), .Y(_9586_) );
NOR2X1 NOR2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_9586_), .B(_9583_), .Y(_9587_) );
NAND3X1 NAND3X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_7778_), .B(_8961_), .C(_7777_), .Y(_9588_) );
NAND3X1 NAND3X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_3839_), .B(_8963_), .C(_3838_), .Y(_9589_) );
NAND2X1 NAND2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_9588_), .B(_9589_), .Y(_9590_) );
NAND3X1 NAND3X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_5853_), .B(_8966_), .C(_5852_), .Y(_9591_) );
NAND3X1 NAND3X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_3759_), .B(_8968_), .C(_3758_), .Y(_9592_) );
NAND2X1 NAND2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_9591_), .B(_9592_), .Y(_9593_) );
NOR2X1 NOR2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_9590_), .B(_9593_), .Y(_9594_) );
NAND2X1 NAND2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_9587_), .B(_9594_), .Y(_9595_) );
NAND3X1 NAND3X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_7960_), .B(_8973_), .C(_7959_), .Y(_9596_) );
NAND3X1 NAND3X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_3463_), .B(_8975_), .C(_3462_), .Y(_9597_) );
NAND2X1 NAND2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_9596_), .B(_9597_), .Y(_9598_) );
NAND3X1 NAND3X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .B(_8978_), .C(_4037_), .Y(_9599_) );
NAND3X1 NAND3X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_4112_), .B(_8980_), .C(_4111_), .Y(_9600_) );
NAND2X1 NAND2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_9600_), .B(_9599_), .Y(_9601_) );
NOR2X1 NOR2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_9598_), .B(_9601_), .Y(_9602_) );
NAND3X1 NAND3X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_5302_), .B(_8984_), .C(_5301_), .Y(_9603_) );
NAND3X1 NAND3X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(_8986_), .C(_5266_), .Y(_9604_) );
NAND2X1 NAND2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_9603_), .B(_9604_), .Y(_9605_) );
NAND3X1 NAND3X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_6564_), .B(_8989_), .C(_6563_), .Y(_9606_) );
NAND3X1 NAND3X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .B(_8991_), .C(_4147_), .Y(_9607_) );
NAND2X1 NAND2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_9606_), .B(_9607_), .Y(_9608_) );
NOR2X1 NOR2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_9605_), .B(_9608_), .Y(_9609_) );
NAND2X1 NAND2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_9602_), .B(_9609_), .Y(_9610_) );
NOR2X1 NOR2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_9595_), .B(_9610_), .Y(_9611_) );
NAND2X1 NAND2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_9580_), .B(_9611_), .Y(_9612_) );
NAND3X1 NAND3X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_8998_), .C(_4886_), .Y(_9613_) );
NAND3X1 NAND3X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_6494_), .B(_9002_), .C(_6493_), .Y(_9614_) );
NAND2X1 NAND2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_9613_), .B(_9614_), .Y(_9615_) );
NAND3X1 NAND3X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_5700_), .B(_9005_), .C(_5699_), .Y(_9616_) );
NAND3X1 NAND3X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .B(_9007_), .C(_4847_), .Y(_9617_) );
NAND2X1 NAND2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_9616_), .B(_9617_), .Y(_9618_) );
NOR2X1 NOR2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_9615_), .B(_9618_), .Y(_9619_) );
NAND3X1 NAND3X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_5738_), .B(_9011_), .C(_5737_), .Y(_9620_) );
NAND3X1 NAND3X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_6780_), .B(_9013_), .C(_6779_), .Y(_9621_) );
NAND2X1 NAND2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_9620_), .B(_9621_), .Y(_9622_) );
NAND3X1 NAND3X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_6741_), .B(_9016_), .C(_6740_), .Y(_9623_) );
NAND3X1 NAND3X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_6882_), .B(_9018_), .C(_6881_), .Y(_9624_) );
NAND2X1 NAND2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_9623_), .B(_9624_), .Y(_9625_) );
NOR2X1 NOR2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_9625_), .B(_9622_), .Y(_9626_) );
NAND2X1 NAND2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_9619_), .B(_9626_), .Y(_9627_) );
NAND3X1 NAND3X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_6264_), .B(_9024_), .C(_6263_), .Y(_9628_) );
NAND3X1 NAND3X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_6336_), .B(_9026_), .C(_6335_), .Y(_9629_) );
NAND2X1 NAND2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_9628_), .B(_9629_), .Y(_9630_) );
NAND3X1 NAND3X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_6041_), .B(_9029_), .C(_6040_), .Y(_9631_) );
NAND3X1 NAND3X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_6099_), .B(_9031_), .C(_6098_), .Y(_9632_) );
NAND2X1 NAND2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_9631_), .B(_9632_), .Y(_9633_) );
NOR2X1 NOR2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_9630_), .B(_9633_), .Y(_9634_) );
NAND3X1 NAND3X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_5659_), .B(_9035_), .C(_5658_), .Y(_9635_) );
NAND3X1 NAND3X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_4655_), .B(_9037_), .C(_4654_), .Y(_9636_) );
NAND2X1 NAND2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_9636_), .B(_9635_), .Y(_9637_) );
NAND3X1 NAND3X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_6300_), .B(_9040_), .C(_6299_), .Y(_9638_) );
NAND3X1 NAND3X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_4317_), .B(_9042_), .C(_4316_), .Y(_9639_) );
NAND2X1 NAND2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_9638_), .B(_9639_), .Y(_9640_) );
NOR2X1 NOR2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_9640_), .B(_9637_), .Y(_9641_) );
NAND2X1 NAND2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_9634_), .B(_9641_), .Y(_9642_) );
NOR2X1 NOR2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_9627_), .B(_9642_), .Y(_9643_) );
NAND3X1 NAND3X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_6188_), .B(_9048_), .C(_6187_), .Y(_9644_) );
NAND3X1 NAND3X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_7923_), .B(_9050_), .C(_7922_), .Y(_9645_) );
NAND2X1 NAND2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_9644_), .B(_9645_), .Y(_9646_) );
NAND3X1 NAND3X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_5472_), .B(_9053_), .C(_5471_), .Y(_9647_) );
NAND3X1 NAND3X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_7886_), .B(_9055_), .C(_7885_), .Y(_9648_) );
NAND2X1 NAND2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_9647_), .B(_9648_), .Y(_9649_) );
NOR2X1 NOR2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_9646_), .B(_9649_), .Y(_9650_) );
NAND3X1 NAND3X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_4438_), .B(_9059_), .C(_4437_), .Y(_9651_) );
NAND3X1 NAND3X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_4398_), .B(_9061_), .C(_4397_), .Y(_9652_) );
NAND2X1 NAND2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_9651_), .B(_9652_), .Y(_9653_) );
NAND3X1 NAND3X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_6226_), .B(_9064_), .C(_6225_), .Y(_9654_) );
NAND3X1 NAND3X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_4358_), .B(_9066_), .C(_4357_), .Y(_9655_) );
NAND2X1 NAND2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_9654_), .B(_9655_), .Y(_9656_) );
NOR2X1 NOR2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_9656_), .B(_9653_), .Y(_9657_) );
NAND2X1 NAND2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_9650_), .B(_9657_), .Y(_9658_) );
NAND3X1 NAND3X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_7582_), .B(_9071_), .C(_7581_), .Y(_9659_) );
NAND3X1 NAND3X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_7546_), .B(_9073_), .C(_7545_), .Y(_9660_) );
NAND2X1 NAND2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_9659_), .B(_9660_), .Y(_9661_) );
NAND3X1 NAND3X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_5776_), .B(_9076_), .C(_5775_), .Y(_9662_) );
NAND3X1 NAND3X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_9078_), .C(_3501_), .Y(_9663_) );
NAND2X1 NAND2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_9662_), .B(_9663_), .Y(_9664_) );
NOR2X1 NOR2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_9661_), .B(_9664_), .Y(_9665_) );
NAND3X1 NAND3X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_5431_), .B(_9082_), .C(_5430_), .Y(_9666_) );
NAND3X1 NAND3X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_3798_), .B(_9084_), .C(_3797_), .Y(_9667_) );
NAND2X1 NAND2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_9667_), .B(_9666_), .Y(_9668_) );
NAND3X1 NAND3X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_6597_), .B(_9087_), .C(_6596_), .Y(_9669_) );
NAND3X1 NAND3X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_3651_), .B(_9089_), .C(_3650_), .Y(_9670_) );
NAND2X1 NAND2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_9669_), .B(_9670_), .Y(_9671_) );
NOR2X1 NOR2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_9668_), .B(_9671_), .Y(_9672_) );
NAND2X1 NAND2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_9665_), .B(_9672_), .Y(_9673_) );
NOR2X1 NOR2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_9658_), .B(_9673_), .Y(_9674_) );
NAND2X1 NAND2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_9643_), .B(_9674_), .Y(_9675_) );
NOR2X1 NOR2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_9612_), .B(_9675_), .Y(_9676_) );
NAND2X1 NAND2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__1_), .Y(_9677_) );
NAND3X1 NAND3X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_3956_), .B(_9099_), .C(_3955_), .Y(_9678_) );
NAND2X1 NAND2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_9677_), .B(_9678_), .Y(_9679_) );
NAND3X1 NAND3X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_5080_), .B(_9102_), .C(_5079_), .Y(_9680_) );
NAND3X1 NAND3X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_6846_), .B(_9104_), .C(_6845_), .Y(_9681_) );
NAND2X1 NAND2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_9681_), .B(_9680_), .Y(_9682_) );
NOR2X1 NOR2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_9679_), .B(_9682_), .Y(_9683_) );
NAND3X1 NAND3X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_15905_), .B(_9109_), .C(_15906_), .Y(_9684_) );
NAND3X1 NAND3X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8369_), .B(_9113_), .C(_8370_), .Y(_9685_) );
NAND3X1 NAND3X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_16115_), .B(_9115_), .C(_16114_), .Y(_9686_) );
NAND3X1 NAND3X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_9684_), .B(_9685_), .C(_9686_), .Y(_9687_) );
NAND3X1 NAND3X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_376_), .C(_377_), .Y(_9688_) );
NAND3X1 NAND3X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_15847_), .B(_9120_), .C(_15848_), .Y(_9689_) );
AND2X2 AND2X2_1563 ( .gnd(gnd), .vdd(vdd), .A(_9689_), .B(_9688_), .Y(_9690_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_201__1_), .B(_9124_), .C(_89__1_), .D(_9123_), .Y(_9691_) );
NAND2X1 NAND2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_9690_), .B(_9691_), .Y(_9692_) );
NAND3X1 NAND3X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_4732_), .B(_9127_), .C(_4733_), .Y(_9693_) );
NAND3X1 NAND3X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_3993_), .B(_9129_), .C(_3994_), .Y(_9694_) );
NAND2X1 NAND2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_9694_), .B(_9693_), .Y(_9695_) );
NOR3X1 NOR3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_9687_), .B(_9695_), .C(_9692_), .Y(_9696_) );
NAND3X1 NAND3X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3404_), .C(_3405_), .Y(_9697_) );
NAND3X1 NAND3X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_5030_), .B(_9135_), .C(_5031_), .Y(_9698_) );
NAND3X1 NAND3X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_6915_), .B(_9137_), .C(_6916_), .Y(_9699_) );
NAND3X1 NAND3X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_9698_), .B(_9699_), .C(_9697_), .Y(_9700_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .B(_9140_), .C(_2__1_), .D(_9141_), .Y(_9701_) );
NAND2X1 NAND2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__1_), .Y(_9702_) );
NAND2X1 NAND2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_200__1_), .Y(_9703_) );
NAND3X1 NAND3X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_9702_), .B(_9703_), .C(_9701_), .Y(_9704_) );
NOR2X1 NOR2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_9700_), .B(_9704_), .Y(_9705_) );
NAND3X1 NAND3X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_9683_), .B(_9705_), .C(_9696_), .Y(_9706_) );
AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_21__1_), .B(_9150_), .C(_185__1_), .D(_9151_), .Y(_9707_) );
AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_243__1_), .B(_9153_), .C(_253__1_), .D(_9154_), .Y(_9708_) );
NAND2X1 NAND2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_9707_), .B(_9708_), .Y(_9709_) );
AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_46__1_), .B(_9158_), .C(_231__1_), .D(_9157_), .Y(_9710_) );
AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .B(_9161_), .C(_244__1_), .D(_9160_), .Y(_9711_) );
NAND2X1 NAND2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_9711_), .B(_9710_), .Y(_9712_) );
NOR2X1 NOR2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_9709_), .B(_9712_), .Y(_9713_) );
NAND2X1 NAND2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_247__1_), .Y(_9714_) );
NAND2X1 NAND2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_9167_), .B(_30__1_), .Y(_9715_) );
AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_218__1_), .B(_9169_), .C(_227__1_), .D(_9170_), .Y(_9716_) );
NAND3X1 NAND3X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_9714_), .B(_9715_), .C(_9716_), .Y(_9717_) );
AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_178__1_), .B(_9173_), .C(_214__1_), .D(_9174_), .Y(_9718_) );
AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_145__1_), .B(_9177_), .C(_29__1_), .D(_9176_), .Y(_9719_) );
NAND2X1 NAND2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_9718_), .B(_9719_), .Y(_9720_) );
NOR2X1 NOR2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_9720_), .B(_9717_), .Y(_9721_) );
NAND2X1 NAND2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_9713_), .B(_9721_), .Y(_9722_) );
AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_234__1_), .B(_9182_), .C(_34__1_), .D(_9183_), .Y(_9723_) );
NAND2X1 NAND2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__1_), .Y(_9724_) );
NAND2X1 NAND2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__1_), .Y(_9725_) );
NAND3X1 NAND3X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_9724_), .B(_9725_), .C(_9723_), .Y(_9726_) );
NAND3X1 NAND3X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_15637_), .B(_9192_), .C(_15638_), .Y(_9727_) );
OAI21X1 OAI21X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_15589_), .B(_9195_), .C(_9727_), .Y(_9728_) );
NAND2X1 NAND2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__1_), .Y(_9729_) );
NAND3X1 NAND3X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_15693_), .B(_9199_), .C(_15694_), .Y(_9730_) );
NAND2X1 NAND2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_9729_), .B(_9730_), .Y(_9731_) );
NOR2X1 NOR2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_9731_), .B(_9728_), .Y(_9732_) );
NAND2X1 NAND2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__1_), .Y(_9733_) );
OAI21X1 OAI21X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_15292_), .B(_9206_), .C(_9733_), .Y(_9734_) );
NAND2X1 NAND2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__1_), .Y(_9735_) );
OAI21X1 OAI21X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_15090_), .B(_9211_), .C(_9735_), .Y(_9736_) );
NOR2X1 NOR2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_9734_), .B(_9736_), .Y(_9737_) );
NOR3X1 NOR3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_15960_), .B(_9215_), .C(_15961_), .Y(_9738_) );
NAND3X1 NAND3X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_15240_), .B(_9217_), .C(_15241_), .Y(_9739_) );
NAND3X1 NAND3X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_15188_), .B(_9219_), .C(_15187_), .Y(_9740_) );
NAND2X1 NAND2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_9740_), .B(_9739_), .Y(_9741_) );
NAND3X1 NAND3X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_15462_), .B(_9222_), .C(_15463_), .Y(_9742_) );
NAND3X1 NAND3X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_15409_), .B(_9224_), .C(_15408_), .Y(_9743_) );
NAND2X1 NAND2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_9742_), .B(_9743_), .Y(_9744_) );
NOR3X1 NOR3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_9738_), .B(_9744_), .C(_9741_), .Y(_9745_) );
NAND3X1 NAND3X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_9737_), .B(_9745_), .C(_9732_), .Y(_9746_) );
NAND3X1 NAND3X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_8478_), .B(_9229_), .C(_8479_), .Y(_9747_) );
NAND3X1 NAND3X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_15520_), .B(_9233_), .C(_15521_), .Y(_9748_) );
NAND2X1 NAND2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .B(_49__1_), .Y(_9749_) );
NAND2X1 NAND2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__1_), .Y(_9750_) );
NAND2X1 NAND2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__1_), .Y(_9751_) );
NAND3X1 NAND3X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_9750_), .B(_9751_), .C(_9749_), .Y(_9752_) );
NAND3X1 NAND3X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_7698_), .B(_9248_), .C(_7700_), .Y(_9753_) );
OAI21X1 OAI21X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_8151_), .B(_9304_), .C(_9753_), .Y(_9754_) );
NAND2X1 NAND2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__1_), .Y(_9755_) );
NAND2X1 NAND2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .B(_186__1_), .Y(_9756_) );
NAND2X1 NAND2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_9755_), .B(_9756_), .Y(_9757_) );
NOR2X1 NOR2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_9757_), .B(_9754_), .Y(_9758_) );
AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_101__1_), .B(_9255_), .C(_197__1_), .D(_9244_), .Y(_9759_) );
AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_65__1_), .B(_9277_), .C(_119__1_), .D(_9268_), .Y(_9760_) );
NAND3X1 NAND3X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_9759_), .B(_9760_), .C(_9758_), .Y(_9761_) );
NOR2X1 NOR2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_9752_), .B(_9761_), .Y(_9762_) );
INVX4 INVX4_67 ( .gnd(gnd), .vdd(vdd), .A(_9281_), .Y(_9763_) );
NOR2X1 NOR2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_9763_), .B(_6413_), .Y(_9764_) );
OR2X2 OR2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_9238_), .B(_9241_), .Y(_9765_) );
NAND3X1 NAND3X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_8219_), .B(_9250_), .C(_8218_), .Y(_9766_) );
OAI21X1 OAI21X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_8699_), .C(_9766_), .Y(_9767_) );
NAND3X1 NAND3X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_7659_), .B(_9321_), .C(_7660_), .Y(_9768_) );
OAI21X1 OAI21X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_5916_), .B(_9323_), .C(_9768_), .Y(_9769_) );
NOR3X1 NOR3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_9764_), .B(_9767_), .C(_9769_), .Y(_9770_) );
NAND2X1 NAND2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_9262_), .B(_137__1_), .Y(_9771_) );
NAND2X1 NAND2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(_154__1_), .Y(_9772_) );
NAND2X1 NAND2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_9771_), .B(_9772_), .Y(_9773_) );
NAND3X1 NAND3X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_7029_), .B(_9266_), .C(_7031_), .Y(_9774_) );
OAI21X1 OAI21X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_4175_), .B(_9254_), .C(_9774_), .Y(_9775_) );
NOR2X1 NOR2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_9775_), .B(_9773_), .Y(_9776_) );
AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_173__1_), .B(_9275_), .C(_187__1_), .D(_9235_), .Y(_9777_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .Y(_9778_) );
AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_182__1_), .B(_9300_), .C(_50__1_), .D(_9778_), .Y(_9779_) );
AND2X2 AND2X2_1564 ( .gnd(gnd), .vdd(vdd), .A(_9777_), .B(_9779_), .Y(_9780_) );
NAND3X1 NAND3X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_9770_), .B(_9776_), .C(_9780_), .Y(_9781_) );
AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_233__1_), .B(_9310_), .C(_251__1_), .D(_9320_), .Y(_9782_) );
OAI21X1 OAI21X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_4206_), .B(_9282_), .C(_9782_), .Y(_9783_) );
AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_252__1_), .B(_9326_), .C(_15__1_), .D(_9313_), .Y(_9784_) );
AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .B(_9274_), .C(_83__1_), .D(_9315_), .Y(_9785_) );
NAND2X1 NAND2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_9785_), .B(_9784_), .Y(_9786_) );
OR2X2 OR2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_9783_), .B(_9786_), .Y(_9787_) );
NOR2X1 NOR2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_9787_), .B(_9781_), .Y(_9788_) );
NAND3X1 NAND3X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_9748_), .B(_9762_), .C(_9788_), .Y(_9789_) );
AOI21X1 AOI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_157__1_), .B(_9232_), .C(_9789_), .Y(_9790_) );
AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_155__1_), .B(_9333_), .C(_172__1_), .D(_9332_), .Y(_9791_) );
NAND3X1 NAND3X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_9747_), .B(_9791_), .C(_9790_), .Y(_9792_) );
NOR3X1 NOR3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_9792_), .B(_9726_), .C(_9746_), .Y(_9793_) );
NAND2X1 NAND2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__1_), .Y(_9794_) );
NAND3X1 NAND3X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_9339_), .C(_431_), .Y(_9795_) );
AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_111__1_), .B(_9342_), .C(_12__1_), .D(_9341_), .Y(_9796_) );
NAND3X1 NAND3X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_9796_), .B(_9794_), .C(_9795_), .Y(_9797_) );
AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_100__1_), .B(_9346_), .C(_212__1_), .D(_9345_), .Y(_9798_) );
AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_245__1_), .B(_9348_), .C(_140__1_), .D(_9349_), .Y(_9799_) );
NAND2X1 NAND2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_9799_), .B(_9798_), .Y(_9800_) );
NOR2X1 NOR2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_9797_), .B(_9800_), .Y(_9801_) );
AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_232__1_), .B(_9354_), .C(_219__1_), .D(_9353_), .Y(_9802_) );
AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_246__1_), .B(_9356_), .C(_226__1_), .D(_9357_), .Y(_9803_) );
NAND2X1 NAND2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_9803_), .B(_9802_), .Y(_9804_) );
NAND3X1 NAND3X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16168_), .C(_16169_), .Y(_9805_) );
OAI21X1 OAI21X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_16218_), .B(_9361_), .C(_9805_), .Y(_9806_) );
NAND3X1 NAND3X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16065_), .C(_16066_), .Y(_9807_) );
NAND3X1 NAND3X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16010_), .C(_16011_), .Y(_9808_) );
NAND2X1 NAND2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_9807_), .B(_9808_), .Y(_9809_) );
NOR2X1 NOR2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_9809_), .B(_9806_), .Y(_9810_) );
NAND3X1 NAND3X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_8652_), .B(_9371_), .C(_8651_), .Y(_9811_) );
NAND3X1 NAND3X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8544_), .C(_8543_), .Y(_9812_) );
NAND2X1 NAND2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_9812_), .B(_9811_), .Y(_9813_) );
NAND3X1 NAND3X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8597_), .C(_8598_), .Y(_9814_) );
NAND3X1 NAND3X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_294_), .C(_295_), .Y(_9815_) );
NAND2X1 NAND2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_9814_), .B(_9815_), .Y(_9816_) );
NOR2X1 NOR2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_9816_), .B(_9813_), .Y(_9817_) );
AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_22__1_), .B(_9382_), .C(_3__1_), .D(_9383_), .Y(_9818_) );
NAND3X1 NAND3X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_9810_), .B(_9817_), .C(_9818_), .Y(_9819_) );
NOR2X1 NOR2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_9819_), .B(_9804_), .Y(_9820_) );
NAND3X1 NAND3X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_9801_), .B(_9820_), .C(_9793_), .Y(_9821_) );
NOR3X1 NOR3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_9706_), .B(_9722_), .C(_9821_), .Y(_9822_) );
NAND3X1 NAND3X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_9549_), .B(_9822_), .C(_9676_), .Y(_9823_) );
NAND2X1 NAND2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__1_), .Y(_9824_) );
NAND2X1 NAND2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__1_), .Y(_9825_) );
NAND2X1 NAND2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_9825_), .B(_9824_), .Y(_9826_) );
NOR3X1 NOR3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_9541_), .B(_9826_), .C(_9823_), .Y(_9827_) );
NOR3X1 NOR3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_9397_), .C(_1843_), .Y(_9828_) );
NAND3X1 NAND3X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1443_), .C(_1442_), .Y(_9829_) );
NAND3X1 NAND3X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_9453_), .B(_1399_), .C(_1397_), .Y(_9830_) );
NAND2X1 NAND2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_9829_), .B(_9830_), .Y(_9831_) );
NAND3X1 NAND3X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1493_), .C(_1492_), .Y(_9832_) );
NAND3X1 NAND3X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1276_), .C(_1275_), .Y(_9833_) );
NAND2X1 NAND2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_9832_), .B(_9833_), .Y(_9834_) );
NOR2X1 NOR2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_9834_), .B(_9831_), .Y(_9835_) );
AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_125__1_), .B(_9411_), .C(_124__1_), .D(_9410_), .Y(_9836_) );
NAND3X1 NAND3X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_9413_), .C(_1084_), .Y(_9837_) );
NAND2X1 NAND2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__1_), .Y(_9838_) );
NAND3X1 NAND3X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_9837_), .B(_9838_), .C(_9836_), .Y(_9839_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_9421_), .C(_799_), .D(_9419_), .Y(_9840_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_9426_), .C(_685_), .D(_9424_), .Y(_9841_) );
NOR2X1 NOR2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_9840_), .B(_9841_), .Y(_9842_) );
NAND3X1 NAND3X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_646_), .C(_647_), .Y(_9843_) );
NAND3X1 NAND3X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_9431_), .C(_524_), .Y(_9844_) );
AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_138__1_), .B(_9434_), .C(_229__1_), .D(_9433_), .Y(_9845_) );
NAND3X1 NAND3X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_9843_), .B(_9844_), .C(_9845_), .Y(_9846_) );
NAND3X1 NAND3X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7399_), .C(_7400_), .Y(_9847_) );
OAI21X1 OAI21X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_9440_), .C(_9847_), .Y(_9848_) );
NOR2X1 NOR2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_9848_), .B(_9846_), .Y(_9849_) );
NAND2X1 NAND2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_9849_), .B(_9842_), .Y(_9850_) );
NAND3X1 NAND3X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_9444_), .C(_1043_), .Y(_9851_) );
NAND2X1 NAND2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__1_), .Y(_9852_) );
AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_130__1_), .B(_9449_), .C(_127__1_), .D(_9448_), .Y(_9853_) );
NAND3X1 NAND3X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_9851_), .B(_9852_), .C(_9853_), .Y(_9854_) );
NOR3X1 NOR3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_9854_), .B(_9839_), .C(_9850_), .Y(_9855_) );
AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_115__1_), .B(_9399_), .C(_114__1_), .D(_9454_), .Y(_9856_) );
NAND3X1 NAND3X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_9856_), .B(_9835_), .C(_9855_), .Y(_9857_) );
NAND3X1 NAND3X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_9457_), .C(_1698_), .Y(_9858_) );
NAND2X1 NAND2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__1_), .Y(_9859_) );
NAND2X1 NAND2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_9859_), .B(_9858_), .Y(_9860_) );
NOR3X1 NOR3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_9860_), .B(_9828_), .C(_9857_), .Y(_9861_) );
NAND3X1 NAND3X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_9534_), .B(_9861_), .C(_9827_), .Y(_9862_) );
NOR2X1 NOR2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_9533_), .B(_9862_), .Y(_9863_) );
NAND3X1 NAND3X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_9522_), .B(_9529_), .C(_9863_), .Y(_9864_) );
NOR3X1 NOR3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_9511_), .B(_9514_), .C(_9864_), .Y(_9865_) );
NAND3X1 NAND3X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_9502_), .B(_9507_), .C(_9865_), .Y(_9866_) );
NAND3X1 NAND3X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_3043_), .B(_9473_), .C(_3044_), .Y(_9867_) );
NAND2X1 NAND2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__1_), .Y(_9868_) );
NAND2X1 NAND2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__1_), .Y(_9869_) );
NAND2X1 NAND2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__1_), .Y(_9870_) );
NAND3X1 NAND3X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_9468_), .C(_2424_), .Y(_9871_) );
NAND3X1 NAND3X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_9869_), .B(_9870_), .C(_9871_), .Y(_9872_) );
AOI21X1 AOI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_68__1_), .B(_9477_), .C(_9872_), .Y(_9873_) );
NAND3X1 NAND3X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_9873_), .B(_9867_), .C(_9868_), .Y(_9874_) );
NOR3X1 NOR3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_9501_), .B(_9874_), .C(_9866_), .Y(_9875_) );
AOI21X1 AOI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_9494_), .B(_9875_), .C(rst), .Y(_0__1_) );
NAND2X1 NAND2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__2_), .Y(_9876_) );
NAND2X1 NAND2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__2_), .Y(_9877_) );
NAND2X1 NAND2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_9876_), .B(_9877_), .Y(_9878_) );
NAND2X1 NAND2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_55__2_), .Y(_9879_) );
NAND2X1 NAND2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__2_), .Y(_9880_) );
NAND2X1 NAND2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_9880_), .B(_9879_), .Y(_9881_) );
NOR2X1 NOR2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_9881_), .B(_9878_), .Y(_9882_) );
NAND3X1 NAND3X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_3151_), .B(_8750_), .C(_3150_), .Y(_9883_) );
NAND3X1 NAND3X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_3097_), .B(_8757_), .C(_3096_), .Y(_9884_) );
NAND2X1 NAND2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_9883_), .B(_9884_), .Y(_9885_) );
NAND3X1 NAND3X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_3264_), .B(_8762_), .C(_3263_), .Y(_9886_) );
NAND3X1 NAND3X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_8774_), .C(_2991_), .Y(_9887_) );
NAND2X1 NAND2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_9886_), .B(_9887_), .Y(_9888_) );
OR2X2 OR2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_9885_), .B(_9888_), .Y(_9889_) );
NAND2X1 NAND2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__2_), .Y(_9890_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .B(_8799_), .C(_2691_), .D(_8792_), .Y(_9891_) );
NAND3X1 NAND3X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_8794_), .C(_2630_), .Y(_9892_) );
NAND3X1 NAND3X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_2799_), .B(_8786_), .C(_2800_), .Y(_9893_) );
NAND2X1 NAND2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_9892_), .B(_9893_), .Y(_9894_) );
NOR2X1 NOR2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_9891_), .B(_9894_), .Y(_9895_) );
AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_77__2_), .B(_9478_), .C(_80__2_), .D(_8805_), .Y(_9896_) );
AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .B(_8806_), .C(_79__2_), .D(_9466_), .Y(_9897_) );
NAND2X1 NAND2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_9897_), .B(_9896_), .Y(_9898_) );
NAND2X1 NAND2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__2_), .Y(_9899_) );
NAND3X1 NAND3X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_2577_), .B(_8803_), .C(_2576_), .Y(_9900_) );
NAND2X1 NAND2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_9900_), .B(_9899_), .Y(_9901_) );
INVX1 INVX1_3867 ( .gnd(gnd), .vdd(vdd), .A(_84__2_), .Y(_9902_) );
NOR2X1 NOR2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_9902_), .Y(_9903_) );
NOR2X1 NOR2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2286_), .Y(_9904_) );
NAND2X1 NAND2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__2_), .Y(_9905_) );
NAND3X1 NAND3X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1898_), .C(_1899_), .Y(_9906_) );
NAND2X1 NAND2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_98__2_), .Y(_9907_) );
NAND3X1 NAND3X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_9906_), .B(_9905_), .C(_9907_), .Y(_9908_) );
NOR3X1 NOR3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_9903_), .B(_9908_), .C(_9904_), .Y(_9909_) );
NAND3X1 NAND3X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .B(_8829_), .C(_2237_), .Y(_9910_) );
NAND3X1 NAND3X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_2130_), .B(_8831_), .C(_2131_), .Y(_9911_) );
NAND2X1 NAND2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_9910_), .B(_9911_), .Y(_9912_) );
NAND3X1 NAND3X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_8834_), .C(_2072_), .Y(_9913_) );
NAND3X1 NAND3X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_2182_), .B(_8836_), .C(_2183_), .Y(_9914_) );
NAND2X1 NAND2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_9913_), .B(_9914_), .Y(_9915_) );
NOR2X1 NOR2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_9915_), .B(_9912_), .Y(_9916_) );
AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_92__2_), .B(_8843_), .C(_91__2_), .D(_8823_), .Y(_9917_) );
AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_94__2_), .B(_8841_), .C(_93__2_), .D(_8840_), .Y(_9918_) );
NAND2X1 NAND2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_9918_), .B(_9917_), .Y(_9919_) );
NAND2X1 NAND2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__2_), .Y(_9920_) );
NAND2X1 NAND2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__2_), .Y(_9921_) );
NAND2X1 NAND2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__2_), .Y(_9922_) );
NAND2X1 NAND2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9921_), .B(_9922_), .Y(_9923_) );
NAND2X1 NAND2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__2_), .Y(_9924_) );
NAND2X1 NAND2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__2_), .Y(_9925_) );
NAND2X1 NAND2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_9925_), .B(_9924_), .Y(_9926_) );
NOR2X1 NOR2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_9926_), .B(_9923_), .Y(_9927_) );
NAND2X1 NAND2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__2_), .Y(_9928_) );
INVX4 INVX4_68 ( .gnd(gnd), .vdd(vdd), .A(_8875_), .Y(_9929_) );
INVX4 INVX4_69 ( .gnd(gnd), .vdd(vdd), .A(_8883_), .Y(_9930_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_7130_), .B(_9930_), .C(_7174_), .D(_9929_), .Y(_9931_) );
INVX4 INVX4_70 ( .gnd(gnd), .vdd(vdd), .A(_8872_), .Y(_9932_) );
NOR2X1 NOR2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7309_), .Y(_9933_) );
INVX4 INVX4_71 ( .gnd(gnd), .vdd(vdd), .A(_8876_), .Y(_9934_) );
NOR2X1 NOR2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7266_), .Y(_9935_) );
NOR3X1 NOR3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_9933_), .B(_9935_), .C(_9931_), .Y(_9936_) );
NAND2X1 NAND2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__2_), .Y(_9937_) );
NAND2X1 NAND2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__2_), .Y(_9938_) );
NAND2X1 NAND2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_9937_), .B(_9938_), .Y(_9939_) );
INVX4 INVX4_72 ( .gnd(gnd), .vdd(vdd), .A(_8873_), .Y(_9940_) );
INVX4 INVX4_73 ( .gnd(gnd), .vdd(vdd), .A(_8884_), .Y(_9941_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_7352_), .B(_9940_), .C(_7220_), .D(_9941_), .Y(_9942_) );
NOR2X1 NOR2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_9942_), .B(_9939_), .Y(_9943_) );
NAND3X1 NAND3X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_9928_), .B(_9936_), .C(_9943_), .Y(_9944_) );
AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_20__2_), .B(_8898_), .C(_236__2_), .D(_8955_), .Y(_9945_) );
AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_237__2_), .B(_8966_), .C(_175__2_), .D(_8904_), .Y(_9946_) );
NAND2X1 NAND2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_9945_), .B(_9946_), .Y(_9947_) );
NAND2X1 NAND2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__2_), .Y(_9948_) );
NAND2X1 NAND2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__2_), .Y(_9949_) );
AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_19__2_), .B(_8914_), .C(_210__2_), .D(_8918_), .Y(_9950_) );
NAND3X1 NAND3X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_9948_), .B(_9949_), .C(_9950_), .Y(_9951_) );
NOR2X1 NOR2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_9947_), .B(_9951_), .Y(_9952_) );
AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_123__2_), .B(_8928_), .C(_9__2_), .D(_8926_), .Y(_9953_) );
NAND2X1 NAND2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__2_), .Y(_9954_) );
NAND2X1 NAND2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_134__2_), .Y(_9955_) );
NAND3X1 NAND3X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_9954_), .B(_9955_), .C(_9953_), .Y(_9956_) );
AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_4__2_), .B(_8937_), .C(_176__2_), .D(_8939_), .Y(_9957_) );
NAND2X1 NAND2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__2_), .Y(_9958_) );
NAND2X1 NAND2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__2_), .Y(_9959_) );
NAND3X1 NAND3X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_9958_), .B(_9959_), .C(_9957_), .Y(_9960_) );
NOR2X1 NOR2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_9960_), .B(_9956_), .Y(_9961_) );
NAND2X1 NAND2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_9952_), .B(_9961_), .Y(_9962_) );
NAND2X1 NAND2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_9082_), .B(_250__2_), .Y(_9963_) );
NAND2X1 NAND2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_47__2_), .Y(_9964_) );
AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_21__2_), .B(_9150_), .C(_185__2_), .D(_9151_), .Y(_9965_) );
NAND3X1 NAND3X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_9963_), .B(_9964_), .C(_9965_), .Y(_9966_) );
AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_246__2_), .B(_9356_), .C(_226__2_), .D(_9357_), .Y(_9967_) );
NAND2X1 NAND2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_9157_), .B(_231__2_), .Y(_9968_) );
NAND2X1 NAND2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_46__2_), .Y(_9969_) );
NAND3X1 NAND3X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_9968_), .B(_9969_), .C(_9967_), .Y(_9970_) );
NOR2X1 NOR2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_9966_), .B(_9970_), .Y(_9971_) );
NAND2X1 NAND2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_178__2_), .Y(_9972_) );
NAND2X1 NAND2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__2_), .Y(_9973_) );
AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_37__2_), .B(_8978_), .C(_35__2_), .D(_8980_), .Y(_9974_) );
NAND3X1 NAND3X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_9972_), .B(_9973_), .C(_9974_), .Y(_9975_) );
NAND2X1 NAND2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .B(_249__2_), .Y(_9976_) );
NAND2X1 NAND2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_253__2_), .Y(_9977_) );
AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_145__2_), .B(_9177_), .C(_213__2_), .D(_8989_), .Y(_9978_) );
NAND3X1 NAND3X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_9976_), .B(_9977_), .C(_9978_), .Y(_9979_) );
NOR2X1 NOR2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_9979_), .B(_9975_), .Y(_9980_) );
NAND2X1 NAND2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_9971_), .B(_9980_), .Y(_9981_) );
NOR2X1 NOR2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_9962_), .B(_9981_), .Y(_9982_) );
NAND2X1 NAND2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__2_), .Y(_9983_) );
NAND2X1 NAND2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__2_), .Y(_9984_) );
AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_13__2_), .B(_9007_), .C(_239__2_), .D(_9076_), .Y(_9985_) );
NAND3X1 NAND3X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_9983_), .B(_9984_), .C(_9985_), .Y(_9986_) );
AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_206__2_), .B(_9013_), .C(_242__2_), .D(_9035_), .Y(_9987_) );
NAND2X1 NAND2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__2_), .Y(_9988_) );
NAND2X1 NAND2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__2_), .Y(_9989_) );
NAND3X1 NAND3X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_9988_), .B(_9989_), .C(_9987_), .Y(_9990_) );
NOR2X1 NOR2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_9986_), .B(_9990_), .Y(_9991_) );
AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_222__2_), .B(_9024_), .C(_220__2_), .D(_9026_), .Y(_9992_) );
NAND2X1 NAND2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__2_), .Y(_9993_) );
NAND2X1 NAND2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__2_), .Y(_9994_) );
NAND3X1 NAND3X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_9993_), .B(_9994_), .C(_9992_), .Y(_9995_) );
AOI22X1 AOI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_18__2_), .B(_9037_), .C(_240__2_), .D(_9011_), .Y(_9996_) );
NAND2X1 NAND2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__2_), .Y(_9997_) );
NAND2X1 NAND2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__2_), .Y(_9998_) );
NAND3X1 NAND3X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_9997_), .B(_9998_), .C(_9996_), .Y(_9999_) );
NOR2X1 NOR2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_9995_), .B(_9999_), .Y(_10000_) );
NAND2X1 NAND2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_9991_), .B(_10000_), .Y(_10001_) );
AOI22X1 AOI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_225__2_), .B(_9048_), .C(_167__2_), .D(_9050_), .Y(_10002_) );
NAND2X1 NAND2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_243__2_), .Y(_10003_) );
NAND2X1 NAND2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__2_), .Y(_10004_) );
NAND3X1 NAND3X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_10003_), .B(_10004_), .C(_10002_), .Y(_10005_) );
NAND2X1 NAND2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__2_), .Y(_10006_) );
NAND2X1 NAND2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__2_), .Y(_10007_) );
AOI22X1 AOI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_224__2_), .B(_9064_), .C(_27__2_), .D(_9066_), .Y(_10008_) );
NAND3X1 NAND3X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_10006_), .B(_10007_), .C(_10008_), .Y(_10009_) );
NOR2X1 NOR2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_10005_), .B(_10009_), .Y(_10010_) );
AOI22X1 AOI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_184__2_), .B(_9073_), .C(_183__2_), .D(_9071_), .Y(_10011_) );
NAND2X1 NAND2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__2_), .Y(_10012_) );
NAND2X1 NAND2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__2_), .Y(_10013_) );
NAND3X1 NAND3X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_10012_), .B(_10013_), .C(_10011_), .Y(_10014_) );
AOI22X1 AOI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_43__2_), .B(_9084_), .C(_244__2_), .D(_9160_), .Y(_10015_) );
NAND2X1 NAND2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__2_), .Y(_10016_) );
NAND2X1 NAND2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__2_), .Y(_10017_) );
NAND3X1 NAND3X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_10016_), .B(_10017_), .C(_10015_), .Y(_10018_) );
NOR2X1 NOR2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_10014_), .B(_10018_), .Y(_10019_) );
NAND2X1 NAND2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_10010_), .B(_10019_), .Y(_10020_) );
NOR2X1 NOR2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_10001_), .B(_10020_), .Y(_10021_) );
NAND3X1 NAND3X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_6817_), .B(_9143_), .C(_6818_), .Y(_10022_) );
NAND3X1 NAND3X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_6963_), .B(_9145_), .C(_6965_), .Y(_10023_) );
NAND2X1 NAND2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_10022_), .B(_10023_), .Y(_10024_) );
NAND3X1 NAND3X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_5033_), .B(_9135_), .C(_5034_), .Y(_10025_) );
NAND3X1 NAND3X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_6918_), .B(_9137_), .C(_6919_), .Y(_10026_) );
NAND2X1 NAND2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_10026_), .B(_10025_), .Y(_10027_) );
NOR2X1 NOR2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_10024_), .B(_10027_), .Y(_10028_) );
NAND3X1 NAND3X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_8308_), .B(_9188_), .C(_8310_), .Y(_10029_) );
NAND3X1 NAND3X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_15908_), .B(_9109_), .C(_15909_), .Y(_10030_) );
NAND3X1 NAND3X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_16117_), .B(_9115_), .C(_16118_), .Y(_10031_) );
NAND3X1 NAND3X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_10030_), .B(_10031_), .C(_10029_), .Y(_10032_) );
AOI22X1 AOI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_234__2_), .B(_9182_), .C(_34__2_), .D(_9183_), .Y(_10033_) );
AOI22X1 AOI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_100__2_), .B(_9346_), .C(_45__2_), .D(_9185_), .Y(_10034_) );
NAND2X1 NAND2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_10034_), .B(_10033_), .Y(_10035_) );
INVX4 INVX4_74 ( .gnd(gnd), .vdd(vdd), .A(_9141_), .Y(_10036_) );
NAND3X1 NAND3X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_9140_), .C(_4692_), .Y(_10037_) );
OAI21X1 OAI21X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_5231_), .B(_10036_), .C(_10037_), .Y(_10038_) );
NOR3X1 NOR3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_10038_), .B(_10032_), .C(_10035_), .Y(_10039_) );
NAND3X1 NAND3X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_3407_), .B(_9133_), .C(_3408_), .Y(_10040_) );
NAND3X1 NAND3X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_4924_), .B(_9097_), .C(_4926_), .Y(_10041_) );
NAND3X1 NAND3X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_9102_), .C(_5083_), .Y(_10042_) );
NAND3X1 NAND3X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_10041_), .B(_10042_), .C(_10040_), .Y(_10043_) );
AOI22X1 AOI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_38__2_), .B(_9129_), .C(_16__2_), .D(_9127_), .Y(_10044_) );
AOI22X1 AOI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_39__2_), .B(_9099_), .C(_204__2_), .D(_9104_), .Y(_10045_) );
NAND2X1 NAND2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_10044_), .B(_10045_), .Y(_10046_) );
NOR2X1 NOR2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_10043_), .B(_10046_), .Y(_10047_) );
NAND3X1 NAND3X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_10028_), .B(_10039_), .C(_10047_), .Y(_10048_) );
AOI22X1 AOI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_227__2_), .B(_9170_), .C(_30__2_), .D(_9167_), .Y(_10049_) );
AOI22X1 AOI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_209__2_), .B(_8957_), .C(_33__2_), .D(_8991_), .Y(_10050_) );
NAND2X1 NAND2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_10049_), .B(_10050_), .Y(_10051_) );
AOI22X1 AOI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_44__2_), .B(_8968_), .C(_42__2_), .D(_8963_), .Y(_10052_) );
AOI22X1 AOI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_238__2_), .B(_8893_), .C(_208__2_), .D(_8950_), .Y(_10053_) );
NAND2X1 NAND2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_10052_), .B(_10053_), .Y(_10054_) );
NOR2X1 NOR2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_10051_), .B(_10054_), .Y(_10055_) );
AOI22X1 AOI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_22__2_), .B(_9382_), .C(_3__2_), .D(_9383_), .Y(_10056_) );
NAND2X1 NAND2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_219__2_), .Y(_10057_) );
NAND2X1 NAND2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(_232__2_), .Y(_10058_) );
NAND3X1 NAND3X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_10057_), .B(_10058_), .C(_10056_), .Y(_10059_) );
AOI22X1 AOI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_255__2_), .B(_8986_), .C(_254__2_), .D(_8984_), .Y(_10060_) );
AOI22X1 AOI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_203__2_), .B(_9018_), .C(_156__2_), .D(_8973_), .Y(_10061_) );
NAND2X1 NAND2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_10060_), .B(_10061_), .Y(_10062_) );
NOR2X1 NOR2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_10059_), .B(_10062_), .Y(_10063_) );
NAND2X1 NAND2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_10055_), .B(_10063_), .Y(_10064_) );
AOI22X1 AOI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_201__2_), .B(_9124_), .C(_212__2_), .D(_9345_), .Y(_10065_) );
NAND3X1 NAND3X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_8423_), .B(_9348_), .C(_8422_), .Y(_10066_) );
NAND3X1 NAND3X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_482_), .C(_484_), .Y(_10067_) );
AND2X2 AND2X2_1565 ( .gnd(gnd), .vdd(vdd), .A(_10067_), .B(_10066_), .Y(_10068_) );
NAND2X1 NAND2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_10065_), .B(_10068_), .Y(_10069_) );
NAND3X1 NAND3X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_15129_), .B(_9208_), .C(_15130_), .Y(_10070_) );
OAI21X1 OAI21X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_15092_), .B(_9211_), .C(_10070_), .Y(_10071_) );
NAND3X1 NAND3X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_15465_), .B(_9222_), .C(_15466_), .Y(_10072_) );
NAND3X1 NAND3X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_15412_), .B(_9224_), .C(_15411_), .Y(_10073_) );
NAND2X1 NAND2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_10072_), .B(_10073_), .Y(_10074_) );
NOR2X1 NOR2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_10074_), .B(_10071_), .Y(_10075_) );
NAND3X1 NAND3X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_15243_), .B(_9217_), .C(_15244_), .Y(_10076_) );
NAND3X1 NAND3X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_15191_), .B(_9219_), .C(_15190_), .Y(_10077_) );
NAND2X1 NAND2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_10077_), .B(_10076_), .Y(_10078_) );
NAND3X1 NAND3X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_15640_), .B(_9192_), .C(_15642_), .Y(_10079_) );
NAND3X1 NAND3X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_15698_), .B(_9199_), .C(_15696_), .Y(_10080_) );
NAND2X1 NAND2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_10080_), .B(_10079_), .Y(_10081_) );
NOR2X1 NOR2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_10081_), .B(_10078_), .Y(_10082_) );
INVX4 INVX4_75 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .Y(_10083_) );
NOR3X1 NOR3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_16170_), .B(_10083_), .C(_16171_), .Y(_10084_) );
INVX4 INVX4_76 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .Y(_10085_) );
NAND3X1 NAND3X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_15294_), .B(_9205_), .C(_15298_), .Y(_10086_) );
OAI21X1 OAI21X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_15338_), .B(_10085_), .C(_10086_), .Y(_10087_) );
NAND3X1 NAND3X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_15523_), .B(_9233_), .C(_15524_), .Y(_10088_) );
NAND3X1 NAND3X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15595_), .C(_15591_), .Y(_10089_) );
NAND2X1 NAND2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_10088_), .B(_10089_), .Y(_10090_) );
NOR3X1 NOR3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_10087_), .B(_10090_), .C(_10084_), .Y(_10091_) );
NAND3X1 NAND3X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_10075_), .B(_10082_), .C(_10091_), .Y(_10092_) );
NAND3X1 NAND3X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_15850_), .B(_9120_), .C(_15852_), .Y(_10093_) );
NAND3X1 NAND3X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_15370_), .B(_9197_), .C(_15371_), .Y(_10094_) );
NAND2X1 NAND2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_9266_), .B(_198__2_), .Y(_10095_) );
AOI22X1 AOI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_137__2_), .B(_9262_), .C(_119__2_), .D(_9268_), .Y(_10096_) );
NAND2X1 NAND2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_10095_), .B(_10096_), .Y(_10097_) );
AOI22X1 AOI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_182__2_), .B(_9300_), .C(_180__2_), .D(_9248_), .Y(_10098_) );
AOI22X1 AOI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_173__2_), .B(_9275_), .C(_78__2_), .D(_9303_), .Y(_10099_) );
NAND2X1 NAND2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_10099_), .B(_10098_), .Y(_10100_) );
NAND2X1 NAND2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_1__2_), .B(_9242_), .Y(_10101_) );
NAND2X1 NAND2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_9244_), .B(_197__2_), .Y(_10102_) );
AOI22X1 AOI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_154__2_), .B(_9292_), .C(_56__2_), .D(_9250_), .Y(_10103_) );
NAND3X1 NAND3X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_10101_), .B(_10102_), .C(_10103_), .Y(_10104_) );
NOR3X1 NOR3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_10097_), .B(_10100_), .C(_10104_), .Y(_10105_) );
NAND2X1 NAND2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .B(_233__2_), .Y(_10106_) );
AOI22X1 AOI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_186__2_), .B(_9298_), .C(_49__2_), .D(_9294_), .Y(_10107_) );
AOI22X1 AOI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .B(_9274_), .C(_31__2_), .D(_9283_), .Y(_10108_) );
NAND3X1 NAND3X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_10106_), .B(_10108_), .C(_10107_), .Y(_10109_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(_9254_), .Y(_10110_) );
AOI22X1 AOI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_32__2_), .B(_10110_), .C(_50__2_), .D(_9778_), .Y(_10111_) );
AOI22X1 AOI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_101__2_), .B(_9255_), .C(_187__2_), .D(_9235_), .Y(_10112_) );
NAND3X1 NAND3X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_8192_), .B(_9286_), .C(_8193_), .Y(_10113_) );
OAI21X1 OAI21X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_6995_), .B(_9288_), .C(_10113_), .Y(_10114_) );
NAND3X1 NAND3X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_2897_), .B(_9277_), .C(_2896_), .Y(_10115_) );
OAI21X1 OAI21X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_6456_), .B(_9259_), .C(_10115_), .Y(_10116_) );
NOR2X1 NOR2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_10116_), .B(_10114_), .Y(_10117_) );
NAND3X1 NAND3X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_10111_), .B(_10112_), .C(_10117_), .Y(_10118_) );
NOR3X1 NOR3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_4767_), .B(_9312_), .C(_4766_), .Y(_10119_) );
NOR3X1 NOR3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_5357_), .B(_9325_), .C(_5359_), .Y(_10120_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .Y(_10121_) );
NOR2X1 NOR2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_10121_), .B(_7665_), .Y(_10122_) );
NOR3X1 NOR3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_10119_), .B(_10122_), .C(_10120_), .Y(_10123_) );
AOI22X1 AOI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_83__2_), .B(_9315_), .C(_251__2_), .D(_9320_), .Y(_10124_) );
AOI22X1 AOI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_217__2_), .B(_9281_), .C(_235__2_), .D(_9324_), .Y(_10125_) );
NAND3X1 NAND3X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_10124_), .B(_10125_), .C(_10123_), .Y(_10126_) );
NOR3X1 NOR3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_10109_), .B(_10118_), .C(_10126_), .Y(_10127_) );
NAND3X1 NAND3X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_10105_), .B(_10094_), .C(_10127_), .Y(_10128_) );
AOI21X1 AOI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_157__2_), .B(_9232_), .C(_10128_), .Y(_10129_) );
AOI22X1 AOI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_155__2_), .B(_9333_), .C(_172__2_), .D(_9332_), .Y(_10130_) );
NAND3X1 NAND3X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_10093_), .B(_10130_), .C(_10129_), .Y(_10131_) );
NOR3X1 NOR3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_10092_), .B(_10131_), .C(_10069_), .Y(_10132_) );
AOI22X1 AOI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(_256__2_), .B(_9113_), .C(_142__2_), .D(_9118_), .Y(_10133_) );
NAND2X1 NAND2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__2_), .Y(_10134_) );
NAND2X1 NAND2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__2_), .Y(_10135_) );
NAND3X1 NAND3X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_10134_), .B(_10135_), .C(_10133_), .Y(_10136_) );
NAND2X1 NAND2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__2_), .Y(_10137_) );
NAND3X1 NAND3X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_9339_), .C(_434_), .Y(_10138_) );
AOI22X1 AOI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(_111__2_), .B(_9342_), .C(_12__2_), .D(_9341_), .Y(_10139_) );
NAND3X1 NAND3X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_10139_), .B(_10137_), .C(_10138_), .Y(_10140_) );
NOR2X1 NOR2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_10136_), .B(_10140_), .Y(_10141_) );
AOI22X1 AOI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_40__2_), .B(_8952_), .C(_29__2_), .D(_9176_), .Y(_10142_) );
AOI22X1 AOI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(_247__2_), .B(_9165_), .C(_218__2_), .D(_9169_), .Y(_10143_) );
NAND2X1 NAND2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_10143_), .B(_10142_), .Y(_10144_) );
NAND3X1 NAND3X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16068_), .C(_16069_), .Y(_10145_) );
NAND3X1 NAND3X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16013_), .C(_16014_), .Y(_10146_) );
NAND2X1 NAND2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_10145_), .B(_10146_), .Y(_10147_) );
NAND3X1 NAND3X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8547_), .C(_8546_), .Y(_10148_) );
OAI21X1 OAI21X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_16221_), .B(_9361_), .C(_10148_), .Y(_10149_) );
NOR2X1 NOR2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_10147_), .B(_10149_), .Y(_10150_) );
NAND2X1 NAND2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_15963_), .B(_15964_), .Y(_10151_) );
NAND3X1 NAND3X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8600_), .C(_8601_), .Y(_10152_) );
OAI21X1 OAI21X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_10151_), .B(_9215_), .C(_10152_), .Y(_10153_) );
NAND3X1 NAND3X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_8655_), .B(_9371_), .C(_8654_), .Y(_10154_) );
NAND3X1 NAND3X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_297_), .C(_298_), .Y(_10155_) );
NAND2X1 NAND2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_10155_), .B(_10154_), .Y(_10156_) );
NOR2X1 NOR2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_10153_), .B(_10156_), .Y(_10157_) );
AOI22X1 AOI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_248__2_), .B(_8901_), .C(_177__2_), .D(_8961_), .Y(_10158_) );
NAND3X1 NAND3X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_10150_), .B(_10157_), .C(_10158_), .Y(_10159_) );
NOR2X1 NOR2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_10144_), .B(_10159_), .Y(_10160_) );
NAND3X1 NAND3X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_10132_), .B(_10141_), .C(_10160_), .Y(_10161_) );
NOR3X1 NOR3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_10048_), .B(_10064_), .C(_10161_), .Y(_10162_) );
NAND3X1 NAND3X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_9982_), .B(_10021_), .C(_10162_), .Y(_10163_) );
NAND3X1 NAND3X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1532_), .C(_1534_), .Y(_10164_) );
NAND3X1 NAND3X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1617_), .C(_1619_), .Y(_10165_) );
NAND2X1 NAND2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_10164_), .B(_10165_), .Y(_10166_) );
NOR3X1 NOR3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_9944_), .B(_10166_), .C(_10163_), .Y(_10167_) );
NAND3X1 NAND3X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_9920_), .B(_9927_), .C(_10167_), .Y(_10168_) );
NAND2X1 NAND2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__2_), .Y(_10169_) );
AOI22X1 AOI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_115__2_), .B(_9399_), .C(_116__2_), .D(_9401_), .Y(_10170_) );
AOI22X1 AOI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_108__2_), .B(_9404_), .C(_109__2_), .D(_9406_), .Y(_10171_) );
NAND2X1 NAND2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_10170_), .B(_10171_), .Y(_10172_) );
NAND2X1 NAND2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_125__2_), .Y(_10173_) );
NAND2X1 NAND2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_122__2_), .Y(_10174_) );
NAND2X1 NAND2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_10173_), .B(_10174_), .Y(_10175_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(_9413_), .Y(_10176_) );
NOR2X1 NOR2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_1089_), .Y(_10177_) );
AND2X2 AND2X2_1566 ( .gnd(gnd), .vdd(vdd), .A(_120__2_), .B(_9415_), .Y(_10178_) );
NOR3X1 NOR3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_10177_), .B(_10178_), .C(_10175_), .Y(_10179_) );
AOI22X1 AOI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_132__2_), .B(_9420_), .C(_131__2_), .D(_9418_), .Y(_10180_) );
NAND2X1 NAND2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__2_), .Y(_10181_) );
NAND2X1 NAND2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__2_), .Y(_10182_) );
NAND3X1 NAND3X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_10181_), .B(_10182_), .C(_10180_), .Y(_10183_) );
NAND3X1 NAND3X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_9431_), .C(_527_), .Y(_10184_) );
NAND2X1 NAND2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__2_), .Y(_10185_) );
NAND2X1 NAND2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__2_), .Y(_10186_) );
NAND3X1 NAND3X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_10186_), .B(_10184_), .C(_10185_), .Y(_10187_) );
AOI21X1 AOI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__2_), .C(_10187_), .Y(_10188_) );
NAND2X1 NAND2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__2_), .Y(_10189_) );
NAND2X1 NAND2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_136__2_), .Y(_10190_) );
NAND3X1 NAND3X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_10189_), .B(_10190_), .C(_10188_), .Y(_10191_) );
NAND3X1 NAND3X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .B(_9410_), .C(_1001_), .Y(_10192_) );
NAND2X1 NAND2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__2_), .Y(_10193_) );
AOI22X1 AOI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_130__2_), .B(_9449_), .C(_127__2_), .D(_9448_), .Y(_10194_) );
NAND3X1 NAND3X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_10192_), .B(_10194_), .C(_10193_), .Y(_10195_) );
NOR3X1 NOR3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_10183_), .B(_10191_), .C(_10195_), .Y(_10196_) );
AOI22X1 AOI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(_110__2_), .B(_9453_), .C(_114__2_), .D(_9454_), .Y(_10197_) );
NAND3X1 NAND3X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_10179_), .B(_10197_), .C(_10196_), .Y(_10198_) );
NOR2X1 NOR2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_10172_), .B(_10198_), .Y(_10199_) );
AOI22X1 AOI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(_102__2_), .B(_9459_), .C(_103__2_), .D(_9457_), .Y(_10200_) );
NAND3X1 NAND3X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_10169_), .B(_10200_), .C(_10199_), .Y(_10201_) );
NOR3X1 NOR3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_9919_), .B(_10201_), .C(_10168_), .Y(_10202_) );
NAND3X1 NAND3X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_9909_), .B(_9916_), .C(_10202_), .Y(_10203_) );
NOR3X1 NOR3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_9898_), .B(_9901_), .C(_10203_), .Y(_10204_) );
NAND3X1 NAND3X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_9890_), .B(_9895_), .C(_10204_), .Y(_10205_) );
NAND3X1 NAND3X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_3046_), .B(_9473_), .C(_3047_), .Y(_10206_) );
NAND2X1 NAND2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__2_), .Y(_10207_) );
NAND3X1 NAND3X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_9468_), .C(_2427_), .Y(_10208_) );
NAND2X1 NAND2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__2_), .Y(_10209_) );
NAND2X1 NAND2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__2_), .Y(_10210_) );
NAND3X1 NAND3X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_10208_), .B(_10210_), .C(_10209_), .Y(_10211_) );
AOI21X1 AOI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_68__2_), .B(_9477_), .C(_10211_), .Y(_10212_) );
NAND3X1 NAND3X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_10206_), .B(_10212_), .C(_10207_), .Y(_10213_) );
NOR3X1 NOR3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_9889_), .B(_10213_), .C(_10205_), .Y(_10214_) );
AOI21X1 AOI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_9882_), .B(_10214_), .C(rst), .Y(_0__2_) );
INVX1 INVX1_3868 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .Y(_10215_) );
NAND2X1 NAND2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_8762_), .B(_54__3_), .Y(_10216_) );
OAI21X1 OAI21X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_3222_), .B(_10215_), .C(_10216_), .Y(_10217_) );
NAND2X1 NAND2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__3_), .Y(_10218_) );
NAND2X1 NAND2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__3_), .Y(_10219_) );
NAND2X1 NAND2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_10219_), .B(_10218_), .Y(_10220_) );
NOR2X1 NOR2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_10217_), .B(_10220_), .Y(_10221_) );
NAND2X1 NAND2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__3_), .Y(_10222_) );
NAND3X1 NAND3X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_8742_), .C(_3129_), .Y(_10223_) );
NAND2X1 NAND2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_10223_), .B(_10222_), .Y(_10224_) );
NAND3X1 NAND3X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_3099_), .C(_3100_), .Y(_10225_) );
NAND2X1 NAND2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_8774_), .B(_62__3_), .Y(_10226_) );
NAND3X1 NAND3X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_9473_), .C(_3050_), .Y(_10227_) );
NAND3X1 NAND3X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_10225_), .B(_10226_), .C(_10227_), .Y(_10228_) );
NAND2X1 NAND2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__3_), .Y(_10229_) );
INVX1 INVX1_3869 ( .gnd(gnd), .vdd(vdd), .A(_84__3_), .Y(_10230_) );
NOR2X1 NOR2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_10230_), .Y(_10231_) );
NOR2X1 NOR2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2288_), .Y(_10232_) );
NAND2X1 NAND2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__3_), .Y(_10233_) );
NAND3X1 NAND3X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1901_), .C(_1902_), .Y(_10234_) );
NAND2X1 NAND2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_98__3_), .Y(_10235_) );
NAND3X1 NAND3X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_10234_), .B(_10233_), .C(_10235_), .Y(_10236_) );
NOR3X1 NOR3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_10231_), .B(_10236_), .C(_10232_), .Y(_10237_) );
NAND3X1 NAND3X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_2239_), .B(_8829_), .C(_2240_), .Y(_10238_) );
NAND3X1 NAND3X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_8831_), .C(_2134_), .Y(_10239_) );
NAND2X1 NAND2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_10238_), .B(_10239_), .Y(_10240_) );
NAND3X1 NAND3X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_2074_), .B(_8834_), .C(_2075_), .Y(_10241_) );
NAND3X1 NAND3X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_2185_), .B(_8836_), .C(_2186_), .Y(_10242_) );
NAND2X1 NAND2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_10241_), .B(_10242_), .Y(_10243_) );
NOR2X1 NOR2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_10243_), .B(_10240_), .Y(_10244_) );
AOI22X1 AOI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_92__3_), .B(_8843_), .C(_91__3_), .D(_8823_), .Y(_10245_) );
NAND2X1 NAND2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(_93__3_), .Y(_10246_) );
NAND2X1 NAND2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_94__3_), .Y(_10247_) );
NAND3X1 NAND3X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_10246_), .B(_10247_), .C(_10245_), .Y(_10248_) );
NAND2X1 NAND2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__3_), .Y(_10249_) );
NAND3X1 NAND3X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1576_), .C(_1577_), .Y(_10250_) );
NAND3X1 NAND3X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_8857_), .C(_1368_), .Y(_10251_) );
NAND2X1 NAND2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_10251_), .B(_10250_), .Y(_10252_) );
NAND3X1 NAND3X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1659_), .C(_1660_), .Y(_10253_) );
NAND3X1 NAND3X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_8862_), .C(_1237_), .Y(_10254_) );
NAND2X1 NAND2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_10253_), .B(_10254_), .Y(_10255_) );
OR2X2 OR2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_10255_), .B(_10252_), .Y(_10256_) );
NOR3X1 NOR3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_8867_), .C(_1205_), .Y(_10257_) );
AOI22X1 AOI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(_191__3_), .B(_8873_), .C(_192__3_), .D(_8872_), .Y(_10258_) );
AOI22X1 AOI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_195__3_), .B(_8875_), .C(_193__3_), .D(_8876_), .Y(_10259_) );
NAND2X1 NAND2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_10258_), .B(_10259_), .Y(_10260_) );
AOI22X1 AOI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(_188__3_), .B(_8879_), .C(_126__3_), .D(_8881_), .Y(_10261_) );
AOI22X1 AOI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_196__3_), .B(_8883_), .C(_194__3_), .D(_8884_), .Y(_10262_) );
NAND2X1 NAND2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_10261_), .B(_10262_), .Y(_10263_) );
NOR3X1 NOR3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_10263_), .B(_10257_), .C(_10260_), .Y(_10264_) );
NAND3X1 NAND3X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_5820_), .B(_8893_), .C(_5819_), .Y(_10265_) );
NAND3X1 NAND3X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_8898_), .C(_4579_), .Y(_10266_) );
NAND2X1 NAND2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_10265_), .B(_10266_), .Y(_10267_) );
NAND3X1 NAND3X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_5517_), .B(_8901_), .C(_5516_), .Y(_10268_) );
NAND3X1 NAND3X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_7855_), .B(_8904_), .C(_7854_), .Y(_10269_) );
NAND2X1 NAND2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_10268_), .B(_10269_), .Y(_10270_) );
NOR2X1 NOR2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_10267_), .B(_10270_), .Y(_10271_) );
NAND3X1 NAND3X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_4080_), .B(_8909_), .C(_4079_), .Y(_10272_) );
NAND3X1 NAND3X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3882_), .C(_3881_), .Y(_10273_) );
NAND2X1 NAND2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_10272_), .B(_10273_), .Y(_10274_) );
NAND3X1 NAND3X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_4621_), .B(_8914_), .C(_4620_), .Y(_10275_) );
NAND3X1 NAND3X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_6642_), .B(_8918_), .C(_6641_), .Y(_10276_) );
NAND2X1 NAND2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_10275_), .B(_10276_), .Y(_10277_) );
NOR2X1 NOR2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_10274_), .B(_10277_), .Y(_10278_) );
NAND2X1 NAND2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_10271_), .B(_10278_), .Y(_10279_) );
NAND3X1 NAND3X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_4961_), .B(_8926_), .C(_4960_), .Y(_10280_) );
NAND3X1 NAND3X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_8029_), .B(_8933_), .C(_8028_), .Y(_10281_) );
NAND2X1 NAND2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_10280_), .B(_10281_), .Y(_10282_) );
NAND3X1 NAND3X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_4483_), .B(_8931_), .C(_4482_), .Y(_10283_) );
NAND3X1 NAND3X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_7993_), .B(_9177_), .C(_7992_), .Y(_10284_) );
NAND2X1 NAND2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_10283_), .B(_10284_), .Y(_10285_) );
NOR2X1 NOR2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_10282_), .B(_10285_), .Y(_10286_) );
NAND3X1 NAND3X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_5175_), .B(_8937_), .C(_5174_), .Y(_10287_) );
NAND3X1 NAND3X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_7817_), .B(_8939_), .C(_7816_), .Y(_10288_) );
NAND2X1 NAND2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_10287_), .B(_10288_), .Y(_10289_) );
NAND3X1 NAND3X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_5137_), .B(_8942_), .C(_5136_), .Y(_10290_) );
NAND3X1 NAND3X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_4999_), .B(_8944_), .C(_4998_), .Y(_10291_) );
NAND2X1 NAND2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_10290_), .B(_10291_), .Y(_10292_) );
NOR2X1 NOR2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_10292_), .B(_10289_), .Y(_10293_) );
NAND2X1 NAND2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_10286_), .B(_10293_), .Y(_10294_) );
NOR2X1 NOR2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_10279_), .B(_10294_), .Y(_10295_) );
NAND3X1 NAND3X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_6713_), .B(_8950_), .C(_6712_), .Y(_10296_) );
NAND3X1 NAND3X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_3923_), .B(_8952_), .C(_3922_), .Y(_10297_) );
NAND2X1 NAND2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_10296_), .B(_10297_), .Y(_10298_) );
NAND3X1 NAND3X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_5892_), .B(_8955_), .C(_5891_), .Y(_10299_) );
NAND3X1 NAND3X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_6681_), .B(_8957_), .C(_6680_), .Y(_10300_) );
NAND2X1 NAND2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_10299_), .B(_10300_), .Y(_10301_) );
NOR2X1 NOR2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_10301_), .B(_10298_), .Y(_10302_) );
NAND3X1 NAND3X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_7783_), .B(_8961_), .C(_7782_), .Y(_10303_) );
NAND3X1 NAND3X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_3844_), .B(_8963_), .C(_3843_), .Y(_10304_) );
NAND2X1 NAND2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_10303_), .B(_10304_), .Y(_10305_) );
NAND3X1 NAND3X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_5858_), .B(_8966_), .C(_5857_), .Y(_10306_) );
NAND3X1 NAND3X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_3764_), .B(_8968_), .C(_3763_), .Y(_10307_) );
NAND2X1 NAND2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_10306_), .B(_10307_), .Y(_10308_) );
NOR2X1 NOR2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_10305_), .B(_10308_), .Y(_10309_) );
NAND2X1 NAND2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_10302_), .B(_10309_), .Y(_10310_) );
NAND3X1 NAND3X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_5272_), .B(_8986_), .C(_5271_), .Y(_10311_) );
NAND3X1 NAND3X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_3468_), .B(_8975_), .C(_3467_), .Y(_10312_) );
NAND2X1 NAND2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_10311_), .B(_10312_), .Y(_10313_) );
NAND3X1 NAND3X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_4043_), .B(_8978_), .C(_4042_), .Y(_10314_) );
NAND3X1 NAND3X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_4117_), .B(_8980_), .C(_4116_), .Y(_10315_) );
NAND2X1 NAND2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_10315_), .B(_10314_), .Y(_10316_) );
NOR2X1 NOR2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_10313_), .B(_10316_), .Y(_10317_) );
NAND3X1 NAND3X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_5307_), .B(_8984_), .C(_5306_), .Y(_10318_) );
NAND3X1 NAND3X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_4153_), .B(_8991_), .C(_4152_), .Y(_10319_) );
NAND2X1 NAND2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_10318_), .B(_10319_), .Y(_10320_) );
NAND3X1 NAND3X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_7965_), .B(_8973_), .C(_7964_), .Y(_10321_) );
NAND3X1 NAND3X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_6887_), .B(_9018_), .C(_6886_), .Y(_10322_) );
NAND2X1 NAND2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_10321_), .B(_10322_), .Y(_10323_) );
NOR2X1 NOR2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_10320_), .B(_10323_), .Y(_10324_) );
NAND2X1 NAND2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_10317_), .B(_10324_), .Y(_10325_) );
NOR2X1 NOR2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_10310_), .B(_10325_), .Y(_10326_) );
NAND2X1 NAND2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_10295_), .B(_10326_), .Y(_10327_) );
NAND3X1 NAND3X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_8998_), .C(_4891_), .Y(_10328_) );
NAND3X1 NAND3X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_6499_), .B(_9002_), .C(_6498_), .Y(_10329_) );
NAND2X1 NAND2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_10328_), .B(_10329_), .Y(_10330_) );
NAND3X1 NAND3X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_5705_), .B(_9005_), .C(_5704_), .Y(_10331_) );
NAND3X1 NAND3X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_4853_), .B(_9007_), .C(_4852_), .Y(_10332_) );
NAND2X1 NAND2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_10331_), .B(_10332_), .Y(_10333_) );
NOR2X1 NOR2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_10330_), .B(_10333_), .Y(_10334_) );
NAND3X1 NAND3X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_5743_), .B(_9011_), .C(_5742_), .Y(_10335_) );
NAND3X1 NAND3X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_6785_), .B(_9013_), .C(_6784_), .Y(_10336_) );
NAND2X1 NAND2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_10335_), .B(_10336_), .Y(_10337_) );
NAND3X1 NAND3X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_6746_), .B(_9016_), .C(_6745_), .Y(_10338_) );
NAND3X1 NAND3X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_6532_), .B(_9174_), .C(_6531_), .Y(_10339_) );
NAND2X1 NAND2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_10338_), .B(_10339_), .Y(_10340_) );
NOR2X1 NOR2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_10340_), .B(_10337_), .Y(_10341_) );
NAND2X1 NAND2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_10334_), .B(_10341_), .Y(_10342_) );
NAND3X1 NAND3X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_6269_), .B(_9024_), .C(_6268_), .Y(_10343_) );
NAND3X1 NAND3X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_6341_), .B(_9026_), .C(_6340_), .Y(_10344_) );
NAND2X1 NAND2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_10343_), .B(_10344_), .Y(_10345_) );
NAND3X1 NAND3X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_6046_), .B(_9029_), .C(_6045_), .Y(_10346_) );
NAND3X1 NAND3X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_6104_), .B(_9031_), .C(_6103_), .Y(_10347_) );
NAND2X1 NAND2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_10346_), .B(_10347_), .Y(_10348_) );
NOR2X1 NOR2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_10345_), .B(_10348_), .Y(_10349_) );
NAND3X1 NAND3X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_5664_), .B(_9035_), .C(_5663_), .Y(_10350_) );
NAND3X1 NAND3X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_4660_), .B(_9037_), .C(_4659_), .Y(_10351_) );
NAND2X1 NAND2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_10351_), .B(_10350_), .Y(_10352_) );
NAND3X1 NAND3X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_6305_), .B(_9040_), .C(_6304_), .Y(_10353_) );
NAND3X1 NAND3X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_4322_), .B(_9042_), .C(_4321_), .Y(_10354_) );
NAND2X1 NAND2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_10353_), .B(_10354_), .Y(_10355_) );
NOR2X1 NOR2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_10355_), .B(_10352_), .Y(_10356_) );
NAND2X1 NAND2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_10349_), .B(_10356_), .Y(_10357_) );
NOR2X1 NOR2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_10342_), .B(_10357_), .Y(_10358_) );
NAND3X1 NAND3X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_6193_), .B(_9048_), .C(_6192_), .Y(_10359_) );
NAND3X1 NAND3X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_7928_), .B(_9050_), .C(_7927_), .Y(_10360_) );
NAND2X1 NAND2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_10359_), .B(_10360_), .Y(_10361_) );
NAND3X1 NAND3X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_5477_), .B(_9053_), .C(_5476_), .Y(_10362_) );
NAND3X1 NAND3X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_7891_), .B(_9055_), .C(_7890_), .Y(_10363_) );
NAND2X1 NAND2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_10362_), .B(_10363_), .Y(_10364_) );
NOR2X1 NOR2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_10361_), .B(_10364_), .Y(_10365_) );
NAND3X1 NAND3X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_4443_), .B(_9059_), .C(_4442_), .Y(_10366_) );
NAND3X1 NAND3X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_4403_), .B(_9061_), .C(_4402_), .Y(_10367_) );
NAND2X1 NAND2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_10366_), .B(_10367_), .Y(_10368_) );
NAND3X1 NAND3X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_6231_), .B(_9064_), .C(_6230_), .Y(_10369_) );
NAND3X1 NAND3X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_4363_), .B(_9066_), .C(_4362_), .Y(_10370_) );
NAND2X1 NAND2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_10369_), .B(_10370_), .Y(_10371_) );
NOR2X1 NOR2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_10371_), .B(_10368_), .Y(_10372_) );
NAND2X1 NAND2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_10365_), .B(_10372_), .Y(_10373_) );
NAND3X1 NAND3X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_7587_), .B(_9071_), .C(_7586_), .Y(_10374_) );
NAND3X1 NAND3X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_7551_), .B(_9073_), .C(_7550_), .Y(_10375_) );
NAND2X1 NAND2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_10374_), .B(_10375_), .Y(_10376_) );
NAND3X1 NAND3X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_5781_), .B(_9076_), .C(_5780_), .Y(_10377_) );
NAND3X1 NAND3X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_3507_), .B(_9078_), .C(_3506_), .Y(_10378_) );
NAND2X1 NAND2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_10377_), .B(_10378_), .Y(_10379_) );
NOR2X1 NOR2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_10376_), .B(_10379_), .Y(_10380_) );
NAND3X1 NAND3X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_5436_), .B(_9082_), .C(_5435_), .Y(_10381_) );
NAND3X1 NAND3X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_3803_), .B(_9084_), .C(_3802_), .Y(_10382_) );
NAND2X1 NAND2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_10382_), .B(_10381_), .Y(_10383_) );
NAND3X1 NAND3X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_6602_), .B(_9087_), .C(_6601_), .Y(_10384_) );
NAND3X1 NAND3X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_3656_), .B(_9089_), .C(_3655_), .Y(_10385_) );
NAND2X1 NAND2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_10384_), .B(_10385_), .Y(_10386_) );
NOR2X1 NOR2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_10383_), .B(_10386_), .Y(_10387_) );
NAND2X1 NAND2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_10380_), .B(_10387_), .Y(_10388_) );
NOR2X1 NOR2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_10373_), .B(_10388_), .Y(_10389_) );
NAND2X1 NAND2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_10358_), .B(_10389_), .Y(_10390_) );
NOR2X1 NOR2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_10327_), .B(_10390_), .Y(_10391_) );
NAND3X1 NAND3X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_6849_), .B(_9104_), .C(_6848_), .Y(_10392_) );
NAND3X1 NAND3X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_3959_), .B(_9099_), .C(_3958_), .Y(_10393_) );
NAND2X1 NAND2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_10393_), .B(_10392_), .Y(_10394_) );
NAND2X1 NAND2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__3_), .Y(_10395_) );
NAND3X1 NAND3X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_5085_), .B(_9102_), .C(_5084_), .Y(_10396_) );
NAND2X1 NAND2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_10395_), .B(_10396_), .Y(_10397_) );
NOR2X1 NOR2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_10397_), .B(_10394_), .Y(_10398_) );
NAND3X1 NAND3X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_15911_), .B(_9109_), .C(_15912_), .Y(_10399_) );
NAND3X1 NAND3X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_8376_), .B(_9113_), .C(_8377_), .Y(_10400_) );
NAND3X1 NAND3X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_16120_), .B(_9115_), .C(_16119_), .Y(_10401_) );
NAND3X1 NAND3X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_10399_), .B(_10400_), .C(_10401_), .Y(_10402_) );
NAND3X1 NAND3X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_382_), .C(_383_), .Y(_10403_) );
NAND3X1 NAND3X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_15854_), .B(_9120_), .C(_15855_), .Y(_10404_) );
AND2X2 AND2X2_1567 ( .gnd(gnd), .vdd(vdd), .A(_10404_), .B(_10403_), .Y(_10405_) );
AOI22X1 AOI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_201__3_), .B(_9124_), .C(_89__3_), .D(_9123_), .Y(_10406_) );
NAND2X1 NAND2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_10405_), .B(_10406_), .Y(_10407_) );
NAND3X1 NAND3X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(_9127_), .C(_4737_), .Y(_10408_) );
NAND3X1 NAND3X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_4001_), .B(_9129_), .C(_4002_), .Y(_10409_) );
NAND2X1 NAND2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_10409_), .B(_10408_), .Y(_10410_) );
NOR3X1 NOR3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_10402_), .B(_10410_), .C(_10407_), .Y(_10411_) );
NAND3X1 NAND3X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3410_), .C(_3411_), .Y(_10412_) );
NAND3X1 NAND3X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_5036_), .B(_9135_), .C(_5037_), .Y(_10413_) );
NAND3X1 NAND3X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_6921_), .B(_9137_), .C(_6922_), .Y(_10414_) );
NAND3X1 NAND3X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_10413_), .B(_10414_), .C(_10412_), .Y(_10415_) );
AOI22X1 AOI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .B(_9140_), .C(_2__3_), .D(_9141_), .Y(_10416_) );
NAND2X1 NAND2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__3_), .Y(_10417_) );
NAND2X1 NAND2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_200__3_), .Y(_10418_) );
NAND3X1 NAND3X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_10417_), .B(_10418_), .C(_10416_), .Y(_10419_) );
NOR2X1 NOR2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_10415_), .B(_10419_), .Y(_10420_) );
NAND3X1 NAND3X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_10398_), .B(_10420_), .C(_10411_), .Y(_10421_) );
AOI22X1 AOI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(_21__3_), .B(_9150_), .C(_185__3_), .D(_9151_), .Y(_10422_) );
AOI22X1 AOI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(_243__3_), .B(_9153_), .C(_253__3_), .D(_9154_), .Y(_10423_) );
NAND2X1 NAND2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_10422_), .B(_10423_), .Y(_10424_) );
AOI22X1 AOI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(_46__3_), .B(_9158_), .C(_231__3_), .D(_9157_), .Y(_10425_) );
AOI22X1 AOI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(_47__3_), .B(_9161_), .C(_244__3_), .D(_9160_), .Y(_10426_) );
NAND2X1 NAND2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_10426_), .B(_10425_), .Y(_10427_) );
NOR2X1 NOR2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_10424_), .B(_10427_), .Y(_10428_) );
NAND2X1 NAND2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_247__3_), .Y(_10429_) );
NAND2X1 NAND2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_9167_), .B(_30__3_), .Y(_10430_) );
AOI22X1 AOI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(_218__3_), .B(_9169_), .C(_227__3_), .D(_9170_), .Y(_10431_) );
NAND3X1 NAND3X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_10429_), .B(_10430_), .C(_10431_), .Y(_10432_) );
AOI22X1 AOI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(_123__3_), .B(_8928_), .C(_213__3_), .D(_8989_), .Y(_10433_) );
AOI22X1 AOI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(_178__3_), .B(_9173_), .C(_29__3_), .D(_9176_), .Y(_10434_) );
NAND2X1 NAND2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_10433_), .B(_10434_), .Y(_10435_) );
NOR2X1 NOR2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_10435_), .B(_10432_), .Y(_10436_) );
NAND2X1 NAND2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_10428_), .B(_10436_), .Y(_10437_) );
AOI22X1 AOI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(_234__3_), .B(_9182_), .C(_34__3_), .D(_9183_), .Y(_10438_) );
NAND2X1 NAND2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__3_), .Y(_10439_) );
NAND2X1 NAND2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__3_), .Y(_10440_) );
NAND3X1 NAND3X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_10439_), .B(_10440_), .C(_10438_), .Y(_10441_) );
NAND3X1 NAND3X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_15644_), .B(_9192_), .C(_15645_), .Y(_10442_) );
OAI21X1 OAI21X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_15597_), .B(_9195_), .C(_10442_), .Y(_10443_) );
NAND2X1 NAND2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__3_), .Y(_10444_) );
NAND3X1 NAND3X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_15700_), .B(_9199_), .C(_15701_), .Y(_10445_) );
NAND2X1 NAND2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_10444_), .B(_10445_), .Y(_10446_) );
NOR2X1 NOR2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_10446_), .B(_10443_), .Y(_10447_) );
NAND2X1 NAND2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__3_), .Y(_10448_) );
OAI21X1 OAI21X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_15300_), .B(_9206_), .C(_10448_), .Y(_10449_) );
NAND2X1 NAND2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__3_), .Y(_10450_) );
OAI21X1 OAI21X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_15094_), .B(_9211_), .C(_10450_), .Y(_10451_) );
NOR2X1 NOR2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_10449_), .B(_10451_), .Y(_10452_) );
NOR3X1 NOR3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_15965_), .B(_9215_), .C(_15966_), .Y(_10453_) );
NAND3X1 NAND3X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_15246_), .B(_9217_), .C(_15247_), .Y(_10454_) );
NAND3X1 NAND3X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_15194_), .B(_9219_), .C(_15193_), .Y(_10455_) );
NAND2X1 NAND2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_10455_), .B(_10454_), .Y(_10456_) );
NAND3X1 NAND3X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_15468_), .B(_9222_), .C(_15469_), .Y(_10457_) );
NAND3X1 NAND3X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_15415_), .B(_9224_), .C(_15414_), .Y(_10458_) );
NAND2X1 NAND2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_10457_), .B(_10458_), .Y(_10459_) );
NOR3X1 NOR3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_10453_), .B(_10459_), .C(_10456_), .Y(_10460_) );
NAND3X1 NAND3X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_10452_), .B(_10460_), .C(_10447_), .Y(_10461_) );
NAND2X1 NAND2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__3_), .Y(_10462_) );
NAND3X1 NAND3X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_15526_), .B(_9233_), .C(_15527_), .Y(_10463_) );
AND2X2 AND2X2_1568 ( .gnd(gnd), .vdd(vdd), .A(_78__3_), .B(_9303_), .Y(_10464_) );
AND2X2 AND2X2_1569 ( .gnd(gnd), .vdd(vdd), .A(_56__3_), .B(_9250_), .Y(_10465_) );
AND2X2 AND2X2_1570 ( .gnd(gnd), .vdd(vdd), .A(_186__3_), .B(_9298_), .Y(_10466_) );
OR2X2 OR2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_10465_), .B(_10466_), .Y(_10467_) );
INVX4 INVX4_77 ( .gnd(gnd), .vdd(vdd), .A(_9277_), .Y(_10468_) );
NAND3X1 NAND3X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_9268_), .C(_1159_), .Y(_10469_) );
OAI21X1 OAI21X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .B(_10468_), .C(_10469_), .Y(_10470_) );
INVX4 INVX4_78 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .Y(_10471_) );
NOR2X1 NOR2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_10471_), .B(_7457_), .Y(_10472_) );
NOR3X1 NOR3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_7080_), .B(_9245_), .C(_7079_), .Y(_10473_) );
NOR3X1 NOR3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_10472_), .B(_10470_), .C(_10473_), .Y(_10474_) );
NAND2X1 NAND2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__3_), .Y(_10475_) );
NAND2X1 NAND2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__3_), .Y(_10476_) );
NAND2X1 NAND2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_10475_), .B(_10476_), .Y(_10477_) );
NAND2X1 NAND2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_1__3_), .B(_9242_), .Y(_10478_) );
OAI21X1 OAI21X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .B(_9295_), .C(_10478_), .Y(_10479_) );
NOR2X1 NOR2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_10477_), .B(_10479_), .Y(_10480_) );
NAND2X1 NAND2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_10474_), .B(_10480_), .Y(_10481_) );
NOR3X1 NOR3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_10464_), .B(_10467_), .C(_10481_), .Y(_10482_) );
NAND3X1 NAND3X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_4209_), .B(_9283_), .C(_4210_), .Y(_10483_) );
NAND3X1 NAND3X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_7703_), .B(_9248_), .C(_7704_), .Y(_10484_) );
NAND3X1 NAND3X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_9262_), .C(_602_), .Y(_10485_) );
NAND3X1 NAND3X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_10483_), .B(_10484_), .C(_10485_), .Y(_10486_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_4805_), .B(_9273_), .C(_5920_), .D(_9323_), .Y(_10487_) );
NOR2X1 NOR2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_10487_), .B(_10486_), .Y(_10488_) );
NAND2X1 NAND2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__3_), .Y(_10489_) );
NAND2X1 NAND2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_173__3_), .Y(_10490_) );
NAND2X1 NAND2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_10489_), .B(_10490_), .Y(_10491_) );
NAND3X1 NAND3X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_15797_), .B(_9292_), .C(_15798_), .Y(_10492_) );
OAI21X1 OAI21X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_7621_), .B(_9301_), .C(_10492_), .Y(_10493_) );
NOR2X1 NOR2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_10493_), .B(_10491_), .Y(_10494_) );
NAND3X1 NAND3X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_7034_), .B(_9266_), .C(_7035_), .Y(_10495_) );
OAI21X1 OAI21X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_3541_), .B(_9306_), .C(_10495_), .Y(_10496_) );
NAND2X1 NAND2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_101__3_), .Y(_10497_) );
OAI21X1 OAI21X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .B(_9254_), .C(_10497_), .Y(_10498_) );
NOR2X1 NOR2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_10496_), .B(_10498_), .Y(_10499_) );
NAND3X1 NAND3X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_10488_), .B(_10499_), .C(_10494_), .Y(_10500_) );
NAND2X1 NAND2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_9320_), .B(_251__3_), .Y(_10501_) );
AOI22X1 AOI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(_252__3_), .B(_9326_), .C(_181__3_), .D(_9321_), .Y(_10502_) );
INVX1 INVX1_3870 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .Y(_10503_) );
NAND3X1 NAND3X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_2345_), .B(_9315_), .C(_2346_), .Y(_10504_) );
OAI21X1 OAI21X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_5953_), .B(_10503_), .C(_10504_), .Y(_10505_) );
NAND3X1 NAND3X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_4769_), .B(_9313_), .C(_4770_), .Y(_10506_) );
OAI21X1 OAI21X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_6417_), .B(_9763_), .C(_10506_), .Y(_10507_) );
NOR2X1 NOR2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_10507_), .B(_10505_), .Y(_10508_) );
NAND3X1 NAND3X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_10501_), .B(_10502_), .C(_10508_), .Y(_10509_) );
NOR2X1 NOR2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_10509_), .B(_10500_), .Y(_10510_) );
NAND3X1 NAND3X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_10463_), .B(_10482_), .C(_10510_), .Y(_10511_) );
AOI21X1 AOI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_157__3_), .B(_9232_), .C(_10511_), .Y(_10512_) );
AOI22X1 AOI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(_155__3_), .B(_9333_), .C(_172__3_), .D(_9332_), .Y(_10513_) );
NAND3X1 NAND3X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_10513_), .B(_10512_), .C(_10462_), .Y(_10514_) );
NOR3X1 NOR3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_10441_), .B(_10514_), .C(_10461_), .Y(_10515_) );
NAND2X1 NAND2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__3_), .Y(_10516_) );
NAND3X1 NAND3X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_9339_), .C(_437_), .Y(_10517_) );
AOI22X1 AOI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(_111__3_), .B(_9342_), .C(_12__3_), .D(_9341_), .Y(_10518_) );
NAND3X1 NAND3X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_10518_), .B(_10516_), .C(_10517_), .Y(_10519_) );
AOI22X1 AOI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(_100__3_), .B(_9346_), .C(_212__3_), .D(_9345_), .Y(_10520_) );
AOI22X1 AOI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(_245__3_), .B(_9348_), .C(_140__3_), .D(_9349_), .Y(_10521_) );
NAND2X1 NAND2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_10521_), .B(_10520_), .Y(_10522_) );
NOR2X1 NOR2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_10519_), .B(_10522_), .Y(_10523_) );
AOI22X1 AOI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(_232__3_), .B(_9354_), .C(_219__3_), .D(_9353_), .Y(_10524_) );
AOI22X1 AOI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(_246__3_), .B(_9356_), .C(_226__3_), .D(_9357_), .Y(_10525_) );
NAND2X1 NAND2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_10525_), .B(_10524_), .Y(_10526_) );
NAND3X1 NAND3X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16173_), .C(_16174_), .Y(_10527_) );
OAI21X1 OAI21X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_16224_), .B(_9361_), .C(_10527_), .Y(_10528_) );
NAND3X1 NAND3X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16071_), .C(_16072_), .Y(_10529_) );
NAND3X1 NAND3X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16016_), .C(_16017_), .Y(_10530_) );
NAND2X1 NAND2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_10529_), .B(_10530_), .Y(_10531_) );
NOR2X1 NOR2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_10531_), .B(_10528_), .Y(_10532_) );
NAND3X1 NAND3X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_8658_), .B(_9371_), .C(_8657_), .Y(_10533_) );
NAND3X1 NAND3X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8550_), .C(_8549_), .Y(_10534_) );
NAND2X1 NAND2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_10534_), .B(_10533_), .Y(_10535_) );
NAND3X1 NAND3X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8603_), .C(_8604_), .Y(_10536_) );
NAND3X1 NAND3X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_300_), .C(_301_), .Y(_10537_) );
NAND2X1 NAND2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_10536_), .B(_10537_), .Y(_10538_) );
NOR2X1 NOR2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_10538_), .B(_10535_), .Y(_10539_) );
AOI22X1 AOI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(_22__3_), .B(_9382_), .C(_3__3_), .D(_9383_), .Y(_10540_) );
NAND3X1 NAND3X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_10532_), .B(_10539_), .C(_10540_), .Y(_10541_) );
NOR2X1 NOR2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_10541_), .B(_10526_), .Y(_10542_) );
NAND3X1 NAND3X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_10523_), .B(_10515_), .C(_10542_), .Y(_10543_) );
NOR3X1 NOR3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_10421_), .B(_10437_), .C(_10543_), .Y(_10544_) );
NAND3X1 NAND3X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_10264_), .B(_10544_), .C(_10391_), .Y(_10545_) );
NAND2X1 NAND2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__3_), .Y(_10546_) );
NAND2X1 NAND2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__3_), .Y(_10547_) );
NAND2X1 NAND2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_10546_), .B(_10547_), .Y(_10548_) );
NOR3X1 NOR3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_10256_), .B(_10548_), .C(_10545_), .Y(_10549_) );
NOR3X1 NOR3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1846_), .B(_9397_), .C(_1847_), .Y(_10550_) );
NAND3X1 NAND3X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_1319_), .C(_1318_), .Y(_10551_) );
NAND3X1 NAND3X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1281_), .C(_1280_), .Y(_10552_) );
NAND2X1 NAND2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_10551_), .B(_10552_), .Y(_10553_) );
NAND3X1 NAND3X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1498_), .C(_1497_), .Y(_10554_) );
NAND3X1 NAND3X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1448_), .C(_1447_), .Y(_10555_) );
NAND2X1 NAND2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_10554_), .B(_10555_), .Y(_10556_) );
NOR2X1 NOR2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_10556_), .B(_10553_), .Y(_10557_) );
AOI22X1 AOI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(_125__3_), .B(_9411_), .C(_124__3_), .D(_9410_), .Y(_10558_) );
NAND3X1 NAND3X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_9413_), .C(_1091_), .Y(_10559_) );
NAND2X1 NAND2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__3_), .Y(_10560_) );
NAND3X1 NAND3X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_10559_), .B(_10560_), .C(_10558_), .Y(_10561_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_9421_), .C(_804_), .D(_9419_), .Y(_10562_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_9426_), .C(_689_), .D(_9424_), .Y(_10563_) );
NOR2X1 NOR2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_10562_), .B(_10563_), .Y(_10564_) );
NAND3X1 NAND3X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_651_), .C(_652_), .Y(_10565_) );
NAND3X1 NAND3X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_9431_), .C(_530_), .Y(_10566_) );
AOI22X1 AOI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(_138__3_), .B(_9434_), .C(_229__3_), .D(_9433_), .Y(_10567_) );
NAND3X1 NAND3X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_10565_), .B(_10566_), .C(_10567_), .Y(_10568_) );
NAND3X1 NAND3X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7404_), .C(_7405_), .Y(_10569_) );
OAI21X1 OAI21X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_9440_), .C(_10569_), .Y(_10570_) );
NOR2X1 NOR2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_10570_), .B(_10568_), .Y(_10571_) );
NAND2X1 NAND2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_10571_), .B(_10564_), .Y(_10572_) );
NAND3X1 NAND3X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_9444_), .C(_1047_), .Y(_10573_) );
NAND2X1 NAND2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__3_), .Y(_10574_) );
AOI22X1 AOI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(_130__3_), .B(_9449_), .C(_127__3_), .D(_9448_), .Y(_10575_) );
NAND3X1 NAND3X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_10573_), .B(_10574_), .C(_10575_), .Y(_10576_) );
NOR3X1 NOR3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_10576_), .B(_10561_), .C(_10572_), .Y(_10577_) );
AOI22X1 AOI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(_114__3_), .B(_9454_), .C(_110__3_), .D(_9453_), .Y(_10578_) );
NAND3X1 NAND3X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_10557_), .B(_10578_), .C(_10577_), .Y(_10579_) );
NAND3X1 NAND3X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(_9457_), .C(_1702_), .Y(_10580_) );
NAND2X1 NAND2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__3_), .Y(_10581_) );
NAND2X1 NAND2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_10581_), .B(_10580_), .Y(_10582_) );
NOR3X1 NOR3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_10582_), .B(_10550_), .C(_10579_), .Y(_10583_) );
NAND3X1 NAND3X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_10249_), .B(_10583_), .C(_10549_), .Y(_10584_) );
NOR2X1 NOR2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_10248_), .B(_10584_), .Y(_10585_) );
NAND3X1 NAND3X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_10237_), .B(_10244_), .C(_10585_), .Y(_10586_) );
NAND2X1 NAND2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__3_), .Y(_10587_) );
NAND2X1 NAND2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__3_), .Y(_10588_) );
AOI22X1 AOI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(_79__3_), .B(_9466_), .C(_80__3_), .D(_8805_), .Y(_10589_) );
NAND3X1 NAND3X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_10587_), .B(_10589_), .C(_10588_), .Y(_10590_) );
NAND3X1 NAND3X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_2632_), .B(_8794_), .C(_2633_), .Y(_10591_) );
NAND3X1 NAND3X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_8806_), .C(_2393_), .Y(_10592_) );
NAND2X1 NAND2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_10592_), .B(_10591_), .Y(_10593_) );
NOR3X1 NOR3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_10590_), .B(_10593_), .C(_10586_), .Y(_10594_) );
INVX1 INVX1_3871 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .Y(_10595_) );
NOR3X1 NOR3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2943_), .B(_10595_), .C(_2939_), .Y(_10596_) );
NAND3X1 NAND3X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_9477_), .C(_2852_), .Y(_10597_) );
AOI22X1 AOI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(_74__3_), .B(_8803_), .C(_73__3_), .D(_9480_), .Y(_10598_) );
AOI22X1 AOI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(_75__3_), .B(_8802_), .C(_81__3_), .D(_9468_), .Y(_10599_) );
NAND3X1 NAND3X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_10597_), .B(_10598_), .C(_10599_), .Y(_10600_) );
NAND3X1 NAND3X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .B(_8798_), .C(_2749_), .Y(_10601_) );
NAND3X1 NAND3X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .B(_8791_), .C(_2693_), .Y(_10602_) );
NAND3X1 NAND3X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_2802_), .B(_8786_), .C(_2804_), .Y(_10603_) );
NAND3X1 NAND3X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_10601_), .B(_10602_), .C(_10603_), .Y(_10604_) );
NOR3X1 NOR3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_10596_), .B(_10604_), .C(_10600_), .Y(_10605_) );
NAND3X1 NAND3X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_10229_), .B(_10605_), .C(_10594_), .Y(_10606_) );
NOR3X1 NOR3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_10224_), .B(_10228_), .C(_10606_), .Y(_10607_) );
AOI21X1 AOI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_10221_), .B(_10607_), .C(rst), .Y(_0__3_) );
NAND2X1 NAND2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__4_), .Y(_10608_) );
NAND2X1 NAND2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__4_), .Y(_10609_) );
NAND2X1 NAND2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_10608_), .B(_10609_), .Y(_10610_) );
NAND2X1 NAND2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_55__4_), .Y(_10611_) );
NAND2X1 NAND2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__4_), .Y(_10612_) );
NAND2X1 NAND2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_10612_), .B(_10611_), .Y(_10613_) );
NOR2X1 NOR2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_10613_), .B(_10610_), .Y(_10614_) );
NAND3X1 NAND3X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .B(_8750_), .C(_3154_), .Y(_10615_) );
NAND3X1 NAND3X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(_8757_), .C(_3102_), .Y(_10616_) );
NAND2X1 NAND2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_10615_), .B(_10616_), .Y(_10617_) );
NAND3X1 NAND3X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_8762_), .C(_3268_), .Y(_10618_) );
NAND3X1 NAND3X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_8774_), .C(_2997_), .Y(_10619_) );
NAND2X1 NAND2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_10618_), .B(_10619_), .Y(_10620_) );
OR2X2 OR2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_10617_), .B(_10620_), .Y(_10621_) );
NAND2X1 NAND2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__4_), .Y(_10622_) );
NAND3X1 NAND3X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_2806_), .B(_8786_), .C(_2807_), .Y(_10623_) );
OAI21X1 OAI21X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .B(_8792_), .C(_10623_), .Y(_10624_) );
NAND3X1 NAND3X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_8794_), .C(_2636_), .Y(_10625_) );
OAI21X1 OAI21X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_8799_), .C(_10625_), .Y(_10626_) );
NOR2X1 NOR2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_10626_), .B(_10624_), .Y(_10627_) );
AOI22X1 AOI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(_76__4_), .B(_9482_), .C(_77__4_), .D(_9478_), .Y(_10628_) );
NAND2X1 NAND2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__4_), .Y(_10629_) );
NAND2X1 NAND2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_82__4_), .Y(_10630_) );
NAND3X1 NAND3X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_10629_), .B(_10630_), .C(_10628_), .Y(_10631_) );
NAND2X1 NAND2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__4_), .Y(_10632_) );
NAND3X1 NAND3X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(_8803_), .C(_2579_), .Y(_10633_) );
NAND2X1 NAND2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_10633_), .B(_10632_), .Y(_10634_) );
INVX1 INVX1_3872 ( .gnd(gnd), .vdd(vdd), .A(_84__4_), .Y(_10635_) );
NOR2X1 NOR2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_10635_), .Y(_10636_) );
NOR2X1 NOR2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2290_), .Y(_10637_) );
NAND2X1 NAND2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__4_), .Y(_10638_) );
NAND3X1 NAND3X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_2001_), .B(_8843_), .C(_2002_), .Y(_10639_) );
NAND3X1 NAND3X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1904_), .C(_1905_), .Y(_10640_) );
NAND3X1 NAND3X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_10640_), .B(_10639_), .C(_10638_), .Y(_10641_) );
NOR3X1 NOR3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_10636_), .B(_10641_), .C(_10637_), .Y(_10642_) );
NAND3X1 NAND3X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_2242_), .B(_8829_), .C(_2243_), .Y(_10643_) );
NAND3X1 NAND3X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_2136_), .B(_8831_), .C(_2137_), .Y(_10644_) );
NAND2X1 NAND2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_10643_), .B(_10644_), .Y(_10645_) );
NAND3X1 NAND3X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_2077_), .B(_8834_), .C(_2078_), .Y(_10646_) );
NAND3X1 NAND3X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .B(_8836_), .C(_2189_), .Y(_10647_) );
NAND2X1 NAND2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_10646_), .B(_10647_), .Y(_10648_) );
NOR2X1 NOR2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_10648_), .B(_10645_), .Y(_10649_) );
AOI22X1 AOI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(_98__4_), .B(_8845_), .C(_93__4_), .D(_8840_), .Y(_10650_) );
NAND2X1 NAND2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_91__4_), .Y(_10651_) );
NAND2X1 NAND2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_94__4_), .Y(_10652_) );
NAND3X1 NAND3X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_10651_), .B(_10652_), .C(_10650_), .Y(_10653_) );
NAND2X1 NAND2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__4_), .Y(_10654_) );
NAND3X1 NAND3X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1537_), .C(_1538_), .Y(_10655_) );
NAND3X1 NAND3X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1622_), .C(_1623_), .Y(_10656_) );
NAND2X1 NAND2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_10655_), .B(_10656_), .Y(_10657_) );
NAND3X1 NAND3X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1662_), .C(_1663_), .Y(_10658_) );
NAND3X1 NAND3X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_8857_), .C(_1371_), .Y(_10659_) );
NAND2X1 NAND2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_10659_), .B(_10658_), .Y(_10660_) );
OR2X2 OR2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_10657_), .B(_10660_), .Y(_10661_) );
NOR3X1 NOR3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_8867_), .C(_1207_), .Y(_10662_) );
AOI22X1 AOI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(_191__4_), .B(_8873_), .C(_192__4_), .D(_8872_), .Y(_10663_) );
AOI22X1 AOI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(_195__4_), .B(_8875_), .C(_193__4_), .D(_8876_), .Y(_10664_) );
NAND2X1 NAND2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_10663_), .B(_10664_), .Y(_10665_) );
AOI22X1 AOI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(_188__4_), .B(_8879_), .C(_126__4_), .D(_8881_), .Y(_10666_) );
AOI22X1 AOI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(_196__4_), .B(_8883_), .C(_194__4_), .D(_8884_), .Y(_10667_) );
NAND2X1 NAND2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_10666_), .B(_10667_), .Y(_10668_) );
NOR3X1 NOR3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_10668_), .B(_10662_), .C(_10665_), .Y(_10669_) );
NAND3X1 NAND3X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_5823_), .B(_8893_), .C(_5822_), .Y(_10670_) );
NAND3X1 NAND3X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_4583_), .B(_8898_), .C(_4582_), .Y(_10671_) );
NAND2X1 NAND2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_10670_), .B(_10671_), .Y(_10672_) );
NAND3X1 NAND3X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_5520_), .B(_8901_), .C(_5519_), .Y(_10673_) );
NAND3X1 NAND3X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_7858_), .B(_8904_), .C(_7857_), .Y(_10674_) );
NAND2X1 NAND2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_10673_), .B(_10674_), .Y(_10675_) );
NOR2X1 NOR2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_10672_), .B(_10675_), .Y(_10676_) );
NAND3X1 NAND3X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_4083_), .B(_8909_), .C(_4082_), .Y(_10677_) );
NAND3X1 NAND3X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3885_), .C(_3884_), .Y(_10678_) );
NAND2X1 NAND2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_10677_), .B(_10678_), .Y(_10679_) );
NAND3X1 NAND3X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_4624_), .B(_8914_), .C(_4623_), .Y(_10680_) );
NAND3X1 NAND3X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_6645_), .B(_8918_), .C(_6644_), .Y(_10681_) );
NAND2X1 NAND2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_10680_), .B(_10681_), .Y(_10682_) );
NOR2X1 NOR2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_10679_), .B(_10682_), .Y(_10683_) );
NAND2X1 NAND2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_10676_), .B(_10683_), .Y(_10684_) );
NAND3X1 NAND3X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_4964_), .B(_8926_), .C(_4963_), .Y(_10685_) );
NAND3X1 NAND3X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_8064_), .B(_8928_), .C(_8063_), .Y(_10686_) );
NAND2X1 NAND2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_10685_), .B(_10686_), .Y(_10687_) );
NAND3X1 NAND3X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_4486_), .B(_8931_), .C(_4485_), .Y(_10688_) );
NAND3X1 NAND3X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_8032_), .B(_8933_), .C(_8031_), .Y(_10689_) );
NAND2X1 NAND2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_10688_), .B(_10689_), .Y(_10690_) );
NOR2X1 NOR2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_10687_), .B(_10690_), .Y(_10691_) );
NAND3X1 NAND3X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_5178_), .B(_8937_), .C(_5177_), .Y(_10692_) );
NAND3X1 NAND3X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_7820_), .B(_8939_), .C(_7819_), .Y(_10693_) );
NAND2X1 NAND2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_10692_), .B(_10693_), .Y(_10694_) );
NAND3X1 NAND3X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_5140_), .B(_8942_), .C(_5139_), .Y(_10695_) );
NAND3X1 NAND3X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_5002_), .B(_8944_), .C(_5001_), .Y(_10696_) );
NAND2X1 NAND2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_10695_), .B(_10696_), .Y(_10697_) );
NOR2X1 NOR2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_10697_), .B(_10694_), .Y(_10698_) );
NAND2X1 NAND2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_10691_), .B(_10698_), .Y(_10699_) );
NOR2X1 NOR2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_10684_), .B(_10699_), .Y(_10700_) );
NAND3X1 NAND3X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_6716_), .B(_8950_), .C(_6715_), .Y(_10701_) );
NAND3X1 NAND3X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_3926_), .B(_8952_), .C(_3925_), .Y(_10702_) );
NAND2X1 NAND2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_10701_), .B(_10702_), .Y(_10703_) );
NAND3X1 NAND3X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_5895_), .B(_8955_), .C(_5894_), .Y(_10704_) );
NAND3X1 NAND3X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_6684_), .B(_8957_), .C(_6683_), .Y(_10705_) );
NAND2X1 NAND2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_10704_), .B(_10705_), .Y(_10706_) );
NOR2X1 NOR2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_10706_), .B(_10703_), .Y(_10707_) );
NAND3X1 NAND3X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_7786_), .B(_8961_), .C(_7785_), .Y(_10708_) );
NAND3X1 NAND3X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .B(_8963_), .C(_3846_), .Y(_10709_) );
NAND2X1 NAND2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_10708_), .B(_10709_), .Y(_10710_) );
NAND3X1 NAND3X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_5861_), .B(_8966_), .C(_5860_), .Y(_10711_) );
NAND3X1 NAND3X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(_8968_), .C(_3766_), .Y(_10712_) );
NAND2X1 NAND2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_10711_), .B(_10712_), .Y(_10713_) );
NOR2X1 NOR2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_10710_), .B(_10713_), .Y(_10714_) );
NAND2X1 NAND2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_10707_), .B(_10714_), .Y(_10715_) );
NAND3X1 NAND3X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_5275_), .B(_8986_), .C(_5274_), .Y(_10716_) );
NAND3X1 NAND3X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_8975_), .C(_3470_), .Y(_10717_) );
NAND2X1 NAND2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_10716_), .B(_10717_), .Y(_10718_) );
NAND3X1 NAND3X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_4046_), .B(_8978_), .C(_4045_), .Y(_10719_) );
NAND3X1 NAND3X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_4120_), .B(_8980_), .C(_4119_), .Y(_10720_) );
NAND2X1 NAND2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_10720_), .B(_10719_), .Y(_10721_) );
NOR2X1 NOR2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_10718_), .B(_10721_), .Y(_10722_) );
NAND3X1 NAND3X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_5310_), .B(_8984_), .C(_5309_), .Y(_10723_) );
NAND3X1 NAND3X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_4156_), .B(_8991_), .C(_4155_), .Y(_10724_) );
NAND2X1 NAND2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_10723_), .B(_10724_), .Y(_10725_) );
NAND3X1 NAND3X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_7968_), .B(_8973_), .C(_7967_), .Y(_10726_) );
NAND3X1 NAND3X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_6890_), .B(_9018_), .C(_6889_), .Y(_10727_) );
NAND2X1 NAND2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_10726_), .B(_10727_), .Y(_10728_) );
NOR2X1 NOR2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_10725_), .B(_10728_), .Y(_10729_) );
NAND2X1 NAND2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_10722_), .B(_10729_), .Y(_10730_) );
NOR2X1 NOR2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_10715_), .B(_10730_), .Y(_10731_) );
NAND2X1 NAND2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_10700_), .B(_10731_), .Y(_10732_) );
NAND3X1 NAND3X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_4895_), .B(_8998_), .C(_4894_), .Y(_10733_) );
NAND3X1 NAND3X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_6502_), .B(_9002_), .C(_6501_), .Y(_10734_) );
NAND2X1 NAND2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_10733_), .B(_10734_), .Y(_10735_) );
NAND3X1 NAND3X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_5708_), .B(_9005_), .C(_5707_), .Y(_10736_) );
NAND3X1 NAND3X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_4856_), .B(_9007_), .C(_4855_), .Y(_10737_) );
NAND2X1 NAND2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_10736_), .B(_10737_), .Y(_10738_) );
NOR2X1 NOR2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_10735_), .B(_10738_), .Y(_10739_) );
NAND3X1 NAND3X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_5746_), .B(_9011_), .C(_5745_), .Y(_10740_) );
NAND3X1 NAND3X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_6788_), .B(_9013_), .C(_6787_), .Y(_10741_) );
NAND2X1 NAND2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_10740_), .B(_10741_), .Y(_10742_) );
NAND3X1 NAND3X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_6749_), .B(_9016_), .C(_6748_), .Y(_10743_) );
NAND3X1 NAND3X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_6535_), .B(_9174_), .C(_6534_), .Y(_10744_) );
NAND2X1 NAND2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_10743_), .B(_10744_), .Y(_10745_) );
NOR2X1 NOR2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_10745_), .B(_10742_), .Y(_10746_) );
NAND2X1 NAND2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_10739_), .B(_10746_), .Y(_10747_) );
NAND3X1 NAND3X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_6272_), .B(_9024_), .C(_6271_), .Y(_10748_) );
NAND3X1 NAND3X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_6344_), .B(_9026_), .C(_6343_), .Y(_10749_) );
NAND2X1 NAND2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_10748_), .B(_10749_), .Y(_10750_) );
NAND3X1 NAND3X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_6049_), .B(_9029_), .C(_6048_), .Y(_10751_) );
NAND3X1 NAND3X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_6107_), .B(_9031_), .C(_6106_), .Y(_10752_) );
NAND2X1 NAND2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_10751_), .B(_10752_), .Y(_10753_) );
NOR2X1 NOR2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_10750_), .B(_10753_), .Y(_10754_) );
NAND3X1 NAND3X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_5667_), .B(_9035_), .C(_5666_), .Y(_10755_) );
NAND3X1 NAND3X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_4663_), .B(_9037_), .C(_4662_), .Y(_10756_) );
NAND2X1 NAND2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_10756_), .B(_10755_), .Y(_10757_) );
NAND3X1 NAND3X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_6308_), .B(_9040_), .C(_6307_), .Y(_10758_) );
NAND3X1 NAND3X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_4325_), .B(_9042_), .C(_4324_), .Y(_10759_) );
NAND2X1 NAND2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_10758_), .B(_10759_), .Y(_10760_) );
NOR2X1 NOR2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_10760_), .B(_10757_), .Y(_10761_) );
NAND2X1 NAND2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_10754_), .B(_10761_), .Y(_10762_) );
NOR2X1 NOR2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_10747_), .B(_10762_), .Y(_10763_) );
NAND3X1 NAND3X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_6196_), .B(_9048_), .C(_6195_), .Y(_10764_) );
NAND3X1 NAND3X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_7931_), .B(_9050_), .C(_7930_), .Y(_10765_) );
NAND2X1 NAND2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_10764_), .B(_10765_), .Y(_10766_) );
NAND3X1 NAND3X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_5480_), .B(_9053_), .C(_5479_), .Y(_10767_) );
NAND3X1 NAND3X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_7894_), .B(_9055_), .C(_7893_), .Y(_10768_) );
NAND2X1 NAND2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_10767_), .B(_10768_), .Y(_10769_) );
NOR2X1 NOR2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_10766_), .B(_10769_), .Y(_10770_) );
NAND3X1 NAND3X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .B(_9059_), .C(_4445_), .Y(_10771_) );
NAND3X1 NAND3X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_9061_), .C(_4405_), .Y(_10772_) );
NAND2X1 NAND2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_10771_), .B(_10772_), .Y(_10773_) );
NAND3X1 NAND3X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_6234_), .B(_9064_), .C(_6233_), .Y(_10774_) );
NAND3X1 NAND3X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_4366_), .B(_9066_), .C(_4365_), .Y(_10775_) );
NAND2X1 NAND2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_10774_), .B(_10775_), .Y(_10776_) );
NOR2X1 NOR2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_10776_), .B(_10773_), .Y(_10777_) );
NAND2X1 NAND2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_10770_), .B(_10777_), .Y(_10778_) );
NAND3X1 NAND3X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_7590_), .B(_9071_), .C(_7589_), .Y(_10779_) );
NAND3X1 NAND3X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_7554_), .B(_9073_), .C(_7553_), .Y(_10780_) );
NAND2X1 NAND2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_10779_), .B(_10780_), .Y(_10781_) );
NAND3X1 NAND3X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_5784_), .B(_9076_), .C(_5783_), .Y(_10782_) );
NAND3X1 NAND3X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_3510_), .B(_9078_), .C(_3509_), .Y(_10783_) );
NAND2X1 NAND2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_10782_), .B(_10783_), .Y(_10784_) );
NOR2X1 NOR2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_10781_), .B(_10784_), .Y(_10785_) );
NAND3X1 NAND3X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_5439_), .B(_9082_), .C(_5438_), .Y(_10786_) );
NAND3X1 NAND3X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_3806_), .B(_9084_), .C(_3805_), .Y(_10787_) );
NAND2X1 NAND2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_10787_), .B(_10786_), .Y(_10788_) );
NAND3X1 NAND3X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_6605_), .B(_9087_), .C(_6604_), .Y(_10789_) );
NAND3X1 NAND3X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_3659_), .B(_9089_), .C(_3658_), .Y(_10790_) );
NAND2X1 NAND2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_10789_), .B(_10790_), .Y(_10791_) );
NOR2X1 NOR2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_10788_), .B(_10791_), .Y(_10792_) );
NAND2X1 NAND2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_10785_), .B(_10792_), .Y(_10793_) );
NOR2X1 NOR2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_10778_), .B(_10793_), .Y(_10794_) );
NAND2X1 NAND2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_10763_), .B(_10794_), .Y(_10795_) );
NOR2X1 NOR2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_10732_), .B(_10795_), .Y(_10796_) );
NAND3X1 NAND3X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_6851_), .B(_9104_), .C(_6850_), .Y(_10797_) );
NAND3X1 NAND3X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_9099_), .C(_3960_), .Y(_10798_) );
NAND2X1 NAND2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_10798_), .B(_10797_), .Y(_10799_) );
NAND2X1 NAND2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__4_), .Y(_10800_) );
NAND3X1 NAND3X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_9102_), .C(_5086_), .Y(_10801_) );
NAND2X1 NAND2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_10800_), .B(_10801_), .Y(_10802_) );
NOR2X1 NOR2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_10802_), .B(_10799_), .Y(_10803_) );
NAND3X1 NAND3X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_15914_), .B(_9109_), .C(_15915_), .Y(_10804_) );
NAND3X1 NAND3X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_8379_), .B(_9113_), .C(_8380_), .Y(_10805_) );
NAND3X1 NAND3X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_16122_), .B(_9115_), .C(_16121_), .Y(_10806_) );
NAND3X1 NAND3X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_10804_), .B(_10805_), .C(_10806_), .Y(_10807_) );
NAND3X1 NAND3X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_385_), .C(_386_), .Y(_10808_) );
NAND3X1 NAND3X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_15857_), .B(_9120_), .C(_15858_), .Y(_10809_) );
AND2X2 AND2X2_1571 ( .gnd(gnd), .vdd(vdd), .A(_10809_), .B(_10808_), .Y(_10810_) );
AOI22X1 AOI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(_201__4_), .B(_9124_), .C(_89__4_), .D(_9123_), .Y(_10811_) );
NAND2X1 NAND2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_10810_), .B(_10811_), .Y(_10812_) );
NAND3X1 NAND3X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_4739_), .B(_9127_), .C(_4740_), .Y(_10813_) );
NAND3X1 NAND3X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_4004_), .B(_9129_), .C(_4005_), .Y(_10814_) );
NAND2X1 NAND2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_10814_), .B(_10813_), .Y(_10815_) );
NOR3X1 NOR3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_10807_), .B(_10815_), .C(_10812_), .Y(_10816_) );
NAND3X1 NAND3X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3413_), .C(_3414_), .Y(_10817_) );
NAND3X1 NAND3X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_5039_), .B(_9135_), .C(_5040_), .Y(_10818_) );
NAND3X1 NAND3X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_6924_), .B(_9137_), .C(_6925_), .Y(_10819_) );
NAND3X1 NAND3X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_10818_), .B(_10819_), .C(_10817_), .Y(_10820_) );
AOI22X1 AOI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(_17__4_), .B(_9140_), .C(_2__4_), .D(_9141_), .Y(_10821_) );
NAND2X1 NAND2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__4_), .Y(_10822_) );
NAND2X1 NAND2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_200__4_), .Y(_10823_) );
NAND3X1 NAND3X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_10822_), .B(_10823_), .C(_10821_), .Y(_10824_) );
NOR2X1 NOR2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_10820_), .B(_10824_), .Y(_10825_) );
NAND3X1 NAND3X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_10803_), .B(_10825_), .C(_10816_), .Y(_10826_) );
AOI22X1 AOI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(_21__4_), .B(_9150_), .C(_185__4_), .D(_9151_), .Y(_10827_) );
AOI22X1 AOI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(_243__4_), .B(_9153_), .C(_253__4_), .D(_9154_), .Y(_10828_) );
NAND2X1 NAND2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_10827_), .B(_10828_), .Y(_10829_) );
AOI22X1 AOI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(_46__4_), .B(_9158_), .C(_231__4_), .D(_9157_), .Y(_10830_) );
AOI22X1 AOI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(_47__4_), .B(_9161_), .C(_244__4_), .D(_9160_), .Y(_10831_) );
NAND2X1 NAND2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_10831_), .B(_10830_), .Y(_10832_) );
NOR2X1 NOR2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_10829_), .B(_10832_), .Y(_10833_) );
NAND2X1 NAND2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_247__4_), .Y(_10834_) );
NAND2X1 NAND2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_9167_), .B(_30__4_), .Y(_10835_) );
AOI22X1 AOI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(_218__4_), .B(_9169_), .C(_227__4_), .D(_9170_), .Y(_10836_) );
NAND3X1 NAND3X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_10834_), .B(_10835_), .C(_10836_), .Y(_10837_) );
AOI22X1 AOI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(_145__4_), .B(_9177_), .C(_213__4_), .D(_8989_), .Y(_10838_) );
AOI22X1 AOI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(_178__4_), .B(_9173_), .C(_29__4_), .D(_9176_), .Y(_10839_) );
NAND2X1 NAND2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_10838_), .B(_10839_), .Y(_10840_) );
NOR2X1 NOR2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_10840_), .B(_10837_), .Y(_10841_) );
NAND2X1 NAND2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_10833_), .B(_10841_), .Y(_10842_) );
AOI22X1 AOI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(_234__4_), .B(_9182_), .C(_34__4_), .D(_9183_), .Y(_10843_) );
NAND2X1 NAND2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__4_), .Y(_10844_) );
NAND2X1 NAND2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__4_), .Y(_10845_) );
NAND3X1 NAND3X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_10844_), .B(_10845_), .C(_10843_), .Y(_10846_) );
NAND3X1 NAND3X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_15647_), .B(_9192_), .C(_15648_), .Y(_10847_) );
OAI21X1 OAI21X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_15599_), .B(_9195_), .C(_10847_), .Y(_10848_) );
NAND2X1 NAND2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__4_), .Y(_10849_) );
NAND3X1 NAND3X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_15703_), .B(_9199_), .C(_15704_), .Y(_10850_) );
NAND2X1 NAND2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_10849_), .B(_10850_), .Y(_10851_) );
NOR2X1 NOR2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_10851_), .B(_10848_), .Y(_10852_) );
NAND2X1 NAND2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__4_), .Y(_10853_) );
OAI21X1 OAI21X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_15302_), .B(_9206_), .C(_10853_), .Y(_10854_) );
NAND2X1 NAND2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__4_), .Y(_10855_) );
OAI21X1 OAI21X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_15096_), .B(_9211_), .C(_10855_), .Y(_10856_) );
NOR2X1 NOR2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_10854_), .B(_10856_), .Y(_10857_) );
NOR3X1 NOR3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_15967_), .B(_9215_), .C(_15968_), .Y(_10858_) );
NAND3X1 NAND3X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_15249_), .B(_9217_), .C(_15250_), .Y(_10859_) );
NAND3X1 NAND3X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_15197_), .B(_9219_), .C(_15196_), .Y(_10860_) );
NAND2X1 NAND2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_10860_), .B(_10859_), .Y(_10861_) );
NAND3X1 NAND3X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_15471_), .B(_9222_), .C(_15472_), .Y(_10862_) );
NAND3X1 NAND3X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_15418_), .B(_9224_), .C(_15417_), .Y(_10863_) );
NAND2X1 NAND2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_10862_), .B(_10863_), .Y(_10864_) );
NOR3X1 NOR3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_10858_), .B(_10864_), .C(_10861_), .Y(_10865_) );
NAND3X1 NAND3X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_10857_), .B(_10865_), .C(_10852_), .Y(_10866_) );
NAND2X1 NAND2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__4_), .Y(_10867_) );
NAND3X1 NAND3X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_15529_), .B(_9233_), .C(_15530_), .Y(_10868_) );
AND2X2 AND2X2_1572 ( .gnd(gnd), .vdd(vdd), .A(_65__4_), .B(_9277_), .Y(_10869_) );
NOR2X1 NOR2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .B(_7624_), .Y(_10870_) );
AND2X2 AND2X2_1573 ( .gnd(gnd), .vdd(vdd), .A(_137__4_), .B(_9262_), .Y(_10871_) );
OR2X2 OR2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_10871_), .B(_10870_), .Y(_10872_) );
NAND3X1 NAND3X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_15800_), .B(_9292_), .C(_15801_), .Y(_10873_) );
OAI21X1 OAI21X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .B(_9306_), .C(_10873_), .Y(_10874_) );
INVX4 INVX4_79 ( .gnd(gnd), .vdd(vdd), .A(_9250_), .Y(_10875_) );
NAND2X1 NAND2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_1__4_), .B(_9242_), .Y(_10876_) );
OAI21X1 OAI21X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_8225_), .B(_10875_), .C(_10876_), .Y(_10877_) );
NOR2X1 NOR2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_10874_), .B(_10877_), .Y(_10878_) );
NAND2X1 NAND2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__4_), .Y(_10879_) );
OAI21X1 OAI21X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_7083_), .B(_9245_), .C(_10879_), .Y(_10880_) );
NAND2X1 NAND2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_173__4_), .Y(_10881_) );
OAI21X1 OAI21X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_4180_), .B(_9254_), .C(_10881_), .Y(_10882_) );
NOR2X1 NOR2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_10880_), .B(_10882_), .Y(_10883_) );
NAND2X1 NAND2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_10883_), .B(_10878_), .Y(_10884_) );
NOR3X1 NOR3X1_281 ( .gnd(gnd), .vdd(vdd), .A(_10869_), .B(_10872_), .C(_10884_), .Y(_10885_) );
NAND3X1 NAND3X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_5393_), .B(_9320_), .C(_5394_), .Y(_10886_) );
NAND2X1 NAND2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__4_), .Y(_10887_) );
NAND3X1 NAND3X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_3592_), .B(_9294_), .C(_3593_), .Y(_10888_) );
NAND3X1 NAND3X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_10887_), .B(_10886_), .C(_10888_), .Y(_10889_) );
NAND3X1 NAND3X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_5955_), .B(_9310_), .C(_5956_), .Y(_10890_) );
OAI21X1 OAI21X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .B(_9325_), .C(_10890_), .Y(_10891_) );
NOR2X1 NOR2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_10891_), .B(_10889_), .Y(_10892_) );
NAND3X1 NAND3X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_6998_), .B(_7000_), .C(_9289_), .Y(_10893_) );
OAI21X1 OAI21X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_7038_), .B(_9267_), .C(_10893_), .Y(_10894_) );
NOR2X1 NOR2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_10471_), .B(_7460_), .Y(_10895_) );
AND2X2 AND2X2_1574 ( .gnd(gnd), .vdd(vdd), .A(_101__4_), .B(_9255_), .Y(_10896_) );
NOR3X1 NOR3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_10896_), .B(_10895_), .C(_10894_), .Y(_10897_) );
NAND2X1 NAND2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .B(_119__4_), .Y(_10898_) );
OAI21X1 OAI21X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_7707_), .B(_9249_), .C(_10898_), .Y(_10899_) );
NAND2X1 NAND2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .B(_186__4_), .Y(_10900_) );
OAI21X1 OAI21X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_8155_), .B(_9304_), .C(_10900_), .Y(_10901_) );
NOR2X1 NOR2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_10899_), .B(_10901_), .Y(_10902_) );
NAND3X1 NAND3X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_10897_), .B(_10892_), .C(_10902_), .Y(_10903_) );
NAND2X1 NAND2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .B(_235__4_), .Y(_10904_) );
AOI22X1 AOI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(_14__4_), .B(_9274_), .C(_217__4_), .D(_9281_), .Y(_10905_) );
AND2X2 AND2X2_1575 ( .gnd(gnd), .vdd(vdd), .A(_10905_), .B(_10904_), .Y(_10906_) );
AOI22X1 AOI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(_31__4_), .B(_9283_), .C(_15__4_), .D(_9313_), .Y(_10907_) );
AOI22X1 AOI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(_181__4_), .B(_9321_), .C(_83__4_), .D(_9315_), .Y(_10908_) );
NAND3X1 NAND3X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_10907_), .B(_10908_), .C(_10906_), .Y(_10909_) );
NOR2X1 NOR2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_10903_), .B(_10909_), .Y(_10910_) );
NAND3X1 NAND3X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_10868_), .B(_10885_), .C(_10910_), .Y(_10911_) );
AOI21X1 AOI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_157__4_), .B(_9232_), .C(_10911_), .Y(_10912_) );
AOI22X1 AOI22X1_179 ( .gnd(gnd), .vdd(vdd), .A(_155__4_), .B(_9333_), .C(_172__4_), .D(_9332_), .Y(_10913_) );
NAND3X1 NAND3X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_10913_), .B(_10867_), .C(_10912_), .Y(_10914_) );
NOR3X1 NOR3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_10846_), .B(_10914_), .C(_10866_), .Y(_10915_) );
NAND2X1 NAND2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__4_), .Y(_10916_) );
NAND3X1 NAND3X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_9339_), .C(_440_), .Y(_10917_) );
AOI22X1 AOI22X1_180 ( .gnd(gnd), .vdd(vdd), .A(_111__4_), .B(_9342_), .C(_12__4_), .D(_9341_), .Y(_10918_) );
NAND3X1 NAND3X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_10918_), .B(_10916_), .C(_10917_), .Y(_10919_) );
AOI22X1 AOI22X1_181 ( .gnd(gnd), .vdd(vdd), .A(_100__4_), .B(_9346_), .C(_212__4_), .D(_9345_), .Y(_10920_) );
AOI22X1 AOI22X1_182 ( .gnd(gnd), .vdd(vdd), .A(_245__4_), .B(_9348_), .C(_140__4_), .D(_9349_), .Y(_10921_) );
NAND2X1 NAND2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_10921_), .B(_10920_), .Y(_10922_) );
NOR2X1 NOR2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_10919_), .B(_10922_), .Y(_10923_) );
AOI22X1 AOI22X1_183 ( .gnd(gnd), .vdd(vdd), .A(_232__4_), .B(_9354_), .C(_219__4_), .D(_9353_), .Y(_10924_) );
AOI22X1 AOI22X1_184 ( .gnd(gnd), .vdd(vdd), .A(_246__4_), .B(_9356_), .C(_226__4_), .D(_9357_), .Y(_10925_) );
NAND2X1 NAND2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_10925_), .B(_10924_), .Y(_10926_) );
NAND3X1 NAND3X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16176_), .C(_16177_), .Y(_10927_) );
OAI21X1 OAI21X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_16227_), .B(_9361_), .C(_10927_), .Y(_10928_) );
NAND3X1 NAND3X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16074_), .C(_16075_), .Y(_10929_) );
NAND3X1 NAND3X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16019_), .C(_16020_), .Y(_10930_) );
NAND2X1 NAND2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_10929_), .B(_10930_), .Y(_10931_) );
NOR2X1 NOR2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_10931_), .B(_10928_), .Y(_10932_) );
NAND3X1 NAND3X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_8661_), .B(_9371_), .C(_8660_), .Y(_10933_) );
NAND3X1 NAND3X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8553_), .C(_8552_), .Y(_10934_) );
NAND2X1 NAND2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_10934_), .B(_10933_), .Y(_10935_) );
NAND3X1 NAND3X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8606_), .C(_8607_), .Y(_10936_) );
NAND3X1 NAND3X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_303_), .C(_304_), .Y(_10937_) );
NAND2X1 NAND2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_10936_), .B(_10937_), .Y(_10938_) );
NOR2X1 NOR2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_10938_), .B(_10935_), .Y(_10939_) );
AOI22X1 AOI22X1_185 ( .gnd(gnd), .vdd(vdd), .A(_22__4_), .B(_9382_), .C(_3__4_), .D(_9383_), .Y(_10940_) );
NAND3X1 NAND3X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_10932_), .B(_10939_), .C(_10940_), .Y(_10941_) );
NOR2X1 NOR2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_10941_), .B(_10926_), .Y(_10942_) );
NAND3X1 NAND3X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_10923_), .B(_10915_), .C(_10942_), .Y(_10943_) );
NOR3X1 NOR3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_10826_), .B(_10842_), .C(_10943_), .Y(_10944_) );
NAND3X1 NAND3X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_10669_), .B(_10944_), .C(_10796_), .Y(_10945_) );
NAND2X1 NAND2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__4_), .Y(_10946_) );
NAND2X1 NAND2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__4_), .Y(_10947_) );
NAND2X1 NAND2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_10947_), .B(_10946_), .Y(_10948_) );
NOR3X1 NOR3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_10661_), .B(_10948_), .C(_10945_), .Y(_10949_) );
NOR3X1 NOR3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_9397_), .C(_1849_), .Y(_10950_) );
NAND3X1 NAND3X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1451_), .C(_1450_), .Y(_10951_) );
NAND3X1 NAND3X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_9453_), .B(_1405_), .C(_1404_), .Y(_10952_) );
NAND2X1 NAND2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_10951_), .B(_10952_), .Y(_10953_) );
NAND3X1 NAND3X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1501_), .C(_1500_), .Y(_10954_) );
NAND3X1 NAND3X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1284_), .C(_1283_), .Y(_10955_) );
NAND2X1 NAND2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_10954_), .B(_10955_), .Y(_10956_) );
NOR2X1 NOR2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_10956_), .B(_10953_), .Y(_10957_) );
AOI22X1 AOI22X1_186 ( .gnd(gnd), .vdd(vdd), .A(_125__4_), .B(_9411_), .C(_124__4_), .D(_9410_), .Y(_10958_) );
NAND3X1 NAND3X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_9413_), .C(_1094_), .Y(_10959_) );
NAND2X1 NAND2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__4_), .Y(_10960_) );
NAND3X1 NAND3X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_10959_), .B(_10960_), .C(_10958_), .Y(_10961_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_9421_), .C(_807_), .D(_9419_), .Y(_10962_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_9426_), .C(_692_), .D(_9424_), .Y(_10963_) );
NOR2X1 NOR2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_10962_), .B(_10963_), .Y(_10964_) );
NAND3X1 NAND3X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_654_), .C(_655_), .Y(_10965_) );
NAND3X1 NAND3X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_9431_), .C(_533_), .Y(_10966_) );
AOI22X1 AOI22X1_187 ( .gnd(gnd), .vdd(vdd), .A(_138__4_), .B(_9434_), .C(_229__4_), .D(_9433_), .Y(_10967_) );
NAND3X1 NAND3X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_10965_), .B(_10966_), .C(_10967_), .Y(_10968_) );
NAND3X1 NAND3X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7407_), .C(_7408_), .Y(_10969_) );
OAI21X1 OAI21X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_9440_), .C(_10969_), .Y(_10970_) );
NOR2X1 NOR2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_10970_), .B(_10968_), .Y(_10971_) );
NAND2X1 NAND2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_10971_), .B(_10964_), .Y(_10972_) );
NAND3X1 NAND3X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_9444_), .C(_1050_), .Y(_10973_) );
NAND2X1 NAND2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__4_), .Y(_10974_) );
AOI22X1 AOI22X1_188 ( .gnd(gnd), .vdd(vdd), .A(_130__4_), .B(_9449_), .C(_127__4_), .D(_9448_), .Y(_10975_) );
NAND3X1 NAND3X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_10973_), .B(_10974_), .C(_10975_), .Y(_10976_) );
NOR3X1 NOR3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_10976_), .B(_10961_), .C(_10972_), .Y(_10977_) );
AOI22X1 AOI22X1_189 ( .gnd(gnd), .vdd(vdd), .A(_115__4_), .B(_9399_), .C(_114__4_), .D(_9454_), .Y(_10978_) );
NAND3X1 NAND3X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_10978_), .B(_10957_), .C(_10977_), .Y(_10979_) );
NAND3X1 NAND3X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .B(_9457_), .C(_1705_), .Y(_10980_) );
NAND2X1 NAND2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__4_), .Y(_10981_) );
NAND2X1 NAND2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_10981_), .B(_10980_), .Y(_10982_) );
NOR3X1 NOR3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_10982_), .B(_10950_), .C(_10979_), .Y(_10983_) );
NAND3X1 NAND3X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_10654_), .B(_10983_), .C(_10949_), .Y(_10984_) );
NOR2X1 NOR2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_10653_), .B(_10984_), .Y(_10985_) );
NAND3X1 NAND3X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_10642_), .B(_10649_), .C(_10985_), .Y(_10986_) );
NOR3X1 NOR3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_10631_), .B(_10634_), .C(_10986_), .Y(_10987_) );
NAND3X1 NAND3X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_10622_), .B(_10627_), .C(_10987_), .Y(_10988_) );
NAND3X1 NAND3X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_3052_), .B(_9473_), .C(_3053_), .Y(_10989_) );
NAND2X1 NAND2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__4_), .Y(_10990_) );
NAND2X1 NAND2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__4_), .Y(_10991_) );
NAND2X1 NAND2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__4_), .Y(_10992_) );
NAND3X1 NAND3X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .B(_9468_), .C(_2431_), .Y(_10993_) );
NAND3X1 NAND3X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_10993_), .B(_10991_), .C(_10992_), .Y(_10994_) );
AOI21X1 AOI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_68__4_), .B(_9477_), .C(_10994_), .Y(_10995_) );
NAND3X1 NAND3X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_10995_), .B(_10989_), .C(_10990_), .Y(_10996_) );
NOR3X1 NOR3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_10621_), .B(_10996_), .C(_10988_), .Y(_10997_) );
AOI21X1 AOI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_10614_), .B(_10997_), .C(rst), .Y(_0__4_) );
NAND2X1 NAND2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__5_), .Y(_10998_) );
NAND2X1 NAND2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__5_), .Y(_10999_) );
NAND2X1 NAND2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_10998_), .B(_10999_), .Y(_11000_) );
NAND2X1 NAND2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__5_), .Y(_11001_) );
NAND2X1 NAND2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__5_), .Y(_11002_) );
NAND2X1 NAND2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_11001_), .B(_11002_), .Y(_11003_) );
NOR2X1 NOR2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_11000_), .B(_11003_), .Y(_11004_) );
NAND3X1 NAND3X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_8762_), .C(_3271_), .Y(_11005_) );
NAND3X1 NAND3X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_8765_), .C(_3225_), .Y(_11006_) );
AND2X2 AND2X2_1576 ( .gnd(gnd), .vdd(vdd), .A(_11006_), .B(_11005_), .Y(_11007_) );
AOI22X1 AOI22X1_190 ( .gnd(gnd), .vdd(vdd), .A(_62__5_), .B(_8774_), .C(_57__5_), .D(_8771_), .Y(_11008_) );
NAND2X1 NAND2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_11007_), .B(_11008_), .Y(_11009_) );
NAND2X1 NAND2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__5_), .Y(_11010_) );
NAND3X1 NAND3X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_2809_), .B(_8786_), .C(_2810_), .Y(_11011_) );
OAI21X1 OAI21X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .B(_8792_), .C(_11011_), .Y(_11012_) );
NAND3X1 NAND3X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_2638_), .B(_8794_), .C(_2639_), .Y(_11013_) );
OAI21X1 OAI21X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_2756_), .B(_8799_), .C(_11013_), .Y(_11014_) );
NOR2X1 NOR2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_11014_), .B(_11012_), .Y(_11015_) );
AOI22X1 AOI22X1_191 ( .gnd(gnd), .vdd(vdd), .A(_75__5_), .B(_8802_), .C(_74__5_), .D(_8803_), .Y(_11016_) );
AOI22X1 AOI22X1_192 ( .gnd(gnd), .vdd(vdd), .A(_80__5_), .B(_8805_), .C(_82__5_), .D(_8806_), .Y(_11017_) );
NAND2X1 NAND2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_11017_), .B(_11016_), .Y(_11018_) );
INVX1 INVX1_3873 ( .gnd(gnd), .vdd(vdd), .A(_84__5_), .Y(_11019_) );
NOR2X1 NOR2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_11019_), .Y(_11020_) );
NOR2X1 NOR2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2292_), .Y(_11021_) );
NAND2X1 NAND2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__5_), .Y(_11022_) );
NAND3X1 NAND3X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_8843_), .C(_2005_), .Y(_11023_) );
NAND3X1 NAND3X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1907_), .C(_1908_), .Y(_11024_) );
NAND3X1 NAND3X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_11024_), .B(_11023_), .C(_11022_), .Y(_11025_) );
NOR3X1 NOR3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_11020_), .B(_11025_), .C(_11021_), .Y(_11026_) );
NAND3X1 NAND3X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_2245_), .B(_8829_), .C(_2246_), .Y(_11027_) );
NAND3X1 NAND3X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_2139_), .B(_8831_), .C(_2140_), .Y(_11028_) );
NAND2X1 NAND2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_11027_), .B(_11028_), .Y(_11029_) );
NAND3X1 NAND3X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_2080_), .B(_8834_), .C(_2081_), .Y(_11030_) );
NAND3X1 NAND3X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_2191_), .B(_8836_), .C(_2192_), .Y(_11031_) );
NAND2X1 NAND2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_11030_), .B(_11031_), .Y(_11032_) );
NOR2X1 NOR2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_11032_), .B(_11029_), .Y(_11033_) );
AOI22X1 AOI22X1_193 ( .gnd(gnd), .vdd(vdd), .A(_98__5_), .B(_8845_), .C(_93__5_), .D(_8840_), .Y(_11034_) );
NAND2X1 NAND2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_91__5_), .Y(_11035_) );
NAND2X1 NAND2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_94__5_), .Y(_11036_) );
NAND3X1 NAND3X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_11035_), .B(_11036_), .C(_11034_), .Y(_11037_) );
NAND2X1 NAND2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__5_), .Y(_11038_) );
NAND3X1 NAND3X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1540_), .C(_1541_), .Y(_11039_) );
NAND3X1 NAND3X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1625_), .C(_1626_), .Y(_11040_) );
NAND2X1 NAND2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_11039_), .B(_11040_), .Y(_11041_) );
NAND3X1 NAND3X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1665_), .C(_1666_), .Y(_11042_) );
NAND3X1 NAND3X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .B(_8857_), .C(_1374_), .Y(_11043_) );
NAND2X1 NAND2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_11043_), .B(_11042_), .Y(_11044_) );
OR2X2 OR2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_11041_), .B(_11044_), .Y(_11045_) );
NOR3X1 NOR3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_8867_), .C(_1209_), .Y(_11046_) );
AOI22X1 AOI22X1_194 ( .gnd(gnd), .vdd(vdd), .A(_191__5_), .B(_8873_), .C(_192__5_), .D(_8872_), .Y(_11047_) );
AOI22X1 AOI22X1_195 ( .gnd(gnd), .vdd(vdd), .A(_195__5_), .B(_8875_), .C(_193__5_), .D(_8876_), .Y(_11048_) );
NAND2X1 NAND2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_11047_), .B(_11048_), .Y(_11049_) );
AOI22X1 AOI22X1_196 ( .gnd(gnd), .vdd(vdd), .A(_188__5_), .B(_8879_), .C(_126__5_), .D(_8881_), .Y(_11050_) );
AOI22X1 AOI22X1_197 ( .gnd(gnd), .vdd(vdd), .A(_196__5_), .B(_8883_), .C(_194__5_), .D(_8884_), .Y(_11051_) );
NAND2X1 NAND2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_11050_), .B(_11051_), .Y(_11052_) );
NOR3X1 NOR3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_11052_), .B(_11046_), .C(_11049_), .Y(_11053_) );
NAND3X1 NAND3X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_5826_), .B(_8893_), .C(_5825_), .Y(_11054_) );
NAND3X1 NAND3X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_8898_), .C(_4585_), .Y(_11055_) );
NAND2X1 NAND2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_11054_), .B(_11055_), .Y(_11056_) );
NAND3X1 NAND3X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_5523_), .B(_8901_), .C(_5522_), .Y(_11057_) );
NAND3X1 NAND3X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_7861_), .B(_8904_), .C(_7860_), .Y(_11058_) );
NAND2X1 NAND2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_11057_), .B(_11058_), .Y(_11059_) );
NOR2X1 NOR2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_11056_), .B(_11059_), .Y(_11060_) );
NAND3X1 NAND3X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_4086_), .B(_8909_), .C(_4085_), .Y(_11061_) );
NAND3X1 NAND3X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3888_), .C(_3887_), .Y(_11062_) );
NAND2X1 NAND2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_11061_), .B(_11062_), .Y(_11063_) );
NAND3X1 NAND3X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_4627_), .B(_8914_), .C(_4626_), .Y(_11064_) );
NAND3X1 NAND3X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_6648_), .B(_8918_), .C(_6647_), .Y(_11065_) );
NAND2X1 NAND2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_11064_), .B(_11065_), .Y(_11066_) );
NOR2X1 NOR2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_11063_), .B(_11066_), .Y(_11067_) );
NAND2X1 NAND2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_11060_), .B(_11067_), .Y(_11068_) );
NAND3X1 NAND3X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_4967_), .B(_8926_), .C(_4966_), .Y(_11069_) );
NAND3X1 NAND3X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_8067_), .B(_8928_), .C(_8066_), .Y(_11070_) );
NAND2X1 NAND2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_11069_), .B(_11070_), .Y(_11071_) );
NAND3X1 NAND3X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_4489_), .B(_8931_), .C(_4488_), .Y(_11072_) );
NAND3X1 NAND3X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_8035_), .B(_8933_), .C(_8034_), .Y(_11073_) );
NAND2X1 NAND2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_11072_), .B(_11073_), .Y(_11074_) );
NOR2X1 NOR2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_11071_), .B(_11074_), .Y(_11075_) );
NAND3X1 NAND3X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_5181_), .B(_8937_), .C(_5180_), .Y(_11076_) );
NAND3X1 NAND3X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_7823_), .B(_8939_), .C(_7822_), .Y(_11077_) );
NAND2X1 NAND2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_11076_), .B(_11077_), .Y(_11078_) );
NAND3X1 NAND3X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_5143_), .B(_8942_), .C(_5142_), .Y(_11079_) );
NAND3X1 NAND3X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_5005_), .B(_8944_), .C(_5004_), .Y(_11080_) );
NAND2X1 NAND2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_11079_), .B(_11080_), .Y(_11081_) );
NOR2X1 NOR2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_11081_), .B(_11078_), .Y(_11082_) );
NAND2X1 NAND2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_11075_), .B(_11082_), .Y(_11083_) );
NOR2X1 NOR2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_11068_), .B(_11083_), .Y(_11084_) );
NAND3X1 NAND3X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_5606_), .B(_9160_), .C(_5605_), .Y(_11085_) );
NAND3X1 NAND3X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_9161_), .C(_3696_), .Y(_11086_) );
NAND2X1 NAND2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_11085_), .B(_11086_), .Y(_11087_) );
NAND3X1 NAND3X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .B(_9150_), .C(_4547_), .Y(_11088_) );
NAND3X1 NAND3X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_7521_), .B(_9151_), .C(_7520_), .Y(_11089_) );
NAND2X1 NAND2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_11088_), .B(_11089_), .Y(_11090_) );
NOR2X1 NOR2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_11087_), .B(_11090_), .Y(_11091_) );
NAND3X1 NAND3X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_5578_), .B(_9356_), .C(_5577_), .Y(_11092_) );
NAND3X1 NAND3X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_6161_), .B(_9357_), .C(_6160_), .Y(_11093_) );
NAND2X1 NAND2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_11092_), .B(_11093_), .Y(_11094_) );
NAND3X1 NAND3X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_6016_), .B(_9157_), .C(_6015_), .Y(_11095_) );
NAND3X1 NAND3X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_9158_), .C(_3730_), .Y(_11096_) );
NAND2X1 NAND2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_11096_), .B(_11095_), .Y(_11097_) );
NOR2X1 NOR2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_11094_), .B(_11097_), .Y(_11098_) );
NAND2X1 NAND2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_11091_), .B(_11098_), .Y(_11099_) );
NAND3X1 NAND3X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_7755_), .B(_9173_), .C(_7754_), .Y(_11100_) );
NAND3X1 NAND3X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(_8975_), .C(_3473_), .Y(_11101_) );
NAND2X1 NAND2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_11100_), .B(_11101_), .Y(_11102_) );
NAND3X1 NAND3X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_4049_), .B(_8978_), .C(_4048_), .Y(_11103_) );
NAND3X1 NAND3X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_4123_), .B(_8980_), .C(_4122_), .Y(_11104_) );
NAND2X1 NAND2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_11104_), .B(_11103_), .Y(_11105_) );
NOR2X1 NOR2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_11102_), .B(_11105_), .Y(_11106_) );
NAND3X1 NAND3X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_5634_), .B(_9153_), .C(_5633_), .Y(_11107_) );
NAND3X1 NAND3X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_5338_), .B(_9154_), .C(_5337_), .Y(_11108_) );
NAND2X1 NAND2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_11107_), .B(_11108_), .Y(_11109_) );
NAND3X1 NAND3X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_7997_), .B(_9177_), .C(_7996_), .Y(_11110_) );
NAND3X1 NAND3X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_6571_), .B(_8989_), .C(_6570_), .Y(_11111_) );
NAND2X1 NAND2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_11111_), .B(_11110_), .Y(_11112_) );
NOR2X1 NOR2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_11109_), .B(_11112_), .Y(_11113_) );
NAND2X1 NAND2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_11106_), .B(_11113_), .Y(_11114_) );
NOR2X1 NOR2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_11099_), .B(_11114_), .Y(_11115_) );
NAND2X1 NAND2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_11084_), .B(_11115_), .Y(_11116_) );
NAND3X1 NAND3X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_8998_), .C(_4897_), .Y(_11117_) );
NAND3X1 NAND3X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_6505_), .B(_9002_), .C(_6504_), .Y(_11118_) );
NAND2X1 NAND2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_11117_), .B(_11118_), .Y(_11119_) );
NAND3X1 NAND3X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_5711_), .B(_9005_), .C(_5710_), .Y(_11120_) );
NAND3X1 NAND3X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_4859_), .B(_9007_), .C(_4858_), .Y(_11121_) );
NAND2X1 NAND2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_11120_), .B(_11121_), .Y(_11122_) );
NOR2X1 NOR2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_11119_), .B(_11122_), .Y(_11123_) );
NAND3X1 NAND3X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_5749_), .B(_9011_), .C(_5748_), .Y(_11124_) );
NAND3X1 NAND3X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_6791_), .B(_9013_), .C(_6790_), .Y(_11125_) );
NAND2X1 NAND2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_11124_), .B(_11125_), .Y(_11126_) );
NAND3X1 NAND3X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_6752_), .B(_9016_), .C(_6751_), .Y(_11127_) );
NAND3X1 NAND3X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_6538_), .B(_9174_), .C(_6537_), .Y(_11128_) );
NAND2X1 NAND2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_11127_), .B(_11128_), .Y(_11129_) );
NOR2X1 NOR2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_11129_), .B(_11126_), .Y(_11130_) );
NAND2X1 NAND2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_11123_), .B(_11130_), .Y(_11131_) );
NAND3X1 NAND3X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_6275_), .B(_9024_), .C(_6274_), .Y(_11132_) );
NAND3X1 NAND3X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_6347_), .B(_9026_), .C(_6346_), .Y(_11133_) );
NAND2X1 NAND2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_11132_), .B(_11133_), .Y(_11134_) );
NAND3X1 NAND3X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_6052_), .B(_9029_), .C(_6051_), .Y(_11135_) );
NAND3X1 NAND3X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_6110_), .B(_9031_), .C(_6109_), .Y(_11136_) );
NAND2X1 NAND2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_11135_), .B(_11136_), .Y(_11137_) );
NOR2X1 NOR2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_11134_), .B(_11137_), .Y(_11138_) );
NAND3X1 NAND3X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_5670_), .B(_9035_), .C(_5669_), .Y(_11139_) );
NAND3X1 NAND3X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_4666_), .B(_9037_), .C(_4665_), .Y(_11140_) );
NAND2X1 NAND2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_11140_), .B(_11139_), .Y(_11141_) );
NAND3X1 NAND3X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_6311_), .B(_9040_), .C(_6310_), .Y(_11142_) );
NAND3X1 NAND3X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_4328_), .B(_9042_), .C(_4327_), .Y(_11143_) );
NAND2X1 NAND2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_11142_), .B(_11143_), .Y(_11144_) );
NOR2X1 NOR2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_11144_), .B(_11141_), .Y(_11145_) );
NAND2X1 NAND2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_11138_), .B(_11145_), .Y(_11146_) );
NOR2X1 NOR2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_11131_), .B(_11146_), .Y(_11147_) );
NAND3X1 NAND3X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_6199_), .B(_9048_), .C(_6198_), .Y(_11148_) );
NAND3X1 NAND3X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_7934_), .B(_9050_), .C(_7933_), .Y(_11149_) );
NAND2X1 NAND2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_11148_), .B(_11149_), .Y(_11150_) );
NAND3X1 NAND3X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_5483_), .B(_9053_), .C(_5482_), .Y(_11151_) );
NAND3X1 NAND3X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_7897_), .B(_9055_), .C(_7896_), .Y(_11152_) );
NAND2X1 NAND2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_11151_), .B(_11152_), .Y(_11153_) );
NOR2X1 NOR2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_11150_), .B(_11153_), .Y(_11154_) );
NAND3X1 NAND3X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_4449_), .B(_9059_), .C(_4448_), .Y(_11155_) );
NAND3X1 NAND3X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_4409_), .B(_9061_), .C(_4408_), .Y(_11156_) );
NAND2X1 NAND2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_11155_), .B(_11156_), .Y(_11157_) );
NAND3X1 NAND3X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_6237_), .B(_9064_), .C(_6236_), .Y(_11158_) );
NAND3X1 NAND3X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_4369_), .B(_9066_), .C(_4368_), .Y(_11159_) );
NAND2X1 NAND2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_11158_), .B(_11159_), .Y(_11160_) );
NOR2X1 NOR2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_11160_), .B(_11157_), .Y(_11161_) );
NAND2X1 NAND2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_11154_), .B(_11161_), .Y(_11162_) );
NAND3X1 NAND3X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_7593_), .B(_9071_), .C(_7592_), .Y(_11163_) );
NAND3X1 NAND3X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_7557_), .B(_9073_), .C(_7556_), .Y(_11164_) );
NAND2X1 NAND2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_11163_), .B(_11164_), .Y(_11165_) );
NAND3X1 NAND3X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_5787_), .B(_9076_), .C(_5786_), .Y(_11166_) );
NAND3X1 NAND3X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_3513_), .B(_9078_), .C(_3512_), .Y(_11167_) );
NAND2X1 NAND2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_11166_), .B(_11167_), .Y(_11168_) );
NOR2X1 NOR2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_11165_), .B(_11168_), .Y(_11169_) );
NAND3X1 NAND3X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_5442_), .B(_9082_), .C(_5441_), .Y(_11170_) );
NAND3X1 NAND3X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_3809_), .B(_9084_), .C(_3808_), .Y(_11171_) );
NAND2X1 NAND2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_11171_), .B(_11170_), .Y(_11172_) );
NAND3X1 NAND3X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_6608_), .B(_9087_), .C(_6607_), .Y(_11173_) );
NAND3X1 NAND3X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_3662_), .B(_9089_), .C(_3661_), .Y(_11174_) );
NAND2X1 NAND2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_11173_), .B(_11174_), .Y(_11175_) );
NOR2X1 NOR2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_11172_), .B(_11175_), .Y(_11176_) );
NAND2X1 NAND2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_11169_), .B(_11176_), .Y(_11177_) );
NOR2X1 NOR2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_11162_), .B(_11177_), .Y(_11178_) );
NAND2X1 NAND2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_11147_), .B(_11178_), .Y(_11179_) );
NOR2X1 NOR2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_11116_), .B(_11179_), .Y(_11180_) );
NAND2X1 NAND2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__5_), .Y(_11181_) );
NAND3X1 NAND3X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_6969_), .B(_9145_), .C(_6968_), .Y(_11182_) );
NAND2X1 NAND2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_11181_), .B(_11182_), .Y(_11183_) );
NAND3X1 NAND3X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_5042_), .B(_9135_), .C(_5043_), .Y(_11184_) );
NAND3X1 NAND3X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_6927_), .B(_9137_), .C(_6926_), .Y(_11185_) );
NAND2X1 NAND2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_11184_), .B(_11185_), .Y(_11186_) );
NOR2X1 NOR2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_11186_), .B(_11183_), .Y(_11187_) );
NAND3X1 NAND3X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_15917_), .B(_9109_), .C(_15918_), .Y(_11188_) );
NAND3X1 NAND3X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_8382_), .B(_9113_), .C(_8383_), .Y(_11189_) );
NAND3X1 NAND3X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_16124_), .B(_9115_), .C(_16123_), .Y(_11190_) );
NAND3X1 NAND3X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_11188_), .B(_11189_), .C(_11190_), .Y(_11191_) );
NAND3X1 NAND3X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_388_), .C(_389_), .Y(_11192_) );
NAND3X1 NAND3X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_15860_), .B(_9120_), .C(_15861_), .Y(_11193_) );
AND2X2 AND2X2_1577 ( .gnd(gnd), .vdd(vdd), .A(_11193_), .B(_11192_), .Y(_11194_) );
AOI22X1 AOI22X1_198 ( .gnd(gnd), .vdd(vdd), .A(_201__5_), .B(_9124_), .C(_89__5_), .D(_9123_), .Y(_11195_) );
NAND2X1 NAND2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_11194_), .B(_11195_), .Y(_11196_) );
NAND3X1 NAND3X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_4697_), .B(_9140_), .C(_4698_), .Y(_11197_) );
OAI21X1 OAI21X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_5236_), .B(_10036_), .C(_11197_), .Y(_11198_) );
NOR3X1 NOR3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_11191_), .B(_11198_), .C(_11196_), .Y(_11199_) );
NAND3X1 NAND3X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3416_), .C(_3417_), .Y(_11200_) );
NAND2X1 NAND2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__5_), .Y(_11201_) );
NAND3X1 NAND3X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_5089_), .B(_9102_), .C(_5090_), .Y(_11202_) );
NAND3X1 NAND3X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_11200_), .B(_11202_), .C(_11201_), .Y(_11203_) );
AOI22X1 AOI22X1_199 ( .gnd(gnd), .vdd(vdd), .A(_38__5_), .B(_9129_), .C(_16__5_), .D(_9127_), .Y(_11204_) );
NAND2X1 NAND2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_9104_), .B(_204__5_), .Y(_11205_) );
NAND2X1 NAND2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_9099_), .B(_39__5_), .Y(_11206_) );
NAND3X1 NAND3X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_11206_), .B(_11205_), .C(_11204_), .Y(_11207_) );
NOR2X1 NOR2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_11203_), .B(_11207_), .Y(_11208_) );
NAND3X1 NAND3X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_11187_), .B(_11208_), .C(_11199_), .Y(_11209_) );
AOI22X1 AOI22X1_200 ( .gnd(gnd), .vdd(vdd), .A(_30__5_), .B(_9167_), .C(_227__5_), .D(_9170_), .Y(_11210_) );
AOI22X1 AOI22X1_201 ( .gnd(gnd), .vdd(vdd), .A(_209__5_), .B(_8957_), .C(_33__5_), .D(_8991_), .Y(_11211_) );
NAND2X1 NAND2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_11210_), .B(_11211_), .Y(_11212_) );
AOI22X1 AOI22X1_202 ( .gnd(gnd), .vdd(vdd), .A(_44__5_), .B(_8968_), .C(_42__5_), .D(_8963_), .Y(_11213_) );
AOI22X1 AOI22X1_203 ( .gnd(gnd), .vdd(vdd), .A(_236__5_), .B(_8955_), .C(_208__5_), .D(_8950_), .Y(_11214_) );
NAND2X1 NAND2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_11213_), .B(_11214_), .Y(_11215_) );
NOR2X1 NOR2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_11212_), .B(_11215_), .Y(_11216_) );
AOI22X1 AOI22X1_204 ( .gnd(gnd), .vdd(vdd), .A(_22__5_), .B(_9382_), .C(_3__5_), .D(_9383_), .Y(_11217_) );
AOI22X1 AOI22X1_205 ( .gnd(gnd), .vdd(vdd), .A(_232__5_), .B(_9354_), .C(_219__5_), .D(_9353_), .Y(_11218_) );
NAND2X1 NAND2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_11217_), .B(_11218_), .Y(_11219_) );
AOI22X1 AOI22X1_206 ( .gnd(gnd), .vdd(vdd), .A(_255__5_), .B(_8986_), .C(_254__5_), .D(_8984_), .Y(_11220_) );
AOI22X1 AOI22X1_207 ( .gnd(gnd), .vdd(vdd), .A(_203__5_), .B(_9018_), .C(_156__5_), .D(_8973_), .Y(_11221_) );
NAND2X1 NAND2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_11221_), .B(_11220_), .Y(_11222_) );
NOR2X1 NOR2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_11219_), .B(_11222_), .Y(_11223_) );
NAND2X1 NAND2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_11216_), .B(_11223_), .Y(_11224_) );
AOI22X1 AOI22X1_208 ( .gnd(gnd), .vdd(vdd), .A(_234__5_), .B(_9182_), .C(_34__5_), .D(_9183_), .Y(_11225_) );
NAND2X1 NAND2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__5_), .Y(_11226_) );
NAND2X1 NAND2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__5_), .Y(_11227_) );
NAND3X1 NAND3X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_11226_), .B(_11227_), .C(_11225_), .Y(_11228_) );
NAND3X1 NAND3X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_15650_), .B(_9192_), .C(_15651_), .Y(_11229_) );
OAI21X1 OAI21X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_15601_), .B(_9195_), .C(_11229_), .Y(_11230_) );
NAND2X1 NAND2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__5_), .Y(_11231_) );
NAND3X1 NAND3X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_15706_), .B(_9199_), .C(_15707_), .Y(_11232_) );
NAND2X1 NAND2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_11231_), .B(_11232_), .Y(_11233_) );
NOR2X1 NOR2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_11233_), .B(_11230_), .Y(_11234_) );
NAND2X1 NAND2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__5_), .Y(_11235_) );
OAI21X1 OAI21X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_15304_), .B(_9206_), .C(_11235_), .Y(_11236_) );
NAND2X1 NAND2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__5_), .Y(_11237_) );
OAI21X1 OAI21X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_15098_), .B(_9211_), .C(_11237_), .Y(_11238_) );
NOR2X1 NOR2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_11236_), .B(_11238_), .Y(_11239_) );
NOR3X1 NOR3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_15969_), .B(_9215_), .C(_15970_), .Y(_11240_) );
NAND3X1 NAND3X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_15252_), .B(_9217_), .C(_15253_), .Y(_11241_) );
NAND3X1 NAND3X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_15200_), .B(_9219_), .C(_15199_), .Y(_11242_) );
NAND2X1 NAND2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_11242_), .B(_11241_), .Y(_11243_) );
NAND3X1 NAND3X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_15474_), .B(_9222_), .C(_15475_), .Y(_11244_) );
NAND3X1 NAND3X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_15421_), .B(_9224_), .C(_15420_), .Y(_11245_) );
NAND2X1 NAND2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_11244_), .B(_11245_), .Y(_11246_) );
NOR3X1 NOR3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_11240_), .B(_11246_), .C(_11243_), .Y(_11247_) );
NAND3X1 NAND3X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_11239_), .B(_11247_), .C(_11234_), .Y(_11248_) );
NAND2X1 NAND2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__5_), .Y(_11249_) );
NAND3X1 NAND3X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_15532_), .B(_9233_), .C(_15533_), .Y(_11250_) );
NOR2X1 NOR2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .B(_7003_), .Y(_11251_) );
NOR2X1 NOR2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_9259_), .B(_6461_), .Y(_11252_) );
AND2X2 AND2X2_1578 ( .gnd(gnd), .vdd(vdd), .A(_186__5_), .B(_9298_), .Y(_11253_) );
NOR3X1 NOR3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_11251_), .B(_11252_), .C(_11253_), .Y(_11254_) );
NAND2X1 NAND2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__5_), .Y(_11255_) );
OAI21X1 OAI21X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_3596_), .B(_9295_), .C(_11255_), .Y(_11256_) );
OAI21X1 OAI21X1_2451 ( .gnd(gnd), .vdd(vdd), .A(IDATA_PROG_data_5_bF_buf1), .B(_8216_), .C(_8227_), .Y(_11257_) );
NAND2X1 NAND2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_173__5_), .Y(_11258_) );
OAI21X1 OAI21X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_11257_), .B(_10875_), .C(_11258_), .Y(_11259_) );
NOR2X1 NOR2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_11256_), .B(_11259_), .Y(_11260_) );
NAND2X1 NAND2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_1__5_), .B(_9242_), .Y(_11261_) );
NAND3X1 NAND3X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_9268_), .C(_1165_), .Y(_11262_) );
NAND2X1 NAND2X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_11262_), .B(_11261_), .Y(_11263_) );
INVX4 INVX4_80 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .Y(_11264_) );
NAND3X1 NAND3X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_1759_), .B(_9255_), .C(_1760_), .Y(_11265_) );
OAI21X1 OAI21X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_15804_), .B(_11264_), .C(_11265_), .Y(_11266_) );
NOR2X1 NOR2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_11266_), .B(_11263_), .Y(_11267_) );
NAND3X1 NAND3X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_11254_), .B(_11267_), .C(_11260_), .Y(_11268_) );
NAND3X1 NAND3X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_7672_), .B(_9321_), .C(_7673_), .Y(_11269_) );
NAND2X1 NAND2X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_9300_), .B(_182__5_), .Y(_11270_) );
NAND3X1 NAND3X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_7085_), .B(_9244_), .C(_7086_), .Y(_11271_) );
NAND3X1 NAND3X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_11270_), .B(_11269_), .C(_11271_), .Y(_11272_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_5924_), .B(_9323_), .C(_6423_), .D(_9763_), .Y(_11273_) );
NOR2X1 NOR2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_11273_), .B(_11272_), .Y(_11274_) );
NAND3X1 NAND3X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_7040_), .B(_9266_), .C(_7041_), .Y(_11275_) );
OAI21X1 OAI21X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_2906_), .B(_10468_), .C(_11275_), .Y(_11276_) );
NOR2X1 NOR2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_10471_), .B(_7463_), .Y(_11277_) );
AND2X2 AND2X2_1579 ( .gnd(gnd), .vdd(vdd), .A(_137__5_), .B(_9262_), .Y(_11278_) );
NOR3X1 NOR3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_11277_), .B(_11278_), .C(_11276_), .Y(_11279_) );
NAND3X1 NAND3X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_7709_), .B(_9248_), .C(_7710_), .Y(_11280_) );
OAI21X1 OAI21X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_4182_), .B(_9254_), .C(_11280_), .Y(_11281_) );
NOR2X1 NOR2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_8158_), .Y(_11282_) );
NOR2X1 NOR2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_9306_), .B(_3547_), .Y(_11283_) );
NOR3X1 NOR3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_11282_), .B(_11283_), .C(_11281_), .Y(_11284_) );
NAND3X1 NAND3X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_11274_), .B(_11279_), .C(_11284_), .Y(_11285_) );
NAND2X1 NAND2X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_9274_), .B(_14__5_), .Y(_11286_) );
AOI22X1 AOI22X1_209 ( .gnd(gnd), .vdd(vdd), .A(_31__5_), .B(_9283_), .C(_251__5_), .D(_9320_), .Y(_11287_) );
NAND3X1 NAND3X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_4775_), .B(_9313_), .C(_4776_), .Y(_11288_) );
OAI21X1 OAI21X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_5366_), .B(_9325_), .C(_11288_), .Y(_11289_) );
NAND3X1 NAND3X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_2351_), .B(_9315_), .C(_2352_), .Y(_11290_) );
OAI21X1 OAI21X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_5959_), .B(_10503_), .C(_11290_), .Y(_11291_) );
NOR2X1 NOR2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_11289_), .B(_11291_), .Y(_11292_) );
NAND3X1 NAND3X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_11286_), .B(_11287_), .C(_11292_), .Y(_11293_) );
NOR3X1 NOR3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_11285_), .B(_11293_), .C(_11268_), .Y(_11294_) );
NAND2X1 NAND2X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_11250_), .B(_11294_), .Y(_11295_) );
AOI21X1 AOI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_157__5_), .B(_9232_), .C(_11295_), .Y(_11296_) );
AOI22X1 AOI22X1_210 ( .gnd(gnd), .vdd(vdd), .A(_155__5_), .B(_9333_), .C(_172__5_), .D(_9332_), .Y(_11297_) );
NAND3X1 NAND3X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_11297_), .B(_11249_), .C(_11296_), .Y(_11298_) );
NOR3X1 NOR3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_11298_), .B(_11228_), .C(_11248_), .Y(_11299_) );
NAND2X1 NAND2X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__5_), .Y(_11300_) );
NAND3X1 NAND3X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_9339_), .C(_443_), .Y(_11301_) );
AOI22X1 AOI22X1_211 ( .gnd(gnd), .vdd(vdd), .A(_111__5_), .B(_9342_), .C(_12__5_), .D(_9341_), .Y(_11302_) );
NAND3X1 NAND3X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_11302_), .B(_11300_), .C(_11301_), .Y(_11303_) );
AOI22X1 AOI22X1_212 ( .gnd(gnd), .vdd(vdd), .A(_100__5_), .B(_9346_), .C(_212__5_), .D(_9345_), .Y(_11304_) );
AOI22X1 AOI22X1_213 ( .gnd(gnd), .vdd(vdd), .A(_245__5_), .B(_9348_), .C(_140__5_), .D(_9349_), .Y(_11305_) );
NAND2X1 NAND2X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_11305_), .B(_11304_), .Y(_11306_) );
NOR2X1 NOR2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_11303_), .B(_11306_), .Y(_11307_) );
AOI22X1 AOI22X1_214 ( .gnd(gnd), .vdd(vdd), .A(_40__5_), .B(_8952_), .C(_29__5_), .D(_9176_), .Y(_11308_) );
AOI22X1 AOI22X1_215 ( .gnd(gnd), .vdd(vdd), .A(_218__5_), .B(_9169_), .C(_247__5_), .D(_9165_), .Y(_11309_) );
NAND2X1 NAND2X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_11309_), .B(_11308_), .Y(_11310_) );
NAND3X1 NAND3X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16179_), .C(_16180_), .Y(_11311_) );
OAI21X1 OAI21X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_16230_), .B(_9361_), .C(_11311_), .Y(_11312_) );
NAND3X1 NAND3X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16077_), .C(_16078_), .Y(_11313_) );
NAND3X1 NAND3X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16022_), .C(_16023_), .Y(_11314_) );
NAND2X1 NAND2X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_11313_), .B(_11314_), .Y(_11315_) );
NOR2X1 NOR2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_11315_), .B(_11312_), .Y(_11316_) );
NAND3X1 NAND3X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_8664_), .B(_9371_), .C(_8663_), .Y(_11317_) );
NAND3X1 NAND3X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8556_), .C(_8555_), .Y(_11318_) );
NAND2X1 NAND2X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_11318_), .B(_11317_), .Y(_11319_) );
NAND3X1 NAND3X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8609_), .C(_8610_), .Y(_11320_) );
NAND3X1 NAND3X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_306_), .C(_307_), .Y(_11321_) );
NAND2X1 NAND2X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_11320_), .B(_11321_), .Y(_11322_) );
NOR2X1 NOR2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_11322_), .B(_11319_), .Y(_11323_) );
AOI22X1 AOI22X1_216 ( .gnd(gnd), .vdd(vdd), .A(_237__5_), .B(_8966_), .C(_177__5_), .D(_8961_), .Y(_11324_) );
NAND3X1 NAND3X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_11316_), .B(_11323_), .C(_11324_), .Y(_11325_) );
NOR2X1 NOR2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_11325_), .B(_11310_), .Y(_11326_) );
NAND3X1 NAND3X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_11307_), .B(_11326_), .C(_11299_), .Y(_11327_) );
NOR3X1 NOR3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_11209_), .B(_11224_), .C(_11327_), .Y(_11328_) );
NAND3X1 NAND3X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_11053_), .B(_11328_), .C(_11180_), .Y(_11329_) );
NAND2X1 NAND2X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__5_), .Y(_11330_) );
NAND2X1 NAND2X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__5_), .Y(_11331_) );
NAND2X1 NAND2X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_11331_), .B(_11330_), .Y(_11332_) );
NOR3X1 NOR3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_11045_), .B(_11332_), .C(_11329_), .Y(_11333_) );
NOR3X1 NOR3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_9397_), .C(_1851_), .Y(_11334_) );
NAND3X1 NAND3X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1454_), .C(_1453_), .Y(_11335_) );
NAND3X1 NAND3X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_9453_), .B(_1408_), .C(_1407_), .Y(_11336_) );
NAND2X1 NAND2X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_11335_), .B(_11336_), .Y(_11337_) );
NAND3X1 NAND3X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1504_), .C(_1503_), .Y(_11338_) );
NAND3X1 NAND3X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1287_), .C(_1286_), .Y(_11339_) );
NAND2X1 NAND2X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_11338_), .B(_11339_), .Y(_11340_) );
NOR2X1 NOR2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_11340_), .B(_11337_), .Y(_11341_) );
AOI22X1 AOI22X1_217 ( .gnd(gnd), .vdd(vdd), .A(_125__5_), .B(_9411_), .C(_122__5_), .D(_9444_), .Y(_11342_) );
NAND3X1 NAND3X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_9413_), .C(_1097_), .Y(_11343_) );
NAND2X1 NAND2X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__5_), .Y(_11344_) );
NAND3X1 NAND3X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_11343_), .B(_11344_), .C(_11342_), .Y(_11345_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_9421_), .C(_810_), .D(_9419_), .Y(_11346_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_9426_), .C(_695_), .D(_9424_), .Y(_11347_) );
NOR2X1 NOR2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_11346_), .B(_11347_), .Y(_11348_) );
NAND3X1 NAND3X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7410_), .C(_7411_), .Y(_11349_) );
NAND3X1 NAND3X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_9431_), .C(_536_), .Y(_11350_) );
AOI22X1 AOI22X1_218 ( .gnd(gnd), .vdd(vdd), .A(_138__5_), .B(_9434_), .C(_229__5_), .D(_9433_), .Y(_11351_) );
NAND3X1 NAND3X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_11350_), .B(_11349_), .C(_11351_), .Y(_11352_) );
NAND3X1 NAND3X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_657_), .C(_658_), .Y(_11353_) );
OAI21X1 OAI21X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_9440_), .C(_11353_), .Y(_11354_) );
NOR2X1 NOR2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_11354_), .B(_11352_), .Y(_11355_) );
NAND2X1 NAND2X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_11355_), .B(_11348_), .Y(_11356_) );
NAND3X1 NAND3X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_9410_), .C(_1006_), .Y(_11357_) );
NAND2X1 NAND2X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__5_), .Y(_11358_) );
AOI22X1 AOI22X1_219 ( .gnd(gnd), .vdd(vdd), .A(_130__5_), .B(_9449_), .C(_127__5_), .D(_9448_), .Y(_11359_) );
NAND3X1 NAND3X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_11357_), .B(_11358_), .C(_11359_), .Y(_11360_) );
NOR3X1 NOR3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_11360_), .B(_11345_), .C(_11356_), .Y(_11361_) );
AOI22X1 AOI22X1_220 ( .gnd(gnd), .vdd(vdd), .A(_115__5_), .B(_9399_), .C(_114__5_), .D(_9454_), .Y(_11362_) );
NAND3X1 NAND3X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_11362_), .B(_11341_), .C(_11361_), .Y(_11363_) );
NAND3X1 NAND3X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(_9457_), .C(_1708_), .Y(_11364_) );
NAND2X1 NAND2X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__5_), .Y(_11365_) );
NAND2X1 NAND2X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_11365_), .B(_11364_), .Y(_11366_) );
NOR3X1 NOR3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_11366_), .B(_11334_), .C(_11363_), .Y(_11367_) );
NAND3X1 NAND3X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_11038_), .B(_11367_), .C(_11333_), .Y(_11368_) );
NOR2X1 NOR2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_11037_), .B(_11368_), .Y(_11369_) );
NAND3X1 NAND3X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_11026_), .B(_11033_), .C(_11369_), .Y(_11370_) );
NAND2X1 NAND2X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__5_), .Y(_11371_) );
NAND3X1 NAND3X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_9468_), .C(_2434_), .Y(_11372_) );
NAND2X1 NAND2X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_11372_), .B(_11371_), .Y(_11373_) );
NOR3X1 NOR3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_11018_), .B(_11373_), .C(_11370_), .Y(_11374_) );
NAND3X1 NAND3X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_11010_), .B(_11015_), .C(_11374_), .Y(_11375_) );
NAND3X1 NAND3X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_9473_), .C(_3056_), .Y(_11376_) );
NAND2X1 NAND2X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__5_), .Y(_11377_) );
NAND2X1 NAND2X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__5_), .Y(_11378_) );
NAND2X1 NAND2X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__5_), .Y(_11379_) );
NAND2X1 NAND2X1_1821 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__5_), .Y(_11380_) );
NAND3X1 NAND3X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_11380_), .B(_11378_), .C(_11379_), .Y(_11381_) );
AOI21X1 AOI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_68__5_), .B(_9477_), .C(_11381_), .Y(_11382_) );
NAND3X1 NAND3X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_11376_), .B(_11382_), .C(_11377_), .Y(_11383_) );
NOR3X1 NOR3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_11009_), .B(_11383_), .C(_11375_), .Y(_11384_) );
AOI21X1 AOI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_11004_), .B(_11384_), .C(rst), .Y(_0__5_) );
NAND2X1 NAND2X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__6_), .Y(_11385_) );
NAND2X1 NAND2X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__6_), .Y(_11386_) );
NAND2X1 NAND2X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_11385_), .B(_11386_), .Y(_11387_) );
NAND2X1 NAND2X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__6_), .Y(_11388_) );
NAND2X1 NAND2X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__6_), .Y(_11389_) );
NAND2X1 NAND2X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_11388_), .B(_11389_), .Y(_11390_) );
NOR2X1 NOR2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_11387_), .B(_11390_), .Y(_11391_) );
NAND3X1 NAND3X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_3275_), .B(_8762_), .C(_3274_), .Y(_11392_) );
NAND3X1 NAND3X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_3229_), .B(_8765_), .C(_3228_), .Y(_11393_) );
AND2X2 AND2X2_1580 ( .gnd(gnd), .vdd(vdd), .A(_11393_), .B(_11392_), .Y(_11394_) );
AOI22X1 AOI22X1_221 ( .gnd(gnd), .vdd(vdd), .A(_62__6_), .B(_8774_), .C(_57__6_), .D(_8771_), .Y(_11395_) );
NAND2X1 NAND2X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_11394_), .B(_11395_), .Y(_11396_) );
NAND2X1 NAND2X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__6_), .Y(_11397_) );
NAND3X1 NAND3X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_2812_), .B(_8786_), .C(_2813_), .Y(_11398_) );
OAI21X1 OAI21X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_2703_), .B(_8792_), .C(_11398_), .Y(_11399_) );
NAND3X1 NAND3X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .B(_8794_), .C(_2642_), .Y(_11400_) );
OAI21X1 OAI21X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_2759_), .B(_8799_), .C(_11400_), .Y(_11401_) );
NOR2X1 NOR2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_11401_), .B(_11399_), .Y(_11402_) );
AOI22X1 AOI22X1_222 ( .gnd(gnd), .vdd(vdd), .A(_76__6_), .B(_9482_), .C(_77__6_), .D(_9478_), .Y(_11403_) );
NAND2X1 NAND2X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__6_), .Y(_11404_) );
NAND2X1 NAND2X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_82__6_), .Y(_11405_) );
NAND3X1 NAND3X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_11404_), .B(_11405_), .C(_11403_), .Y(_11406_) );
NAND2X1 NAND2X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__6_), .Y(_11407_) );
NAND3X1 NAND3X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_2583_), .B(_8803_), .C(_2582_), .Y(_11408_) );
NAND2X1 NAND2X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_11408_), .B(_11407_), .Y(_11409_) );
INVX1 INVX1_3874 ( .gnd(gnd), .vdd(vdd), .A(_84__6_), .Y(_11410_) );
NOR2X1 NOR2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_11410_), .Y(_11411_) );
NOR2X1 NOR2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2294_), .Y(_11412_) );
NAND2X1 NAND2X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__6_), .Y(_11413_) );
NAND3X1 NAND3X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_2043_), .B(_8823_), .C(_2044_), .Y(_11414_) );
NAND3X1 NAND3X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1910_), .C(_1911_), .Y(_11415_) );
NAND3X1 NAND3X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_11415_), .B(_11414_), .C(_11413_), .Y(_11416_) );
NOR3X1 NOR3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_11411_), .B(_11416_), .C(_11412_), .Y(_11417_) );
NAND3X1 NAND3X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_2248_), .B(_8829_), .C(_2249_), .Y(_11418_) );
NAND3X1 NAND3X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_8831_), .C(_2143_), .Y(_11419_) );
NAND2X1 NAND2X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_11418_), .B(_11419_), .Y(_11420_) );
NAND3X1 NAND3X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_8834_), .C(_2084_), .Y(_11421_) );
NAND3X1 NAND3X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_2194_), .B(_8836_), .C(_2195_), .Y(_11422_) );
NAND2X1 NAND2X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_11421_), .B(_11422_), .Y(_11423_) );
NOR2X1 NOR2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_11423_), .B(_11420_), .Y(_11424_) );
AOI22X1 AOI22X1_223 ( .gnd(gnd), .vdd(vdd), .A(_94__6_), .B(_8841_), .C(_93__6_), .D(_8840_), .Y(_11425_) );
AOI22X1 AOI22X1_224 ( .gnd(gnd), .vdd(vdd), .A(_98__6_), .B(_8845_), .C(_92__6_), .D(_8843_), .Y(_11426_) );
NAND2X1 NAND2X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_11426_), .B(_11425_), .Y(_11427_) );
NAND2X1 NAND2X1_1838 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__6_), .Y(_11428_) );
NAND2X1 NAND2X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__6_), .Y(_11429_) );
NAND2X1 NAND2X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__6_), .Y(_11430_) );
NAND2X1 NAND2X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_11429_), .B(_11430_), .Y(_11431_) );
NAND2X1 NAND2X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__6_), .Y(_11432_) );
NAND2X1 NAND2X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__6_), .Y(_11433_) );
NAND2X1 NAND2X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_11433_), .B(_11432_), .Y(_11434_) );
NOR2X1 NOR2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_11434_), .B(_11431_), .Y(_11435_) );
NAND2X1 NAND2X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__6_), .Y(_11436_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_7139_), .B(_9930_), .C(_7183_), .D(_9929_), .Y(_11437_) );
NOR2X1 NOR2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7318_), .Y(_11438_) );
NOR2X1 NOR2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7275_), .Y(_11439_) );
NOR3X1 NOR3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_11438_), .B(_11439_), .C(_11437_), .Y(_11440_) );
NAND2X1 NAND2X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__6_), .Y(_11441_) );
NAND2X1 NAND2X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__6_), .Y(_11442_) );
NAND2X1 NAND2X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_11441_), .B(_11442_), .Y(_11443_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_7361_), .B(_9940_), .C(_7229_), .D(_9941_), .Y(_11444_) );
NOR2X1 NOR2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_11444_), .B(_11443_), .Y(_11445_) );
NAND3X1 NAND3X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_11436_), .B(_11440_), .C(_11445_), .Y(_11446_) );
AOI22X1 AOI22X1_225 ( .gnd(gnd), .vdd(vdd), .A(_20__6_), .B(_8898_), .C(_236__6_), .D(_8955_), .Y(_11447_) );
AOI22X1 AOI22X1_226 ( .gnd(gnd), .vdd(vdd), .A(_237__6_), .B(_8966_), .C(_175__6_), .D(_8904_), .Y(_11448_) );
NAND2X1 NAND2X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_11447_), .B(_11448_), .Y(_11449_) );
NAND2X1 NAND2X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__6_), .Y(_11450_) );
NAND2X1 NAND2X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__6_), .Y(_11451_) );
AOI22X1 AOI22X1_227 ( .gnd(gnd), .vdd(vdd), .A(_19__6_), .B(_8914_), .C(_210__6_), .D(_8918_), .Y(_11452_) );
NAND3X1 NAND3X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_11450_), .B(_11451_), .C(_11452_), .Y(_11453_) );
NOR2X1 NOR2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_11449_), .B(_11453_), .Y(_11454_) );
AOI22X1 AOI22X1_228 ( .gnd(gnd), .vdd(vdd), .A(_123__6_), .B(_8928_), .C(_9__6_), .D(_8926_), .Y(_11455_) );
NAND2X1 NAND2X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__6_), .Y(_11456_) );
NAND2X1 NAND2X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_134__6_), .Y(_11457_) );
NAND3X1 NAND3X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_11456_), .B(_11457_), .C(_11455_), .Y(_11458_) );
AOI22X1 AOI22X1_229 ( .gnd(gnd), .vdd(vdd), .A(_4__6_), .B(_8937_), .C(_176__6_), .D(_8939_), .Y(_11459_) );
NAND2X1 NAND2X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__6_), .Y(_11460_) );
NAND2X1 NAND2X1_1855 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__6_), .Y(_11461_) );
NAND3X1 NAND3X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_11460_), .B(_11461_), .C(_11459_), .Y(_11462_) );
NOR2X1 NOR2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_11462_), .B(_11458_), .Y(_11463_) );
NAND2X1 NAND2X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_11454_), .B(_11463_), .Y(_11464_) );
NAND2X1 NAND2X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_9082_), .B(_250__6_), .Y(_11465_) );
NAND2X1 NAND2X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_47__6_), .Y(_11466_) );
AOI22X1 AOI22X1_230 ( .gnd(gnd), .vdd(vdd), .A(_21__6_), .B(_9150_), .C(_185__6_), .D(_9151_), .Y(_11467_) );
NAND3X1 NAND3X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_11465_), .B(_11466_), .C(_11467_), .Y(_11468_) );
AOI22X1 AOI22X1_231 ( .gnd(gnd), .vdd(vdd), .A(_246__6_), .B(_9356_), .C(_226__6_), .D(_9357_), .Y(_11469_) );
NAND2X1 NAND2X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_9157_), .B(_231__6_), .Y(_11470_) );
NAND2X1 NAND2X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_46__6_), .Y(_11471_) );
NAND3X1 NAND3X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_11470_), .B(_11471_), .C(_11469_), .Y(_11472_) );
NOR2X1 NOR2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_11468_), .B(_11472_), .Y(_11473_) );
NAND2X1 NAND2X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_178__6_), .Y(_11474_) );
NAND2X1 NAND2X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__6_), .Y(_11475_) );
AOI22X1 AOI22X1_232 ( .gnd(gnd), .vdd(vdd), .A(_37__6_), .B(_8978_), .C(_35__6_), .D(_8980_), .Y(_11476_) );
NAND3X1 NAND3X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_11474_), .B(_11475_), .C(_11476_), .Y(_11477_) );
NAND2X1 NAND2X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .B(_249__6_), .Y(_11478_) );
NAND2X1 NAND2X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_253__6_), .Y(_11479_) );
AOI22X1 AOI22X1_233 ( .gnd(gnd), .vdd(vdd), .A(_145__6_), .B(_9177_), .C(_213__6_), .D(_8989_), .Y(_11480_) );
NAND3X1 NAND3X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_11478_), .B(_11479_), .C(_11480_), .Y(_11481_) );
NOR2X1 NOR2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_11481_), .B(_11477_), .Y(_11482_) );
NAND2X1 NAND2X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_11473_), .B(_11482_), .Y(_11483_) );
NOR2X1 NOR2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_11464_), .B(_11483_), .Y(_11484_) );
NAND2X1 NAND2X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__6_), .Y(_11485_) );
NAND2X1 NAND2X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__6_), .Y(_11486_) );
AOI22X1 AOI22X1_234 ( .gnd(gnd), .vdd(vdd), .A(_13__6_), .B(_9007_), .C(_239__6_), .D(_9076_), .Y(_11487_) );
NAND3X1 NAND3X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_11485_), .B(_11486_), .C(_11487_), .Y(_11488_) );
AOI22X1 AOI22X1_235 ( .gnd(gnd), .vdd(vdd), .A(_206__6_), .B(_9013_), .C(_242__6_), .D(_9035_), .Y(_11489_) );
NAND2X1 NAND2X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__6_), .Y(_11490_) );
NAND2X1 NAND2X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__6_), .Y(_11491_) );
NAND3X1 NAND3X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_11490_), .B(_11491_), .C(_11489_), .Y(_11492_) );
NOR2X1 NOR2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_11488_), .B(_11492_), .Y(_11493_) );
AOI22X1 AOI22X1_236 ( .gnd(gnd), .vdd(vdd), .A(_222__6_), .B(_9024_), .C(_220__6_), .D(_9026_), .Y(_11494_) );
NAND2X1 NAND2X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__6_), .Y(_11495_) );
NAND2X1 NAND2X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__6_), .Y(_11496_) );
NAND3X1 NAND3X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_11495_), .B(_11496_), .C(_11494_), .Y(_11497_) );
AOI22X1 AOI22X1_237 ( .gnd(gnd), .vdd(vdd), .A(_18__6_), .B(_9037_), .C(_240__6_), .D(_9011_), .Y(_11498_) );
NAND2X1 NAND2X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__6_), .Y(_11499_) );
NAND2X1 NAND2X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__6_), .Y(_11500_) );
NAND3X1 NAND3X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_11499_), .B(_11500_), .C(_11498_), .Y(_11501_) );
NOR2X1 NOR2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_11497_), .B(_11501_), .Y(_11502_) );
NAND2X1 NAND2X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_11493_), .B(_11502_), .Y(_11503_) );
AOI22X1 AOI22X1_238 ( .gnd(gnd), .vdd(vdd), .A(_225__6_), .B(_9048_), .C(_167__6_), .D(_9050_), .Y(_11504_) );
NAND2X1 NAND2X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_243__6_), .Y(_11505_) );
NAND2X1 NAND2X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__6_), .Y(_11506_) );
NAND3X1 NAND3X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_11505_), .B(_11506_), .C(_11504_), .Y(_11507_) );
NAND2X1 NAND2X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__6_), .Y(_11508_) );
NAND2X1 NAND2X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__6_), .Y(_11509_) );
AOI22X1 AOI22X1_239 ( .gnd(gnd), .vdd(vdd), .A(_224__6_), .B(_9064_), .C(_27__6_), .D(_9066_), .Y(_11510_) );
NAND3X1 NAND3X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_11508_), .B(_11509_), .C(_11510_), .Y(_11511_) );
NOR2X1 NOR2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_11507_), .B(_11511_), .Y(_11512_) );
AOI22X1 AOI22X1_240 ( .gnd(gnd), .vdd(vdd), .A(_184__6_), .B(_9073_), .C(_183__6_), .D(_9071_), .Y(_11513_) );
NAND2X1 NAND2X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__6_), .Y(_11514_) );
NAND2X1 NAND2X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__6_), .Y(_11515_) );
NAND3X1 NAND3X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_11514_), .B(_11515_), .C(_11513_), .Y(_11516_) );
AOI22X1 AOI22X1_241 ( .gnd(gnd), .vdd(vdd), .A(_43__6_), .B(_9084_), .C(_244__6_), .D(_9160_), .Y(_11517_) );
NAND2X1 NAND2X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__6_), .Y(_11518_) );
NAND2X1 NAND2X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__6_), .Y(_11519_) );
NAND3X1 NAND3X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_11518_), .B(_11519_), .C(_11517_), .Y(_11520_) );
NOR2X1 NOR2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_11516_), .B(_11520_), .Y(_11521_) );
NAND2X1 NAND2X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_11512_), .B(_11521_), .Y(_11522_) );
NOR2X1 NOR2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_11503_), .B(_11522_), .Y(_11523_) );
NAND3X1 NAND3X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_6823_), .B(_9143_), .C(_6824_), .Y(_11524_) );
NAND3X1 NAND3X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_6971_), .B(_9145_), .C(_6972_), .Y(_11525_) );
NAND2X1 NAND2X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_11524_), .B(_11525_), .Y(_11526_) );
NAND3X1 NAND3X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_5045_), .B(_9135_), .C(_5046_), .Y(_11527_) );
NAND3X1 NAND3X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_6929_), .B(_9137_), .C(_6930_), .Y(_11528_) );
NAND2X1 NAND2X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_11528_), .B(_11527_), .Y(_11529_) );
NOR2X1 NOR2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_11526_), .B(_11529_), .Y(_11530_) );
NAND3X1 NAND3X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_8315_), .B(_9188_), .C(_8316_), .Y(_11531_) );
NAND3X1 NAND3X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_15920_), .B(_9109_), .C(_15921_), .Y(_11532_) );
NAND3X1 NAND3X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_16126_), .B(_9115_), .C(_16127_), .Y(_11533_) );
NAND3X1 NAND3X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_11532_), .B(_11533_), .C(_11531_), .Y(_11534_) );
AOI22X1 AOI22X1_242 ( .gnd(gnd), .vdd(vdd), .A(_234__6_), .B(_9182_), .C(_34__6_), .D(_9183_), .Y(_11535_) );
AOI22X1 AOI22X1_243 ( .gnd(gnd), .vdd(vdd), .A(_100__6_), .B(_9346_), .C(_45__6_), .D(_9185_), .Y(_11536_) );
NAND2X1 NAND2X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_11536_), .B(_11535_), .Y(_11537_) );
NAND3X1 NAND3X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(_9140_), .C(_4700_), .Y(_11538_) );
OAI21X1 OAI21X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_5239_), .B(_10036_), .C(_11538_), .Y(_11539_) );
NOR3X1 NOR3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_11539_), .B(_11534_), .C(_11537_), .Y(_11540_) );
NAND3X1 NAND3X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_9133_), .C(_3420_), .Y(_11541_) );
NAND3X1 NAND3X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(_9097_), .C(_4932_), .Y(_11542_) );
NAND3X1 NAND3X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .B(_9102_), .C(_5093_), .Y(_11543_) );
NAND3X1 NAND3X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_11542_), .B(_11543_), .C(_11541_), .Y(_11544_) );
AOI22X1 AOI22X1_244 ( .gnd(gnd), .vdd(vdd), .A(_38__6_), .B(_9129_), .C(_16__6_), .D(_9127_), .Y(_11545_) );
AOI22X1 AOI22X1_245 ( .gnd(gnd), .vdd(vdd), .A(_39__6_), .B(_9099_), .C(_204__6_), .D(_9104_), .Y(_11546_) );
NAND2X1 NAND2X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_11545_), .B(_11546_), .Y(_11547_) );
NOR2X1 NOR2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_11544_), .B(_11547_), .Y(_11548_) );
NAND3X1 NAND3X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_11530_), .B(_11540_), .C(_11548_), .Y(_11549_) );
AOI22X1 AOI22X1_246 ( .gnd(gnd), .vdd(vdd), .A(_227__6_), .B(_9170_), .C(_30__6_), .D(_9167_), .Y(_11550_) );
AOI22X1 AOI22X1_247 ( .gnd(gnd), .vdd(vdd), .A(_209__6_), .B(_8957_), .C(_33__6_), .D(_8991_), .Y(_11551_) );
NAND2X1 NAND2X1_1888 ( .gnd(gnd), .vdd(vdd), .A(_11550_), .B(_11551_), .Y(_11552_) );
AOI22X1 AOI22X1_248 ( .gnd(gnd), .vdd(vdd), .A(_44__6_), .B(_8968_), .C(_42__6_), .D(_8963_), .Y(_11553_) );
AOI22X1 AOI22X1_249 ( .gnd(gnd), .vdd(vdd), .A(_238__6_), .B(_8893_), .C(_208__6_), .D(_8950_), .Y(_11554_) );
NAND2X1 NAND2X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_11553_), .B(_11554_), .Y(_11555_) );
NOR2X1 NOR2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_11552_), .B(_11555_), .Y(_11556_) );
AOI22X1 AOI22X1_250 ( .gnd(gnd), .vdd(vdd), .A(_22__6_), .B(_9382_), .C(_3__6_), .D(_9383_), .Y(_11557_) );
NAND2X1 NAND2X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_219__6_), .Y(_11558_) );
NAND2X1 NAND2X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(_232__6_), .Y(_11559_) );
NAND3X1 NAND3X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_11558_), .B(_11559_), .C(_11557_), .Y(_11560_) );
AOI22X1 AOI22X1_251 ( .gnd(gnd), .vdd(vdd), .A(_255__6_), .B(_8986_), .C(_254__6_), .D(_8984_), .Y(_11561_) );
AOI22X1 AOI22X1_252 ( .gnd(gnd), .vdd(vdd), .A(_203__6_), .B(_9018_), .C(_156__6_), .D(_8973_), .Y(_11562_) );
NAND2X1 NAND2X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_11561_), .B(_11562_), .Y(_11563_) );
NOR2X1 NOR2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_11560_), .B(_11563_), .Y(_11564_) );
NAND2X1 NAND2X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_11556_), .B(_11564_), .Y(_11565_) );
AOI22X1 AOI22X1_253 ( .gnd(gnd), .vdd(vdd), .A(_201__6_), .B(_9124_), .C(_212__6_), .D(_9345_), .Y(_11566_) );
NAND3X1 NAND3X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_8429_), .B(_9348_), .C(_8428_), .Y(_11567_) );
NAND3X1 NAND3X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_489_), .C(_490_), .Y(_11568_) );
AND2X2 AND2X2_1581 ( .gnd(gnd), .vdd(vdd), .A(_11568_), .B(_11567_), .Y(_11569_) );
NAND2X1 NAND2X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_11566_), .B(_11569_), .Y(_11570_) );
NAND3X1 NAND3X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_15135_), .B(_9208_), .C(_15136_), .Y(_11571_) );
OAI21X1 OAI21X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_15100_), .B(_9211_), .C(_11571_), .Y(_11572_) );
NAND3X1 NAND3X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_15477_), .B(_9222_), .C(_15478_), .Y(_11573_) );
NAND3X1 NAND3X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_15424_), .B(_9224_), .C(_15423_), .Y(_11574_) );
NAND2X1 NAND2X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_11573_), .B(_11574_), .Y(_11575_) );
NOR2X1 NOR2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_11575_), .B(_11572_), .Y(_11576_) );
NAND3X1 NAND3X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_15255_), .B(_9217_), .C(_15256_), .Y(_11577_) );
NAND3X1 NAND3X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_15203_), .B(_9219_), .C(_15202_), .Y(_11578_) );
NAND2X1 NAND2X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_11578_), .B(_11577_), .Y(_11579_) );
NAND3X1 NAND3X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_15653_), .B(_9192_), .C(_15654_), .Y(_11580_) );
NAND3X1 NAND3X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_15710_), .B(_9199_), .C(_15709_), .Y(_11581_) );
NAND2X1 NAND2X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_11581_), .B(_11580_), .Y(_11582_) );
NOR2X1 NOR2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_11582_), .B(_11579_), .Y(_11583_) );
NOR3X1 NOR3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_16181_), .B(_10083_), .C(_16182_), .Y(_11584_) );
NAND3X1 NAND3X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_15306_), .B(_9205_), .C(_15307_), .Y(_11585_) );
OAI21X1 OAI21X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_15343_), .B(_10085_), .C(_11585_), .Y(_11586_) );
NAND3X1 NAND3X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_15535_), .B(_9233_), .C(_15536_), .Y(_11587_) );
NAND3X1 NAND3X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15604_), .C(_15603_), .Y(_11588_) );
NAND2X1 NAND2X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_11587_), .B(_11588_), .Y(_11589_) );
NOR3X1 NOR3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_11586_), .B(_11589_), .C(_11584_), .Y(_11590_) );
NAND3X1 NAND3X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_11576_), .B(_11583_), .C(_11590_), .Y(_11591_) );
NAND3X1 NAND3X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_15863_), .B(_9120_), .C(_15864_), .Y(_11592_) );
NAND3X1 NAND3X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_15376_), .B(_9197_), .C(_15377_), .Y(_11593_) );
NAND3X1 NAND3X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_7089_), .B(_9244_), .C(_7088_), .Y(_11594_) );
OAI21X1 OAI21X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_8706_), .C(_11594_), .Y(_11595_) );
AOI21X1 AOI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .B(_187__6_), .C(_11595_), .Y(_11596_) );
NAND3X1 NAND3X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_7713_), .B(_9248_), .C(_7712_), .Y(_11597_) );
OAI21X1 OAI21X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_8161_), .B(_9304_), .C(_11597_), .Y(_11598_) );
NAND3X1 NAND3X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_1762_), .B(_9255_), .C(_1763_), .Y(_11599_) );
OAI21X1 OAI21X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_4184_), .B(_9254_), .C(_11599_), .Y(_11600_) );
NOR2X1 NOR2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_11598_), .B(_11600_), .Y(_11601_) );
NAND3X1 NAND3X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_9262_), .C(_606_), .Y(_11602_) );
OAI21X1 OAI21X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_6464_), .B(_9259_), .C(_11602_), .Y(_11603_) );
NAND3X1 NAND3X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_9268_), .C(_1167_), .Y(_11604_) );
OAI21X1 OAI21X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_7044_), .B(_9267_), .C(_11604_), .Y(_11605_) );
NOR2X1 NOR2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_11603_), .B(_11605_), .Y(_11606_) );
NAND3X1 NAND3X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_11596_), .B(_11606_), .C(_11601_), .Y(_11607_) );
NOR2X1 NOR2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .B(_4812_), .Y(_11608_) );
NAND3X1 NAND3X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_9277_), .C(_2908_), .Y(_11609_) );
OAI21X1 OAI21X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_14907_), .B(_9276_), .C(_11609_), .Y(_11610_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_4218_), .B(_9282_), .C(_6426_), .D(_9763_), .Y(_11611_) );
NOR3X1 NOR3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_11608_), .B(_11610_), .C(_11611_), .Y(_11612_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .Y(_11613_) );
NAND2X1 NAND2X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__6_), .Y(_11614_) );
OAI21X1 OAI21X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_7492_), .B(_11613_), .C(_11614_), .Y(_11615_) );
NAND3X1 NAND3X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_15806_), .B(_9292_), .C(_15807_), .Y(_11616_) );
OAI21X1 OAI21X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_3599_), .B(_9295_), .C(_11616_), .Y(_11617_) );
NOR2X1 NOR2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_11615_), .B(_11617_), .Y(_11618_) );
NAND3X1 NAND3X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_8230_), .B(_9250_), .C(_8231_), .Y(_11619_) );
OAI21X1 OAI21X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_7628_), .B(_9301_), .C(_11619_), .Y(_11620_) );
NAND2X1 NAND2X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__6_), .Y(_11621_) );
OAI21X1 OAI21X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_3550_), .B(_9306_), .C(_11621_), .Y(_11622_) );
NOR2X1 NOR2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_11622_), .B(_11620_), .Y(_11623_) );
NAND3X1 NAND3X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_11612_), .B(_11618_), .C(_11623_), .Y(_11624_) );
NAND3X1 NAND3X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_5961_), .B(_9310_), .C(_5962_), .Y(_11625_) );
NAND3X1 NAND3X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_4778_), .B(_9313_), .C(_4779_), .Y(_11626_) );
NAND3X1 NAND3X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_9315_), .C(_2355_), .Y(_11627_) );
NAND3X1 NAND3X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_11626_), .B(_11627_), .C(_11625_), .Y(_11628_) );
INVX1 INVX1_3875 ( .gnd(gnd), .vdd(vdd), .A(_11628_), .Y(_11629_) );
AOI22X1 AOI22X1_254 ( .gnd(gnd), .vdd(vdd), .A(_181__6_), .B(_9321_), .C(_251__6_), .D(_9320_), .Y(_11630_) );
AOI22X1 AOI22X1_255 ( .gnd(gnd), .vdd(vdd), .A(_252__6_), .B(_9326_), .C(_235__6_), .D(_9324_), .Y(_11631_) );
NAND3X1 NAND3X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_11630_), .B(_11631_), .C(_11629_), .Y(_11632_) );
NOR3X1 NOR3X1_315 ( .gnd(gnd), .vdd(vdd), .A(_11607_), .B(_11632_), .C(_11624_), .Y(_11633_) );
NAND2X1 NAND2X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_11593_), .B(_11633_), .Y(_11634_) );
AOI21X1 AOI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_157__6_), .B(_9232_), .C(_11634_), .Y(_11635_) );
AOI22X1 AOI22X1_256 ( .gnd(gnd), .vdd(vdd), .A(_155__6_), .B(_9333_), .C(_172__6_), .D(_9332_), .Y(_11636_) );
NAND3X1 NAND3X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_11592_), .B(_11636_), .C(_11635_), .Y(_11637_) );
NOR3X1 NOR3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_11591_), .B(_11637_), .C(_11570_), .Y(_11638_) );
AOI22X1 AOI22X1_257 ( .gnd(gnd), .vdd(vdd), .A(_256__6_), .B(_9113_), .C(_142__6_), .D(_9118_), .Y(_11639_) );
NAND2X1 NAND2X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__6_), .Y(_11640_) );
NAND2X1 NAND2X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__6_), .Y(_11641_) );
NAND3X1 NAND3X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_11640_), .B(_11641_), .C(_11639_), .Y(_11642_) );
NAND2X1 NAND2X1_1904 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__6_), .Y(_11643_) );
NAND3X1 NAND3X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_9339_), .C(_446_), .Y(_11644_) );
AOI22X1 AOI22X1_258 ( .gnd(gnd), .vdd(vdd), .A(_111__6_), .B(_9342_), .C(_12__6_), .D(_9341_), .Y(_11645_) );
NAND3X1 NAND3X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_11645_), .B(_11643_), .C(_11644_), .Y(_11646_) );
NOR2X1 NOR2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_11642_), .B(_11646_), .Y(_11647_) );
AOI22X1 AOI22X1_259 ( .gnd(gnd), .vdd(vdd), .A(_40__6_), .B(_8952_), .C(_29__6_), .D(_9176_), .Y(_11648_) );
AOI22X1 AOI22X1_260 ( .gnd(gnd), .vdd(vdd), .A(_247__6_), .B(_9165_), .C(_218__6_), .D(_9169_), .Y(_11649_) );
NAND2X1 NAND2X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_11649_), .B(_11648_), .Y(_11650_) );
NAND3X1 NAND3X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16080_), .C(_16081_), .Y(_11651_) );
NAND3X1 NAND3X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16025_), .C(_16026_), .Y(_11652_) );
NAND2X1 NAND2X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_11651_), .B(_11652_), .Y(_11653_) );
NAND3X1 NAND3X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8559_), .C(_8558_), .Y(_11654_) );
OAI21X1 OAI21X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_9361_), .C(_11654_), .Y(_11655_) );
NOR2X1 NOR2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_11653_), .B(_11655_), .Y(_11656_) );
NAND2X1 NAND2X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_15972_), .B(_15973_), .Y(_11657_) );
NAND3X1 NAND3X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8612_), .C(_8613_), .Y(_11658_) );
OAI21X1 OAI21X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_11657_), .B(_9215_), .C(_11658_), .Y(_11659_) );
NAND3X1 NAND3X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_8667_), .B(_9371_), .C(_8666_), .Y(_11660_) );
NAND3X1 NAND3X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_309_), .C(_310_), .Y(_11661_) );
NAND2X1 NAND2X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_11661_), .B(_11660_), .Y(_11662_) );
NOR2X1 NOR2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_11659_), .B(_11662_), .Y(_11663_) );
AOI22X1 AOI22X1_261 ( .gnd(gnd), .vdd(vdd), .A(_248__6_), .B(_8901_), .C(_177__6_), .D(_8961_), .Y(_11664_) );
NAND3X1 NAND3X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_11656_), .B(_11663_), .C(_11664_), .Y(_11665_) );
NOR2X1 NOR2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_11650_), .B(_11665_), .Y(_11666_) );
NAND3X1 NAND3X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_11638_), .B(_11647_), .C(_11666_), .Y(_11667_) );
NOR3X1 NOR3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_11549_), .B(_11565_), .C(_11667_), .Y(_11668_) );
NAND3X1 NAND3X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_11484_), .B(_11523_), .C(_11668_), .Y(_11669_) );
NAND3X1 NAND3X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1543_), .C(_1544_), .Y(_11670_) );
NAND3X1 NAND3X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1628_), .C(_1629_), .Y(_11671_) );
NAND2X1 NAND2X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_11670_), .B(_11671_), .Y(_11672_) );
NOR3X1 NOR3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_11446_), .B(_11672_), .C(_11669_), .Y(_11673_) );
NAND3X1 NAND3X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_11428_), .B(_11435_), .C(_11673_), .Y(_11674_) );
NAND2X1 NAND2X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__6_), .Y(_11675_) );
AOI22X1 AOI22X1_262 ( .gnd(gnd), .vdd(vdd), .A(_115__6_), .B(_9399_), .C(_116__6_), .D(_9401_), .Y(_11676_) );
AOI22X1 AOI22X1_263 ( .gnd(gnd), .vdd(vdd), .A(_108__6_), .B(_9404_), .C(_109__6_), .D(_9406_), .Y(_11677_) );
NAND2X1 NAND2X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_11676_), .B(_11677_), .Y(_11678_) );
NAND2X1 NAND2X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_125__6_), .Y(_11679_) );
NAND2X1 NAND2X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_122__6_), .Y(_11680_) );
NAND2X1 NAND2X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_11679_), .B(_11680_), .Y(_11681_) );
NOR2X1 NOR2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_1101_), .Y(_11682_) );
AND2X2 AND2X2_1582 ( .gnd(gnd), .vdd(vdd), .A(_120__6_), .B(_9415_), .Y(_11683_) );
NOR3X1 NOR3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_11682_), .B(_11683_), .C(_11681_), .Y(_11684_) );
AOI22X1 AOI22X1_264 ( .gnd(gnd), .vdd(vdd), .A(_132__6_), .B(_9420_), .C(_131__6_), .D(_9418_), .Y(_11685_) );
NAND2X1 NAND2X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__6_), .Y(_11686_) );
NAND2X1 NAND2X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__6_), .Y(_11687_) );
NAND3X1 NAND3X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_11686_), .B(_11687_), .C(_11685_), .Y(_11688_) );
NAND3X1 NAND3X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_9431_), .C(_539_), .Y(_11689_) );
NAND2X1 NAND2X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__6_), .Y(_11690_) );
NAND2X1 NAND2X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__6_), .Y(_11691_) );
NAND3X1 NAND3X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_11691_), .B(_11689_), .C(_11690_), .Y(_11692_) );
AOI21X1 AOI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__6_), .C(_11692_), .Y(_11693_) );
NAND2X1 NAND2X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__6_), .Y(_11694_) );
NAND2X1 NAND2X1_1920 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_136__6_), .Y(_11695_) );
NAND3X1 NAND3X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_11694_), .B(_11695_), .C(_11693_), .Y(_11696_) );
NAND3X1 NAND3X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_9410_), .C(_1009_), .Y(_11697_) );
NAND2X1 NAND2X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__6_), .Y(_11698_) );
AOI22X1 AOI22X1_265 ( .gnd(gnd), .vdd(vdd), .A(_130__6_), .B(_9449_), .C(_127__6_), .D(_9448_), .Y(_11699_) );
NAND3X1 NAND3X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_11697_), .B(_11699_), .C(_11698_), .Y(_11700_) );
NOR3X1 NOR3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_11688_), .B(_11696_), .C(_11700_), .Y(_11701_) );
AOI22X1 AOI22X1_266 ( .gnd(gnd), .vdd(vdd), .A(_110__6_), .B(_9453_), .C(_114__6_), .D(_9454_), .Y(_11702_) );
NAND3X1 NAND3X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_11684_), .B(_11702_), .C(_11701_), .Y(_11703_) );
NOR2X1 NOR2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_11678_), .B(_11703_), .Y(_11704_) );
AOI22X1 AOI22X1_267 ( .gnd(gnd), .vdd(vdd), .A(_102__6_), .B(_9459_), .C(_103__6_), .D(_9457_), .Y(_11705_) );
NAND3X1 NAND3X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_11675_), .B(_11705_), .C(_11704_), .Y(_11706_) );
NOR3X1 NOR3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_11427_), .B(_11706_), .C(_11674_), .Y(_11707_) );
NAND3X1 NAND3X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_11417_), .B(_11424_), .C(_11707_), .Y(_11708_) );
NOR3X1 NOR3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_11406_), .B(_11409_), .C(_11708_), .Y(_11709_) );
NAND3X1 NAND3X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_11397_), .B(_11402_), .C(_11709_), .Y(_11710_) );
NAND3X1 NAND3X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(_9473_), .C(_3059_), .Y(_11711_) );
NAND2X1 NAND2X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__6_), .Y(_11712_) );
NAND2X1 NAND2X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__6_), .Y(_11713_) );
NAND2X1 NAND2X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__6_), .Y(_11714_) );
NAND3X1 NAND3X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_2436_), .B(_9468_), .C(_2437_), .Y(_11715_) );
NAND3X1 NAND3X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_11715_), .B(_11713_), .C(_11714_), .Y(_11716_) );
AOI21X1 AOI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_68__6_), .B(_9477_), .C(_11716_), .Y(_11717_) );
NAND3X1 NAND3X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_11717_), .B(_11711_), .C(_11712_), .Y(_11718_) );
NOR3X1 NOR3X1_323 ( .gnd(gnd), .vdd(vdd), .A(_11396_), .B(_11718_), .C(_11710_), .Y(_11719_) );
AOI21X1 AOI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_11391_), .B(_11719_), .C(rst), .Y(_0__6_) );
NAND2X1 NAND2X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__7_), .Y(_11720_) );
NAND2X1 NAND2X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__7_), .Y(_11721_) );
NAND2X1 NAND2X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_11720_), .B(_11721_), .Y(_11722_) );
NAND2X1 NAND2X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__7_), .Y(_11723_) );
NAND2X1 NAND2X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__7_), .Y(_11724_) );
NAND2X1 NAND2X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_11723_), .B(_11724_), .Y(_11725_) );
NOR2X1 NOR2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_11722_), .B(_11725_), .Y(_11726_) );
NAND3X1 NAND3X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(_8762_), .C(_3277_), .Y(_11727_) );
NAND3X1 NAND3X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(_8765_), .C(_3231_), .Y(_11728_) );
AND2X2 AND2X2_1583 ( .gnd(gnd), .vdd(vdd), .A(_11728_), .B(_11727_), .Y(_11729_) );
AOI22X1 AOI22X1_268 ( .gnd(gnd), .vdd(vdd), .A(_62__7_), .B(_8774_), .C(_57__7_), .D(_8771_), .Y(_11730_) );
NAND2X1 NAND2X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_11729_), .B(_11730_), .Y(_11731_) );
NAND2X1 NAND2X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__7_), .Y(_11732_) );
NAND3X1 NAND3X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(_8794_), .C(_2645_), .Y(_11733_) );
OAI21X1 OAI21X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_2706_), .B(_8792_), .C(_11733_), .Y(_11734_) );
NAND3X1 NAND3X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_2815_), .B(_8786_), .C(_2816_), .Y(_11735_) );
OAI21X1 OAI21X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_8799_), .C(_11735_), .Y(_11736_) );
NOR2X1 NOR2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_11734_), .B(_11736_), .Y(_11737_) );
AOI22X1 AOI22X1_269 ( .gnd(gnd), .vdd(vdd), .A(_73__7_), .B(_9480_), .C(_74__7_), .D(_8803_), .Y(_11738_) );
AOI22X1 AOI22X1_270 ( .gnd(gnd), .vdd(vdd), .A(_76__7_), .B(_9482_), .C(_81__7_), .D(_9468_), .Y(_11739_) );
NAND2X1 NAND2X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_11739_), .B(_11738_), .Y(_11740_) );
INVX1 INVX1_3876 ( .gnd(gnd), .vdd(vdd), .A(_84__7_), .Y(_11741_) );
NOR2X1 NOR2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_11741_), .Y(_11742_) );
NOR2X1 NOR2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2296_), .Y(_11743_) );
NAND2X1 NAND2X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__7_), .Y(_11744_) );
NAND3X1 NAND3X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_8843_), .C(_2010_), .Y(_11745_) );
NAND3X1 NAND3X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1913_), .C(_1914_), .Y(_11746_) );
NAND3X1 NAND3X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_11746_), .B(_11745_), .C(_11744_), .Y(_11747_) );
NOR3X1 NOR3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_11742_), .B(_11747_), .C(_11743_), .Y(_11748_) );
NAND3X1 NAND3X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_2251_), .B(_8829_), .C(_2252_), .Y(_11749_) );
NAND3X1 NAND3X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(_8831_), .C(_2146_), .Y(_11750_) );
NAND2X1 NAND2X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_11749_), .B(_11750_), .Y(_11751_) );
NAND3X1 NAND3X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_8834_), .C(_2087_), .Y(_11752_) );
NAND3X1 NAND3X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_2197_), .B(_8836_), .C(_2198_), .Y(_11753_) );
NAND2X1 NAND2X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_11752_), .B(_11753_), .Y(_11754_) );
NOR2X1 NOR2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_11754_), .B(_11751_), .Y(_11755_) );
AOI22X1 AOI22X1_271 ( .gnd(gnd), .vdd(vdd), .A(_98__7_), .B(_8845_), .C(_93__7_), .D(_8840_), .Y(_11756_) );
NAND2X1 NAND2X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_8823_), .B(_91__7_), .Y(_11757_) );
NAND2X1 NAND2X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_94__7_), .Y(_11758_) );
NAND3X1 NAND3X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_11757_), .B(_11758_), .C(_11756_), .Y(_11759_) );
NAND2X1 NAND2X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__7_), .Y(_11760_) );
NAND3X1 NAND3X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1546_), .C(_1547_), .Y(_11761_) );
NAND3X1 NAND3X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1631_), .C(_1632_), .Y(_11762_) );
NAND2X1 NAND2X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_11761_), .B(_11762_), .Y(_11763_) );
NAND3X1 NAND3X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1669_), .C(_1670_), .Y(_11764_) );
NAND3X1 NAND3X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .B(_8857_), .C(_1378_), .Y(_11765_) );
NAND2X1 NAND2X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_11765_), .B(_11764_), .Y(_11766_) );
OR2X2 OR2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_11763_), .B(_11766_), .Y(_11767_) );
NOR3X1 NOR3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_8867_), .C(_1212_), .Y(_11768_) );
AOI22X1 AOI22X1_272 ( .gnd(gnd), .vdd(vdd), .A(_191__7_), .B(_8873_), .C(_192__7_), .D(_8872_), .Y(_11769_) );
AOI22X1 AOI22X1_273 ( .gnd(gnd), .vdd(vdd), .A(_195__7_), .B(_8875_), .C(_193__7_), .D(_8876_), .Y(_11770_) );
NAND2X1 NAND2X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_11769_), .B(_11770_), .Y(_11771_) );
AOI22X1 AOI22X1_274 ( .gnd(gnd), .vdd(vdd), .A(_188__7_), .B(_8879_), .C(_126__7_), .D(_8881_), .Y(_11772_) );
AOI22X1 AOI22X1_275 ( .gnd(gnd), .vdd(vdd), .A(_196__7_), .B(_8883_), .C(_194__7_), .D(_8884_), .Y(_11773_) );
NAND2X1 NAND2X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_11772_), .B(_11773_), .Y(_11774_) );
NOR3X1 NOR3X1_326 ( .gnd(gnd), .vdd(vdd), .A(_11774_), .B(_11768_), .C(_11771_), .Y(_11775_) );
NAND3X1 NAND3X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_5638_), .B(_9153_), .C(_5637_), .Y(_11776_) );
NAND3X1 NAND3X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_4590_), .B(_8898_), .C(_4589_), .Y(_11777_) );
NAND2X1 NAND2X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_11776_), .B(_11777_), .Y(_11778_) );
NAND3X1 NAND3X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_5610_), .B(_9160_), .C(_5609_), .Y(_11779_) );
NAND3X1 NAND3X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_7865_), .B(_8904_), .C(_7864_), .Y(_11780_) );
NAND2X1 NAND2X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_11779_), .B(_11780_), .Y(_11781_) );
NOR2X1 NOR2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_11778_), .B(_11781_), .Y(_11782_) );
NAND3X1 NAND3X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_3478_), .B(_8975_), .C(_3477_), .Y(_11783_) );
NAND3X1 NAND3X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3892_), .C(_3891_), .Y(_11784_) );
NAND2X1 NAND2X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_11783_), .B(_11784_), .Y(_11785_) );
NAND3X1 NAND3X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_8914_), .C(_4630_), .Y(_11786_) );
NAND3X1 NAND3X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_6652_), .B(_8918_), .C(_6651_), .Y(_11787_) );
NAND2X1 NAND2X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_11786_), .B(_11787_), .Y(_11788_) );
NOR2X1 NOR2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_11785_), .B(_11788_), .Y(_11789_) );
NAND2X1 NAND2X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_11782_), .B(_11789_), .Y(_11790_) );
NAND3X1 NAND3X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_4971_), .B(_8926_), .C(_4970_), .Y(_11791_) );
NAND3X1 NAND3X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_8071_), .B(_8928_), .C(_8070_), .Y(_11792_) );
NAND2X1 NAND2X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_11791_), .B(_11792_), .Y(_11793_) );
NAND3X1 NAND3X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_4493_), .B(_8931_), .C(_4492_), .Y(_11794_) );
NAND3X1 NAND3X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_8039_), .B(_8933_), .C(_8038_), .Y(_11795_) );
NAND2X1 NAND2X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_11794_), .B(_11795_), .Y(_11796_) );
NOR2X1 NOR2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_11793_), .B(_11796_), .Y(_11797_) );
NAND3X1 NAND3X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_5185_), .B(_8937_), .C(_5184_), .Y(_11798_) );
NAND3X1 NAND3X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_7827_), .B(_8939_), .C(_7826_), .Y(_11799_) );
NAND2X1 NAND2X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_11798_), .B(_11799_), .Y(_11800_) );
NAND3X1 NAND3X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_5147_), .B(_8942_), .C(_5146_), .Y(_11801_) );
NAND3X1 NAND3X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_5009_), .B(_8944_), .C(_5008_), .Y(_11802_) );
NAND2X1 NAND2X1_1952 ( .gnd(gnd), .vdd(vdd), .A(_11801_), .B(_11802_), .Y(_11803_) );
NOR2X1 NOR2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_11803_), .B(_11800_), .Y(_11804_) );
NAND2X1 NAND2X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_11797_), .B(_11804_), .Y(_11805_) );
NOR2X1 NOR2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_11790_), .B(_11805_), .Y(_11806_) );
NAND3X1 NAND3X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_5527_), .B(_8901_), .C(_5526_), .Y(_11807_) );
NAND3X1 NAND3X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_3701_), .B(_9161_), .C(_3700_), .Y(_11808_) );
NAND2X1 NAND2X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_11807_), .B(_11808_), .Y(_11809_) );
NAND3X1 NAND3X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_4552_), .B(_9150_), .C(_4551_), .Y(_11810_) );
NAND3X1 NAND3X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_7525_), .B(_9151_), .C(_7524_), .Y(_11811_) );
NAND2X1 NAND2X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_11810_), .B(_11811_), .Y(_11812_) );
NOR2X1 NOR2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_11809_), .B(_11812_), .Y(_11813_) );
NAND3X1 NAND3X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_5582_), .B(_9356_), .C(_5581_), .Y(_11814_) );
NAND3X1 NAND3X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_6165_), .B(_9357_), .C(_6164_), .Y(_11815_) );
NAND2X1 NAND2X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_11814_), .B(_11815_), .Y(_11816_) );
NAND3X1 NAND3X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_6020_), .B(_9157_), .C(_6019_), .Y(_11817_) );
NAND3X1 NAND3X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .B(_9158_), .C(_3734_), .Y(_11818_) );
NAND2X1 NAND2X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_11818_), .B(_11817_), .Y(_11819_) );
NOR2X1 NOR2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_11816_), .B(_11819_), .Y(_11820_) );
NAND2X1 NAND2X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_11813_), .B(_11820_), .Y(_11821_) );
NAND3X1 NAND3X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_7759_), .B(_9173_), .C(_7758_), .Y(_11822_) );
NAND3X1 NAND3X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_9084_), .C(_3812_), .Y(_11823_) );
NAND2X1 NAND2X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_11822_), .B(_11823_), .Y(_11824_) );
NAND3X1 NAND3X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_5830_), .B(_8893_), .C(_5829_), .Y(_11825_) );
NAND3X1 NAND3X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_3666_), .B(_9089_), .C(_3665_), .Y(_11826_) );
NAND2X1 NAND2X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_11825_), .B(_11826_), .Y(_11827_) );
NOR2X1 NOR2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_11824_), .B(_11827_), .Y(_11828_) );
NAND3X1 NAND3X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_5900_), .B(_8955_), .C(_5899_), .Y(_11829_) );
NAND3X1 NAND3X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_5342_), .B(_9154_), .C(_5341_), .Y(_11830_) );
NAND2X1 NAND2X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_11829_), .B(_11830_), .Y(_11831_) );
NAND3X1 NAND3X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_8001_), .B(_9177_), .C(_8000_), .Y(_11832_) );
NAND3X1 NAND3X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_6575_), .B(_8989_), .C(_6574_), .Y(_11833_) );
NAND2X1 NAND2X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_11833_), .B(_11832_), .Y(_11834_) );
NOR2X1 NOR2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_11831_), .B(_11834_), .Y(_11835_) );
NAND2X1 NAND2X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_11828_), .B(_11835_), .Y(_11836_) );
NOR2X1 NOR2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_11821_), .B(_11836_), .Y(_11837_) );
NAND2X1 NAND2X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_11806_), .B(_11837_), .Y(_11838_) );
NAND3X1 NAND3X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_4902_), .B(_8998_), .C(_4901_), .Y(_11839_) );
NAND3X1 NAND3X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_6509_), .B(_9002_), .C(_6508_), .Y(_11840_) );
NAND2X1 NAND2X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_11839_), .B(_11840_), .Y(_11841_) );
NAND3X1 NAND3X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_5715_), .B(_9005_), .C(_5714_), .Y(_11842_) );
NAND3X1 NAND3X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_4863_), .B(_9007_), .C(_4862_), .Y(_11843_) );
NAND2X1 NAND2X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_11842_), .B(_11843_), .Y(_11844_) );
NOR2X1 NOR2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_11841_), .B(_11844_), .Y(_11845_) );
NAND3X1 NAND3X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_5753_), .B(_9011_), .C(_5752_), .Y(_11846_) );
NAND3X1 NAND3X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_6795_), .B(_9013_), .C(_6794_), .Y(_11847_) );
NAND2X1 NAND2X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_11846_), .B(_11847_), .Y(_11848_) );
NAND3X1 NAND3X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_6756_), .B(_9016_), .C(_6755_), .Y(_11849_) );
NAND3X1 NAND3X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_6542_), .B(_9174_), .C(_6541_), .Y(_11850_) );
NAND2X1 NAND2X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_11849_), .B(_11850_), .Y(_11851_) );
NOR2X1 NOR2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_11851_), .B(_11848_), .Y(_11852_) );
NAND2X1 NAND2X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_11845_), .B(_11852_), .Y(_11853_) );
NAND3X1 NAND3X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_6279_), .B(_9024_), .C(_6278_), .Y(_11854_) );
NAND3X1 NAND3X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_6351_), .B(_9026_), .C(_6350_), .Y(_11855_) );
NAND2X1 NAND2X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_11854_), .B(_11855_), .Y(_11856_) );
NAND3X1 NAND3X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_6056_), .B(_9029_), .C(_6055_), .Y(_11857_) );
NAND3X1 NAND3X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_6114_), .B(_9031_), .C(_6113_), .Y(_11858_) );
NAND2X1 NAND2X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_11857_), .B(_11858_), .Y(_11859_) );
NOR2X1 NOR2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_11856_), .B(_11859_), .Y(_11860_) );
NAND3X1 NAND3X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_5674_), .B(_9035_), .C(_5673_), .Y(_11861_) );
NAND3X1 NAND3X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_4670_), .B(_9037_), .C(_4669_), .Y(_11862_) );
NAND2X1 NAND2X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_11862_), .B(_11861_), .Y(_11863_) );
NAND3X1 NAND3X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_6315_), .B(_9040_), .C(_6314_), .Y(_11864_) );
NAND3X1 NAND3X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_9042_), .C(_4331_), .Y(_11865_) );
NAND2X1 NAND2X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_11864_), .B(_11865_), .Y(_11866_) );
NOR2X1 NOR2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_11866_), .B(_11863_), .Y(_11867_) );
NAND2X1 NAND2X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_11860_), .B(_11867_), .Y(_11868_) );
NOR2X1 NOR2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_11853_), .B(_11868_), .Y(_11869_) );
NAND3X1 NAND3X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_6203_), .B(_9048_), .C(_6202_), .Y(_11870_) );
NAND3X1 NAND3X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_7938_), .B(_9050_), .C(_7937_), .Y(_11871_) );
NAND2X1 NAND2X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_11870_), .B(_11871_), .Y(_11872_) );
NAND3X1 NAND3X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_7901_), .B(_9055_), .C(_7900_), .Y(_11873_) );
NAND3X1 NAND3X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_4127_), .B(_8980_), .C(_4126_), .Y(_11874_) );
NAND2X1 NAND2X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_11873_), .B(_11874_), .Y(_11875_) );
NOR2X1 NOR2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_11872_), .B(_11875_), .Y(_11876_) );
NAND3X1 NAND3X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_4453_), .B(_9059_), .C(_4452_), .Y(_11877_) );
NAND3X1 NAND3X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_4413_), .B(_9061_), .C(_4412_), .Y(_11878_) );
NAND2X1 NAND2X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_11877_), .B(_11878_), .Y(_11879_) );
NAND3X1 NAND3X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_6241_), .B(_9064_), .C(_6240_), .Y(_11880_) );
NAND3X1 NAND3X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_4373_), .B(_9066_), .C(_4372_), .Y(_11881_) );
NAND2X1 NAND2X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_11880_), .B(_11881_), .Y(_11882_) );
NOR2X1 NOR2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_11882_), .B(_11879_), .Y(_11883_) );
NAND2X1 NAND2X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_11876_), .B(_11883_), .Y(_11884_) );
NAND3X1 NAND3X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_7597_), .B(_9071_), .C(_7596_), .Y(_11885_) );
NAND3X1 NAND3X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_7561_), .B(_9073_), .C(_7560_), .Y(_11886_) );
NAND2X1 NAND2X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_11885_), .B(_11886_), .Y(_11887_) );
NAND3X1 NAND3X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_5791_), .B(_9076_), .C(_5790_), .Y(_11888_) );
NAND3X1 NAND3X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_3517_), .B(_9078_), .C(_3516_), .Y(_11889_) );
NAND2X1 NAND2X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_11888_), .B(_11889_), .Y(_11890_) );
NOR2X1 NOR2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_11887_), .B(_11890_), .Y(_11891_) );
NAND3X1 NAND3X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_5867_), .B(_8966_), .C(_5866_), .Y(_11892_) );
NAND3X1 NAND3X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_4090_), .B(_8909_), .C(_4089_), .Y(_11893_) );
NAND2X1 NAND2X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_11892_), .B(_11893_), .Y(_11894_) );
NAND3X1 NAND3X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_6612_), .B(_9087_), .C(_6611_), .Y(_11895_) );
NAND3X1 NAND3X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_4053_), .B(_8978_), .C(_4052_), .Y(_11896_) );
NAND2X1 NAND2X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_11895_), .B(_11896_), .Y(_11897_) );
NOR2X1 NOR2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_11894_), .B(_11897_), .Y(_11898_) );
NAND2X1 NAND2X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_11891_), .B(_11898_), .Y(_11899_) );
NOR2X1 NOR2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_11884_), .B(_11899_), .Y(_11900_) );
NAND2X1 NAND2X1_1985 ( .gnd(gnd), .vdd(vdd), .A(_11869_), .B(_11900_), .Y(_11901_) );
NOR2X1 NOR2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_11838_), .B(_11901_), .Y(_11902_) );
NAND2X1 NAND2X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__7_), .Y(_11903_) );
NAND3X1 NAND3X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_6974_), .B(_9145_), .C(_6973_), .Y(_11904_) );
NAND2X1 NAND2X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_11903_), .B(_11904_), .Y(_11905_) );
NAND3X1 NAND3X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_5048_), .B(_9135_), .C(_5049_), .Y(_11906_) );
NAND3X1 NAND3X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_6932_), .B(_9137_), .C(_6931_), .Y(_11907_) );
NAND2X1 NAND2X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_11906_), .B(_11907_), .Y(_11908_) );
NOR2X1 NOR2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_11908_), .B(_11905_), .Y(_11909_) );
NAND3X1 NAND3X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_16129_), .B(_9115_), .C(_16130_), .Y(_11910_) );
NAND3X1 NAND3X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_8388_), .B(_9113_), .C(_8389_), .Y(_11911_) );
NAND3X1 NAND3X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_15923_), .B(_9109_), .C(_15924_), .Y(_11912_) );
NAND3X1 NAND3X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_11910_), .B(_11912_), .C(_11911_), .Y(_11913_) );
NAND3X1 NAND3X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_394_), .C(_395_), .Y(_11914_) );
NAND3X1 NAND3X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_15866_), .B(_9120_), .C(_15867_), .Y(_11915_) );
AND2X2 AND2X2_1584 ( .gnd(gnd), .vdd(vdd), .A(_11915_), .B(_11914_), .Y(_11916_) );
AOI22X1 AOI22X1_276 ( .gnd(gnd), .vdd(vdd), .A(_201__7_), .B(_9124_), .C(_89__7_), .D(_9123_), .Y(_11917_) );
NAND2X1 NAND2X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_11916_), .B(_11917_), .Y(_11918_) );
NAND3X1 NAND3X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_4703_), .B(_9140_), .C(_4704_), .Y(_11919_) );
OAI21X1 OAI21X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_5242_), .B(_10036_), .C(_11919_), .Y(_11920_) );
NOR3X1 NOR3X1_327 ( .gnd(gnd), .vdd(vdd), .A(_11913_), .B(_11920_), .C(_11918_), .Y(_11921_) );
NAND3X1 NAND3X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3422_), .C(_3423_), .Y(_11922_) );
NAND2X1 NAND2X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__7_), .Y(_11923_) );
NAND3X1 NAND3X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_9102_), .C(_5096_), .Y(_11924_) );
NAND3X1 NAND3X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_11922_), .B(_11924_), .C(_11923_), .Y(_11925_) );
AOI22X1 AOI22X1_277 ( .gnd(gnd), .vdd(vdd), .A(_38__7_), .B(_9129_), .C(_16__7_), .D(_9127_), .Y(_11926_) );
NAND2X1 NAND2X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_9104_), .B(_204__7_), .Y(_11927_) );
NAND2X1 NAND2X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_9099_), .B(_39__7_), .Y(_11928_) );
NAND3X1 NAND3X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_11928_), .B(_11927_), .C(_11926_), .Y(_11929_) );
NOR2X1 NOR2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_11925_), .B(_11929_), .Y(_11930_) );
NAND3X1 NAND3X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_11909_), .B(_11930_), .C(_11921_), .Y(_11931_) );
AOI22X1 AOI22X1_278 ( .gnd(gnd), .vdd(vdd), .A(_30__7_), .B(_9167_), .C(_227__7_), .D(_9170_), .Y(_11932_) );
AOI22X1 AOI22X1_279 ( .gnd(gnd), .vdd(vdd), .A(_209__7_), .B(_8957_), .C(_33__7_), .D(_8991_), .Y(_11933_) );
NAND2X1 NAND2X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_11932_), .B(_11933_), .Y(_11934_) );
AOI22X1 AOI22X1_280 ( .gnd(gnd), .vdd(vdd), .A(_44__7_), .B(_8968_), .C(_42__7_), .D(_8963_), .Y(_11935_) );
AOI22X1 AOI22X1_281 ( .gnd(gnd), .vdd(vdd), .A(_249__7_), .B(_9053_), .C(_208__7_), .D(_8950_), .Y(_11936_) );
NAND2X1 NAND2X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_11935_), .B(_11936_), .Y(_11937_) );
NOR2X1 NOR2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_11934_), .B(_11937_), .Y(_11938_) );
AOI22X1 AOI22X1_282 ( .gnd(gnd), .vdd(vdd), .A(_22__7_), .B(_9382_), .C(_3__7_), .D(_9383_), .Y(_11939_) );
AOI22X1 AOI22X1_283 ( .gnd(gnd), .vdd(vdd), .A(_232__7_), .B(_9354_), .C(_219__7_), .D(_9353_), .Y(_11940_) );
NAND2X1 NAND2X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_11939_), .B(_11940_), .Y(_11941_) );
AOI22X1 AOI22X1_284 ( .gnd(gnd), .vdd(vdd), .A(_255__7_), .B(_8986_), .C(_254__7_), .D(_8984_), .Y(_11942_) );
AOI22X1 AOI22X1_285 ( .gnd(gnd), .vdd(vdd), .A(_203__7_), .B(_9018_), .C(_156__7_), .D(_8973_), .Y(_11943_) );
NAND2X1 NAND2X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_11943_), .B(_11942_), .Y(_11944_) );
NOR2X1 NOR2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_11941_), .B(_11944_), .Y(_11945_) );
NAND2X1 NAND2X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_11938_), .B(_11945_), .Y(_11946_) );
AOI22X1 AOI22X1_286 ( .gnd(gnd), .vdd(vdd), .A(_234__7_), .B(_9182_), .C(_34__7_), .D(_9183_), .Y(_11947_) );
NAND2X1 NAND2X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__7_), .Y(_11948_) );
NAND2X1 NAND2X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__7_), .Y(_11949_) );
NAND3X1 NAND3X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_11948_), .B(_11949_), .C(_11947_), .Y(_11950_) );
NAND3X1 NAND3X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_15656_), .B(_9192_), .C(_15657_), .Y(_11951_) );
OAI21X1 OAI21X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_15606_), .B(_9195_), .C(_11951_), .Y(_11952_) );
NAND2X1 NAND2X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__7_), .Y(_11953_) );
NAND3X1 NAND3X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_15712_), .B(_9199_), .C(_15713_), .Y(_11954_) );
NAND2X1 NAND2X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_11953_), .B(_11954_), .Y(_11955_) );
NOR2X1 NOR2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_11955_), .B(_11952_), .Y(_11956_) );
NAND2X1 NAND2X1_2002 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__7_), .Y(_11957_) );
OAI21X1 OAI21X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_15309_), .B(_9206_), .C(_11957_), .Y(_11958_) );
NAND2X1 NAND2X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__7_), .Y(_11959_) );
OAI21X1 OAI21X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_15102_), .B(_9211_), .C(_11959_), .Y(_11960_) );
NOR2X1 NOR2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_11958_), .B(_11960_), .Y(_11961_) );
NOR3X1 NOR3X1_328 ( .gnd(gnd), .vdd(vdd), .A(_15974_), .B(_9215_), .C(_15975_), .Y(_11962_) );
NAND3X1 NAND3X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_15258_), .B(_9217_), .C(_15259_), .Y(_11963_) );
NAND3X1 NAND3X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_15206_), .B(_9219_), .C(_15205_), .Y(_11964_) );
NAND2X1 NAND2X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_11964_), .B(_11963_), .Y(_11965_) );
NAND3X1 NAND3X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_15480_), .B(_9222_), .C(_15481_), .Y(_11966_) );
NAND3X1 NAND3X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_15427_), .B(_9224_), .C(_15426_), .Y(_11967_) );
NAND2X1 NAND2X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_11966_), .B(_11967_), .Y(_11968_) );
NOR3X1 NOR3X1_329 ( .gnd(gnd), .vdd(vdd), .A(_11962_), .B(_11968_), .C(_11965_), .Y(_11969_) );
NAND3X1 NAND3X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_11961_), .B(_11969_), .C(_11956_), .Y(_11970_) );
NAND2X1 NAND2X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__7_), .Y(_11971_) );
NAND3X1 NAND3X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_15538_), .B(_9233_), .C(_15539_), .Y(_11972_) );
NOR2X1 NOR2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_10471_), .B(_7468_), .Y(_11973_) );
AND2X2 AND2X2_1585 ( .gnd(gnd), .vdd(vdd), .A(_186__7_), .B(_9298_), .Y(_11974_) );
NOR2X1 NOR2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_11974_), .B(_11973_), .Y(_11975_) );
OAI21X1 OAI21X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_7007_), .B(_9288_), .C(_11975_), .Y(_11976_) );
NAND2X1 NAND2X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__7_), .Y(_11977_) );
OAI21X1 OAI21X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_8234_), .B(_10875_), .C(_11977_), .Y(_11978_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_7047_), .B(_9267_), .C(_7092_), .D(_9245_), .Y(_11979_) );
NOR2X1 NOR2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_11979_), .B(_11978_), .Y(_11980_) );
NAND3X1 NAND3X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_7715_), .B(_9248_), .C(_7716_), .Y(_11981_) );
OAI21X1 OAI21X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_9306_), .C(_11981_), .Y(_11982_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_8164_), .B(_9304_), .C(_7631_), .D(_9301_), .Y(_11983_) );
NOR2X1 NOR2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_11983_), .B(_11982_), .Y(_11984_) );
NAND2X1 NAND2X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_11980_), .B(_11984_), .Y(_11985_) );
NOR2X1 NOR2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_11976_), .B(_11985_), .Y(_11986_) );
NOR2X1 NOR2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_9763_), .B(_6429_), .Y(_11987_) );
NAND3X1 NAND3X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_9262_), .C(_609_), .Y(_11988_) );
OAI21X1 OAI21X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_10468_), .C(_11988_), .Y(_11989_) );
NAND3X1 NAND3X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_2357_), .B(_9315_), .C(_2358_), .Y(_11990_) );
OAI21X1 OAI21X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_5400_), .B(_9319_), .C(_11990_), .Y(_11991_) );
NOR3X1 NOR3X1_330 ( .gnd(gnd), .vdd(vdd), .A(_11989_), .B(_11987_), .C(_11991_), .Y(_11992_) );
NAND2X1 NAND2X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_1__7_), .B(_9242_), .Y(_11993_) );
NAND2X1 NAND2X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_101__7_), .Y(_11994_) );
NAND2X1 NAND2X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_11993_), .B(_11994_), .Y(_11995_) );
NAND2X1 NAND2X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_9292_), .B(_154__7_), .Y(_11996_) );
OAI21X1 OAI21X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_4186_), .B(_9254_), .C(_11996_), .Y(_11997_) );
NOR2X1 NOR2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_11995_), .B(_11997_), .Y(_11998_) );
NAND2X1 NAND2X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__7_), .Y(_11999_) );
OAI21X1 OAI21X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .B(_9295_), .C(_11999_), .Y(_12000_) );
NAND2X1 NAND2X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_9268_), .B(_119__7_), .Y(_12001_) );
NAND2X1 NAND2X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_173__7_), .Y(_12002_) );
NAND2X1 NAND2X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_12001_), .B(_12002_), .Y(_12003_) );
NOR2X1 NOR2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_12000_), .B(_12003_), .Y(_12004_) );
NAND3X1 NAND3X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_11992_), .B(_11998_), .C(_12004_), .Y(_12005_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4219_), .B(_9282_), .C(_4780_), .D(_9312_), .Y(_12006_) );
AOI21X1 AOI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_9324_), .B(_235__7_), .C(_12006_), .Y(_12007_) );
AOI22X1 AOI22X1_287 ( .gnd(gnd), .vdd(vdd), .A(_181__7_), .B(_9321_), .C(_252__7_), .D(_9326_), .Y(_12008_) );
AOI22X1 AOI22X1_288 ( .gnd(gnd), .vdd(vdd), .A(_14__7_), .B(_9274_), .C(_233__7_), .D(_9310_), .Y(_12009_) );
NAND3X1 NAND3X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_12007_), .B(_12009_), .C(_12008_), .Y(_12010_) );
NOR2X1 NOR2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_12010_), .B(_12005_), .Y(_12011_) );
NAND3X1 NAND3X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_11972_), .B(_11986_), .C(_12011_), .Y(_12012_) );
AOI21X1 AOI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_157__7_), .B(_9232_), .C(_12012_), .Y(_12013_) );
AOI22X1 AOI22X1_289 ( .gnd(gnd), .vdd(vdd), .A(_155__7_), .B(_9333_), .C(_172__7_), .D(_9332_), .Y(_12014_) );
NAND3X1 NAND3X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_12014_), .B(_12013_), .C(_11971_), .Y(_12015_) );
NOR3X1 NOR3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_11950_), .B(_12015_), .C(_11970_), .Y(_12016_) );
NAND2X1 NAND2X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__7_), .Y(_12017_) );
NAND3X1 NAND3X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_9339_), .C(_449_), .Y(_12018_) );
AOI22X1 AOI22X1_290 ( .gnd(gnd), .vdd(vdd), .A(_111__7_), .B(_9342_), .C(_12__7_), .D(_9341_), .Y(_12019_) );
NAND3X1 NAND3X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_12019_), .B(_12017_), .C(_12018_), .Y(_12020_) );
AOI22X1 AOI22X1_291 ( .gnd(gnd), .vdd(vdd), .A(_100__7_), .B(_9346_), .C(_212__7_), .D(_9345_), .Y(_12021_) );
AOI22X1 AOI22X1_292 ( .gnd(gnd), .vdd(vdd), .A(_245__7_), .B(_9348_), .C(_140__7_), .D(_9349_), .Y(_12022_) );
NAND2X1 NAND2X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_12022_), .B(_12021_), .Y(_12023_) );
NOR2X1 NOR2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_12020_), .B(_12023_), .Y(_12024_) );
AOI22X1 AOI22X1_293 ( .gnd(gnd), .vdd(vdd), .A(_40__7_), .B(_8952_), .C(_29__7_), .D(_9176_), .Y(_12025_) );
AOI22X1 AOI22X1_294 ( .gnd(gnd), .vdd(vdd), .A(_218__7_), .B(_9169_), .C(_247__7_), .D(_9165_), .Y(_12026_) );
NAND2X1 NAND2X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_12026_), .B(_12025_), .Y(_12027_) );
NAND3X1 NAND3X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16184_), .C(_16185_), .Y(_12028_) );
OAI21X1 OAI21X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_9361_), .C(_12028_), .Y(_12029_) );
NAND3X1 NAND3X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16083_), .C(_16084_), .Y(_12030_) );
NAND3X1 NAND3X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16028_), .C(_16029_), .Y(_12031_) );
NAND2X1 NAND2X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_12030_), .B(_12031_), .Y(_12032_) );
NOR2X1 NOR2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_12032_), .B(_12029_), .Y(_12033_) );
NAND3X1 NAND3X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_8670_), .B(_9371_), .C(_8669_), .Y(_12034_) );
NAND3X1 NAND3X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8562_), .C(_8561_), .Y(_12035_) );
NAND2X1 NAND2X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_12035_), .B(_12034_), .Y(_12036_) );
NAND3X1 NAND3X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8615_), .C(_8616_), .Y(_12037_) );
NAND3X1 NAND3X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_312_), .C(_313_), .Y(_12038_) );
NAND2X1 NAND2X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_12037_), .B(_12038_), .Y(_12039_) );
NOR2X1 NOR2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_12039_), .B(_12036_), .Y(_12040_) );
AOI22X1 AOI22X1_295 ( .gnd(gnd), .vdd(vdd), .A(_250__7_), .B(_9082_), .C(_177__7_), .D(_8961_), .Y(_12041_) );
NAND3X1 NAND3X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_12033_), .B(_12040_), .C(_12041_), .Y(_12042_) );
NOR2X1 NOR2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_12042_), .B(_12027_), .Y(_12043_) );
NAND3X1 NAND3X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_12024_), .B(_12016_), .C(_12043_), .Y(_12044_) );
NOR3X1 NOR3X1_332 ( .gnd(gnd), .vdd(vdd), .A(_11931_), .B(_11946_), .C(_12044_), .Y(_12045_) );
NAND3X1 NAND3X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_11775_), .B(_12045_), .C(_11902_), .Y(_12046_) );
NAND2X1 NAND2X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__7_), .Y(_12047_) );
NAND2X1 NAND2X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__7_), .Y(_12048_) );
NAND2X1 NAND2X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_12048_), .B(_12047_), .Y(_12049_) );
NOR3X1 NOR3X1_333 ( .gnd(gnd), .vdd(vdd), .A(_11767_), .B(_12049_), .C(_12046_), .Y(_12050_) );
NOR3X1 NOR3X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_9397_), .C(_1854_), .Y(_12051_) );
NAND3X1 NAND3X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1458_), .C(_1457_), .Y(_12052_) );
NAND3X1 NAND3X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_9453_), .B(_1412_), .C(_1411_), .Y(_12053_) );
NAND2X1 NAND2X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_12052_), .B(_12053_), .Y(_12054_) );
NAND3X1 NAND3X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1508_), .C(_1507_), .Y(_12055_) );
NAND3X1 NAND3X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1291_), .C(_1290_), .Y(_12056_) );
NAND2X1 NAND2X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_12055_), .B(_12056_), .Y(_12057_) );
NOR2X1 NOR2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_12057_), .B(_12054_), .Y(_12058_) );
AOI22X1 AOI22X1_296 ( .gnd(gnd), .vdd(vdd), .A(_125__7_), .B(_9411_), .C(_122__7_), .D(_9444_), .Y(_12059_) );
NAND3X1 NAND3X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_9413_), .C(_1103_), .Y(_12060_) );
NAND2X1 NAND2X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__7_), .Y(_12061_) );
NAND3X1 NAND3X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_12060_), .B(_12061_), .C(_12059_), .Y(_12062_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_776_), .B(_9421_), .C(_814_), .D(_9419_), .Y(_12063_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_9426_), .C(_699_), .D(_9424_), .Y(_12064_) );
NOR2X1 NOR2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_12063_), .B(_12064_), .Y(_12065_) );
NAND3X1 NAND3X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7414_), .C(_7415_), .Y(_12066_) );
NAND2X1 NAND2X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__7_), .Y(_12067_) );
AOI22X1 AOI22X1_297 ( .gnd(gnd), .vdd(vdd), .A(_229__7_), .B(_9433_), .C(_139__7_), .D(_9431_), .Y(_12068_) );
NAND3X1 NAND3X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_12067_), .B(_12066_), .C(_12068_), .Y(_12069_) );
NAND3X1 NAND3X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_661_), .C(_662_), .Y(_12070_) );
OAI21X1 OAI21X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_9440_), .C(_12070_), .Y(_12071_) );
NOR2X1 NOR2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_12071_), .B(_12069_), .Y(_12072_) );
NAND2X1 NAND2X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_12072_), .B(_12065_), .Y(_12073_) );
NAND3X1 NAND3X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_9410_), .C(_1012_), .Y(_12074_) );
NAND2X1 NAND2X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__7_), .Y(_12075_) );
AOI22X1 AOI22X1_298 ( .gnd(gnd), .vdd(vdd), .A(_130__7_), .B(_9449_), .C(_127__7_), .D(_9448_), .Y(_12076_) );
NAND3X1 NAND3X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_12074_), .B(_12075_), .C(_12076_), .Y(_12077_) );
NOR3X1 NOR3X1_335 ( .gnd(gnd), .vdd(vdd), .A(_12077_), .B(_12062_), .C(_12073_), .Y(_12078_) );
AOI22X1 AOI22X1_299 ( .gnd(gnd), .vdd(vdd), .A(_115__7_), .B(_9399_), .C(_114__7_), .D(_9454_), .Y(_12079_) );
NAND3X1 NAND3X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_12079_), .B(_12058_), .C(_12078_), .Y(_12080_) );
NAND3X1 NAND3X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_9457_), .C(_1712_), .Y(_12081_) );
NAND2X1 NAND2X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__7_), .Y(_12082_) );
NAND2X1 NAND2X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_12082_), .B(_12081_), .Y(_12083_) );
NOR3X1 NOR3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_12083_), .B(_12051_), .C(_12080_), .Y(_12084_) );
NAND3X1 NAND3X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_11760_), .B(_12084_), .C(_12050_), .Y(_12085_) );
NOR2X1 NOR2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_11759_), .B(_12085_), .Y(_12086_) );
NAND3X1 NAND3X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_11748_), .B(_11755_), .C(_12086_), .Y(_12087_) );
NAND2X1 NAND2X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__7_), .Y(_12088_) );
NAND3X1 NAND3X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .B(_8806_), .C(_2399_), .Y(_12089_) );
NAND2X1 NAND2X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_12089_), .B(_12088_), .Y(_12090_) );
NOR3X1 NOR3X1_337 ( .gnd(gnd), .vdd(vdd), .A(_11740_), .B(_12090_), .C(_12087_), .Y(_12091_) );
NAND3X1 NAND3X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_11732_), .B(_11737_), .C(_12091_), .Y(_12092_) );
NAND3X1 NAND3X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_3061_), .B(_9473_), .C(_3062_), .Y(_12093_) );
NAND2X1 NAND2X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__7_), .Y(_12094_) );
NAND2X1 NAND2X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__7_), .Y(_12095_) );
NAND2X1 NAND2X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__7_), .Y(_12096_) );
NAND2X1 NAND2X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__7_), .Y(_12097_) );
NAND3X1 NAND3X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_12095_), .B(_12096_), .C(_12097_), .Y(_12098_) );
AOI21X1 AOI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_68__7_), .B(_9477_), .C(_12098_), .Y(_12099_) );
NAND3X1 NAND3X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_12093_), .B(_12099_), .C(_12094_), .Y(_12100_) );
NOR3X1 NOR3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_11731_), .B(_12100_), .C(_12092_), .Y(_12101_) );
AOI21X1 AOI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_11726_), .B(_12101_), .C(rst), .Y(_0__7_) );
NAND2X1 NAND2X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__8_), .Y(_12102_) );
NAND2X1 NAND2X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__8_), .Y(_12103_) );
NAND2X1 NAND2X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_12102_), .B(_12103_), .Y(_12104_) );
NAND2X1 NAND2X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__8_), .Y(_12105_) );
NAND2X1 NAND2X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__8_), .Y(_12106_) );
NAND2X1 NAND2X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_12105_), .B(_12106_), .Y(_12107_) );
NOR2X1 NOR2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_12104_), .B(_12107_), .Y(_12108_) );
NAND3X1 NAND3X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_3281_), .B(_8762_), .C(_3280_), .Y(_12109_) );
NAND3X1 NAND3X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_3235_), .B(_8765_), .C(_3234_), .Y(_12110_) );
AND2X2 AND2X2_1586 ( .gnd(gnd), .vdd(vdd), .A(_12110_), .B(_12109_), .Y(_12111_) );
AOI22X1 AOI22X1_300 ( .gnd(gnd), .vdd(vdd), .A(_62__8_), .B(_8774_), .C(_57__8_), .D(_8771_), .Y(_12112_) );
NAND2X1 NAND2X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_12111_), .B(_12112_), .Y(_12113_) );
NAND2X1 NAND2X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__8_), .Y(_12114_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_2765_), .B(_8799_), .C(_2709_), .D(_8792_), .Y(_12115_) );
NAND3X1 NAND3X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .B(_8794_), .C(_2648_), .Y(_12116_) );
NAND3X1 NAND3X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_2818_), .B(_8786_), .C(_2819_), .Y(_12117_) );
NAND2X1 NAND2X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_12116_), .B(_12117_), .Y(_12118_) );
NOR2X1 NOR2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_12115_), .B(_12118_), .Y(_12119_) );
AOI22X1 AOI22X1_301 ( .gnd(gnd), .vdd(vdd), .A(_80__8_), .B(_8805_), .C(_79__8_), .D(_9466_), .Y(_12120_) );
AOI22X1 AOI22X1_302 ( .gnd(gnd), .vdd(vdd), .A(_75__8_), .B(_8802_), .C(_81__8_), .D(_9468_), .Y(_12121_) );
NAND2X1 NAND2X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_12120_), .B(_12121_), .Y(_12122_) );
NAND2X1 NAND2X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__8_), .Y(_12123_) );
NAND2X1 NAND2X1_2051 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__8_), .Y(_12124_) );
NAND2X1 NAND2X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_12123_), .B(_12124_), .Y(_12125_) );
INVX1 INVX1_3877 ( .gnd(gnd), .vdd(vdd), .A(_84__8_), .Y(_12126_) );
NOR2X1 NOR2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_12126_), .Y(_12127_) );
NOR2X1 NOR2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2298_), .Y(_12128_) );
NAND2X1 NAND2X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__8_), .Y(_12129_) );
NAND3X1 NAND3X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .B(_8840_), .C(_1973_), .Y(_12130_) );
NAND3X1 NAND3X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1916_), .C(_1917_), .Y(_12131_) );
NAND3X1 NAND3X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_12131_), .B(_12130_), .C(_12129_), .Y(_12132_) );
NOR3X1 NOR3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_12127_), .B(_12132_), .C(_12128_), .Y(_12133_) );
NAND3X1 NAND3X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_2254_), .B(_8829_), .C(_2255_), .Y(_12134_) );
NAND3X1 NAND3X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_2148_), .B(_8831_), .C(_2149_), .Y(_12135_) );
NAND2X1 NAND2X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_12134_), .B(_12135_), .Y(_12136_) );
NAND3X1 NAND3X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .B(_8834_), .C(_2090_), .Y(_12137_) );
NAND3X1 NAND3X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .B(_8836_), .C(_2201_), .Y(_12138_) );
NAND2X1 NAND2X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_12137_), .B(_12138_), .Y(_12139_) );
NOR2X1 NOR2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_12139_), .B(_12136_), .Y(_12140_) );
AOI22X1 AOI22X1_303 ( .gnd(gnd), .vdd(vdd), .A(_94__8_), .B(_8841_), .C(_91__8_), .D(_8823_), .Y(_12141_) );
AOI22X1 AOI22X1_304 ( .gnd(gnd), .vdd(vdd), .A(_98__8_), .B(_8845_), .C(_92__8_), .D(_8843_), .Y(_12142_) );
NAND2X1 NAND2X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_12142_), .B(_12141_), .Y(_12143_) );
NAND2X1 NAND2X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__8_), .Y(_12144_) );
NAND2X1 NAND2X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__8_), .Y(_12145_) );
NAND2X1 NAND2X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__8_), .Y(_12146_) );
NAND2X1 NAND2X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_12145_), .B(_12146_), .Y(_12147_) );
NAND2X1 NAND2X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__8_), .Y(_12148_) );
NAND2X1 NAND2X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__8_), .Y(_12149_) );
NAND2X1 NAND2X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_12148_), .B(_12149_), .Y(_12150_) );
NOR2X1 NOR2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_12147_), .B(_12150_), .Y(_12151_) );
NAND2X1 NAND2X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__8_), .Y(_12152_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_7144_), .B(_9930_), .C(_7188_), .D(_9929_), .Y(_12153_) );
NOR2X1 NOR2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7323_), .Y(_12154_) );
NOR2X1 NOR2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7280_), .Y(_12155_) );
NOR3X1 NOR3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_12154_), .B(_12155_), .C(_12153_), .Y(_12156_) );
NAND2X1 NAND2X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__8_), .Y(_12157_) );
NAND2X1 NAND2X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__8_), .Y(_12158_) );
NAND2X1 NAND2X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_12157_), .B(_12158_), .Y(_12159_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_7366_), .B(_9940_), .C(_7234_), .D(_9941_), .Y(_12160_) );
NOR2X1 NOR2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_12160_), .B(_12159_), .Y(_12161_) );
NAND3X1 NAND3X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_12152_), .B(_12156_), .C(_12161_), .Y(_12162_) );
AOI22X1 AOI22X1_305 ( .gnd(gnd), .vdd(vdd), .A(_20__8_), .B(_8898_), .C(_236__8_), .D(_8955_), .Y(_12163_) );
AOI22X1 AOI22X1_306 ( .gnd(gnd), .vdd(vdd), .A(_237__8_), .B(_8966_), .C(_175__8_), .D(_8904_), .Y(_12164_) );
NAND2X1 NAND2X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_12163_), .B(_12164_), .Y(_12165_) );
NAND2X1 NAND2X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__8_), .Y(_12166_) );
NAND2X1 NAND2X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__8_), .Y(_12167_) );
AOI22X1 AOI22X1_307 ( .gnd(gnd), .vdd(vdd), .A(_19__8_), .B(_8914_), .C(_210__8_), .D(_8918_), .Y(_12168_) );
NAND3X1 NAND3X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_12166_), .B(_12167_), .C(_12168_), .Y(_12169_) );
NOR2X1 NOR2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_12165_), .B(_12169_), .Y(_12170_) );
AOI22X1 AOI22X1_308 ( .gnd(gnd), .vdd(vdd), .A(_123__8_), .B(_8928_), .C(_9__8_), .D(_8926_), .Y(_12171_) );
NAND2X1 NAND2X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__8_), .Y(_12172_) );
NAND2X1 NAND2X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_134__8_), .Y(_12173_) );
NAND3X1 NAND3X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_12172_), .B(_12173_), .C(_12171_), .Y(_12174_) );
AOI22X1 AOI22X1_309 ( .gnd(gnd), .vdd(vdd), .A(_4__8_), .B(_8937_), .C(_176__8_), .D(_8939_), .Y(_12175_) );
NAND2X1 NAND2X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__8_), .Y(_12176_) );
NAND2X1 NAND2X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__8_), .Y(_12177_) );
NAND3X1 NAND3X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_12176_), .B(_12177_), .C(_12175_), .Y(_12178_) );
NOR2X1 NOR2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_12178_), .B(_12174_), .Y(_12179_) );
NAND2X1 NAND2X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_12170_), .B(_12179_), .Y(_12180_) );
NAND2X1 NAND2X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_9082_), .B(_250__8_), .Y(_12181_) );
NAND2X1 NAND2X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_9161_), .B(_47__8_), .Y(_12182_) );
AOI22X1 AOI22X1_310 ( .gnd(gnd), .vdd(vdd), .A(_21__8_), .B(_9150_), .C(_185__8_), .D(_9151_), .Y(_12183_) );
NAND3X1 NAND3X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_12181_), .B(_12182_), .C(_12183_), .Y(_12184_) );
AOI22X1 AOI22X1_311 ( .gnd(gnd), .vdd(vdd), .A(_246__8_), .B(_9356_), .C(_226__8_), .D(_9357_), .Y(_12185_) );
NAND2X1 NAND2X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_9157_), .B(_231__8_), .Y(_12186_) );
NAND2X1 NAND2X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_46__8_), .Y(_12187_) );
NAND3X1 NAND3X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_12186_), .B(_12187_), .C(_12185_), .Y(_12188_) );
NOR2X1 NOR2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_12184_), .B(_12188_), .Y(_12189_) );
NAND2X1 NAND2X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_145__8_), .Y(_12190_) );
NAND2X1 NAND2X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__8_), .Y(_12191_) );
AOI22X1 AOI22X1_312 ( .gnd(gnd), .vdd(vdd), .A(_37__8_), .B(_8978_), .C(_35__8_), .D(_8980_), .Y(_12192_) );
NAND3X1 NAND3X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_12190_), .B(_12191_), .C(_12192_), .Y(_12193_) );
NAND2X1 NAND2X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_9053_), .B(_249__8_), .Y(_12194_) );
NAND2X1 NAND2X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_253__8_), .Y(_12195_) );
AOI22X1 AOI22X1_313 ( .gnd(gnd), .vdd(vdd), .A(_178__8_), .B(_9173_), .C(_214__8_), .D(_9174_), .Y(_12196_) );
NAND3X1 NAND3X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_12194_), .B(_12195_), .C(_12196_), .Y(_12197_) );
NOR2X1 NOR2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_12193_), .B(_12197_), .Y(_12198_) );
NAND2X1 NAND2X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_12189_), .B(_12198_), .Y(_12199_) );
NOR2X1 NOR2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_12180_), .B(_12199_), .Y(_12200_) );
NAND2X1 NAND2X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__8_), .Y(_12201_) );
NAND2X1 NAND2X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__8_), .Y(_12202_) );
AOI22X1 AOI22X1_314 ( .gnd(gnd), .vdd(vdd), .A(_13__8_), .B(_9007_), .C(_239__8_), .D(_9076_), .Y(_12203_) );
NAND3X1 NAND3X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_12201_), .B(_12202_), .C(_12203_), .Y(_12204_) );
AOI22X1 AOI22X1_315 ( .gnd(gnd), .vdd(vdd), .A(_206__8_), .B(_9013_), .C(_242__8_), .D(_9035_), .Y(_12205_) );
NAND2X1 NAND2X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__8_), .Y(_12206_) );
NAND2X1 NAND2X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_9018_), .B(_203__8_), .Y(_12207_) );
NAND3X1 NAND3X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_12206_), .B(_12207_), .C(_12205_), .Y(_12208_) );
NOR2X1 NOR2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_12204_), .B(_12208_), .Y(_12209_) );
AOI22X1 AOI22X1_316 ( .gnd(gnd), .vdd(vdd), .A(_222__8_), .B(_9024_), .C(_220__8_), .D(_9026_), .Y(_12210_) );
NAND2X1 NAND2X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__8_), .Y(_12211_) );
NAND2X1 NAND2X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__8_), .Y(_12212_) );
NAND3X1 NAND3X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_12211_), .B(_12212_), .C(_12210_), .Y(_12213_) );
AOI22X1 AOI22X1_317 ( .gnd(gnd), .vdd(vdd), .A(_18__8_), .B(_9037_), .C(_240__8_), .D(_9011_), .Y(_12214_) );
NAND2X1 NAND2X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__8_), .Y(_12215_) );
NAND2X1 NAND2X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__8_), .Y(_12216_) );
NAND3X1 NAND3X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_12215_), .B(_12216_), .C(_12214_), .Y(_12217_) );
NOR2X1 NOR2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_12213_), .B(_12217_), .Y(_12218_) );
NAND2X1 NAND2X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_12209_), .B(_12218_), .Y(_12219_) );
AOI22X1 AOI22X1_318 ( .gnd(gnd), .vdd(vdd), .A(_225__8_), .B(_9048_), .C(_167__8_), .D(_9050_), .Y(_12220_) );
NAND2X1 NAND2X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_243__8_), .Y(_12221_) );
NAND2X1 NAND2X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__8_), .Y(_12222_) );
NAND3X1 NAND3X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_12221_), .B(_12222_), .C(_12220_), .Y(_12223_) );
NAND2X1 NAND2X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__8_), .Y(_12224_) );
NAND2X1 NAND2X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__8_), .Y(_12225_) );
AOI22X1 AOI22X1_319 ( .gnd(gnd), .vdd(vdd), .A(_224__8_), .B(_9064_), .C(_27__8_), .D(_9066_), .Y(_12226_) );
NAND3X1 NAND3X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_12224_), .B(_12225_), .C(_12226_), .Y(_12227_) );
NOR2X1 NOR2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_12223_), .B(_12227_), .Y(_12228_) );
AOI22X1 AOI22X1_320 ( .gnd(gnd), .vdd(vdd), .A(_184__8_), .B(_9073_), .C(_183__8_), .D(_9071_), .Y(_12229_) );
NAND2X1 NAND2X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__8_), .Y(_12230_) );
NAND2X1 NAND2X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__8_), .Y(_12231_) );
NAND3X1 NAND3X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_12230_), .B(_12231_), .C(_12229_), .Y(_12232_) );
AOI22X1 AOI22X1_321 ( .gnd(gnd), .vdd(vdd), .A(_43__8_), .B(_9084_), .C(_244__8_), .D(_9160_), .Y(_12233_) );
NAND2X1 NAND2X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__8_), .Y(_12234_) );
NAND2X1 NAND2X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__8_), .Y(_12235_) );
NAND3X1 NAND3X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_12234_), .B(_12235_), .C(_12233_), .Y(_12236_) );
NOR2X1 NOR2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_12232_), .B(_12236_), .Y(_12237_) );
NAND2X1 NAND2X1_2102 ( .gnd(gnd), .vdd(vdd), .A(_12228_), .B(_12237_), .Y(_12238_) );
NOR2X1 NOR2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_12219_), .B(_12238_), .Y(_12239_) );
NAND3X1 NAND3X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_6976_), .B(_9145_), .C(_6977_), .Y(_12240_) );
NAND3X1 NAND3X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_6934_), .B(_9137_), .C(_6935_), .Y(_12241_) );
NAND2X1 NAND2X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_12240_), .B(_12241_), .Y(_12242_) );
NAND3X1 NAND3X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_9135_), .C(_5052_), .Y(_12243_) );
NAND2X1 NAND2X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__8_), .Y(_12244_) );
NAND2X1 NAND2X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_12243_), .B(_12244_), .Y(_12245_) );
NOR2X1 NOR2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_12242_), .B(_12245_), .Y(_12246_) );
NAND3X1 NAND3X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_15926_), .B(_9109_), .C(_15927_), .Y(_12247_) );
NAND3X1 NAND3X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_8319_), .B(_9188_), .C(_8320_), .Y(_12248_) );
NAND3X1 NAND3X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_16132_), .B(_9115_), .C(_16133_), .Y(_12249_) );
NAND3X1 NAND3X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_12247_), .B(_12249_), .C(_12248_), .Y(_12250_) );
AOI22X1 AOI22X1_322 ( .gnd(gnd), .vdd(vdd), .A(_234__8_), .B(_9182_), .C(_34__8_), .D(_9183_), .Y(_12251_) );
AOI22X1 AOI22X1_323 ( .gnd(gnd), .vdd(vdd), .A(_100__8_), .B(_9346_), .C(_45__8_), .D(_9185_), .Y(_12252_) );
NAND2X1 NAND2X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_12252_), .B(_12251_), .Y(_12253_) );
NAND3X1 NAND3X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_4707_), .B(_9140_), .C(_4706_), .Y(_12254_) );
OAI21X1 OAI21X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_5245_), .B(_10036_), .C(_12254_), .Y(_12255_) );
NOR3X1 NOR3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_12255_), .B(_12250_), .C(_12253_), .Y(_12256_) );
NAND3X1 NAND3X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_3425_), .B(_9133_), .C(_3426_), .Y(_12257_) );
NAND3X1 NAND3X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .B(_9102_), .C(_5099_), .Y(_12258_) );
NAND3X1 NAND3X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_6857_), .B(_9104_), .C(_6858_), .Y(_12259_) );
NAND3X1 NAND3X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_12258_), .B(_12259_), .C(_12257_), .Y(_12260_) );
AOI22X1 AOI22X1_324 ( .gnd(gnd), .vdd(vdd), .A(_38__8_), .B(_9129_), .C(_16__8_), .D(_9127_), .Y(_12261_) );
AOI22X1 AOI22X1_325 ( .gnd(gnd), .vdd(vdd), .A(_39__8_), .B(_9099_), .C(_10__8_), .D(_9097_), .Y(_12262_) );
NAND2X1 NAND2X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_12261_), .B(_12262_), .Y(_12263_) );
NOR2X1 NOR2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_12260_), .B(_12263_), .Y(_12264_) );
NAND3X1 NAND3X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_12246_), .B(_12256_), .C(_12264_), .Y(_12265_) );
AOI22X1 AOI22X1_326 ( .gnd(gnd), .vdd(vdd), .A(_227__8_), .B(_9170_), .C(_30__8_), .D(_9167_), .Y(_12266_) );
AOI22X1 AOI22X1_327 ( .gnd(gnd), .vdd(vdd), .A(_33__8_), .B(_8991_), .C(_213__8_), .D(_8989_), .Y(_12267_) );
NAND2X1 NAND2X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_12266_), .B(_12267_), .Y(_12268_) );
AOI22X1 AOI22X1_328 ( .gnd(gnd), .vdd(vdd), .A(_44__8_), .B(_8968_), .C(_42__8_), .D(_8963_), .Y(_12269_) );
AOI22X1 AOI22X1_329 ( .gnd(gnd), .vdd(vdd), .A(_238__8_), .B(_8893_), .C(_208__8_), .D(_8950_), .Y(_12270_) );
NAND2X1 NAND2X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_12269_), .B(_12270_), .Y(_12271_) );
NOR2X1 NOR2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_12268_), .B(_12271_), .Y(_12272_) );
AOI22X1 AOI22X1_330 ( .gnd(gnd), .vdd(vdd), .A(_22__8_), .B(_9382_), .C(_3__8_), .D(_9383_), .Y(_12273_) );
NAND2X1 NAND2X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_219__8_), .Y(_12274_) );
NAND2X1 NAND2X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(_232__8_), .Y(_12275_) );
NAND3X1 NAND3X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_12274_), .B(_12275_), .C(_12273_), .Y(_12276_) );
AOI22X1 AOI22X1_331 ( .gnd(gnd), .vdd(vdd), .A(_209__8_), .B(_8957_), .C(_254__8_), .D(_8984_), .Y(_12277_) );
AOI22X1 AOI22X1_332 ( .gnd(gnd), .vdd(vdd), .A(_255__8_), .B(_8986_), .C(_156__8_), .D(_8973_), .Y(_12278_) );
NAND2X1 NAND2X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_12277_), .B(_12278_), .Y(_12279_) );
NOR2X1 NOR2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_12276_), .B(_12279_), .Y(_12280_) );
NAND2X1 NAND2X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_12272_), .B(_12280_), .Y(_12281_) );
AOI22X1 AOI22X1_333 ( .gnd(gnd), .vdd(vdd), .A(_201__8_), .B(_9124_), .C(_212__8_), .D(_9345_), .Y(_12282_) );
NAND3X1 NAND3X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_8433_), .B(_9348_), .C(_8432_), .Y(_12283_) );
NAND3X1 NAND3X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_493_), .C(_494_), .Y(_12284_) );
AND2X2 AND2X2_1587 ( .gnd(gnd), .vdd(vdd), .A(_12284_), .B(_12283_), .Y(_12285_) );
NAND2X1 NAND2X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_12282_), .B(_12285_), .Y(_12286_) );
NAND3X1 NAND3X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_15139_), .B(_9208_), .C(_15140_), .Y(_12287_) );
OAI21X1 OAI21X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_15104_), .B(_9211_), .C(_12287_), .Y(_12288_) );
NAND3X1 NAND3X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_15483_), .B(_9222_), .C(_15484_), .Y(_12289_) );
NAND3X1 NAND3X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_15430_), .B(_9224_), .C(_15429_), .Y(_12290_) );
NAND2X1 NAND2X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_12289_), .B(_12290_), .Y(_12291_) );
NOR2X1 NOR2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_12291_), .B(_12288_), .Y(_12292_) );
NAND3X1 NAND3X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_15261_), .B(_9217_), .C(_15262_), .Y(_12293_) );
NAND3X1 NAND3X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_15209_), .B(_9219_), .C(_15208_), .Y(_12294_) );
NAND2X1 NAND2X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_12294_), .B(_12293_), .Y(_12295_) );
NAND3X1 NAND3X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_15659_), .B(_9192_), .C(_15660_), .Y(_12296_) );
NAND3X1 NAND3X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_15716_), .B(_9199_), .C(_15715_), .Y(_12297_) );
NAND2X1 NAND2X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_12297_), .B(_12296_), .Y(_12298_) );
NOR2X1 NOR2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_12298_), .B(_12295_), .Y(_12299_) );
NOR3X1 NOR3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_16186_), .B(_10083_), .C(_16187_), .Y(_12300_) );
NAND3X1 NAND3X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_15311_), .B(_9205_), .C(_15312_), .Y(_12301_) );
OAI21X1 OAI21X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_15346_), .B(_10085_), .C(_12301_), .Y(_12302_) );
NAND3X1 NAND3X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_15541_), .B(_9233_), .C(_15542_), .Y(_12303_) );
NAND3X1 NAND3X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15609_), .C(_15608_), .Y(_12304_) );
NAND2X1 NAND2X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_12303_), .B(_12304_), .Y(_12305_) );
NOR3X1 NOR3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_12302_), .B(_12305_), .C(_12300_), .Y(_12306_) );
NAND3X1 NAND3X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_12292_), .B(_12299_), .C(_12306_), .Y(_12307_) );
NAND3X1 NAND3X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_15869_), .B(_9120_), .C(_15870_), .Y(_12308_) );
NAND3X1 NAND3X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_15380_), .B(_9197_), .C(_15381_), .Y(_12309_) );
NOR2X1 NOR2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_9267_), .B(_7050_), .Y(_12310_) );
AND2X2 AND2X2_1588 ( .gnd(gnd), .vdd(vdd), .A(_187__8_), .B(_9235_), .Y(_12311_) );
NOR2X1 NOR2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_11264_), .B(_15811_), .Y(_12312_) );
OR2X2 OR2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_12311_), .B(_12312_), .Y(_12313_) );
NAND3X1 NAND3X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_7009_), .B(_7010_), .C(_9289_), .Y(_12314_) );
OAI21X1 OAI21X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_8710_), .C(_12314_), .Y(_12315_) );
NAND3X1 NAND3X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_7095_), .B(_9244_), .C(_7094_), .Y(_12316_) );
OAI21X1 OAI21X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_14912_), .B(_9276_), .C(_12316_), .Y(_12317_) );
NOR2X1 NOR2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_12317_), .B(_12315_), .Y(_12318_) );
NOR2X1 NOR2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_8167_), .Y(_12319_) );
NOR2X1 NOR2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_11613_), .B(_7496_), .Y(_12320_) );
NAND3X1 NAND3X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_8200_), .B(_9286_), .C(_8201_), .Y(_12321_) );
NAND3X1 NAND3X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(_9268_), .C(_1171_), .Y(_12322_) );
NAND2X1 NAND2X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_12322_), .B(_12321_), .Y(_12323_) );
NOR3X1 NOR3X1_344 ( .gnd(gnd), .vdd(vdd), .A(_12319_), .B(_12320_), .C(_12323_), .Y(_12324_) );
NAND2X1 NAND2X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_12318_), .B(_12324_), .Y(_12325_) );
NOR3X1 NOR3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_12310_), .B(_12313_), .C(_12325_), .Y(_12326_) );
NAND3X1 NAND3X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_9310_), .B(_5965_), .C(_5966_), .Y(_12327_) );
NAND3X1 NAND3X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_6467_), .B(_6468_), .C(_9260_), .Y(_12328_) );
NAND3X1 NAND3X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_3604_), .B(_9294_), .C(_3605_), .Y(_12329_) );
NAND3X1 NAND3X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_12328_), .B(_12327_), .C(_12329_), .Y(_12330_) );
NAND3X1 NAND3X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_7677_), .B(_9321_), .C(_7678_), .Y(_12331_) );
OAI21X1 OAI21X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_5403_), .B(_9319_), .C(_12331_), .Y(_12332_) );
NOR2X1 NOR2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_12332_), .B(_12330_), .Y(_12333_) );
NAND3X1 NAND3X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_8236_), .B(_9250_), .C(_8237_), .Y(_12334_) );
OAI21X1 OAI21X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_3556_), .B(_9306_), .C(_12334_), .Y(_12335_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_7634_), .B(_9301_), .C(_4188_), .D(_9254_), .Y(_12336_) );
NOR2X1 NOR2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_12336_), .B(_12335_), .Y(_12337_) );
NAND3X1 NAND3X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_7718_), .B(_9248_), .C(_7719_), .Y(_12338_) );
OAI21X1 OAI21X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_9263_), .C(_12338_), .Y(_12339_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .Y(_12340_) );
NAND3X1 NAND3X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_2914_), .B(_9277_), .C(_2915_), .Y(_12341_) );
OAI21X1 OAI21X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(_12340_), .C(_12341_), .Y(_12342_) );
NOR2X1 NOR2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_12339_), .B(_12342_), .Y(_12343_) );
NAND3X1 NAND3X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_12337_), .B(_12343_), .C(_12333_), .Y(_12344_) );
NAND2X1 NAND2X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_9326_), .B(_252__8_), .Y(_12345_) );
AOI22X1 AOI22X1_334 ( .gnd(gnd), .vdd(vdd), .A(_15__8_), .B(_9313_), .C(_235__8_), .D(_9324_), .Y(_12346_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_4222_), .B(_9282_), .C(_4816_), .D(_9273_), .Y(_12347_) );
NAND3X1 NAND3X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_2360_), .B(_9315_), .C(_2361_), .Y(_12348_) );
OAI21X1 OAI21X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_6432_), .B(_9763_), .C(_12348_), .Y(_12349_) );
NOR2X1 NOR2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_12347_), .B(_12349_), .Y(_12350_) );
NAND3X1 NAND3X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_12345_), .B(_12346_), .C(_12350_), .Y(_12351_) );
NOR2X1 NOR2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_12351_), .B(_12344_), .Y(_12352_) );
NAND3X1 NAND3X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_12309_), .B(_12326_), .C(_12352_), .Y(_12353_) );
AOI21X1 AOI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_157__8_), .B(_9232_), .C(_12353_), .Y(_12354_) );
AOI22X1 AOI22X1_335 ( .gnd(gnd), .vdd(vdd), .A(_155__8_), .B(_9333_), .C(_172__8_), .D(_9332_), .Y(_12355_) );
NAND3X1 NAND3X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_12308_), .B(_12355_), .C(_12354_), .Y(_12356_) );
NOR3X1 NOR3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_12307_), .B(_12356_), .C(_12286_), .Y(_12357_) );
AOI22X1 AOI22X1_336 ( .gnd(gnd), .vdd(vdd), .A(_256__8_), .B(_9113_), .C(_142__8_), .D(_9118_), .Y(_12358_) );
NAND2X1 NAND2X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__8_), .Y(_12359_) );
NAND2X1 NAND2X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__8_), .Y(_12360_) );
NAND3X1 NAND3X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_12359_), .B(_12360_), .C(_12358_), .Y(_12361_) );
NAND2X1 NAND2X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__8_), .Y(_12362_) );
NAND3X1 NAND3X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_9339_), .C(_452_), .Y(_12363_) );
AOI22X1 AOI22X1_337 ( .gnd(gnd), .vdd(vdd), .A(_111__8_), .B(_9342_), .C(_12__8_), .D(_9341_), .Y(_12364_) );
NAND3X1 NAND3X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_12364_), .B(_12362_), .C(_12363_), .Y(_12365_) );
NOR2X1 NOR2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_12361_), .B(_12365_), .Y(_12366_) );
AOI22X1 AOI22X1_338 ( .gnd(gnd), .vdd(vdd), .A(_40__8_), .B(_8952_), .C(_29__8_), .D(_9176_), .Y(_12367_) );
AOI22X1 AOI22X1_339 ( .gnd(gnd), .vdd(vdd), .A(_247__8_), .B(_9165_), .C(_218__8_), .D(_9169_), .Y(_12368_) );
NAND2X1 NAND2X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_12368_), .B(_12367_), .Y(_12369_) );
NAND3X1 NAND3X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16086_), .C(_16087_), .Y(_12370_) );
NAND3X1 NAND3X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16031_), .C(_16032_), .Y(_12371_) );
NAND2X1 NAND2X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_12370_), .B(_12371_), .Y(_12372_) );
NAND3X1 NAND3X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8565_), .C(_8564_), .Y(_12373_) );
OAI21X1 OAI21X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_9361_), .C(_12373_), .Y(_12374_) );
NOR2X1 NOR2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_12372_), .B(_12374_), .Y(_12375_) );
NAND2X1 NAND2X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_15977_), .B(_15978_), .Y(_12376_) );
NAND3X1 NAND3X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8618_), .C(_8619_), .Y(_12377_) );
OAI21X1 OAI21X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_12376_), .B(_9215_), .C(_12377_), .Y(_12378_) );
NAND3X1 NAND3X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_8673_), .B(_9371_), .C(_8672_), .Y(_12379_) );
NAND3X1 NAND3X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_315_), .C(_316_), .Y(_12380_) );
NAND2X1 NAND2X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_12380_), .B(_12379_), .Y(_12381_) );
NOR2X1 NOR2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_12378_), .B(_12381_), .Y(_12382_) );
AOI22X1 AOI22X1_340 ( .gnd(gnd), .vdd(vdd), .A(_248__8_), .B(_8901_), .C(_177__8_), .D(_8961_), .Y(_12383_) );
NAND3X1 NAND3X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_12375_), .B(_12382_), .C(_12383_), .Y(_12384_) );
NOR2X1 NOR2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_12369_), .B(_12384_), .Y(_12385_) );
NAND3X1 NAND3X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_12357_), .B(_12366_), .C(_12385_), .Y(_12386_) );
NOR3X1 NOR3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_12265_), .B(_12281_), .C(_12386_), .Y(_12387_) );
NAND3X1 NAND3X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_12200_), .B(_12239_), .C(_12387_), .Y(_12388_) );
NAND3X1 NAND3X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1583_), .C(_1585_), .Y(_12389_) );
NAND3X1 NAND3X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_8862_), .C(_1246_), .Y(_12390_) );
NAND2X1 NAND2X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_12389_), .B(_12390_), .Y(_12391_) );
NOR3X1 NOR3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_12162_), .B(_12391_), .C(_12388_), .Y(_12392_) );
NAND3X1 NAND3X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_12144_), .B(_12151_), .C(_12392_), .Y(_12393_) );
NAND2X1 NAND2X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__8_), .Y(_12394_) );
NAND3X1 NAND3X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_9406_), .C(_1461_), .Y(_12395_) );
NAND3X1 NAND3X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_9453_), .C(_1415_), .Y(_12396_) );
AND2X2 AND2X2_1589 ( .gnd(gnd), .vdd(vdd), .A(_12395_), .B(_12396_), .Y(_12397_) );
NAND2X1 NAND2X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_108__8_), .Y(_12398_) );
NAND2X1 NAND2X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_116__8_), .Y(_12399_) );
NAND3X1 NAND3X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_12398_), .B(_12399_), .C(_12397_), .Y(_12400_) );
NAND2X1 NAND2X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_125__8_), .Y(_12401_) );
NAND2X1 NAND2X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_122__8_), .Y(_12402_) );
NAND2X1 NAND2X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_12401_), .B(_12402_), .Y(_12403_) );
NOR2X1 NOR2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_1107_), .Y(_12404_) );
AND2X2 AND2X2_1590 ( .gnd(gnd), .vdd(vdd), .A(_120__8_), .B(_9415_), .Y(_12405_) );
NOR3X1 NOR3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_12404_), .B(_12405_), .C(_12403_), .Y(_12406_) );
AOI22X1 AOI22X1_341 ( .gnd(gnd), .vdd(vdd), .A(_132__8_), .B(_9420_), .C(_131__8_), .D(_9418_), .Y(_12407_) );
NAND2X1 NAND2X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__8_), .Y(_12408_) );
NAND2X1 NAND2X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__8_), .Y(_12409_) );
NAND3X1 NAND3X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_12408_), .B(_12409_), .C(_12407_), .Y(_12410_) );
NAND3X1 NAND3X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_9431_), .C(_547_), .Y(_12411_) );
NAND2X1 NAND2X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__8_), .Y(_12412_) );
NAND2X1 NAND2X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__8_), .Y(_12413_) );
NAND3X1 NAND3X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_12413_), .B(_12411_), .C(_12412_), .Y(_12414_) );
AOI21X1 AOI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__8_), .C(_12414_), .Y(_12415_) );
NAND2X1 NAND2X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__8_), .Y(_12416_) );
NAND2X1 NAND2X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_136__8_), .Y(_12417_) );
NAND3X1 NAND3X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_12416_), .B(_12417_), .C(_12415_), .Y(_12418_) );
NAND3X1 NAND3X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_9410_), .C(_1015_), .Y(_12419_) );
NAND2X1 NAND2X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__8_), .Y(_12420_) );
AOI22X1 AOI22X1_342 ( .gnd(gnd), .vdd(vdd), .A(_130__8_), .B(_9449_), .C(_127__8_), .D(_9448_), .Y(_12421_) );
NAND3X1 NAND3X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_12419_), .B(_12421_), .C(_12420_), .Y(_12422_) );
NOR3X1 NOR3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_12410_), .B(_12418_), .C(_12422_), .Y(_12423_) );
AOI22X1 AOI22X1_343 ( .gnd(gnd), .vdd(vdd), .A(_115__8_), .B(_9399_), .C(_114__8_), .D(_9454_), .Y(_12424_) );
NAND3X1 NAND3X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_12406_), .B(_12424_), .C(_12423_), .Y(_12425_) );
NOR2X1 NOR2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_12400_), .B(_12425_), .Y(_12426_) );
AOI22X1 AOI22X1_344 ( .gnd(gnd), .vdd(vdd), .A(_102__8_), .B(_9459_), .C(_103__8_), .D(_9457_), .Y(_12427_) );
NAND3X1 NAND3X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_12394_), .B(_12427_), .C(_12426_), .Y(_12428_) );
NOR3X1 NOR3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_12143_), .B(_12428_), .C(_12393_), .Y(_12429_) );
NAND3X1 NAND3X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_12133_), .B(_12140_), .C(_12429_), .Y(_12430_) );
NOR3X1 NOR3X1_352 ( .gnd(gnd), .vdd(vdd), .A(_12122_), .B(_12125_), .C(_12430_), .Y(_12431_) );
NAND3X1 NAND3X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_12114_), .B(_12119_), .C(_12431_), .Y(_12432_) );
NAND3X1 NAND3X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_9473_), .C(_3065_), .Y(_12433_) );
NAND2X1 NAND2X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__8_), .Y(_12434_) );
NAND3X1 NAND3X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_2586_), .B(_8803_), .C(_2585_), .Y(_12435_) );
NAND2X1 NAND2X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__8_), .Y(_12436_) );
NAND3X1 NAND3X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_2401_), .B(_8806_), .C(_2402_), .Y(_12437_) );
NAND3X1 NAND3X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_12435_), .B(_12437_), .C(_12436_), .Y(_12438_) );
AOI21X1 AOI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_68__8_), .B(_9477_), .C(_12438_), .Y(_12439_) );
NAND3X1 NAND3X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_12433_), .B(_12439_), .C(_12434_), .Y(_12440_) );
NOR3X1 NOR3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_12113_), .B(_12440_), .C(_12432_), .Y(_12441_) );
AOI21X1 AOI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_12108_), .B(_12441_), .C(rst), .Y(_0__8_) );
NAND2X1 NAND2X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__9_), .Y(_12442_) );
NAND2X1 NAND2X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__9_), .Y(_12443_) );
NAND2X1 NAND2X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_12442_), .B(_12443_), .Y(_12444_) );
NAND2X1 NAND2X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_55__9_), .Y(_12445_) );
NAND2X1 NAND2X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__9_), .Y(_12446_) );
NAND2X1 NAND2X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_12446_), .B(_12445_), .Y(_12447_) );
NOR2X1 NOR2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_12447_), .B(_12444_), .Y(_12448_) );
NAND3X1 NAND3X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_3162_), .B(_8750_), .C(_3161_), .Y(_12449_) );
NAND3X1 NAND3X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .B(_8757_), .C(_3109_), .Y(_12450_) );
NAND2X1 NAND2X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_12449_), .B(_12450_), .Y(_12451_) );
NAND3X1 NAND3X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(_8762_), .C(_3283_), .Y(_12452_) );
NAND3X1 NAND3X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_8774_), .C(_3012_), .Y(_12453_) );
NAND2X1 NAND2X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_12452_), .B(_12453_), .Y(_12454_) );
OR2X2 OR2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_12451_), .B(_12454_), .Y(_12455_) );
NAND2X1 NAND2X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__9_), .Y(_12456_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_8799_), .C(_2712_), .D(_8792_), .Y(_12457_) );
NAND3X1 NAND3X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(_8794_), .C(_2651_), .Y(_12458_) );
NAND3X1 NAND3X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_8786_), .C(_2822_), .Y(_12459_) );
NAND2X1 NAND2X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_12458_), .B(_12459_), .Y(_12460_) );
NOR2X1 NOR2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_12457_), .B(_12460_), .Y(_12461_) );
AOI22X1 AOI22X1_345 ( .gnd(gnd), .vdd(vdd), .A(_73__9_), .B(_9480_), .C(_74__9_), .D(_8803_), .Y(_12462_) );
AOI22X1 AOI22X1_346 ( .gnd(gnd), .vdd(vdd), .A(_79__9_), .B(_9466_), .C(_81__9_), .D(_9468_), .Y(_12463_) );
NAND2X1 NAND2X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_12463_), .B(_12462_), .Y(_12464_) );
INVX1 INVX1_3878 ( .gnd(gnd), .vdd(vdd), .A(_84__9_), .Y(_12465_) );
NOR2X1 NOR2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_12465_), .Y(_12466_) );
NOR2X1 NOR2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2300_), .Y(_12467_) );
NAND2X1 NAND2X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__9_), .Y(_12468_) );
NAND3X1 NAND3X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_8843_), .C(_2015_), .Y(_12469_) );
NAND3X1 NAND3X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1919_), .C(_1920_), .Y(_12470_) );
NAND3X1 NAND3X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_12470_), .B(_12469_), .C(_12468_), .Y(_12471_) );
NOR3X1 NOR3X1_354 ( .gnd(gnd), .vdd(vdd), .A(_12466_), .B(_12471_), .C(_12467_), .Y(_12472_) );
NAND3X1 NAND3X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_2257_), .B(_8829_), .C(_2258_), .Y(_12473_) );
NAND3X1 NAND3X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(_8831_), .C(_2152_), .Y(_12474_) );
NAND2X1 NAND2X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_12473_), .B(_12474_), .Y(_12475_) );
NAND3X1 NAND3X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_2092_), .B(_8834_), .C(_2093_), .Y(_12476_) );
NAND3X1 NAND3X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_2203_), .B(_8836_), .C(_2204_), .Y(_12477_) );
NAND2X1 NAND2X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_12476_), .B(_12477_), .Y(_12478_) );
NOR2X1 NOR2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_12478_), .B(_12475_), .Y(_12479_) );
AOI22X1 AOI22X1_347 ( .gnd(gnd), .vdd(vdd), .A(_98__9_), .B(_8845_), .C(_93__9_), .D(_8840_), .Y(_12480_) );
AOI22X1 AOI22X1_348 ( .gnd(gnd), .vdd(vdd), .A(_94__9_), .B(_8841_), .C(_91__9_), .D(_8823_), .Y(_12481_) );
NAND2X1 NAND2X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_12480_), .B(_12481_), .Y(_12482_) );
NAND2X1 NAND2X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__9_), .Y(_12483_) );
NAND2X1 NAND2X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__9_), .Y(_12484_) );
NAND2X1 NAND2X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__9_), .Y(_12485_) );
NAND2X1 NAND2X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_12484_), .B(_12485_), .Y(_12486_) );
NAND2X1 NAND2X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__9_), .Y(_12487_) );
NAND2X1 NAND2X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__9_), .Y(_12488_) );
NAND2X1 NAND2X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_12487_), .B(_12488_), .Y(_12489_) );
NOR2X1 NOR2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_12486_), .B(_12489_), .Y(_12490_) );
NAND2X1 NAND2X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__9_), .Y(_12491_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_7147_), .B(_9930_), .C(_7191_), .D(_9929_), .Y(_12492_) );
NOR2X1 NOR2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7326_), .Y(_12493_) );
NOR2X1 NOR2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7283_), .Y(_12494_) );
NOR3X1 NOR3X1_355 ( .gnd(gnd), .vdd(vdd), .A(_12493_), .B(_12494_), .C(_12492_), .Y(_12495_) );
NAND2X1 NAND2X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__9_), .Y(_12496_) );
NAND2X1 NAND2X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__9_), .Y(_12497_) );
NAND2X1 NAND2X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_12496_), .B(_12497_), .Y(_12498_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_7369_), .B(_9940_), .C(_7237_), .D(_9941_), .Y(_12499_) );
NOR2X1 NOR2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_12499_), .B(_12498_), .Y(_12500_) );
NAND3X1 NAND3X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_12491_), .B(_12495_), .C(_12500_), .Y(_12501_) );
AOI22X1 AOI22X1_349 ( .gnd(gnd), .vdd(vdd), .A(_20__9_), .B(_8898_), .C(_236__9_), .D(_8955_), .Y(_12502_) );
AOI22X1 AOI22X1_350 ( .gnd(gnd), .vdd(vdd), .A(_237__9_), .B(_8966_), .C(_175__9_), .D(_8904_), .Y(_12503_) );
NAND2X1 NAND2X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_12502_), .B(_12503_), .Y(_12504_) );
NAND2X1 NAND2X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__9_), .Y(_12505_) );
NAND2X1 NAND2X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__9_), .Y(_12506_) );
AOI22X1 AOI22X1_351 ( .gnd(gnd), .vdd(vdd), .A(_19__9_), .B(_8914_), .C(_210__9_), .D(_8918_), .Y(_12507_) );
NAND3X1 NAND3X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_12505_), .B(_12506_), .C(_12507_), .Y(_12508_) );
NOR2X1 NOR2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_12504_), .B(_12508_), .Y(_12509_) );
AOI22X1 AOI22X1_352 ( .gnd(gnd), .vdd(vdd), .A(_123__9_), .B(_8928_), .C(_9__9_), .D(_8926_), .Y(_12510_) );
NAND2X1 NAND2X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__9_), .Y(_12511_) );
NAND2X1 NAND2X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_134__9_), .Y(_12512_) );
NAND3X1 NAND3X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_12511_), .B(_12512_), .C(_12510_), .Y(_12513_) );
AOI22X1 AOI22X1_353 ( .gnd(gnd), .vdd(vdd), .A(_4__9_), .B(_8937_), .C(_176__9_), .D(_8939_), .Y(_12514_) );
NAND2X1 NAND2X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__9_), .Y(_12515_) );
NAND2X1 NAND2X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__9_), .Y(_12516_) );
NAND3X1 NAND3X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_12515_), .B(_12516_), .C(_12514_), .Y(_12517_) );
NOR2X1 NOR2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_12517_), .B(_12513_), .Y(_12518_) );
NAND2X1 NAND2X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_12509_), .B(_12518_), .Y(_12519_) );
NAND2X1 NAND2X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_208__9_), .Y(_12520_) );
NAND2X1 NAND2X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_8952_), .B(_40__9_), .Y(_12521_) );
AOI22X1 AOI22X1_354 ( .gnd(gnd), .vdd(vdd), .A(_238__9_), .B(_8893_), .C(_209__9_), .D(_8957_), .Y(_12522_) );
NAND3X1 NAND3X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_12520_), .B(_12521_), .C(_12522_), .Y(_12523_) );
AOI22X1 AOI22X1_355 ( .gnd(gnd), .vdd(vdd), .A(_42__9_), .B(_8963_), .C(_177__9_), .D(_8961_), .Y(_12524_) );
NAND2X1 NAND2X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_8901_), .B(_248__9_), .Y(_12525_) );
NAND2X1 NAND2X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_8968_), .B(_44__9_), .Y(_12526_) );
NAND3X1 NAND3X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_12525_), .B(_12526_), .C(_12524_), .Y(_12527_) );
NOR2X1 NOR2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_12523_), .B(_12527_), .Y(_12528_) );
NAND2X1 NAND2X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_8986_), .B(_255__9_), .Y(_12529_) );
NAND2X1 NAND2X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_9084_), .B(_43__9_), .Y(_12530_) );
AOI22X1 AOI22X1_356 ( .gnd(gnd), .vdd(vdd), .A(_48__9_), .B(_9089_), .C(_244__9_), .D(_9160_), .Y(_12531_) );
NAND3X1 NAND3X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_12529_), .B(_12530_), .C(_12531_), .Y(_12532_) );
NAND2X1 NAND2X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_8984_), .B(_254__9_), .Y(_12533_) );
NAND2X1 NAND2X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(_33__9_), .Y(_12534_) );
AOI22X1 AOI22X1_357 ( .gnd(gnd), .vdd(vdd), .A(_203__9_), .B(_9018_), .C(_156__9_), .D(_8973_), .Y(_12535_) );
NAND3X1 NAND3X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_12533_), .B(_12534_), .C(_12535_), .Y(_12536_) );
NOR2X1 NOR2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_12532_), .B(_12536_), .Y(_12537_) );
NAND2X1 NAND2X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_12528_), .B(_12537_), .Y(_12538_) );
NOR2X1 NOR2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_12519_), .B(_12538_), .Y(_12539_) );
NAND2X1 NAND2X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__9_), .Y(_12540_) );
NAND2X1 NAND2X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__9_), .Y(_12541_) );
AOI22X1 AOI22X1_358 ( .gnd(gnd), .vdd(vdd), .A(_13__9_), .B(_9007_), .C(_239__9_), .D(_9076_), .Y(_12542_) );
NAND3X1 NAND3X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_12540_), .B(_12541_), .C(_12542_), .Y(_12543_) );
AOI22X1 AOI22X1_359 ( .gnd(gnd), .vdd(vdd), .A(_206__9_), .B(_9013_), .C(_242__9_), .D(_9035_), .Y(_12544_) );
NAND2X1 NAND2X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__9_), .Y(_12545_) );
NAND2X1 NAND2X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__9_), .Y(_12546_) );
NAND3X1 NAND3X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_12545_), .B(_12546_), .C(_12544_), .Y(_12547_) );
NOR2X1 NOR2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_12543_), .B(_12547_), .Y(_12548_) );
AOI22X1 AOI22X1_360 ( .gnd(gnd), .vdd(vdd), .A(_222__9_), .B(_9024_), .C(_220__9_), .D(_9026_), .Y(_12549_) );
NAND2X1 NAND2X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__9_), .Y(_12550_) );
NAND2X1 NAND2X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__9_), .Y(_12551_) );
NAND3X1 NAND3X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_12550_), .B(_12551_), .C(_12549_), .Y(_12552_) );
AOI22X1 AOI22X1_361 ( .gnd(gnd), .vdd(vdd), .A(_18__9_), .B(_9037_), .C(_240__9_), .D(_9011_), .Y(_12553_) );
NAND2X1 NAND2X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__9_), .Y(_12554_) );
NAND2X1 NAND2X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__9_), .Y(_12555_) );
NAND3X1 NAND3X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_12554_), .B(_12555_), .C(_12553_), .Y(_12556_) );
NOR2X1 NOR2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_12552_), .B(_12556_), .Y(_12557_) );
NAND2X1 NAND2X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_12548_), .B(_12557_), .Y(_12558_) );
AOI22X1 AOI22X1_362 ( .gnd(gnd), .vdd(vdd), .A(_225__9_), .B(_9048_), .C(_167__9_), .D(_9050_), .Y(_12559_) );
NAND2X1 NAND2X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__9_), .Y(_12560_) );
NAND2X1 NAND2X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_8980_), .B(_35__9_), .Y(_12561_) );
NAND3X1 NAND3X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_12560_), .B(_12561_), .C(_12559_), .Y(_12562_) );
NAND2X1 NAND2X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__9_), .Y(_12563_) );
NAND2X1 NAND2X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__9_), .Y(_12564_) );
AOI22X1 AOI22X1_363 ( .gnd(gnd), .vdd(vdd), .A(_224__9_), .B(_9064_), .C(_27__9_), .D(_9066_), .Y(_12565_) );
NAND3X1 NAND3X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_12563_), .B(_12564_), .C(_12565_), .Y(_12566_) );
NOR2X1 NOR2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_12562_), .B(_12566_), .Y(_12567_) );
AOI22X1 AOI22X1_364 ( .gnd(gnd), .vdd(vdd), .A(_184__9_), .B(_9073_), .C(_183__9_), .D(_9071_), .Y(_12568_) );
NAND2X1 NAND2X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__9_), .Y(_12569_) );
NAND2X1 NAND2X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__9_), .Y(_12570_) );
NAND3X1 NAND3X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_12569_), .B(_12570_), .C(_12568_), .Y(_12571_) );
AOI22X1 AOI22X1_365 ( .gnd(gnd), .vdd(vdd), .A(_243__9_), .B(_9153_), .C(_36__9_), .D(_8909_), .Y(_12572_) );
NAND2X1 NAND2X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__9_), .Y(_12573_) );
NAND2X1 NAND2X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_8978_), .B(_37__9_), .Y(_12574_) );
NAND3X1 NAND3X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_12573_), .B(_12574_), .C(_12572_), .Y(_12575_) );
NOR2X1 NOR2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_12571_), .B(_12575_), .Y(_12576_) );
NAND2X1 NAND2X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_12567_), .B(_12576_), .Y(_12577_) );
NOR2X1 NOR2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_12558_), .B(_12577_), .Y(_12578_) );
NAND3X1 NAND3X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_6860_), .B(_9104_), .C(_6861_), .Y(_12579_) );
NAND3X1 NAND3X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_9099_), .C(_3969_), .Y(_12580_) );
NAND2X1 NAND2X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_12579_), .B(_12580_), .Y(_12581_) );
NAND2X1 NAND2X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__9_), .Y(_12582_) );
NAND3X1 NAND3X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_5101_), .B(_9102_), .C(_5102_), .Y(_12583_) );
NAND2X1 NAND2X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_12583_), .B(_12582_), .Y(_12584_) );
NOR2X1 NOR2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_12581_), .B(_12584_), .Y(_12585_) );
NAND3X1 NAND3X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_8322_), .B(_9188_), .C(_8323_), .Y(_12586_) );
NAND3X1 NAND3X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_15929_), .B(_9109_), .C(_15930_), .Y(_12587_) );
NAND3X1 NAND3X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_16135_), .B(_9115_), .C(_16136_), .Y(_12588_) );
NAND3X1 NAND3X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_12587_), .B(_12588_), .C(_12586_), .Y(_12589_) );
AOI22X1 AOI22X1_366 ( .gnd(gnd), .vdd(vdd), .A(_234__9_), .B(_9182_), .C(_34__9_), .D(_9183_), .Y(_12590_) );
AOI22X1 AOI22X1_367 ( .gnd(gnd), .vdd(vdd), .A(_100__9_), .B(_9346_), .C(_45__9_), .D(_9185_), .Y(_12591_) );
NAND2X1 NAND2X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_12591_), .B(_12590_), .Y(_12592_) );
NAND3X1 NAND3X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(_9127_), .C(_4746_), .Y(_12593_) );
NAND3X1 NAND3X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_4011_), .B(_9129_), .C(_4012_), .Y(_12594_) );
NAND2X1 NAND2X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_12593_), .B(_12594_), .Y(_12595_) );
NOR3X1 NOR3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_12589_), .B(_12595_), .C(_12592_), .Y(_12596_) );
NAND3X1 NAND3X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_3428_), .B(_9133_), .C(_3429_), .Y(_12597_) );
NAND3X1 NAND3X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_5054_), .B(_9135_), .C(_5055_), .Y(_12598_) );
NAND3X1 NAND3X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_6937_), .B(_9137_), .C(_6938_), .Y(_12599_) );
NAND3X1 NAND3X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_12598_), .B(_12599_), .C(_12597_), .Y(_12600_) );
AOI22X1 AOI22X1_368 ( .gnd(gnd), .vdd(vdd), .A(_17__9_), .B(_9140_), .C(_2__9_), .D(_9141_), .Y(_12601_) );
AOI22X1 AOI22X1_369 ( .gnd(gnd), .vdd(vdd), .A(_205__9_), .B(_9143_), .C(_200__9_), .D(_9145_), .Y(_12602_) );
NAND2X1 NAND2X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_12601_), .B(_12602_), .Y(_12603_) );
NOR2X1 NOR2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_12600_), .B(_12603_), .Y(_12604_) );
NAND3X1 NAND3X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_12585_), .B(_12596_), .C(_12604_), .Y(_12605_) );
AOI22X1 AOI22X1_370 ( .gnd(gnd), .vdd(vdd), .A(_21__9_), .B(_9150_), .C(_185__9_), .D(_9151_), .Y(_12606_) );
AOI22X1 AOI22X1_371 ( .gnd(gnd), .vdd(vdd), .A(_249__9_), .B(_9053_), .C(_253__9_), .D(_9154_), .Y(_12607_) );
NAND2X1 NAND2X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_12606_), .B(_12607_), .Y(_12608_) );
AOI22X1 AOI22X1_372 ( .gnd(gnd), .vdd(vdd), .A(_46__9_), .B(_9158_), .C(_231__9_), .D(_9157_), .Y(_12609_) );
AOI22X1 AOI22X1_373 ( .gnd(gnd), .vdd(vdd), .A(_47__9_), .B(_9161_), .C(_250__9_), .D(_9082_), .Y(_12610_) );
NAND2X1 NAND2X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_12610_), .B(_12609_), .Y(_12611_) );
NOR2X1 NOR2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_12608_), .B(_12611_), .Y(_12612_) );
AOI22X1 AOI22X1_374 ( .gnd(gnd), .vdd(vdd), .A(_247__9_), .B(_9165_), .C(_30__9_), .D(_9167_), .Y(_12613_) );
AOI22X1 AOI22X1_375 ( .gnd(gnd), .vdd(vdd), .A(_227__9_), .B(_9170_), .C(_218__9_), .D(_9169_), .Y(_12614_) );
NAND2X1 NAND2X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_12613_), .B(_12614_), .Y(_12615_) );
AOI22X1 AOI22X1_376 ( .gnd(gnd), .vdd(vdd), .A(_145__9_), .B(_9177_), .C(_213__9_), .D(_8989_), .Y(_12616_) );
AOI22X1 AOI22X1_377 ( .gnd(gnd), .vdd(vdd), .A(_29__9_), .B(_9176_), .C(_178__9_), .D(_9173_), .Y(_12617_) );
NAND2X1 NAND2X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_12616_), .B(_12617_), .Y(_12618_) );
NOR2X1 NOR2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_12615_), .B(_12618_), .Y(_12619_) );
NAND2X1 NAND2X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_12612_), .B(_12619_), .Y(_12620_) );
AOI22X1 AOI22X1_378 ( .gnd(gnd), .vdd(vdd), .A(_201__9_), .B(_9124_), .C(_212__9_), .D(_9345_), .Y(_12621_) );
NAND3X1 NAND3X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_8436_), .B(_9348_), .C(_8435_), .Y(_12622_) );
NAND3X1 NAND3X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_496_), .C(_497_), .Y(_12623_) );
AND2X2 AND2X2_1591 ( .gnd(gnd), .vdd(vdd), .A(_12623_), .B(_12622_), .Y(_12624_) );
NAND2X1 NAND2X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_12621_), .B(_12624_), .Y(_12625_) );
NAND3X1 NAND3X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_15142_), .B(_9208_), .C(_15143_), .Y(_12626_) );
OAI21X1 OAI21X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_15106_), .B(_9211_), .C(_12626_), .Y(_12627_) );
NAND3X1 NAND3X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_15486_), .B(_9222_), .C(_15487_), .Y(_12628_) );
NAND3X1 NAND3X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_15433_), .B(_9224_), .C(_15432_), .Y(_12629_) );
NAND2X1 NAND2X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_12628_), .B(_12629_), .Y(_12630_) );
NOR2X1 NOR2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_12630_), .B(_12627_), .Y(_12631_) );
NAND3X1 NAND3X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_15264_), .B(_9217_), .C(_15265_), .Y(_12632_) );
NAND3X1 NAND3X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_15212_), .B(_9219_), .C(_15211_), .Y(_12633_) );
NAND2X1 NAND2X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_12633_), .B(_12632_), .Y(_12634_) );
NAND3X1 NAND3X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_15662_), .B(_9192_), .C(_15663_), .Y(_12635_) );
NAND3X1 NAND3X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_15719_), .B(_9199_), .C(_15718_), .Y(_12636_) );
NAND2X1 NAND2X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_12636_), .B(_12635_), .Y(_12637_) );
NOR2X1 NOR2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_12637_), .B(_12634_), .Y(_12638_) );
NOR3X1 NOR3X1_357 ( .gnd(gnd), .vdd(vdd), .A(_16188_), .B(_10083_), .C(_16189_), .Y(_12639_) );
NAND3X1 NAND3X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_15314_), .B(_9205_), .C(_15315_), .Y(_12640_) );
OAI21X1 OAI21X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_15348_), .B(_10085_), .C(_12640_), .Y(_12641_) );
NAND3X1 NAND3X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_15544_), .B(_9233_), .C(_15545_), .Y(_12642_) );
NAND3X1 NAND3X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15612_), .C(_15611_), .Y(_12643_) );
NAND2X1 NAND2X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_12642_), .B(_12643_), .Y(_12644_) );
NOR3X1 NOR3X1_358 ( .gnd(gnd), .vdd(vdd), .A(_12641_), .B(_12644_), .C(_12639_), .Y(_12645_) );
NAND3X1 NAND3X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_12631_), .B(_12638_), .C(_12645_), .Y(_12646_) );
NAND3X1 NAND3X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_15872_), .B(_9120_), .C(_15873_), .Y(_12647_) );
NAND3X1 NAND3X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_15383_), .B(_9197_), .C(_15384_), .Y(_12648_) );
NAND2X1 NAND2X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__9_), .Y(_12649_) );
NAND2X1 NAND2X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__9_), .Y(_12650_) );
NAND2X1 NAND2X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .B(_186__9_), .Y(_12651_) );
NAND3X1 NAND3X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_12651_), .B(_12650_), .C(_12649_), .Y(_12652_) );
NAND2X1 NAND2X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__9_), .Y(_12653_) );
NAND2X1 NAND2X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_9294_), .B(_49__9_), .Y(_12654_) );
AOI22X1 AOI22X1_379 ( .gnd(gnd), .vdd(vdd), .A(_198__9_), .B(_9266_), .C(_119__9_), .D(_9268_), .Y(_12655_) );
NAND3X1 NAND3X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_12653_), .B(_12654_), .C(_12655_), .Y(_12656_) );
NAND2X1 NAND2X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_9250_), .B(_56__9_), .Y(_12657_) );
NAND2X1 NAND2X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_101__9_), .Y(_12658_) );
AOI22X1 AOI22X1_380 ( .gnd(gnd), .vdd(vdd), .A(_173__9_), .B(_9275_), .C(_137__9_), .D(_9262_), .Y(_12659_) );
NAND3X1 NAND3X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_12657_), .B(_12658_), .C(_12659_), .Y(_12660_) );
NOR3X1 NOR3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_12660_), .B(_12652_), .C(_12656_), .Y(_12661_) );
NAND2X1 NAND2X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_181__9_), .Y(_12662_) );
AOI22X1 AOI22X1_381 ( .gnd(gnd), .vdd(vdd), .A(_32__9_), .B(_10110_), .C(_187__9_), .D(_9235_), .Y(_12663_) );
AOI22X1 AOI22X1_382 ( .gnd(gnd), .vdd(vdd), .A(_83__9_), .B(_9315_), .C(_235__9_), .D(_9324_), .Y(_12664_) );
NAND3X1 NAND3X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_12662_), .B(_12663_), .C(_12664_), .Y(_12665_) );
NAND3X1 NAND3X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_7722_), .B(_9248_), .C(_7721_), .Y(_12666_) );
OAI21X1 OAI21X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_8170_), .B(_9304_), .C(_12666_), .Y(_12667_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_7637_), .B(_9301_), .C(_9765_), .D(_8713_), .Y(_12668_) );
NOR2X1 NOR2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_12667_), .B(_12668_), .Y(_12669_) );
AOI22X1 AOI22X1_383 ( .gnd(gnd), .vdd(vdd), .A(_154__9_), .B(_9292_), .C(_50__9_), .D(_9778_), .Y(_12670_) );
AOI22X1 AOI22X1_384 ( .gnd(gnd), .vdd(vdd), .A(_65__9_), .B(_9277_), .C(_197__9_), .D(_9244_), .Y(_12671_) );
NAND3X1 NAND3X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_12670_), .B(_12671_), .C(_12669_), .Y(_12672_) );
NOR2X1 NOR2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .B(_4819_), .Y(_12673_) );
NOR2X1 NOR2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_9319_), .B(_5406_), .Y(_12674_) );
NOR2X1 NOR2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .B(_4225_), .Y(_12675_) );
NOR3X1 NOR3X1_360 ( .gnd(gnd), .vdd(vdd), .A(_12673_), .B(_12675_), .C(_12674_), .Y(_12676_) );
AOI22X1 AOI22X1_385 ( .gnd(gnd), .vdd(vdd), .A(_217__9_), .B(_9281_), .C(_252__9_), .D(_9326_), .Y(_12677_) );
AOI22X1 AOI22X1_386 ( .gnd(gnd), .vdd(vdd), .A(_15__9_), .B(_9313_), .C(_233__9_), .D(_9310_), .Y(_12678_) );
NAND3X1 NAND3X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_12676_), .B(_12677_), .C(_12678_), .Y(_12679_) );
NOR3X1 NOR3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_12672_), .B(_12665_), .C(_12679_), .Y(_12680_) );
NAND3X1 NAND3X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_12661_), .B(_12648_), .C(_12680_), .Y(_12681_) );
AOI21X1 AOI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_157__9_), .B(_9232_), .C(_12681_), .Y(_12682_) );
AOI22X1 AOI22X1_387 ( .gnd(gnd), .vdd(vdd), .A(_155__9_), .B(_9333_), .C(_172__9_), .D(_9332_), .Y(_12683_) );
NAND3X1 NAND3X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_12647_), .B(_12683_), .C(_12682_), .Y(_12684_) );
NOR3X1 NOR3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_12646_), .B(_12684_), .C(_12625_), .Y(_12685_) );
AOI22X1 AOI22X1_388 ( .gnd(gnd), .vdd(vdd), .A(_256__9_), .B(_9113_), .C(_142__9_), .D(_9118_), .Y(_12686_) );
NAND2X1 NAND2X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__9_), .Y(_12687_) );
NAND2X1 NAND2X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__9_), .Y(_12688_) );
NAND3X1 NAND3X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_12687_), .B(_12688_), .C(_12686_), .Y(_12689_) );
NAND2X1 NAND2X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__9_), .Y(_12690_) );
NAND3X1 NAND3X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_9339_), .C(_455_), .Y(_12691_) );
AOI22X1 AOI22X1_389 ( .gnd(gnd), .vdd(vdd), .A(_111__9_), .B(_9342_), .C(_12__9_), .D(_9341_), .Y(_12692_) );
NAND3X1 NAND3X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_12692_), .B(_12690_), .C(_12691_), .Y(_12693_) );
NOR2X1 NOR2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_12689_), .B(_12693_), .Y(_12694_) );
AOI22X1 AOI22X1_390 ( .gnd(gnd), .vdd(vdd), .A(_232__9_), .B(_9354_), .C(_219__9_), .D(_9353_), .Y(_12695_) );
AOI22X1 AOI22X1_391 ( .gnd(gnd), .vdd(vdd), .A(_246__9_), .B(_9356_), .C(_226__9_), .D(_9357_), .Y(_12696_) );
NAND2X1 NAND2X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_12695_), .B(_12696_), .Y(_12697_) );
NAND3X1 NAND3X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16089_), .C(_16090_), .Y(_12698_) );
NAND3X1 NAND3X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16034_), .C(_16035_), .Y(_12699_) );
NAND2X1 NAND2X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_12698_), .B(_12699_), .Y(_12700_) );
NAND3X1 NAND3X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8568_), .C(_8567_), .Y(_12701_) );
OAI21X1 OAI21X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_9361_), .C(_12701_), .Y(_12702_) );
NOR2X1 NOR2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_12700_), .B(_12702_), .Y(_12703_) );
NAND2X1 NAND2X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_15980_), .B(_15981_), .Y(_12704_) );
NAND3X1 NAND3X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8621_), .C(_8622_), .Y(_12705_) );
OAI21X1 OAI21X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_12704_), .B(_9215_), .C(_12705_), .Y(_12706_) );
NAND3X1 NAND3X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_8676_), .B(_9371_), .C(_8675_), .Y(_12707_) );
NAND3X1 NAND3X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_318_), .C(_319_), .Y(_12708_) );
NAND2X1 NAND2X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_12708_), .B(_12707_), .Y(_12709_) );
NOR2X1 NOR2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_12706_), .B(_12709_), .Y(_12710_) );
AOI22X1 AOI22X1_392 ( .gnd(gnd), .vdd(vdd), .A(_22__9_), .B(_9382_), .C(_3__9_), .D(_9383_), .Y(_12711_) );
NAND3X1 NAND3X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_12703_), .B(_12710_), .C(_12711_), .Y(_12712_) );
NOR2X1 NOR2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_12697_), .B(_12712_), .Y(_12713_) );
NAND3X1 NAND3X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_12685_), .B(_12694_), .C(_12713_), .Y(_12714_) );
NOR3X1 NOR3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_12605_), .B(_12620_), .C(_12714_), .Y(_12715_) );
NAND3X1 NAND3X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_12539_), .B(_12578_), .C(_12715_), .Y(_12716_) );
NAND3X1 NAND3X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1587_), .C(_1588_), .Y(_12717_) );
NAND3X1 NAND3X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_8862_), .C(_1249_), .Y(_12718_) );
NAND2X1 NAND2X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_12717_), .B(_12718_), .Y(_12719_) );
NOR3X1 NOR3X1_364 ( .gnd(gnd), .vdd(vdd), .A(_12501_), .B(_12719_), .C(_12716_), .Y(_12720_) );
NAND3X1 NAND3X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_12483_), .B(_12490_), .C(_12720_), .Y(_12721_) );
NAND2X1 NAND2X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__9_), .Y(_12722_) );
NAND3X1 NAND3X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_9406_), .C(_1464_), .Y(_12723_) );
NAND3X1 NAND3X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_9453_), .C(_1418_), .Y(_12724_) );
AND2X2 AND2X2_1592 ( .gnd(gnd), .vdd(vdd), .A(_12723_), .B(_12724_), .Y(_12725_) );
NAND2X1 NAND2X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_108__9_), .Y(_12726_) );
NAND2X1 NAND2X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_116__9_), .Y(_12727_) );
NAND3X1 NAND3X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_12726_), .B(_12727_), .C(_12725_), .Y(_12728_) );
AOI22X1 AOI22X1_393 ( .gnd(gnd), .vdd(vdd), .A(_125__9_), .B(_9411_), .C(_124__9_), .D(_9410_), .Y(_12729_) );
AOI22X1 AOI22X1_394 ( .gnd(gnd), .vdd(vdd), .A(_120__9_), .B(_9415_), .C(_121__9_), .D(_9413_), .Y(_12730_) );
AND2X2 AND2X2_1593 ( .gnd(gnd), .vdd(vdd), .A(_12730_), .B(_12729_), .Y(_12731_) );
AOI22X1 AOI22X1_395 ( .gnd(gnd), .vdd(vdd), .A(_132__9_), .B(_9420_), .C(_131__9_), .D(_9418_), .Y(_12732_) );
NAND2X1 NAND2X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__9_), .Y(_12733_) );
NAND2X1 NAND2X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__9_), .Y(_12734_) );
NAND3X1 NAND3X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_12733_), .B(_12734_), .C(_12732_), .Y(_12735_) );
NAND3X1 NAND3X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_9431_), .C(_550_), .Y(_12736_) );
NAND2X1 NAND2X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__9_), .Y(_12737_) );
NAND2X1 NAND2X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__9_), .Y(_12738_) );
NAND3X1 NAND3X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_12738_), .B(_12736_), .C(_12737_), .Y(_12739_) );
AOI21X1 AOI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_136__9_), .B(_9429_), .C(_12739_), .Y(_12740_) );
NAND2X1 NAND2X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__9_), .Y(_12741_) );
NAND2X1 NAND2X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__9_), .Y(_12742_) );
NAND3X1 NAND3X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_12741_), .B(_12742_), .C(_12740_), .Y(_12743_) );
NAND3X1 NAND3X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_9444_), .C(_1057_), .Y(_12744_) );
NAND2X1 NAND2X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__9_), .Y(_12745_) );
AOI22X1 AOI22X1_396 ( .gnd(gnd), .vdd(vdd), .A(_130__9_), .B(_9449_), .C(_127__9_), .D(_9448_), .Y(_12746_) );
NAND3X1 NAND3X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_12744_), .B(_12746_), .C(_12745_), .Y(_12747_) );
NOR3X1 NOR3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_12735_), .B(_12743_), .C(_12747_), .Y(_12748_) );
AOI22X1 AOI22X1_397 ( .gnd(gnd), .vdd(vdd), .A(_115__9_), .B(_9399_), .C(_114__9_), .D(_9454_), .Y(_12749_) );
NAND3X1 NAND3X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_12749_), .B(_12731_), .C(_12748_), .Y(_12750_) );
NOR2X1 NOR2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_12728_), .B(_12750_), .Y(_12751_) );
AOI22X1 AOI22X1_398 ( .gnd(gnd), .vdd(vdd), .A(_102__9_), .B(_9459_), .C(_103__9_), .D(_9457_), .Y(_12752_) );
NAND3X1 NAND3X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_12722_), .B(_12752_), .C(_12751_), .Y(_12753_) );
NOR3X1 NOR3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_12482_), .B(_12753_), .C(_12721_), .Y(_12754_) );
NAND3X1 NAND3X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_12472_), .B(_12479_), .C(_12754_), .Y(_12755_) );
NAND2X1 NAND2X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__9_), .Y(_12756_) );
NAND3X1 NAND3X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .B(_8806_), .C(_2405_), .Y(_12757_) );
NAND2X1 NAND2X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_12757_), .B(_12756_), .Y(_12758_) );
NOR3X1 NOR3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_12464_), .B(_12758_), .C(_12755_), .Y(_12759_) );
NAND3X1 NAND3X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_12456_), .B(_12461_), .C(_12759_), .Y(_12760_) );
NAND3X1 NAND3X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_3067_), .B(_9473_), .C(_3068_), .Y(_12761_) );
NAND2X1 NAND2X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__9_), .Y(_12762_) );
NAND2X1 NAND2X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__9_), .Y(_12763_) );
NAND2X1 NAND2X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__9_), .Y(_12764_) );
NAND2X1 NAND2X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__9_), .Y(_12765_) );
NAND3X1 NAND3X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_12763_), .B(_12764_), .C(_12765_), .Y(_12766_) );
AOI21X1 AOI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_68__9_), .B(_9477_), .C(_12766_), .Y(_12767_) );
NAND3X1 NAND3X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_12761_), .B(_12767_), .C(_12762_), .Y(_12768_) );
NOR3X1 NOR3X1_368 ( .gnd(gnd), .vdd(vdd), .A(_12455_), .B(_12768_), .C(_12760_), .Y(_12769_) );
AOI21X1 AOI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_12448_), .B(_12769_), .C(rst), .Y(_0__9_) );
NAND2X1 NAND2X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__10_), .Y(_12770_) );
NAND2X1 NAND2X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__10_), .Y(_12771_) );
NAND2X1 NAND2X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_12770_), .B(_12771_), .Y(_12772_) );
NAND2X1 NAND2X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__10_), .Y(_12773_) );
NAND2X1 NAND2X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__10_), .Y(_12774_) );
NAND2X1 NAND2X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_12773_), .B(_12774_), .Y(_12775_) );
NOR2X1 NOR2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_12772_), .B(_12775_), .Y(_12776_) );
NAND3X1 NAND3X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_3287_), .B(_8762_), .C(_3286_), .Y(_12777_) );
NAND3X1 NAND3X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_3239_), .B(_8765_), .C(_3238_), .Y(_12778_) );
AND2X2 AND2X2_1594 ( .gnd(gnd), .vdd(vdd), .A(_12778_), .B(_12777_), .Y(_12779_) );
AOI22X1 AOI22X1_399 ( .gnd(gnd), .vdd(vdd), .A(_62__10_), .B(_8774_), .C(_57__10_), .D(_8771_), .Y(_12780_) );
NAND2X1 NAND2X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_12779_), .B(_12780_), .Y(_12781_) );
NAND2X1 NAND2X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__10_), .Y(_12782_) );
NAND3X1 NAND3X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(_8786_), .C(_2825_), .Y(_12783_) );
OAI21X1 OAI21X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_8792_), .C(_12783_), .Y(_12784_) );
NAND3X1 NAND3X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_8794_), .C(_2654_), .Y(_12785_) );
OAI21X1 OAI21X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_8799_), .C(_12785_), .Y(_12786_) );
NOR2X1 NOR2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_12786_), .B(_12784_), .Y(_12787_) );
AOI22X1 AOI22X1_400 ( .gnd(gnd), .vdd(vdd), .A(_76__10_), .B(_9482_), .C(_77__10_), .D(_9478_), .Y(_12788_) );
NAND2X1 NAND2X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__10_), .Y(_12789_) );
NAND2X1 NAND2X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_82__10_), .Y(_12790_) );
NAND3X1 NAND3X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_12789_), .B(_12790_), .C(_12788_), .Y(_12791_) );
NAND2X1 NAND2X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__10_), .Y(_12792_) );
NAND3X1 NAND3X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .B(_8803_), .C(_2588_), .Y(_12793_) );
NAND2X1 NAND2X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_12793_), .B(_12792_), .Y(_12794_) );
INVX1 INVX1_3879 ( .gnd(gnd), .vdd(vdd), .A(_84__10_), .Y(_12795_) );
NOR2X1 NOR2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_12795_), .Y(_12796_) );
NOR2X1 NOR2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2302_), .Y(_12797_) );
NAND2X1 NAND2X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__10_), .Y(_12798_) );
NAND3X1 NAND3X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_8843_), .C(_2018_), .Y(_12799_) );
NAND3X1 NAND3X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1922_), .C(_1923_), .Y(_12800_) );
NAND3X1 NAND3X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_12800_), .B(_12799_), .C(_12798_), .Y(_12801_) );
NOR3X1 NOR3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_12796_), .B(_12801_), .C(_12797_), .Y(_12802_) );
NAND3X1 NAND3X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_2260_), .B(_8829_), .C(_2261_), .Y(_12803_) );
NAND3X1 NAND3X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_2154_), .B(_8831_), .C(_2155_), .Y(_12804_) );
NAND2X1 NAND2X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_12803_), .B(_12804_), .Y(_12805_) );
NAND3X1 NAND3X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_2095_), .B(_8834_), .C(_2096_), .Y(_12806_) );
NAND3X1 NAND3X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_2206_), .B(_8836_), .C(_2207_), .Y(_12807_) );
NAND2X1 NAND2X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_12806_), .B(_12807_), .Y(_12808_) );
NOR2X1 NOR2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_12808_), .B(_12805_), .Y(_12809_) );
AOI22X1 AOI22X1_401 ( .gnd(gnd), .vdd(vdd), .A(_98__10_), .B(_8845_), .C(_93__10_), .D(_8840_), .Y(_12810_) );
AOI22X1 AOI22X1_402 ( .gnd(gnd), .vdd(vdd), .A(_94__10_), .B(_8841_), .C(_91__10_), .D(_8823_), .Y(_12811_) );
NAND2X1 NAND2X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_12810_), .B(_12811_), .Y(_12812_) );
NAND2X1 NAND2X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__10_), .Y(_12813_) );
NAND2X1 NAND2X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__10_), .Y(_12814_) );
NAND2X1 NAND2X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__10_), .Y(_12815_) );
NAND2X1 NAND2X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_12814_), .B(_12815_), .Y(_12816_) );
NAND2X1 NAND2X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__10_), .Y(_12817_) );
NAND2X1 NAND2X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__10_), .Y(_12818_) );
NAND2X1 NAND2X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_12817_), .B(_12818_), .Y(_12819_) );
NOR2X1 NOR2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_12816_), .B(_12819_), .Y(_12820_) );
NAND2X1 NAND2X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__10_), .Y(_12821_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_7150_), .B(_9930_), .C(_7194_), .D(_9929_), .Y(_12822_) );
NOR2X1 NOR2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7329_), .Y(_12823_) );
NOR2X1 NOR2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7286_), .Y(_12824_) );
NOR3X1 NOR3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_12823_), .B(_12824_), .C(_12822_), .Y(_12825_) );
NAND2X1 NAND2X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__10_), .Y(_12826_) );
NAND2X1 NAND2X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__10_), .Y(_12827_) );
NAND2X1 NAND2X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_12826_), .B(_12827_), .Y(_12828_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_7372_), .B(_9940_), .C(_7240_), .D(_9941_), .Y(_12829_) );
NOR2X1 NOR2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_12829_), .B(_12828_), .Y(_12830_) );
NAND3X1 NAND3X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_12821_), .B(_12825_), .C(_12830_), .Y(_12831_) );
AOI22X1 AOI22X1_403 ( .gnd(gnd), .vdd(vdd), .A(_20__10_), .B(_8898_), .C(_236__10_), .D(_8955_), .Y(_12832_) );
AOI22X1 AOI22X1_404 ( .gnd(gnd), .vdd(vdd), .A(_237__10_), .B(_8966_), .C(_175__10_), .D(_8904_), .Y(_12833_) );
NAND2X1 NAND2X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_12832_), .B(_12833_), .Y(_12834_) );
NAND2X1 NAND2X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__10_), .Y(_12835_) );
NAND2X1 NAND2X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__10_), .Y(_12836_) );
AOI22X1 AOI22X1_405 ( .gnd(gnd), .vdd(vdd), .A(_19__10_), .B(_8914_), .C(_210__10_), .D(_8918_), .Y(_12837_) );
NAND3X1 NAND3X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_12835_), .B(_12836_), .C(_12837_), .Y(_12838_) );
NOR2X1 NOR2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_12834_), .B(_12838_), .Y(_12839_) );
AOI22X1 AOI22X1_406 ( .gnd(gnd), .vdd(vdd), .A(_123__10_), .B(_8928_), .C(_9__10_), .D(_8926_), .Y(_12840_) );
NAND2X1 NAND2X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__10_), .Y(_12841_) );
NAND2X1 NAND2X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_134__10_), .Y(_12842_) );
NAND3X1 NAND3X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_12841_), .B(_12842_), .C(_12840_), .Y(_12843_) );
AOI22X1 AOI22X1_407 ( .gnd(gnd), .vdd(vdd), .A(_4__10_), .B(_8937_), .C(_176__10_), .D(_8939_), .Y(_12844_) );
NAND2X1 NAND2X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__10_), .Y(_12845_) );
NAND2X1 NAND2X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__10_), .Y(_12846_) );
NAND3X1 NAND3X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_12845_), .B(_12846_), .C(_12844_), .Y(_12847_) );
NOR2X1 NOR2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_12847_), .B(_12843_), .Y(_12848_) );
NAND2X1 NAND2X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_12839_), .B(_12848_), .Y(_12849_) );
NAND2X1 NAND2X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_208__10_), .Y(_12850_) );
NAND2X1 NAND2X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_8952_), .B(_40__10_), .Y(_12851_) );
AOI22X1 AOI22X1_408 ( .gnd(gnd), .vdd(vdd), .A(_238__10_), .B(_8893_), .C(_209__10_), .D(_8957_), .Y(_12852_) );
NAND3X1 NAND3X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_12850_), .B(_12851_), .C(_12852_), .Y(_12853_) );
AOI22X1 AOI22X1_409 ( .gnd(gnd), .vdd(vdd), .A(_42__10_), .B(_8963_), .C(_177__10_), .D(_8961_), .Y(_12854_) );
NAND2X1 NAND2X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_8901_), .B(_248__10_), .Y(_12855_) );
NAND2X1 NAND2X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_8968_), .B(_44__10_), .Y(_12856_) );
NAND3X1 NAND3X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_12855_), .B(_12856_), .C(_12854_), .Y(_12857_) );
NOR2X1 NOR2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_12853_), .B(_12857_), .Y(_12858_) );
NAND2X1 NAND2X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_8986_), .B(_255__10_), .Y(_12859_) );
NAND2X1 NAND2X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__10_), .Y(_12860_) );
AOI22X1 AOI22X1_410 ( .gnd(gnd), .vdd(vdd), .A(_37__10_), .B(_8978_), .C(_35__10_), .D(_8980_), .Y(_12861_) );
NAND3X1 NAND3X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_12859_), .B(_12860_), .C(_12861_), .Y(_12862_) );
NAND2X1 NAND2X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_8984_), .B(_254__10_), .Y(_12863_) );
NAND2X1 NAND2X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(_33__10_), .Y(_12864_) );
AOI22X1 AOI22X1_411 ( .gnd(gnd), .vdd(vdd), .A(_203__10_), .B(_9018_), .C(_156__10_), .D(_8973_), .Y(_12865_) );
NAND3X1 NAND3X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_12863_), .B(_12864_), .C(_12865_), .Y(_12866_) );
NOR2X1 NOR2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_12866_), .B(_12862_), .Y(_12867_) );
NAND2X1 NAND2X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_12858_), .B(_12867_), .Y(_12868_) );
NOR2X1 NOR2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_12849_), .B(_12868_), .Y(_12869_) );
NAND2X1 NAND2X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__10_), .Y(_12870_) );
NAND2X1 NAND2X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__10_), .Y(_12871_) );
AOI22X1 AOI22X1_412 ( .gnd(gnd), .vdd(vdd), .A(_13__10_), .B(_9007_), .C(_239__10_), .D(_9076_), .Y(_12872_) );
NAND3X1 NAND3X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_12870_), .B(_12871_), .C(_12872_), .Y(_12873_) );
AOI22X1 AOI22X1_413 ( .gnd(gnd), .vdd(vdd), .A(_206__10_), .B(_9013_), .C(_242__10_), .D(_9035_), .Y(_12874_) );
NAND2X1 NAND2X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__10_), .Y(_12875_) );
NAND2X1 NAND2X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__10_), .Y(_12876_) );
NAND3X1 NAND3X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_12875_), .B(_12876_), .C(_12874_), .Y(_12877_) );
NOR2X1 NOR2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_12873_), .B(_12877_), .Y(_12878_) );
AOI22X1 AOI22X1_414 ( .gnd(gnd), .vdd(vdd), .A(_222__10_), .B(_9024_), .C(_220__10_), .D(_9026_), .Y(_12879_) );
NAND2X1 NAND2X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__10_), .Y(_12880_) );
NAND2X1 NAND2X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__10_), .Y(_12881_) );
NAND3X1 NAND3X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_12880_), .B(_12881_), .C(_12879_), .Y(_12882_) );
AOI22X1 AOI22X1_415 ( .gnd(gnd), .vdd(vdd), .A(_18__10_), .B(_9037_), .C(_240__10_), .D(_9011_), .Y(_12883_) );
NAND2X1 NAND2X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__10_), .Y(_12884_) );
NAND2X1 NAND2X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__10_), .Y(_12885_) );
NAND3X1 NAND3X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_12884_), .B(_12885_), .C(_12883_), .Y(_12886_) );
NOR2X1 NOR2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_12882_), .B(_12886_), .Y(_12887_) );
NAND2X1 NAND2X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_12878_), .B(_12887_), .Y(_12888_) );
AOI22X1 AOI22X1_416 ( .gnd(gnd), .vdd(vdd), .A(_225__10_), .B(_9048_), .C(_167__10_), .D(_9050_), .Y(_12889_) );
NAND2X1 NAND2X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_9153_), .B(_243__10_), .Y(_12890_) );
NAND2X1 NAND2X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__10_), .Y(_12891_) );
NAND3X1 NAND3X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_12890_), .B(_12891_), .C(_12889_), .Y(_12892_) );
NAND2X1 NAND2X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__10_), .Y(_12893_) );
NAND2X1 NAND2X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__10_), .Y(_12894_) );
AOI22X1 AOI22X1_417 ( .gnd(gnd), .vdd(vdd), .A(_224__10_), .B(_9064_), .C(_27__10_), .D(_9066_), .Y(_12895_) );
NAND3X1 NAND3X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_12893_), .B(_12894_), .C(_12895_), .Y(_12896_) );
NOR2X1 NOR2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_12892_), .B(_12896_), .Y(_12897_) );
AOI22X1 AOI22X1_418 ( .gnd(gnd), .vdd(vdd), .A(_184__10_), .B(_9073_), .C(_183__10_), .D(_9071_), .Y(_12898_) );
NAND2X1 NAND2X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__10_), .Y(_12899_) );
NAND2X1 NAND2X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__10_), .Y(_12900_) );
NAND3X1 NAND3X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_12899_), .B(_12900_), .C(_12898_), .Y(_12901_) );
AOI22X1 AOI22X1_419 ( .gnd(gnd), .vdd(vdd), .A(_43__10_), .B(_9084_), .C(_244__10_), .D(_9160_), .Y(_12902_) );
NAND2X1 NAND2X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__10_), .Y(_12903_) );
NAND2X1 NAND2X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__10_), .Y(_12904_) );
NAND3X1 NAND3X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_12903_), .B(_12904_), .C(_12902_), .Y(_12905_) );
NOR2X1 NOR2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_12901_), .B(_12905_), .Y(_12906_) );
NAND2X1 NAND2X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_12897_), .B(_12906_), .Y(_12907_) );
NOR2X1 NOR2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_12888_), .B(_12907_), .Y(_12908_) );
NAND3X1 NAND3X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_6863_), .B(_9104_), .C(_6864_), .Y(_12909_) );
NAND3X1 NAND3X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_3971_), .B(_9099_), .C(_3972_), .Y(_12910_) );
NAND2X1 NAND2X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_12909_), .B(_12910_), .Y(_12911_) );
NAND2X1 NAND2X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__10_), .Y(_12912_) );
NAND3X1 NAND3X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .B(_9102_), .C(_5105_), .Y(_12913_) );
NAND2X1 NAND2X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_12913_), .B(_12912_), .Y(_12914_) );
NOR2X1 NOR2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_12911_), .B(_12914_), .Y(_12915_) );
NAND3X1 NAND3X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_8325_), .B(_9188_), .C(_8326_), .Y(_12916_) );
NAND3X1 NAND3X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_15932_), .B(_9109_), .C(_15933_), .Y(_12917_) );
NAND3X1 NAND3X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_16138_), .B(_9115_), .C(_16139_), .Y(_12918_) );
NAND3X1 NAND3X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_12917_), .B(_12918_), .C(_12916_), .Y(_12919_) );
AOI22X1 AOI22X1_420 ( .gnd(gnd), .vdd(vdd), .A(_234__10_), .B(_9182_), .C(_34__10_), .D(_9183_), .Y(_12920_) );
AOI22X1 AOI22X1_421 ( .gnd(gnd), .vdd(vdd), .A(_100__10_), .B(_9346_), .C(_45__10_), .D(_9185_), .Y(_12921_) );
NAND2X1 NAND2X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_12921_), .B(_12920_), .Y(_12922_) );
NAND3X1 NAND3X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_4750_), .B(_9127_), .C(_4749_), .Y(_12923_) );
NAND3X1 NAND3X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_9129_), .C(_4015_), .Y(_12924_) );
NAND2X1 NAND2X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_12923_), .B(_12924_), .Y(_12925_) );
NOR3X1 NOR3X1_371 ( .gnd(gnd), .vdd(vdd), .A(_12919_), .B(_12925_), .C(_12922_), .Y(_12926_) );
NAND3X1 NAND3X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .B(_9133_), .C(_3432_), .Y(_12927_) );
NAND3X1 NAND3X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_5057_), .B(_9135_), .C(_5058_), .Y(_12928_) );
NAND3X1 NAND3X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_6940_), .B(_9137_), .C(_6941_), .Y(_12929_) );
NAND3X1 NAND3X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_12928_), .B(_12929_), .C(_12927_), .Y(_12930_) );
AOI22X1 AOI22X1_422 ( .gnd(gnd), .vdd(vdd), .A(_17__10_), .B(_9140_), .C(_2__10_), .D(_9141_), .Y(_12931_) );
AOI22X1 AOI22X1_423 ( .gnd(gnd), .vdd(vdd), .A(_205__10_), .B(_9143_), .C(_200__10_), .D(_9145_), .Y(_12932_) );
NAND2X1 NAND2X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_12931_), .B(_12932_), .Y(_12933_) );
NOR2X1 NOR2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_12930_), .B(_12933_), .Y(_12934_) );
NAND3X1 NAND3X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_12915_), .B(_12926_), .C(_12934_), .Y(_12935_) );
AOI22X1 AOI22X1_424 ( .gnd(gnd), .vdd(vdd), .A(_21__10_), .B(_9150_), .C(_185__10_), .D(_9151_), .Y(_12936_) );
AOI22X1 AOI22X1_425 ( .gnd(gnd), .vdd(vdd), .A(_249__10_), .B(_9053_), .C(_253__10_), .D(_9154_), .Y(_12937_) );
NAND2X1 NAND2X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_12936_), .B(_12937_), .Y(_12938_) );
AOI22X1 AOI22X1_426 ( .gnd(gnd), .vdd(vdd), .A(_46__10_), .B(_9158_), .C(_231__10_), .D(_9157_), .Y(_12939_) );
AOI22X1 AOI22X1_427 ( .gnd(gnd), .vdd(vdd), .A(_47__10_), .B(_9161_), .C(_250__10_), .D(_9082_), .Y(_12940_) );
NAND2X1 NAND2X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_12940_), .B(_12939_), .Y(_12941_) );
NOR2X1 NOR2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_12938_), .B(_12941_), .Y(_12942_) );
AOI22X1 AOI22X1_428 ( .gnd(gnd), .vdd(vdd), .A(_247__10_), .B(_9165_), .C(_30__10_), .D(_9167_), .Y(_12943_) );
AOI22X1 AOI22X1_429 ( .gnd(gnd), .vdd(vdd), .A(_227__10_), .B(_9170_), .C(_218__10_), .D(_9169_), .Y(_12944_) );
NAND2X1 NAND2X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_12943_), .B(_12944_), .Y(_12945_) );
AOI22X1 AOI22X1_430 ( .gnd(gnd), .vdd(vdd), .A(_145__10_), .B(_9177_), .C(_213__10_), .D(_8989_), .Y(_12946_) );
AOI22X1 AOI22X1_431 ( .gnd(gnd), .vdd(vdd), .A(_29__10_), .B(_9176_), .C(_178__10_), .D(_9173_), .Y(_12947_) );
NAND2X1 NAND2X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_12946_), .B(_12947_), .Y(_12948_) );
NOR2X1 NOR2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_12945_), .B(_12948_), .Y(_12949_) );
NAND2X1 NAND2X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_12942_), .B(_12949_), .Y(_12950_) );
AOI22X1 AOI22X1_432 ( .gnd(gnd), .vdd(vdd), .A(_201__10_), .B(_9124_), .C(_212__10_), .D(_9345_), .Y(_12951_) );
NAND3X1 NAND3X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_8439_), .B(_9348_), .C(_8438_), .Y(_12952_) );
NAND3X1 NAND3X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_499_), .C(_500_), .Y(_12953_) );
AND2X2 AND2X2_1595 ( .gnd(gnd), .vdd(vdd), .A(_12953_), .B(_12952_), .Y(_12954_) );
NAND2X1 NAND2X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_12951_), .B(_12954_), .Y(_12955_) );
NAND3X1 NAND3X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_15145_), .B(_9208_), .C(_15146_), .Y(_12956_) );
OAI21X1 OAI21X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_15108_), .B(_9211_), .C(_12956_), .Y(_12957_) );
NAND3X1 NAND3X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_15489_), .B(_9222_), .C(_15490_), .Y(_12958_) );
NAND3X1 NAND3X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_15436_), .B(_9224_), .C(_15435_), .Y(_12959_) );
NAND2X1 NAND2X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_12958_), .B(_12959_), .Y(_12960_) );
NOR2X1 NOR2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_12960_), .B(_12957_), .Y(_12961_) );
NAND3X1 NAND3X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_15267_), .B(_9217_), .C(_15268_), .Y(_12962_) );
NAND3X1 NAND3X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_15215_), .B(_9219_), .C(_15214_), .Y(_12963_) );
NAND2X1 NAND2X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_12963_), .B(_12962_), .Y(_12964_) );
NAND3X1 NAND3X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_15665_), .B(_9192_), .C(_15666_), .Y(_12965_) );
NAND3X1 NAND3X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_15722_), .B(_9199_), .C(_15721_), .Y(_12966_) );
NAND2X1 NAND2X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_12966_), .B(_12965_), .Y(_12967_) );
NOR2X1 NOR2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_12967_), .B(_12964_), .Y(_12968_) );
NOR3X1 NOR3X1_372 ( .gnd(gnd), .vdd(vdd), .A(_16190_), .B(_10083_), .C(_16191_), .Y(_12969_) );
NAND3X1 NAND3X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_15317_), .B(_9205_), .C(_15318_), .Y(_12970_) );
OAI21X1 OAI21X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_15350_), .B(_10085_), .C(_12970_), .Y(_12971_) );
NAND3X1 NAND3X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_15547_), .B(_9233_), .C(_15548_), .Y(_12972_) );
NAND3X1 NAND3X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15615_), .C(_15614_), .Y(_12973_) );
NAND2X1 NAND2X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_12972_), .B(_12973_), .Y(_12974_) );
NOR3X1 NOR3X1_373 ( .gnd(gnd), .vdd(vdd), .A(_12971_), .B(_12974_), .C(_12969_), .Y(_12975_) );
NAND3X1 NAND3X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_12961_), .B(_12968_), .C(_12975_), .Y(_12976_) );
NAND3X1 NAND3X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_15875_), .B(_9120_), .C(_15876_), .Y(_12977_) );
NAND3X1 NAND3X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_15386_), .B(_9197_), .C(_15387_), .Y(_12978_) );
NOR2X1 NOR2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_9276_), .B(_14917_), .Y(_12979_) );
NOR3X1 NOR3X1_374 ( .gnd(gnd), .vdd(vdd), .A(_4190_), .B(_9254_), .C(_4192_), .Y(_12980_) );
NOR2X1 NOR2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_12340_), .B(_1771_), .Y(_12981_) );
NOR3X1 NOR3X1_375 ( .gnd(gnd), .vdd(vdd), .A(_12979_), .B(_12981_), .C(_12980_), .Y(_12982_) );
AND2X2 AND2X2_1596 ( .gnd(gnd), .vdd(vdd), .A(_186__10_), .B(_9298_), .Y(_12983_) );
NOR3X1 NOR3X1_376 ( .gnd(gnd), .vdd(vdd), .A(_7472_), .B(_10471_), .C(_7473_), .Y(_12984_) );
NAND3X1 NAND3X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_8241_), .B(_9250_), .C(_8240_), .Y(_12985_) );
OAI21X1 OAI21X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_8716_), .C(_12985_), .Y(_12986_) );
NOR3X1 NOR3X1_377 ( .gnd(gnd), .vdd(vdd), .A(_12984_), .B(_12983_), .C(_12986_), .Y(_12987_) );
NAND3X1 NAND3X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_7099_), .B(_9244_), .C(_7098_), .Y(_12988_) );
OAI21X1 OAI21X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .B(_9306_), .C(_12988_), .Y(_12989_) );
NAND3X1 NAND3X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_15817_), .B(_9292_), .C(_15816_), .Y(_12990_) );
OAI21X1 OAI21X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_7640_), .B(_9301_), .C(_12990_), .Y(_12991_) );
NOR2X1 NOR2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_12991_), .B(_12989_), .Y(_12992_) );
NAND3X1 NAND3X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_12982_), .B(_12992_), .C(_12987_), .Y(_12993_) );
NOR3X1 NOR3X1_378 ( .gnd(gnd), .vdd(vdd), .A(_6435_), .B(_9763_), .C(_6436_), .Y(_12994_) );
NAND3X1 NAND3X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_7054_), .B(_9266_), .C(_7053_), .Y(_12995_) );
OAI21X1 OAI21X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_7725_), .B(_9249_), .C(_12995_), .Y(_12996_) );
NAND3X1 NAND3X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_9321_), .B(_7681_), .C(_7682_), .Y(_12997_) );
OAI21X1 OAI21X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .B(_9273_), .C(_12997_), .Y(_12998_) );
NOR3X1 NOR3X1_379 ( .gnd(gnd), .vdd(vdd), .A(_12998_), .B(_12996_), .C(_12994_), .Y(_12999_) );
NAND2X1 NAND2X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__10_), .Y(_13000_) );
OAI21X1 OAI21X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_8173_), .B(_9304_), .C(_13000_), .Y(_13001_) );
NAND3X1 NAND3X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_8204_), .B(_9286_), .C(_8205_), .Y(_13002_) );
NAND3X1 NAND3X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_9268_), .C(_1176_), .Y(_13003_) );
NAND2X1 NAND2X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_13002_), .B(_13003_), .Y(_13004_) );
NOR2X1 NOR2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_13001_), .B(_13004_), .Y(_13005_) );
NAND3X1 NAND3X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .B(_9277_), .C(_2919_), .Y(_13006_) );
OAI21X1 OAI21X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_3609_), .B(_9295_), .C(_13006_), .Y(_13007_) );
NAND2X1 NAND2X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__10_), .Y(_13008_) );
OAI21X1 OAI21X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_9263_), .C(_13008_), .Y(_13009_) );
NOR2X1 NOR2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_13009_), .B(_13007_), .Y(_13010_) );
NAND3X1 NAND3X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_12999_), .B(_13005_), .C(_13010_), .Y(_13011_) );
NOR2X1 NOR2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_9325_), .B(_5374_), .Y(_13012_) );
NOR3X1 NOR3X1_380 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(_9312_), .C(_4784_), .Y(_13013_) );
NOR2X1 NOR2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .B(_4228_), .Y(_13014_) );
NOR3X1 NOR3X1_381 ( .gnd(gnd), .vdd(vdd), .A(_13012_), .B(_13014_), .C(_13013_), .Y(_13015_) );
AOI22X1 AOI22X1_433 ( .gnd(gnd), .vdd(vdd), .A(_83__10_), .B(_9315_), .C(_235__10_), .D(_9324_), .Y(_13016_) );
AOI22X1 AOI22X1_434 ( .gnd(gnd), .vdd(vdd), .A(_233__10_), .B(_9310_), .C(_251__10_), .D(_9320_), .Y(_13017_) );
NAND3X1 NAND3X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_13015_), .B(_13016_), .C(_13017_), .Y(_13018_) );
NOR3X1 NOR3X1_382 ( .gnd(gnd), .vdd(vdd), .A(_13011_), .B(_13018_), .C(_12993_), .Y(_13019_) );
NAND2X1 NAND2X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_12978_), .B(_13019_), .Y(_13020_) );
AOI21X1 AOI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_157__10_), .B(_9232_), .C(_13020_), .Y(_13021_) );
AOI22X1 AOI22X1_435 ( .gnd(gnd), .vdd(vdd), .A(_155__10_), .B(_9333_), .C(_172__10_), .D(_9332_), .Y(_13022_) );
NAND3X1 NAND3X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_12977_), .B(_13022_), .C(_13021_), .Y(_13023_) );
NOR3X1 NOR3X1_383 ( .gnd(gnd), .vdd(vdd), .A(_12976_), .B(_13023_), .C(_12955_), .Y(_13024_) );
AOI22X1 AOI22X1_436 ( .gnd(gnd), .vdd(vdd), .A(_256__10_), .B(_9113_), .C(_142__10_), .D(_9118_), .Y(_13025_) );
NAND2X1 NAND2X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__10_), .Y(_13026_) );
NAND2X1 NAND2X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__10_), .Y(_13027_) );
NAND3X1 NAND3X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_13026_), .B(_13027_), .C(_13025_), .Y(_13028_) );
NAND2X1 NAND2X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__10_), .Y(_13029_) );
NAND3X1 NAND3X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_9339_), .C(_458_), .Y(_13030_) );
AOI22X1 AOI22X1_437 ( .gnd(gnd), .vdd(vdd), .A(_111__10_), .B(_9342_), .C(_12__10_), .D(_9341_), .Y(_13031_) );
NAND3X1 NAND3X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_13031_), .B(_13029_), .C(_13030_), .Y(_13032_) );
NOR2X1 NOR2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_13028_), .B(_13032_), .Y(_13033_) );
AOI22X1 AOI22X1_438 ( .gnd(gnd), .vdd(vdd), .A(_232__10_), .B(_9354_), .C(_219__10_), .D(_9353_), .Y(_13034_) );
AOI22X1 AOI22X1_439 ( .gnd(gnd), .vdd(vdd), .A(_246__10_), .B(_9356_), .C(_226__10_), .D(_9357_), .Y(_13035_) );
NAND2X1 NAND2X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_13034_), .B(_13035_), .Y(_13036_) );
NAND3X1 NAND3X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16092_), .C(_16093_), .Y(_13037_) );
NAND3X1 NAND3X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16037_), .C(_16038_), .Y(_13038_) );
NAND2X1 NAND2X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_13037_), .B(_13038_), .Y(_13039_) );
NAND3X1 NAND3X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8571_), .C(_8570_), .Y(_13040_) );
OAI21X1 OAI21X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_9361_), .C(_13040_), .Y(_13041_) );
NOR2X1 NOR2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_13039_), .B(_13041_), .Y(_13042_) );
NAND2X1 NAND2X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_15983_), .B(_15984_), .Y(_13043_) );
NAND3X1 NAND3X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8624_), .C(_8625_), .Y(_13044_) );
OAI21X1 OAI21X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_13043_), .B(_9215_), .C(_13044_), .Y(_13045_) );
NAND3X1 NAND3X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_8679_), .B(_9371_), .C(_8678_), .Y(_13046_) );
NAND3X1 NAND3X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_321_), .C(_322_), .Y(_13047_) );
NAND2X1 NAND2X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_13047_), .B(_13046_), .Y(_13048_) );
NOR2X1 NOR2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_13045_), .B(_13048_), .Y(_13049_) );
AOI22X1 AOI22X1_440 ( .gnd(gnd), .vdd(vdd), .A(_22__10_), .B(_9382_), .C(_3__10_), .D(_9383_), .Y(_13050_) );
NAND3X1 NAND3X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_13042_), .B(_13049_), .C(_13050_), .Y(_13051_) );
NOR2X1 NOR2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_13036_), .B(_13051_), .Y(_13052_) );
NAND3X1 NAND3X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_13024_), .B(_13033_), .C(_13052_), .Y(_13053_) );
NOR3X1 NOR3X1_384 ( .gnd(gnd), .vdd(vdd), .A(_12935_), .B(_12950_), .C(_13053_), .Y(_13054_) );
NAND3X1 NAND3X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_12869_), .B(_12908_), .C(_13054_), .Y(_13055_) );
NAND3X1 NAND3X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1590_), .C(_1591_), .Y(_13056_) );
NAND3X1 NAND3X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_1251_), .B(_8862_), .C(_1252_), .Y(_13057_) );
NAND2X1 NAND2X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_13056_), .B(_13057_), .Y(_13058_) );
NOR3X1 NOR3X1_385 ( .gnd(gnd), .vdd(vdd), .A(_12831_), .B(_13058_), .C(_13055_), .Y(_13059_) );
NAND3X1 NAND3X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_12813_), .B(_12820_), .C(_13059_), .Y(_13060_) );
NAND2X1 NAND2X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__10_), .Y(_13061_) );
NAND3X1 NAND3X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_9406_), .C(_1467_), .Y(_13062_) );
NAND3X1 NAND3X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_9453_), .C(_1421_), .Y(_13063_) );
AND2X2 AND2X2_1597 ( .gnd(gnd), .vdd(vdd), .A(_13062_), .B(_13063_), .Y(_13064_) );
NAND2X1 NAND2X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_108__10_), .Y(_13065_) );
NAND2X1 NAND2X1_2346 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_116__10_), .Y(_13066_) );
NAND3X1 NAND3X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_13065_), .B(_13066_), .C(_13064_), .Y(_13067_) );
AOI22X1 AOI22X1_441 ( .gnd(gnd), .vdd(vdd), .A(_125__10_), .B(_9411_), .C(_124__10_), .D(_9410_), .Y(_13068_) );
AOI22X1 AOI22X1_442 ( .gnd(gnd), .vdd(vdd), .A(_120__10_), .B(_9415_), .C(_121__10_), .D(_9413_), .Y(_13069_) );
AND2X2 AND2X2_1598 ( .gnd(gnd), .vdd(vdd), .A(_13069_), .B(_13068_), .Y(_13070_) );
AOI22X1 AOI22X1_443 ( .gnd(gnd), .vdd(vdd), .A(_132__10_), .B(_9420_), .C(_131__10_), .D(_9418_), .Y(_13071_) );
NAND2X1 NAND2X1_2347 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__10_), .Y(_13072_) );
NAND2X1 NAND2X1_2348 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__10_), .Y(_13073_) );
NAND3X1 NAND3X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_13072_), .B(_13073_), .C(_13071_), .Y(_13074_) );
NAND3X1 NAND3X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_9431_), .C(_553_), .Y(_13075_) );
NAND2X1 NAND2X1_2349 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__10_), .Y(_13076_) );
NAND2X1 NAND2X1_2350 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__10_), .Y(_13077_) );
NAND3X1 NAND3X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_13077_), .B(_13075_), .C(_13076_), .Y(_13078_) );
AOI21X1 AOI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_136__10_), .B(_9429_), .C(_13078_), .Y(_13079_) );
NAND2X1 NAND2X1_2351 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__10_), .Y(_13080_) );
NAND2X1 NAND2X1_2352 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__10_), .Y(_13081_) );
NAND3X1 NAND3X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_13080_), .B(_13081_), .C(_13079_), .Y(_13082_) );
NAND3X1 NAND3X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_9444_), .C(_1060_), .Y(_13083_) );
NAND2X1 NAND2X1_2353 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__10_), .Y(_13084_) );
AOI22X1 AOI22X1_444 ( .gnd(gnd), .vdd(vdd), .A(_130__10_), .B(_9449_), .C(_127__10_), .D(_9448_), .Y(_13085_) );
NAND3X1 NAND3X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_13083_), .B(_13085_), .C(_13084_), .Y(_13086_) );
NOR3X1 NOR3X1_386 ( .gnd(gnd), .vdd(vdd), .A(_13074_), .B(_13082_), .C(_13086_), .Y(_13087_) );
AOI22X1 AOI22X1_445 ( .gnd(gnd), .vdd(vdd), .A(_115__10_), .B(_9399_), .C(_114__10_), .D(_9454_), .Y(_13088_) );
NAND3X1 NAND3X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_13088_), .B(_13070_), .C(_13087_), .Y(_13089_) );
NOR2X1 NOR2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_13067_), .B(_13089_), .Y(_13090_) );
AOI22X1 AOI22X1_446 ( .gnd(gnd), .vdd(vdd), .A(_102__10_), .B(_9459_), .C(_103__10_), .D(_9457_), .Y(_13091_) );
NAND3X1 NAND3X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_13061_), .B(_13091_), .C(_13090_), .Y(_13092_) );
NOR3X1 NOR3X1_387 ( .gnd(gnd), .vdd(vdd), .A(_12812_), .B(_13092_), .C(_13060_), .Y(_13093_) );
NAND3X1 NAND3X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_12802_), .B(_12809_), .C(_13093_), .Y(_13094_) );
NOR3X1 NOR3X1_388 ( .gnd(gnd), .vdd(vdd), .A(_12791_), .B(_12794_), .C(_13094_), .Y(_13095_) );
NAND3X1 NAND3X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_12782_), .B(_12787_), .C(_13095_), .Y(_13096_) );
NAND3X1 NAND3X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_3070_), .B(_9473_), .C(_3071_), .Y(_13097_) );
NAND2X1 NAND2X1_2354 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__10_), .Y(_13098_) );
NAND2X1 NAND2X1_2355 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__10_), .Y(_13099_) );
NAND2X1 NAND2X1_2356 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__10_), .Y(_13100_) );
NAND3X1 NAND3X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_2442_), .B(_9468_), .C(_2443_), .Y(_13101_) );
NAND3X1 NAND3X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_13101_), .B(_13099_), .C(_13100_), .Y(_13102_) );
AOI21X1 AOI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_68__10_), .B(_9477_), .C(_13102_), .Y(_13103_) );
NAND3X1 NAND3X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_13103_), .B(_13097_), .C(_13098_), .Y(_13104_) );
NOR3X1 NOR3X1_389 ( .gnd(gnd), .vdd(vdd), .A(_12781_), .B(_13104_), .C(_13096_), .Y(_13105_) );
AOI21X1 AOI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_12776_), .B(_13105_), .C(rst), .Y(_0__10_) );
NAND2X1 NAND2X1_2357 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__11_), .Y(_13106_) );
NAND2X1 NAND2X1_2358 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__11_), .Y(_13107_) );
NAND2X1 NAND2X1_2359 ( .gnd(gnd), .vdd(vdd), .A(_13106_), .B(_13107_), .Y(_13108_) );
NAND2X1 NAND2X1_2360 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_55__11_), .Y(_13109_) );
NAND2X1 NAND2X1_2361 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__11_), .Y(_13110_) );
NAND2X1 NAND2X1_2362 ( .gnd(gnd), .vdd(vdd), .A(_13110_), .B(_13109_), .Y(_13111_) );
NOR2X1 NOR2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_13111_), .B(_13108_), .Y(_13112_) );
NAND3X1 NAND3X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_8750_), .C(_3165_), .Y(_13113_) );
NAND3X1 NAND3X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_3114_), .B(_8757_), .C(_3113_), .Y(_13114_) );
NAND2X1 NAND2X1_2363 ( .gnd(gnd), .vdd(vdd), .A(_13113_), .B(_13114_), .Y(_13115_) );
NAND3X1 NAND3X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_3290_), .B(_8762_), .C(_3289_), .Y(_13116_) );
NAND3X1 NAND3X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_8774_), .C(_3018_), .Y(_13117_) );
NAND2X1 NAND2X1_2364 ( .gnd(gnd), .vdd(vdd), .A(_13116_), .B(_13117_), .Y(_13118_) );
OR2X2 OR2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_13115_), .B(_13118_), .Y(_13119_) );
NAND2X1 NAND2X1_2365 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__11_), .Y(_13120_) );
NAND3X1 NAND3X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_2827_), .B(_8786_), .C(_2828_), .Y(_13121_) );
OAI21X1 OAI21X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_2718_), .B(_8792_), .C(_13121_), .Y(_13122_) );
NAND3X1 NAND3X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_2656_), .B(_8794_), .C(_2657_), .Y(_13123_) );
OAI21X1 OAI21X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_2774_), .B(_8799_), .C(_13123_), .Y(_13124_) );
NOR2X1 NOR2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_13124_), .B(_13122_), .Y(_13125_) );
AOI22X1 AOI22X1_447 ( .gnd(gnd), .vdd(vdd), .A(_76__11_), .B(_9482_), .C(_77__11_), .D(_9478_), .Y(_13126_) );
NAND2X1 NAND2X1_2366 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__11_), .Y(_13127_) );
NAND2X1 NAND2X1_2367 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_82__11_), .Y(_13128_) );
NAND3X1 NAND3X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_13127_), .B(_13128_), .C(_13126_), .Y(_13129_) );
NAND2X1 NAND2X1_2368 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__11_), .Y(_13130_) );
NAND3X1 NAND3X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_2591_), .B(_8803_), .C(_2590_), .Y(_13131_) );
NAND2X1 NAND2X1_2369 ( .gnd(gnd), .vdd(vdd), .A(_13131_), .B(_13130_), .Y(_13132_) );
INVX1 INVX1_3880 ( .gnd(gnd), .vdd(vdd), .A(_84__11_), .Y(_13133_) );
NOR2X1 NOR2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_13133_), .Y(_13134_) );
NOR2X1 NOR2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2304_), .Y(_13135_) );
NAND2X1 NAND2X1_2370 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__11_), .Y(_13136_) );
NAND3X1 NAND3X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_1979_), .B(_8840_), .C(_1980_), .Y(_13137_) );
NAND3X1 NAND3X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1925_), .C(_1926_), .Y(_13138_) );
NAND3X1 NAND3X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_13138_), .B(_13137_), .C(_13136_), .Y(_13139_) );
NOR3X1 NOR3X1_390 ( .gnd(gnd), .vdd(vdd), .A(_13134_), .B(_13139_), .C(_13135_), .Y(_13140_) );
NAND3X1 NAND3X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_2263_), .B(_8829_), .C(_2264_), .Y(_13141_) );
NAND3X1 NAND3X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(_8831_), .C(_2158_), .Y(_13142_) );
NAND2X1 NAND2X1_2371 ( .gnd(gnd), .vdd(vdd), .A(_13141_), .B(_13142_), .Y(_13143_) );
NAND3X1 NAND3X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_8834_), .C(_2099_), .Y(_13144_) );
NAND3X1 NAND3X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_2209_), .B(_8836_), .C(_2210_), .Y(_13145_) );
NAND2X1 NAND2X1_2372 ( .gnd(gnd), .vdd(vdd), .A(_13144_), .B(_13145_), .Y(_13146_) );
NOR2X1 NOR2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_13146_), .B(_13143_), .Y(_13147_) );
AOI22X1 AOI22X1_448 ( .gnd(gnd), .vdd(vdd), .A(_94__11_), .B(_8841_), .C(_91__11_), .D(_8823_), .Y(_13148_) );
NAND2X1 NAND2X1_2373 ( .gnd(gnd), .vdd(vdd), .A(_8843_), .B(_92__11_), .Y(_13149_) );
NAND2X1 NAND2X1_2374 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_98__11_), .Y(_13150_) );
NAND3X1 NAND3X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_13149_), .B(_13150_), .C(_13148_), .Y(_13151_) );
NAND2X1 NAND2X1_2375 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__11_), .Y(_13152_) );
NAND3X1 NAND3X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1552_), .C(_1553_), .Y(_13153_) );
NAND3X1 NAND3X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1637_), .C(_1638_), .Y(_13154_) );
NAND2X1 NAND2X1_2376 ( .gnd(gnd), .vdd(vdd), .A(_13153_), .B(_13154_), .Y(_13155_) );
NAND3X1 NAND3X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1675_), .C(_1676_), .Y(_13156_) );
NAND3X1 NAND3X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_8857_), .C(_1384_), .Y(_13157_) );
NAND2X1 NAND2X1_2377 ( .gnd(gnd), .vdd(vdd), .A(_13157_), .B(_13156_), .Y(_13158_) );
OR2X2 OR2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_13155_), .B(_13158_), .Y(_13159_) );
NOR3X1 NOR3X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1216_), .B(_8867_), .C(_1217_), .Y(_13160_) );
AOI22X1 AOI22X1_449 ( .gnd(gnd), .vdd(vdd), .A(_191__11_), .B(_8873_), .C(_192__11_), .D(_8872_), .Y(_13161_) );
AOI22X1 AOI22X1_450 ( .gnd(gnd), .vdd(vdd), .A(_195__11_), .B(_8875_), .C(_193__11_), .D(_8876_), .Y(_13162_) );
NAND2X1 NAND2X1_2378 ( .gnd(gnd), .vdd(vdd), .A(_13161_), .B(_13162_), .Y(_13163_) );
AOI22X1 AOI22X1_451 ( .gnd(gnd), .vdd(vdd), .A(_188__11_), .B(_8879_), .C(_126__11_), .D(_8881_), .Y(_13164_) );
AOI22X1 AOI22X1_452 ( .gnd(gnd), .vdd(vdd), .A(_196__11_), .B(_8883_), .C(_194__11_), .D(_8884_), .Y(_13165_) );
NAND2X1 NAND2X1_2379 ( .gnd(gnd), .vdd(vdd), .A(_13164_), .B(_13165_), .Y(_13166_) );
NOR3X1 NOR3X1_392 ( .gnd(gnd), .vdd(vdd), .A(_13166_), .B(_13160_), .C(_13163_), .Y(_13167_) );
NAND3X1 NAND3X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_5837_), .B(_8893_), .C(_5836_), .Y(_13168_) );
NAND3X1 NAND3X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_4596_), .B(_8898_), .C(_4595_), .Y(_13169_) );
NAND2X1 NAND2X1_2380 ( .gnd(gnd), .vdd(vdd), .A(_13168_), .B(_13169_), .Y(_13170_) );
NAND3X1 NAND3X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_5534_), .B(_8901_), .C(_5533_), .Y(_13171_) );
NAND3X1 NAND3X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_7871_), .B(_8904_), .C(_7870_), .Y(_13172_) );
NAND2X1 NAND2X1_2381 ( .gnd(gnd), .vdd(vdd), .A(_13171_), .B(_13172_), .Y(_13173_) );
NOR2X1 NOR2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_13170_), .B(_13173_), .Y(_13174_) );
NAND3X1 NAND3X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_4096_), .B(_8909_), .C(_4095_), .Y(_13175_) );
NAND3X1 NAND3X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3898_), .C(_3897_), .Y(_13176_) );
NAND2X1 NAND2X1_2382 ( .gnd(gnd), .vdd(vdd), .A(_13175_), .B(_13176_), .Y(_13177_) );
NAND3X1 NAND3X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_4637_), .B(_8914_), .C(_4636_), .Y(_13178_) );
NAND3X1 NAND3X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_6658_), .B(_8918_), .C(_6657_), .Y(_13179_) );
NAND2X1 NAND2X1_2383 ( .gnd(gnd), .vdd(vdd), .A(_13178_), .B(_13179_), .Y(_13180_) );
NOR2X1 NOR2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_13177_), .B(_13180_), .Y(_13181_) );
NAND2X1 NAND2X1_2384 ( .gnd(gnd), .vdd(vdd), .A(_13174_), .B(_13181_), .Y(_13182_) );
NAND3X1 NAND3X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_4977_), .B(_8926_), .C(_4976_), .Y(_13183_) );
NAND3X1 NAND3X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_8045_), .B(_8933_), .C(_8044_), .Y(_13184_) );
NAND2X1 NAND2X1_2385 ( .gnd(gnd), .vdd(vdd), .A(_13183_), .B(_13184_), .Y(_13185_) );
NAND3X1 NAND3X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_4499_), .B(_8931_), .C(_4498_), .Y(_13186_) );
NAND3X1 NAND3X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_8008_), .B(_9177_), .C(_8007_), .Y(_13187_) );
NAND2X1 NAND2X1_2386 ( .gnd(gnd), .vdd(vdd), .A(_13186_), .B(_13187_), .Y(_13188_) );
NOR2X1 NOR2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_13185_), .B(_13188_), .Y(_13189_) );
NAND3X1 NAND3X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_5191_), .B(_8937_), .C(_5190_), .Y(_13190_) );
NAND3X1 NAND3X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_7833_), .B(_8939_), .C(_7832_), .Y(_13191_) );
NAND2X1 NAND2X1_2387 ( .gnd(gnd), .vdd(vdd), .A(_13190_), .B(_13191_), .Y(_13192_) );
NAND3X1 NAND3X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_5153_), .B(_8942_), .C(_5152_), .Y(_13193_) );
NAND3X1 NAND3X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_5015_), .B(_8944_), .C(_5014_), .Y(_13194_) );
NAND2X1 NAND2X1_2388 ( .gnd(gnd), .vdd(vdd), .A(_13193_), .B(_13194_), .Y(_13195_) );
NOR2X1 NOR2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_13195_), .B(_13192_), .Y(_13196_) );
NAND2X1 NAND2X1_2389 ( .gnd(gnd), .vdd(vdd), .A(_13189_), .B(_13196_), .Y(_13197_) );
NOR2X1 NOR2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_13182_), .B(_13197_), .Y(_13198_) );
NAND3X1 NAND3X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_6726_), .B(_8950_), .C(_6725_), .Y(_13199_) );
NAND3X1 NAND3X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_3936_), .B(_8952_), .C(_3935_), .Y(_13200_) );
NAND2X1 NAND2X1_2390 ( .gnd(gnd), .vdd(vdd), .A(_13199_), .B(_13200_), .Y(_13201_) );
NAND3X1 NAND3X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_5906_), .B(_8955_), .C(_5905_), .Y(_13202_) );
NAND3X1 NAND3X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_6694_), .B(_8957_), .C(_6693_), .Y(_13203_) );
NAND2X1 NAND2X1_2391 ( .gnd(gnd), .vdd(vdd), .A(_13202_), .B(_13203_), .Y(_13204_) );
NOR2X1 NOR2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_13204_), .B(_13201_), .Y(_13205_) );
NAND3X1 NAND3X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_7796_), .B(_8961_), .C(_7795_), .Y(_13206_) );
NAND3X1 NAND3X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_3857_), .B(_8963_), .C(_3856_), .Y(_13207_) );
NAND2X1 NAND2X1_2392 ( .gnd(gnd), .vdd(vdd), .A(_13206_), .B(_13207_), .Y(_13208_) );
NAND3X1 NAND3X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_5873_), .B(_8966_), .C(_5872_), .Y(_13209_) );
NAND3X1 NAND3X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_3777_), .B(_8968_), .C(_3776_), .Y(_13210_) );
NAND2X1 NAND2X1_2393 ( .gnd(gnd), .vdd(vdd), .A(_13209_), .B(_13210_), .Y(_13211_) );
NOR2X1 NOR2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_13208_), .B(_13211_), .Y(_13212_) );
NAND2X1 NAND2X1_2394 ( .gnd(gnd), .vdd(vdd), .A(_13205_), .B(_13212_), .Y(_13213_) );
NAND3X1 NAND3X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_5285_), .B(_8986_), .C(_5284_), .Y(_13214_) );
NAND3X1 NAND3X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .B(_8975_), .C(_3483_), .Y(_13215_) );
NAND2X1 NAND2X1_2395 ( .gnd(gnd), .vdd(vdd), .A(_13214_), .B(_13215_), .Y(_13216_) );
NAND3X1 NAND3X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_4059_), .B(_8978_), .C(_4058_), .Y(_13217_) );
NAND3X1 NAND3X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_4133_), .B(_8980_), .C(_4132_), .Y(_13218_) );
NAND2X1 NAND2X1_2396 ( .gnd(gnd), .vdd(vdd), .A(_13218_), .B(_13217_), .Y(_13219_) );
NOR2X1 NOR2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_13216_), .B(_13219_), .Y(_13220_) );
NAND3X1 NAND3X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_5320_), .B(_8984_), .C(_5319_), .Y(_13221_) );
NAND3X1 NAND3X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_4166_), .B(_8991_), .C(_4165_), .Y(_13222_) );
NAND2X1 NAND2X1_2397 ( .gnd(gnd), .vdd(vdd), .A(_13221_), .B(_13222_), .Y(_13223_) );
NAND3X1 NAND3X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_7977_), .B(_8973_), .C(_7976_), .Y(_13224_) );
NAND3X1 NAND3X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_6900_), .B(_9018_), .C(_6899_), .Y(_13225_) );
NAND2X1 NAND2X1_2398 ( .gnd(gnd), .vdd(vdd), .A(_13224_), .B(_13225_), .Y(_13226_) );
NOR2X1 NOR2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_13223_), .B(_13226_), .Y(_13227_) );
NAND2X1 NAND2X1_2399 ( .gnd(gnd), .vdd(vdd), .A(_13220_), .B(_13227_), .Y(_13228_) );
NOR2X1 NOR2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_13213_), .B(_13228_), .Y(_13229_) );
NAND2X1 NAND2X1_2400 ( .gnd(gnd), .vdd(vdd), .A(_13198_), .B(_13229_), .Y(_13230_) );
NAND3X1 NAND3X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_4908_), .B(_8998_), .C(_4907_), .Y(_13231_) );
NAND3X1 NAND3X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_6515_), .B(_9002_), .C(_6514_), .Y(_13232_) );
NAND2X1 NAND2X1_2401 ( .gnd(gnd), .vdd(vdd), .A(_13231_), .B(_13232_), .Y(_13233_) );
NAND3X1 NAND3X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_5721_), .B(_9005_), .C(_5720_), .Y(_13234_) );
NAND3X1 NAND3X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(_9007_), .C(_4868_), .Y(_13235_) );
NAND2X1 NAND2X1_2402 ( .gnd(gnd), .vdd(vdd), .A(_13234_), .B(_13235_), .Y(_13236_) );
NOR2X1 NOR2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_13233_), .B(_13236_), .Y(_13237_) );
NAND3X1 NAND3X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_5759_), .B(_9011_), .C(_5758_), .Y(_13238_) );
NAND3X1 NAND3X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_6801_), .B(_9013_), .C(_6800_), .Y(_13239_) );
NAND2X1 NAND2X1_2403 ( .gnd(gnd), .vdd(vdd), .A(_13238_), .B(_13239_), .Y(_13240_) );
NAND3X1 NAND3X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_6762_), .B(_9016_), .C(_6761_), .Y(_13241_) );
NAND3X1 NAND3X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_6548_), .B(_9174_), .C(_6547_), .Y(_13242_) );
NAND2X1 NAND2X1_2404 ( .gnd(gnd), .vdd(vdd), .A(_13241_), .B(_13242_), .Y(_13243_) );
NOR2X1 NOR2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_13243_), .B(_13240_), .Y(_13244_) );
NAND2X1 NAND2X1_2405 ( .gnd(gnd), .vdd(vdd), .A(_13237_), .B(_13244_), .Y(_13245_) );
NAND3X1 NAND3X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_6285_), .B(_9024_), .C(_6284_), .Y(_13246_) );
NAND3X1 NAND3X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_6357_), .B(_9026_), .C(_6356_), .Y(_13247_) );
NAND2X1 NAND2X1_2406 ( .gnd(gnd), .vdd(vdd), .A(_13246_), .B(_13247_), .Y(_13248_) );
NAND3X1 NAND3X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_6062_), .B(_9029_), .C(_6061_), .Y(_13249_) );
NAND3X1 NAND3X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_6120_), .B(_9031_), .C(_6119_), .Y(_13250_) );
NAND2X1 NAND2X1_2407 ( .gnd(gnd), .vdd(vdd), .A(_13249_), .B(_13250_), .Y(_13251_) );
NOR2X1 NOR2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_13248_), .B(_13251_), .Y(_13252_) );
NAND3X1 NAND3X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_5680_), .B(_9035_), .C(_5679_), .Y(_13253_) );
NAND3X1 NAND3X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_9037_), .C(_4675_), .Y(_13254_) );
NAND2X1 NAND2X1_2408 ( .gnd(gnd), .vdd(vdd), .A(_13254_), .B(_13253_), .Y(_13255_) );
NAND3X1 NAND3X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_6321_), .B(_9040_), .C(_6320_), .Y(_13256_) );
NAND3X1 NAND3X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_4338_), .B(_9042_), .C(_4337_), .Y(_13257_) );
NAND2X1 NAND2X1_2409 ( .gnd(gnd), .vdd(vdd), .A(_13256_), .B(_13257_), .Y(_13258_) );
NOR2X1 NOR2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_13258_), .B(_13255_), .Y(_13259_) );
NAND2X1 NAND2X1_2410 ( .gnd(gnd), .vdd(vdd), .A(_13252_), .B(_13259_), .Y(_13260_) );
NOR2X1 NOR2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_13245_), .B(_13260_), .Y(_13261_) );
NAND3X1 NAND3X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_6209_), .B(_9048_), .C(_6208_), .Y(_13262_) );
NAND3X1 NAND3X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_7944_), .B(_9050_), .C(_7943_), .Y(_13263_) );
NAND2X1 NAND2X1_2411 ( .gnd(gnd), .vdd(vdd), .A(_13262_), .B(_13263_), .Y(_13264_) );
NAND3X1 NAND3X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_5492_), .B(_9053_), .C(_5491_), .Y(_13265_) );
NAND3X1 NAND3X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_7907_), .B(_9055_), .C(_7906_), .Y(_13266_) );
NAND2X1 NAND2X1_2412 ( .gnd(gnd), .vdd(vdd), .A(_13265_), .B(_13266_), .Y(_13267_) );
NOR2X1 NOR2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_13264_), .B(_13267_), .Y(_13268_) );
NAND3X1 NAND3X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_4459_), .B(_9059_), .C(_4458_), .Y(_13269_) );
NAND3X1 NAND3X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_4419_), .B(_9061_), .C(_4418_), .Y(_13270_) );
NAND2X1 NAND2X1_2413 ( .gnd(gnd), .vdd(vdd), .A(_13269_), .B(_13270_), .Y(_13271_) );
NAND3X1 NAND3X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_6247_), .B(_9064_), .C(_6246_), .Y(_13272_) );
NAND3X1 NAND3X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_4379_), .B(_9066_), .C(_4378_), .Y(_13273_) );
NAND2X1 NAND2X1_2414 ( .gnd(gnd), .vdd(vdd), .A(_13272_), .B(_13273_), .Y(_13274_) );
NOR2X1 NOR2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_13274_), .B(_13271_), .Y(_13275_) );
NAND2X1 NAND2X1_2415 ( .gnd(gnd), .vdd(vdd), .A(_13268_), .B(_13275_), .Y(_13276_) );
NAND3X1 NAND3X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_7603_), .B(_9071_), .C(_7602_), .Y(_13277_) );
NAND3X1 NAND3X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_7567_), .B(_9073_), .C(_7566_), .Y(_13278_) );
NAND2X1 NAND2X1_2416 ( .gnd(gnd), .vdd(vdd), .A(_13277_), .B(_13278_), .Y(_13279_) );
NAND3X1 NAND3X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_5797_), .B(_9076_), .C(_5796_), .Y(_13280_) );
NAND3X1 NAND3X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_9078_), .C(_3522_), .Y(_13281_) );
NAND2X1 NAND2X1_2417 ( .gnd(gnd), .vdd(vdd), .A(_13280_), .B(_13281_), .Y(_13282_) );
NOR2X1 NOR2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_13279_), .B(_13282_), .Y(_13283_) );
NAND3X1 NAND3X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_5451_), .B(_9082_), .C(_5450_), .Y(_13284_) );
NAND3X1 NAND3X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_3819_), .B(_9084_), .C(_3818_), .Y(_13285_) );
NAND2X1 NAND2X1_2418 ( .gnd(gnd), .vdd(vdd), .A(_13285_), .B(_13284_), .Y(_13286_) );
NAND3X1 NAND3X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_6618_), .B(_9087_), .C(_6617_), .Y(_13287_) );
NAND3X1 NAND3X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .B(_9089_), .C(_3671_), .Y(_13288_) );
NAND2X1 NAND2X1_2419 ( .gnd(gnd), .vdd(vdd), .A(_13287_), .B(_13288_), .Y(_13289_) );
NOR2X1 NOR2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_13286_), .B(_13289_), .Y(_13290_) );
NAND2X1 NAND2X1_2420 ( .gnd(gnd), .vdd(vdd), .A(_13283_), .B(_13290_), .Y(_13291_) );
NOR2X1 NOR2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_13276_), .B(_13291_), .Y(_13292_) );
NAND2X1 NAND2X1_2421 ( .gnd(gnd), .vdd(vdd), .A(_13261_), .B(_13292_), .Y(_13293_) );
NOR2X1 NOR2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_13230_), .B(_13293_), .Y(_13294_) );
NAND3X1 NAND3X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_6866_), .B(_9104_), .C(_6865_), .Y(_13295_) );
NAND3X1 NAND3X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_3974_), .B(_9099_), .C(_3973_), .Y(_13296_) );
NAND2X1 NAND2X1_2422 ( .gnd(gnd), .vdd(vdd), .A(_13296_), .B(_13295_), .Y(_13297_) );
NAND2X1 NAND2X1_2423 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__11_), .Y(_13298_) );
NAND3X1 NAND3X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_5107_), .B(_9102_), .C(_5106_), .Y(_13299_) );
NAND2X1 NAND2X1_2424 ( .gnd(gnd), .vdd(vdd), .A(_13298_), .B(_13299_), .Y(_13300_) );
NOR2X1 NOR2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_13300_), .B(_13297_), .Y(_13301_) );
NAND3X1 NAND3X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_15935_), .B(_9109_), .C(_15936_), .Y(_13302_) );
NAND3X1 NAND3X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_8400_), .B(_9113_), .C(_8401_), .Y(_13303_) );
NAND3X1 NAND3X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_16141_), .B(_9115_), .C(_16140_), .Y(_13304_) );
NAND3X1 NAND3X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_13302_), .B(_13303_), .C(_13304_), .Y(_13305_) );
NAND3X1 NAND3X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_406_), .C(_407_), .Y(_13306_) );
NAND3X1 NAND3X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_15878_), .B(_9120_), .C(_15879_), .Y(_13307_) );
AND2X2 AND2X2_1599 ( .gnd(gnd), .vdd(vdd), .A(_13307_), .B(_13306_), .Y(_13308_) );
AOI22X1 AOI22X1_453 ( .gnd(gnd), .vdd(vdd), .A(_201__11_), .B(_9124_), .C(_89__11_), .D(_9123_), .Y(_13309_) );
NAND2X1 NAND2X1_2425 ( .gnd(gnd), .vdd(vdd), .A(_13308_), .B(_13309_), .Y(_13310_) );
NAND3X1 NAND3X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_4752_), .B(_9127_), .C(_4753_), .Y(_13311_) );
NAND3X1 NAND3X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_4017_), .B(_9129_), .C(_4018_), .Y(_13312_) );
NAND2X1 NAND2X1_2426 ( .gnd(gnd), .vdd(vdd), .A(_13312_), .B(_13311_), .Y(_13313_) );
NOR3X1 NOR3X1_393 ( .gnd(gnd), .vdd(vdd), .A(_13305_), .B(_13313_), .C(_13310_), .Y(_13314_) );
NAND3X1 NAND3X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3434_), .C(_3435_), .Y(_13315_) );
NAND3X1 NAND3X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_5060_), .B(_9135_), .C(_5061_), .Y(_13316_) );
NAND3X1 NAND3X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_6943_), .B(_9137_), .C(_6944_), .Y(_13317_) );
NAND3X1 NAND3X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_13316_), .B(_13317_), .C(_13315_), .Y(_13318_) );
AOI22X1 AOI22X1_454 ( .gnd(gnd), .vdd(vdd), .A(_17__11_), .B(_9140_), .C(_2__11_), .D(_9141_), .Y(_13319_) );
NAND2X1 NAND2X1_2427 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__11_), .Y(_13320_) );
NAND2X1 NAND2X1_2428 ( .gnd(gnd), .vdd(vdd), .A(_9145_), .B(_200__11_), .Y(_13321_) );
NAND3X1 NAND3X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_13320_), .B(_13321_), .C(_13319_), .Y(_13322_) );
NOR2X1 NOR2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_13318_), .B(_13322_), .Y(_13323_) );
NAND3X1 NAND3X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_13301_), .B(_13323_), .C(_13314_), .Y(_13324_) );
AOI22X1 AOI22X1_455 ( .gnd(gnd), .vdd(vdd), .A(_21__11_), .B(_9150_), .C(_185__11_), .D(_9151_), .Y(_13325_) );
AOI22X1 AOI22X1_456 ( .gnd(gnd), .vdd(vdd), .A(_243__11_), .B(_9153_), .C(_253__11_), .D(_9154_), .Y(_13326_) );
NAND2X1 NAND2X1_2429 ( .gnd(gnd), .vdd(vdd), .A(_13325_), .B(_13326_), .Y(_13327_) );
AOI22X1 AOI22X1_457 ( .gnd(gnd), .vdd(vdd), .A(_46__11_), .B(_9158_), .C(_231__11_), .D(_9157_), .Y(_13328_) );
AOI22X1 AOI22X1_458 ( .gnd(gnd), .vdd(vdd), .A(_47__11_), .B(_9161_), .C(_244__11_), .D(_9160_), .Y(_13329_) );
NAND2X1 NAND2X1_2430 ( .gnd(gnd), .vdd(vdd), .A(_13329_), .B(_13328_), .Y(_13330_) );
NOR2X1 NOR2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_13327_), .B(_13330_), .Y(_13331_) );
NAND2X1 NAND2X1_2431 ( .gnd(gnd), .vdd(vdd), .A(_9165_), .B(_247__11_), .Y(_13332_) );
NAND2X1 NAND2X1_2432 ( .gnd(gnd), .vdd(vdd), .A(_9167_), .B(_30__11_), .Y(_13333_) );
AOI22X1 AOI22X1_459 ( .gnd(gnd), .vdd(vdd), .A(_218__11_), .B(_9169_), .C(_227__11_), .D(_9170_), .Y(_13334_) );
NAND3X1 NAND3X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_13332_), .B(_13333_), .C(_13334_), .Y(_13335_) );
AOI22X1 AOI22X1_460 ( .gnd(gnd), .vdd(vdd), .A(_123__11_), .B(_8928_), .C(_213__11_), .D(_8989_), .Y(_13336_) );
AOI22X1 AOI22X1_461 ( .gnd(gnd), .vdd(vdd), .A(_178__11_), .B(_9173_), .C(_29__11_), .D(_9176_), .Y(_13337_) );
NAND2X1 NAND2X1_2433 ( .gnd(gnd), .vdd(vdd), .A(_13336_), .B(_13337_), .Y(_13338_) );
NOR2X1 NOR2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_13338_), .B(_13335_), .Y(_13339_) );
NAND2X1 NAND2X1_2434 ( .gnd(gnd), .vdd(vdd), .A(_13331_), .B(_13339_), .Y(_13340_) );
AOI22X1 AOI22X1_462 ( .gnd(gnd), .vdd(vdd), .A(_234__11_), .B(_9182_), .C(_34__11_), .D(_9183_), .Y(_13341_) );
NAND2X1 NAND2X1_2435 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__11_), .Y(_13342_) );
NAND2X1 NAND2X1_2436 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__11_), .Y(_13343_) );
NAND3X1 NAND3X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_13342_), .B(_13343_), .C(_13341_), .Y(_13344_) );
NAND3X1 NAND3X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_15668_), .B(_9192_), .C(_15669_), .Y(_13345_) );
OAI21X1 OAI21X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_15617_), .B(_9195_), .C(_13345_), .Y(_13346_) );
NAND2X1 NAND2X1_2437 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__11_), .Y(_13347_) );
NAND3X1 NAND3X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_15724_), .B(_9199_), .C(_15725_), .Y(_13348_) );
NAND2X1 NAND2X1_2438 ( .gnd(gnd), .vdd(vdd), .A(_13347_), .B(_13348_), .Y(_13349_) );
NOR2X1 NOR2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_13349_), .B(_13346_), .Y(_13350_) );
NAND2X1 NAND2X1_2439 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__11_), .Y(_13351_) );
OAI21X1 OAI21X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_15320_), .B(_9206_), .C(_13351_), .Y(_13352_) );
NAND2X1 NAND2X1_2440 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__11_), .Y(_13353_) );
OAI21X1 OAI21X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_15110_), .B(_9211_), .C(_13353_), .Y(_13354_) );
NOR2X1 NOR2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(_13352_), .B(_13354_), .Y(_13355_) );
NOR3X1 NOR3X1_394 ( .gnd(gnd), .vdd(vdd), .A(_15985_), .B(_9215_), .C(_15986_), .Y(_13356_) );
NAND3X1 NAND3X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_15270_), .B(_9217_), .C(_15271_), .Y(_13357_) );
NAND3X1 NAND3X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_15218_), .B(_9219_), .C(_15217_), .Y(_13358_) );
NAND2X1 NAND2X1_2441 ( .gnd(gnd), .vdd(vdd), .A(_13358_), .B(_13357_), .Y(_13359_) );
NAND3X1 NAND3X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_15492_), .B(_9222_), .C(_15493_), .Y(_13360_) );
NAND3X1 NAND3X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_15439_), .B(_9224_), .C(_15438_), .Y(_13361_) );
NAND2X1 NAND2X1_2442 ( .gnd(gnd), .vdd(vdd), .A(_13360_), .B(_13361_), .Y(_13362_) );
NOR3X1 NOR3X1_395 ( .gnd(gnd), .vdd(vdd), .A(_13356_), .B(_13362_), .C(_13359_), .Y(_13363_) );
NAND3X1 NAND3X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_13355_), .B(_13363_), .C(_13350_), .Y(_13364_) );
NAND2X1 NAND2X1_2443 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__11_), .Y(_13365_) );
NAND3X1 NAND3X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_15550_), .B(_9233_), .C(_15551_), .Y(_13366_) );
AND2X2 AND2X2_1600 ( .gnd(gnd), .vdd(vdd), .A(_32__11_), .B(_10110_), .Y(_13367_) );
AND2X2 AND2X2_1601 ( .gnd(gnd), .vdd(vdd), .A(_186__11_), .B(_9298_), .Y(_13368_) );
AND2X2 AND2X2_1602 ( .gnd(gnd), .vdd(vdd), .A(_65__11_), .B(_9277_), .Y(_13369_) );
OR2X2 OR2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_13369_), .B(_13368_), .Y(_13370_) );
NOR3X1 NOR3X1_396 ( .gnd(gnd), .vdd(vdd), .A(_7474_), .B(_10471_), .C(_7475_), .Y(_13371_) );
NOR2X1 NOR2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_9267_), .B(_7057_), .Y(_13372_) );
NAND3X1 NAND3X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_8244_), .B(_9250_), .C(_8243_), .Y(_13373_) );
OAI21X1 OAI21X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_7015_), .B(_9288_), .C(_13373_), .Y(_13374_) );
NOR3X1 NOR3X1_397 ( .gnd(gnd), .vdd(vdd), .A(_13372_), .B(_13374_), .C(_13371_), .Y(_13375_) );
NAND3X1 NAND3X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_9268_), .C(_1179_), .Y(_13376_) );
OAI21X1 OAI21X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_15820_), .B(_11264_), .C(_13376_), .Y(_13377_) );
NAND2X1 NAND2X1_2444 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__11_), .Y(_13378_) );
OAI21X1 OAI21X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_7643_), .B(_9301_), .C(_13378_), .Y(_13379_) );
NOR2X1 NOR2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_13379_), .B(_13377_), .Y(_13380_) );
NAND2X1 NAND2X1_2445 ( .gnd(gnd), .vdd(vdd), .A(_13375_), .B(_13380_), .Y(_13381_) );
NOR3X1 NOR3X1_398 ( .gnd(gnd), .vdd(vdd), .A(_13367_), .B(_13370_), .C(_13381_), .Y(_13382_) );
NOR2X1 NOR2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .B(_5933_), .Y(_13383_) );
NAND3X1 NAND3X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_7102_), .B(_9244_), .C(_7101_), .Y(_13384_) );
OAI21X1 OAI21X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_12340_), .C(_13384_), .Y(_13385_) );
NAND3X1 NAND3X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_7684_), .B(_9321_), .C(_7685_), .Y(_13386_) );
OAI21X1 OAI21X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_4825_), .B(_9273_), .C(_13386_), .Y(_13387_) );
NOR3X1 NOR3X1_399 ( .gnd(gnd), .vdd(vdd), .A(_13385_), .B(_13383_), .C(_13387_), .Y(_13388_) );
NAND2X1 NAND2X1_2446 ( .gnd(gnd), .vdd(vdd), .A(_9260_), .B(_216__11_), .Y(_13389_) );
NAND2X1 NAND2X1_2447 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_173__11_), .Y(_13390_) );
NAND2X1 NAND2X1_2448 ( .gnd(gnd), .vdd(vdd), .A(_13389_), .B(_13390_), .Y(_13391_) );
NAND3X1 NAND3X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_3611_), .B(_9294_), .C(_3612_), .Y(_13392_) );
OAI21X1 OAI21X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .B(_9306_), .C(_13392_), .Y(_13393_) );
NOR2X1 NOR2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_13393_), .B(_13391_), .Y(_13394_) );
NAND3X1 NAND3X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_7727_), .B(_9248_), .C(_7728_), .Y(_13395_) );
OAI21X1 OAI21X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_8176_), .B(_9304_), .C(_13395_), .Y(_13396_) );
NAND2X1 NAND2X1_2449 ( .gnd(gnd), .vdd(vdd), .A(_1__11_), .B(_9242_), .Y(_13397_) );
NAND2X1 NAND2X1_2450 ( .gnd(gnd), .vdd(vdd), .A(_9262_), .B(_137__11_), .Y(_13398_) );
NAND2X1 NAND2X1_2451 ( .gnd(gnd), .vdd(vdd), .A(_13397_), .B(_13398_), .Y(_13399_) );
NOR2X1 NOR2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_13396_), .B(_13399_), .Y(_13400_) );
NAND3X1 NAND3X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_13400_), .B(_13388_), .C(_13394_), .Y(_13401_) );
NOR2X1 NOR2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_9312_), .B(_4788_), .Y(_13402_) );
NOR2X1 NOR2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_9763_), .B(_6439_), .Y(_13403_) );
AND2X2 AND2X2_1603 ( .gnd(gnd), .vdd(vdd), .A(_252__11_), .B(_9326_), .Y(_13404_) );
NOR3X1 NOR3X1_400 ( .gnd(gnd), .vdd(vdd), .A(_13402_), .B(_13403_), .C(_13404_), .Y(_13405_) );
AOI22X1 AOI22X1_463 ( .gnd(gnd), .vdd(vdd), .A(_233__11_), .B(_9310_), .C(_251__11_), .D(_9320_), .Y(_13406_) );
AOI22X1 AOI22X1_464 ( .gnd(gnd), .vdd(vdd), .A(_83__11_), .B(_9315_), .C(_31__11_), .D(_9283_), .Y(_13407_) );
NAND3X1 NAND3X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_13406_), .B(_13407_), .C(_13405_), .Y(_13408_) );
NOR2X1 NOR2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_13408_), .B(_13401_), .Y(_13409_) );
NAND3X1 NAND3X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_13366_), .B(_13382_), .C(_13409_), .Y(_13410_) );
AOI21X1 AOI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_157__11_), .B(_9232_), .C(_13410_), .Y(_13411_) );
AOI22X1 AOI22X1_465 ( .gnd(gnd), .vdd(vdd), .A(_155__11_), .B(_9333_), .C(_172__11_), .D(_9332_), .Y(_13412_) );
NAND3X1 NAND3X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_13412_), .B(_13411_), .C(_13365_), .Y(_13413_) );
NOR3X1 NOR3X1_401 ( .gnd(gnd), .vdd(vdd), .A(_13344_), .B(_13413_), .C(_13364_), .Y(_13414_) );
NAND2X1 NAND2X1_2452 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__11_), .Y(_13415_) );
NAND3X1 NAND3X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_9339_), .C(_461_), .Y(_13416_) );
AOI22X1 AOI22X1_466 ( .gnd(gnd), .vdd(vdd), .A(_111__11_), .B(_9342_), .C(_12__11_), .D(_9341_), .Y(_13417_) );
NAND3X1 NAND3X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_13417_), .B(_13415_), .C(_13416_), .Y(_13418_) );
AOI22X1 AOI22X1_467 ( .gnd(gnd), .vdd(vdd), .A(_100__11_), .B(_9346_), .C(_212__11_), .D(_9345_), .Y(_13419_) );
AOI22X1 AOI22X1_468 ( .gnd(gnd), .vdd(vdd), .A(_245__11_), .B(_9348_), .C(_140__11_), .D(_9349_), .Y(_13420_) );
NAND2X1 NAND2X1_2453 ( .gnd(gnd), .vdd(vdd), .A(_13420_), .B(_13419_), .Y(_13421_) );
NOR2X1 NOR2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_13418_), .B(_13421_), .Y(_13422_) );
AOI22X1 AOI22X1_469 ( .gnd(gnd), .vdd(vdd), .A(_232__11_), .B(_9354_), .C(_219__11_), .D(_9353_), .Y(_13423_) );
AOI22X1 AOI22X1_470 ( .gnd(gnd), .vdd(vdd), .A(_246__11_), .B(_9356_), .C(_226__11_), .D(_9357_), .Y(_13424_) );
NAND2X1 NAND2X1_2454 ( .gnd(gnd), .vdd(vdd), .A(_13424_), .B(_13423_), .Y(_13425_) );
NAND3X1 NAND3X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16193_), .C(_16194_), .Y(_13426_) );
OAI21X1 OAI21X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_9361_), .C(_13426_), .Y(_13427_) );
NAND3X1 NAND3X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16095_), .C(_16096_), .Y(_13428_) );
NAND3X1 NAND3X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16040_), .C(_16041_), .Y(_13429_) );
NAND2X1 NAND2X1_2455 ( .gnd(gnd), .vdd(vdd), .A(_13428_), .B(_13429_), .Y(_13430_) );
NOR2X1 NOR2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_13430_), .B(_13427_), .Y(_13431_) );
NAND3X1 NAND3X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_8682_), .B(_9371_), .C(_8681_), .Y(_13432_) );
NAND3X1 NAND3X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8574_), .C(_8573_), .Y(_13433_) );
NAND2X1 NAND2X1_2456 ( .gnd(gnd), .vdd(vdd), .A(_13433_), .B(_13432_), .Y(_13434_) );
NAND3X1 NAND3X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8627_), .C(_8628_), .Y(_13435_) );
NAND3X1 NAND3X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_324_), .C(_325_), .Y(_13436_) );
NAND2X1 NAND2X1_2457 ( .gnd(gnd), .vdd(vdd), .A(_13435_), .B(_13436_), .Y(_13437_) );
NOR2X1 NOR2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_13437_), .B(_13434_), .Y(_13438_) );
AOI22X1 AOI22X1_471 ( .gnd(gnd), .vdd(vdd), .A(_22__11_), .B(_9382_), .C(_3__11_), .D(_9383_), .Y(_13439_) );
NAND3X1 NAND3X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_13431_), .B(_13438_), .C(_13439_), .Y(_13440_) );
NOR2X1 NOR2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_13440_), .B(_13425_), .Y(_13441_) );
NAND3X1 NAND3X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_13422_), .B(_13414_), .C(_13441_), .Y(_13442_) );
NOR3X1 NOR3X1_402 ( .gnd(gnd), .vdd(vdd), .A(_13324_), .B(_13340_), .C(_13442_), .Y(_13443_) );
NAND3X1 NAND3X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_13167_), .B(_13443_), .C(_13294_), .Y(_13444_) );
NAND2X1 NAND2X1_2458 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__11_), .Y(_13445_) );
NAND2X1 NAND2X1_2459 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__11_), .Y(_13446_) );
NAND2X1 NAND2X1_2460 ( .gnd(gnd), .vdd(vdd), .A(_13446_), .B(_13445_), .Y(_13447_) );
NOR3X1 NOR3X1_403 ( .gnd(gnd), .vdd(vdd), .A(_13159_), .B(_13447_), .C(_13444_), .Y(_13448_) );
NOR3X1 NOR3X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1858_), .B(_9397_), .C(_1859_), .Y(_13449_) );
NAND3X1 NAND3X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1470_), .C(_1469_), .Y(_13450_) );
NAND3X1 NAND3X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_9453_), .B(_1424_), .C(_1423_), .Y(_13451_) );
NAND2X1 NAND2X1_2461 ( .gnd(gnd), .vdd(vdd), .A(_13450_), .B(_13451_), .Y(_13452_) );
NAND3X1 NAND3X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1514_), .C(_1513_), .Y(_13453_) );
NAND3X1 NAND3X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1297_), .C(_1296_), .Y(_13454_) );
NAND2X1 NAND2X1_2462 ( .gnd(gnd), .vdd(vdd), .A(_13453_), .B(_13454_), .Y(_13455_) );
NOR2X1 NOR2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_13455_), .B(_13452_), .Y(_13456_) );
AOI22X1 AOI22X1_472 ( .gnd(gnd), .vdd(vdd), .A(_125__11_), .B(_9411_), .C(_124__11_), .D(_9410_), .Y(_13457_) );
NAND3X1 NAND3X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_9413_), .C(_1115_), .Y(_13458_) );
NAND2X1 NAND2X1_2463 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__11_), .Y(_13459_) );
NAND3X1 NAND3X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_13458_), .B(_13459_), .C(_13457_), .Y(_13460_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_9421_), .C(_820_), .D(_9419_), .Y(_13461_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_9426_), .C(_705_), .D(_9424_), .Y(_13462_) );
NOR2X1 NOR2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_13461_), .B(_13462_), .Y(_13463_) );
NAND3X1 NAND3X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_667_), .C(_668_), .Y(_13464_) );
NAND3X1 NAND3X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_9431_), .C(_556_), .Y(_13465_) );
AOI22X1 AOI22X1_473 ( .gnd(gnd), .vdd(vdd), .A(_138__11_), .B(_9434_), .C(_229__11_), .D(_9433_), .Y(_13466_) );
NAND3X1 NAND3X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_13464_), .B(_13465_), .C(_13466_), .Y(_13467_) );
NAND3X1 NAND3X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7420_), .C(_7421_), .Y(_13468_) );
OAI21X1 OAI21X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_9440_), .C(_13468_), .Y(_13469_) );
NOR2X1 NOR2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_13469_), .B(_13467_), .Y(_13470_) );
NAND2X1 NAND2X1_2464 ( .gnd(gnd), .vdd(vdd), .A(_13470_), .B(_13463_), .Y(_13471_) );
NAND3X1 NAND3X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_1064_), .B(_9444_), .C(_1063_), .Y(_13472_) );
NAND2X1 NAND2X1_2465 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__11_), .Y(_13473_) );
AOI22X1 AOI22X1_474 ( .gnd(gnd), .vdd(vdd), .A(_130__11_), .B(_9449_), .C(_127__11_), .D(_9448_), .Y(_13474_) );
NAND3X1 NAND3X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_13472_), .B(_13473_), .C(_13474_), .Y(_13475_) );
NOR3X1 NOR3X1_405 ( .gnd(gnd), .vdd(vdd), .A(_13475_), .B(_13460_), .C(_13471_), .Y(_13476_) );
AOI22X1 AOI22X1_475 ( .gnd(gnd), .vdd(vdd), .A(_115__11_), .B(_9399_), .C(_114__11_), .D(_9454_), .Y(_13477_) );
NAND3X1 NAND3X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_13477_), .B(_13456_), .C(_13476_), .Y(_13478_) );
NAND3X1 NAND3X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(_9457_), .C(_1718_), .Y(_13479_) );
NAND2X1 NAND2X1_2466 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__11_), .Y(_13480_) );
NAND2X1 NAND2X1_2467 ( .gnd(gnd), .vdd(vdd), .A(_13480_), .B(_13479_), .Y(_13481_) );
NOR3X1 NOR3X1_406 ( .gnd(gnd), .vdd(vdd), .A(_13481_), .B(_13449_), .C(_13478_), .Y(_13482_) );
NAND3X1 NAND3X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_13152_), .B(_13482_), .C(_13448_), .Y(_13483_) );
NOR2X1 NOR2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_13151_), .B(_13483_), .Y(_13484_) );
NAND3X1 NAND3X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_13140_), .B(_13147_), .C(_13484_), .Y(_13485_) );
NOR3X1 NOR3X1_407 ( .gnd(gnd), .vdd(vdd), .A(_13129_), .B(_13132_), .C(_13485_), .Y(_13486_) );
NAND3X1 NAND3X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_13120_), .B(_13125_), .C(_13486_), .Y(_13487_) );
NAND3X1 NAND3X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_3073_), .B(_9473_), .C(_3074_), .Y(_13488_) );
NAND2X1 NAND2X1_2468 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__11_), .Y(_13489_) );
NAND2X1 NAND2X1_2469 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__11_), .Y(_13490_) );
NAND2X1 NAND2X1_2470 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__11_), .Y(_13491_) );
NAND3X1 NAND3X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_2445_), .B(_9468_), .C(_2446_), .Y(_13492_) );
NAND3X1 NAND3X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_13492_), .B(_13490_), .C(_13491_), .Y(_13493_) );
AOI21X1 AOI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_68__11_), .B(_9477_), .C(_13493_), .Y(_13494_) );
NAND3X1 NAND3X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_13494_), .B(_13488_), .C(_13489_), .Y(_13495_) );
NOR3X1 NOR3X1_408 ( .gnd(gnd), .vdd(vdd), .A(_13119_), .B(_13495_), .C(_13487_), .Y(_13496_) );
AOI21X1 AOI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_13112_), .B(_13496_), .C(rst), .Y(_0__11_) );
NAND2X1 NAND2X1_2471 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__12_), .Y(_13497_) );
NAND2X1 NAND2X1_2472 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__12_), .Y(_13498_) );
NAND2X1 NAND2X1_2473 ( .gnd(gnd), .vdd(vdd), .A(_13497_), .B(_13498_), .Y(_13499_) );
NAND2X1 NAND2X1_2474 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__12_), .Y(_13500_) );
NAND2X1 NAND2X1_2475 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__12_), .Y(_13501_) );
NAND2X1 NAND2X1_2476 ( .gnd(gnd), .vdd(vdd), .A(_13500_), .B(_13501_), .Y(_13502_) );
NOR2X1 NOR2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(_13499_), .B(_13502_), .Y(_13503_) );
NAND3X1 NAND3X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_3293_), .B(_8762_), .C(_3292_), .Y(_13504_) );
NAND3X1 NAND3X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_8765_), .C(_3242_), .Y(_13505_) );
AND2X2 AND2X2_1604 ( .gnd(gnd), .vdd(vdd), .A(_13505_), .B(_13504_), .Y(_13506_) );
AOI22X1 AOI22X1_476 ( .gnd(gnd), .vdd(vdd), .A(_62__12_), .B(_8774_), .C(_57__12_), .D(_8771_), .Y(_13507_) );
NAND2X1 NAND2X1_2477 ( .gnd(gnd), .vdd(vdd), .A(_13506_), .B(_13507_), .Y(_13508_) );
NAND2X1 NAND2X1_2478 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__12_), .Y(_13509_) );
NAND3X1 NAND3X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_2830_), .B(_8786_), .C(_2831_), .Y(_13510_) );
OAI21X1 OAI21X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_2721_), .B(_8792_), .C(_13510_), .Y(_13511_) );
NAND3X1 NAND3X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .B(_8794_), .C(_2660_), .Y(_13512_) );
OAI21X1 OAI21X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_2777_), .B(_8799_), .C(_13512_), .Y(_13513_) );
NOR2X1 NOR2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_13513_), .B(_13511_), .Y(_13514_) );
AOI22X1 AOI22X1_477 ( .gnd(gnd), .vdd(vdd), .A(_75__12_), .B(_8802_), .C(_74__12_), .D(_8803_), .Y(_13515_) );
AOI22X1 AOI22X1_478 ( .gnd(gnd), .vdd(vdd), .A(_80__12_), .B(_8805_), .C(_82__12_), .D(_8806_), .Y(_13516_) );
NAND2X1 NAND2X1_2479 ( .gnd(gnd), .vdd(vdd), .A(_13516_), .B(_13515_), .Y(_13517_) );
INVX1 INVX1_3881 ( .gnd(gnd), .vdd(vdd), .A(_84__12_), .Y(_13518_) );
NOR2X1 NOR2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_13518_), .Y(_13519_) );
NOR2X1 NOR2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2306_), .Y(_13520_) );
NAND2X1 NAND2X1_2480 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__12_), .Y(_13521_) );
NAND3X1 NAND3X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1928_), .C(_1929_), .Y(_13522_) );
NAND2X1 NAND2X1_2481 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_98__12_), .Y(_13523_) );
NAND3X1 NAND3X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_13522_), .B(_13521_), .C(_13523_), .Y(_13524_) );
NOR3X1 NOR3X1_409 ( .gnd(gnd), .vdd(vdd), .A(_13519_), .B(_13524_), .C(_13520_), .Y(_13525_) );
NAND3X1 NAND3X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_2266_), .B(_8829_), .C(_2267_), .Y(_13526_) );
NAND3X1 NAND3X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_2160_), .B(_8831_), .C(_2161_), .Y(_13527_) );
NAND2X1 NAND2X1_2482 ( .gnd(gnd), .vdd(vdd), .A(_13526_), .B(_13527_), .Y(_13528_) );
NAND3X1 NAND3X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .B(_8834_), .C(_2102_), .Y(_13529_) );
NAND3X1 NAND3X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_2212_), .B(_8836_), .C(_2213_), .Y(_13530_) );
NAND2X1 NAND2X1_2483 ( .gnd(gnd), .vdd(vdd), .A(_13529_), .B(_13530_), .Y(_13531_) );
NOR2X1 NOR2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_13531_), .B(_13528_), .Y(_13532_) );
AOI22X1 AOI22X1_479 ( .gnd(gnd), .vdd(vdd), .A(_92__12_), .B(_8843_), .C(_91__12_), .D(_8823_), .Y(_13533_) );
NAND2X1 NAND2X1_2484 ( .gnd(gnd), .vdd(vdd), .A(_8840_), .B(_93__12_), .Y(_13534_) );
NAND2X1 NAND2X1_2485 ( .gnd(gnd), .vdd(vdd), .A(_8841_), .B(_94__12_), .Y(_13535_) );
NAND3X1 NAND3X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_13534_), .B(_13535_), .C(_13533_), .Y(_13536_) );
NAND2X1 NAND2X1_2486 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__12_), .Y(_13537_) );
NAND3X1 NAND3X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1594_), .C(_1595_), .Y(_13538_) );
NAND3X1 NAND3X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_1388_), .B(_8857_), .C(_1387_), .Y(_13539_) );
NAND2X1 NAND2X1_2487 ( .gnd(gnd), .vdd(vdd), .A(_13539_), .B(_13538_), .Y(_13540_) );
NAND3X1 NAND3X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_1678_), .C(_1679_), .Y(_13541_) );
NAND3X1 NAND3X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_8862_), .C(_1255_), .Y(_13542_) );
NAND2X1 NAND2X1_2488 ( .gnd(gnd), .vdd(vdd), .A(_13541_), .B(_13542_), .Y(_13543_) );
OR2X2 OR2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_13543_), .B(_13540_), .Y(_13544_) );
NOR3X1 NOR3X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1218_), .B(_8867_), .C(_1219_), .Y(_13545_) );
AOI22X1 AOI22X1_480 ( .gnd(gnd), .vdd(vdd), .A(_191__12_), .B(_8873_), .C(_192__12_), .D(_8872_), .Y(_13546_) );
AOI22X1 AOI22X1_481 ( .gnd(gnd), .vdd(vdd), .A(_195__12_), .B(_8875_), .C(_193__12_), .D(_8876_), .Y(_13547_) );
NAND2X1 NAND2X1_2489 ( .gnd(gnd), .vdd(vdd), .A(_13546_), .B(_13547_), .Y(_13548_) );
AOI22X1 AOI22X1_482 ( .gnd(gnd), .vdd(vdd), .A(_188__12_), .B(_8879_), .C(_126__12_), .D(_8881_), .Y(_13549_) );
AOI22X1 AOI22X1_483 ( .gnd(gnd), .vdd(vdd), .A(_196__12_), .B(_8883_), .C(_194__12_), .D(_8884_), .Y(_13550_) );
NAND2X1 NAND2X1_2490 ( .gnd(gnd), .vdd(vdd), .A(_13549_), .B(_13550_), .Y(_13551_) );
NOR3X1 NOR3X1_411 ( .gnd(gnd), .vdd(vdd), .A(_13551_), .B(_13545_), .C(_13548_), .Y(_13552_) );
NAND3X1 NAND3X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_5840_), .B(_8893_), .C(_5839_), .Y(_13553_) );
NAND3X1 NAND3X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_4599_), .B(_8898_), .C(_4598_), .Y(_13554_) );
NAND2X1 NAND2X1_2491 ( .gnd(gnd), .vdd(vdd), .A(_13553_), .B(_13554_), .Y(_13555_) );
NAND3X1 NAND3X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_5537_), .B(_8901_), .C(_5536_), .Y(_13556_) );
NAND3X1 NAND3X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_7874_), .B(_8904_), .C(_7873_), .Y(_13557_) );
NAND2X1 NAND2X1_2492 ( .gnd(gnd), .vdd(vdd), .A(_13556_), .B(_13557_), .Y(_13558_) );
NOR2X1 NOR2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_13555_), .B(_13558_), .Y(_13559_) );
NAND3X1 NAND3X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_4099_), .B(_8909_), .C(_4098_), .Y(_13560_) );
NAND3X1 NAND3X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_3901_), .C(_3900_), .Y(_13561_) );
NAND2X1 NAND2X1_2493 ( .gnd(gnd), .vdd(vdd), .A(_13560_), .B(_13561_), .Y(_13562_) );
NAND3X1 NAND3X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_4640_), .B(_8914_), .C(_4639_), .Y(_13563_) );
NAND3X1 NAND3X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_6661_), .B(_8918_), .C(_6660_), .Y(_13564_) );
NAND2X1 NAND2X1_2494 ( .gnd(gnd), .vdd(vdd), .A(_13563_), .B(_13564_), .Y(_13565_) );
NOR2X1 NOR2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_13562_), .B(_13565_), .Y(_13566_) );
NAND2X1 NAND2X1_2495 ( .gnd(gnd), .vdd(vdd), .A(_13559_), .B(_13566_), .Y(_13567_) );
NAND3X1 NAND3X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_4980_), .B(_8926_), .C(_4979_), .Y(_13568_) );
NAND3X1 NAND3X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_8078_), .B(_8928_), .C(_8077_), .Y(_13569_) );
NAND2X1 NAND2X1_2496 ( .gnd(gnd), .vdd(vdd), .A(_13568_), .B(_13569_), .Y(_13570_) );
NAND3X1 NAND3X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_4502_), .B(_8931_), .C(_4501_), .Y(_13571_) );
NAND3X1 NAND3X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_8048_), .B(_8933_), .C(_8047_), .Y(_13572_) );
NAND2X1 NAND2X1_2497 ( .gnd(gnd), .vdd(vdd), .A(_13571_), .B(_13572_), .Y(_13573_) );
NOR2X1 NOR2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_13570_), .B(_13573_), .Y(_13574_) );
NAND3X1 NAND3X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_5194_), .B(_8937_), .C(_5193_), .Y(_13575_) );
NAND3X1 NAND3X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_7836_), .B(_8939_), .C(_7835_), .Y(_13576_) );
NAND2X1 NAND2X1_2498 ( .gnd(gnd), .vdd(vdd), .A(_13575_), .B(_13576_), .Y(_13577_) );
NAND3X1 NAND3X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_5156_), .B(_8942_), .C(_5155_), .Y(_13578_) );
NAND3X1 NAND3X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_5018_), .B(_8944_), .C(_5017_), .Y(_13579_) );
NAND2X1 NAND2X1_2499 ( .gnd(gnd), .vdd(vdd), .A(_13578_), .B(_13579_), .Y(_13580_) );
NOR2X1 NOR2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_13580_), .B(_13577_), .Y(_13581_) );
NAND2X1 NAND2X1_2500 ( .gnd(gnd), .vdd(vdd), .A(_13574_), .B(_13581_), .Y(_13582_) );
NOR2X1 NOR2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_13567_), .B(_13582_), .Y(_13583_) );
NAND3X1 NAND3X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_5617_), .B(_9160_), .C(_5616_), .Y(_13584_) );
NAND3X1 NAND3X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_3709_), .B(_9161_), .C(_3708_), .Y(_13585_) );
NAND2X1 NAND2X1_2501 ( .gnd(gnd), .vdd(vdd), .A(_13584_), .B(_13585_), .Y(_13586_) );
NAND3X1 NAND3X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_4560_), .B(_9150_), .C(_4559_), .Y(_13587_) );
NAND3X1 NAND3X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_7533_), .B(_9151_), .C(_7532_), .Y(_13588_) );
NAND2X1 NAND2X1_2502 ( .gnd(gnd), .vdd(vdd), .A(_13587_), .B(_13588_), .Y(_13589_) );
NOR2X1 NOR2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_13586_), .B(_13589_), .Y(_13590_) );
NAND3X1 NAND3X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_5590_), .B(_9356_), .C(_5589_), .Y(_13591_) );
NAND3X1 NAND3X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_6173_), .B(_9357_), .C(_6172_), .Y(_13592_) );
NAND2X1 NAND2X1_2503 ( .gnd(gnd), .vdd(vdd), .A(_13591_), .B(_13592_), .Y(_13593_) );
NAND3X1 NAND3X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_6028_), .B(_9157_), .C(_6027_), .Y(_13594_) );
NAND3X1 NAND3X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_3743_), .B(_9158_), .C(_3742_), .Y(_13595_) );
NAND2X1 NAND2X1_2504 ( .gnd(gnd), .vdd(vdd), .A(_13595_), .B(_13594_), .Y(_13596_) );
NOR2X1 NOR2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_13593_), .B(_13596_), .Y(_13597_) );
NAND2X1 NAND2X1_2505 ( .gnd(gnd), .vdd(vdd), .A(_13590_), .B(_13597_), .Y(_13598_) );
NAND3X1 NAND3X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_7766_), .B(_9173_), .C(_7765_), .Y(_13599_) );
NAND3X1 NAND3X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_3487_), .B(_8975_), .C(_3486_), .Y(_13600_) );
NAND2X1 NAND2X1_2506 ( .gnd(gnd), .vdd(vdd), .A(_13599_), .B(_13600_), .Y(_13601_) );
NAND3X1 NAND3X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_4062_), .B(_8978_), .C(_4061_), .Y(_13602_) );
NAND3X1 NAND3X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_8980_), .C(_4135_), .Y(_13603_) );
NAND2X1 NAND2X1_2507 ( .gnd(gnd), .vdd(vdd), .A(_13603_), .B(_13602_), .Y(_13604_) );
NOR2X1 NOR2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_13601_), .B(_13604_), .Y(_13605_) );
NAND3X1 NAND3X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_5645_), .B(_9153_), .C(_5644_), .Y(_13606_) );
NAND3X1 NAND3X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_5350_), .B(_9154_), .C(_5349_), .Y(_13607_) );
NAND2X1 NAND2X1_2508 ( .gnd(gnd), .vdd(vdd), .A(_13606_), .B(_13607_), .Y(_13608_) );
NAND3X1 NAND3X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_8011_), .B(_9177_), .C(_8010_), .Y(_13609_) );
NAND3X1 NAND3X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_6583_), .B(_8989_), .C(_6582_), .Y(_13610_) );
NAND2X1 NAND2X1_2509 ( .gnd(gnd), .vdd(vdd), .A(_13610_), .B(_13609_), .Y(_13611_) );
NOR2X1 NOR2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_13608_), .B(_13611_), .Y(_13612_) );
NAND2X1 NAND2X1_2510 ( .gnd(gnd), .vdd(vdd), .A(_13605_), .B(_13612_), .Y(_13613_) );
NOR2X1 NOR2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_13598_), .B(_13613_), .Y(_13614_) );
NAND2X1 NAND2X1_2511 ( .gnd(gnd), .vdd(vdd), .A(_13583_), .B(_13614_), .Y(_13615_) );
NAND3X1 NAND3X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .B(_8998_), .C(_4910_), .Y(_13616_) );
NAND3X1 NAND3X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_6518_), .B(_9002_), .C(_6517_), .Y(_13617_) );
NAND2X1 NAND2X1_2512 ( .gnd(gnd), .vdd(vdd), .A(_13616_), .B(_13617_), .Y(_13618_) );
NAND3X1 NAND3X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_5724_), .B(_9005_), .C(_5723_), .Y(_13619_) );
NAND3X1 NAND3X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_4872_), .B(_9007_), .C(_4871_), .Y(_13620_) );
NAND2X1 NAND2X1_2513 ( .gnd(gnd), .vdd(vdd), .A(_13619_), .B(_13620_), .Y(_13621_) );
NOR2X1 NOR2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_13618_), .B(_13621_), .Y(_13622_) );
NAND3X1 NAND3X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_5762_), .B(_9011_), .C(_5761_), .Y(_13623_) );
NAND3X1 NAND3X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_6804_), .B(_9013_), .C(_6803_), .Y(_13624_) );
NAND2X1 NAND2X1_2514 ( .gnd(gnd), .vdd(vdd), .A(_13623_), .B(_13624_), .Y(_13625_) );
NAND3X1 NAND3X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_6765_), .B(_9016_), .C(_6764_), .Y(_13626_) );
NAND3X1 NAND3X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_6551_), .B(_9174_), .C(_6550_), .Y(_13627_) );
NAND2X1 NAND2X1_2515 ( .gnd(gnd), .vdd(vdd), .A(_13626_), .B(_13627_), .Y(_13628_) );
NOR2X1 NOR2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_13628_), .B(_13625_), .Y(_13629_) );
NAND2X1 NAND2X1_2516 ( .gnd(gnd), .vdd(vdd), .A(_13622_), .B(_13629_), .Y(_13630_) );
NAND3X1 NAND3X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_6288_), .B(_9024_), .C(_6287_), .Y(_13631_) );
NAND3X1 NAND3X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_6360_), .B(_9026_), .C(_6359_), .Y(_13632_) );
NAND2X1 NAND2X1_2517 ( .gnd(gnd), .vdd(vdd), .A(_13631_), .B(_13632_), .Y(_13633_) );
NAND3X1 NAND3X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_6065_), .B(_9029_), .C(_6064_), .Y(_13634_) );
NAND3X1 NAND3X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_6123_), .B(_9031_), .C(_6122_), .Y(_13635_) );
NAND2X1 NAND2X1_2518 ( .gnd(gnd), .vdd(vdd), .A(_13634_), .B(_13635_), .Y(_13636_) );
NOR2X1 NOR2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_13633_), .B(_13636_), .Y(_13637_) );
NAND3X1 NAND3X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_5683_), .B(_9035_), .C(_5682_), .Y(_13638_) );
NAND3X1 NAND3X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_4679_), .B(_9037_), .C(_4678_), .Y(_13639_) );
NAND2X1 NAND2X1_2519 ( .gnd(gnd), .vdd(vdd), .A(_13639_), .B(_13638_), .Y(_13640_) );
NAND3X1 NAND3X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_6324_), .B(_9040_), .C(_6323_), .Y(_13641_) );
NAND3X1 NAND3X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_4341_), .B(_9042_), .C(_4340_), .Y(_13642_) );
NAND2X1 NAND2X1_2520 ( .gnd(gnd), .vdd(vdd), .A(_13641_), .B(_13642_), .Y(_13643_) );
NOR2X1 NOR2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_13643_), .B(_13640_), .Y(_13644_) );
NAND2X1 NAND2X1_2521 ( .gnd(gnd), .vdd(vdd), .A(_13637_), .B(_13644_), .Y(_13645_) );
NOR2X1 NOR2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_13630_), .B(_13645_), .Y(_13646_) );
NAND3X1 NAND3X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_6212_), .B(_9048_), .C(_6211_), .Y(_13647_) );
NAND3X1 NAND3X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_7947_), .B(_9050_), .C(_7946_), .Y(_13648_) );
NAND2X1 NAND2X1_2522 ( .gnd(gnd), .vdd(vdd), .A(_13647_), .B(_13648_), .Y(_13649_) );
NAND3X1 NAND3X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_5495_), .B(_9053_), .C(_5494_), .Y(_13650_) );
NAND3X1 NAND3X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_7910_), .B(_9055_), .C(_7909_), .Y(_13651_) );
NAND2X1 NAND2X1_2523 ( .gnd(gnd), .vdd(vdd), .A(_13650_), .B(_13651_), .Y(_13652_) );
NOR2X1 NOR2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_13649_), .B(_13652_), .Y(_13653_) );
NAND3X1 NAND3X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_4462_), .B(_9059_), .C(_4461_), .Y(_13654_) );
NAND3X1 NAND3X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_4422_), .B(_9061_), .C(_4421_), .Y(_13655_) );
NAND2X1 NAND2X1_2524 ( .gnd(gnd), .vdd(vdd), .A(_13654_), .B(_13655_), .Y(_13656_) );
NAND3X1 NAND3X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_6250_), .B(_9064_), .C(_6249_), .Y(_13657_) );
NAND3X1 NAND3X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_4382_), .B(_9066_), .C(_4381_), .Y(_13658_) );
NAND2X1 NAND2X1_2525 ( .gnd(gnd), .vdd(vdd), .A(_13657_), .B(_13658_), .Y(_13659_) );
NOR2X1 NOR2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_13659_), .B(_13656_), .Y(_13660_) );
NAND2X1 NAND2X1_2526 ( .gnd(gnd), .vdd(vdd), .A(_13653_), .B(_13660_), .Y(_13661_) );
NAND3X1 NAND3X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_7606_), .B(_9071_), .C(_7605_), .Y(_13662_) );
NAND3X1 NAND3X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_7570_), .B(_9073_), .C(_7569_), .Y(_13663_) );
NAND2X1 NAND2X1_2527 ( .gnd(gnd), .vdd(vdd), .A(_13662_), .B(_13663_), .Y(_13664_) );
NAND3X1 NAND3X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_5800_), .B(_9076_), .C(_5799_), .Y(_13665_) );
NAND3X1 NAND3X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_9078_), .C(_3525_), .Y(_13666_) );
NAND2X1 NAND2X1_2528 ( .gnd(gnd), .vdd(vdd), .A(_13665_), .B(_13666_), .Y(_13667_) );
NOR2X1 NOR2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_13664_), .B(_13667_), .Y(_13668_) );
NAND3X1 NAND3X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_5454_), .B(_9082_), .C(_5453_), .Y(_13669_) );
NAND3X1 NAND3X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_3822_), .B(_9084_), .C(_3821_), .Y(_13670_) );
NAND2X1 NAND2X1_2529 ( .gnd(gnd), .vdd(vdd), .A(_13670_), .B(_13669_), .Y(_13671_) );
NAND3X1 NAND3X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_6621_), .B(_9087_), .C(_6620_), .Y(_13672_) );
NAND3X1 NAND3X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(_9089_), .C(_3674_), .Y(_13673_) );
NAND2X1 NAND2X1_2530 ( .gnd(gnd), .vdd(vdd), .A(_13672_), .B(_13673_), .Y(_13674_) );
NOR2X1 NOR2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_13671_), .B(_13674_), .Y(_13675_) );
NAND2X1 NAND2X1_2531 ( .gnd(gnd), .vdd(vdd), .A(_13668_), .B(_13675_), .Y(_13676_) );
NOR2X1 NOR2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_13661_), .B(_13676_), .Y(_13677_) );
NAND2X1 NAND2X1_2532 ( .gnd(gnd), .vdd(vdd), .A(_13646_), .B(_13677_), .Y(_13678_) );
NOR2X1 NOR2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_13615_), .B(_13678_), .Y(_13679_) );
NAND2X1 NAND2X1_2533 ( .gnd(gnd), .vdd(vdd), .A(_9143_), .B(_205__12_), .Y(_13680_) );
NAND3X1 NAND3X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_6982_), .B(_9145_), .C(_6981_), .Y(_13681_) );
NAND2X1 NAND2X1_2534 ( .gnd(gnd), .vdd(vdd), .A(_13680_), .B(_13681_), .Y(_13682_) );
NAND3X1 NAND3X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_5063_), .B(_9135_), .C(_5064_), .Y(_13683_) );
NAND3X1 NAND3X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_6946_), .B(_9137_), .C(_6945_), .Y(_13684_) );
NAND2X1 NAND2X1_2535 ( .gnd(gnd), .vdd(vdd), .A(_13683_), .B(_13684_), .Y(_13685_) );
NOR2X1 NOR2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_13685_), .B(_13682_), .Y(_13686_) );
NAND3X1 NAND3X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_16143_), .B(_9115_), .C(_16144_), .Y(_13687_) );
NAND3X1 NAND3X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_8403_), .B(_9113_), .C(_8404_), .Y(_13688_) );
NAND3X1 NAND3X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_15938_), .B(_9109_), .C(_15939_), .Y(_13689_) );
NAND3X1 NAND3X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_13687_), .B(_13689_), .C(_13688_), .Y(_13690_) );
NAND3X1 NAND3X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_9118_), .B(_409_), .C(_410_), .Y(_13691_) );
NAND3X1 NAND3X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_15881_), .B(_9120_), .C(_15882_), .Y(_13692_) );
AND2X2 AND2X2_1605 ( .gnd(gnd), .vdd(vdd), .A(_13692_), .B(_13691_), .Y(_13693_) );
AOI22X1 AOI22X1_484 ( .gnd(gnd), .vdd(vdd), .A(_201__12_), .B(_9124_), .C(_89__12_), .D(_9123_), .Y(_13694_) );
NAND2X1 NAND2X1_2536 ( .gnd(gnd), .vdd(vdd), .A(_13693_), .B(_13694_), .Y(_13695_) );
NAND3X1 NAND3X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_4712_), .B(_9140_), .C(_4713_), .Y(_13696_) );
OAI21X1 OAI21X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_5251_), .B(_10036_), .C(_13696_), .Y(_13697_) );
NOR3X1 NOR3X1_412 ( .gnd(gnd), .vdd(vdd), .A(_13690_), .B(_13697_), .C(_13695_), .Y(_13698_) );
NAND3X1 NAND3X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_9133_), .B(_3437_), .C(_3438_), .Y(_13699_) );
NAND2X1 NAND2X1_2537 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__12_), .Y(_13700_) );
NAND3X1 NAND3X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .B(_9102_), .C(_5110_), .Y(_13701_) );
NAND3X1 NAND3X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_13699_), .B(_13701_), .C(_13700_), .Y(_13702_) );
AOI22X1 AOI22X1_485 ( .gnd(gnd), .vdd(vdd), .A(_38__12_), .B(_9129_), .C(_16__12_), .D(_9127_), .Y(_13703_) );
NAND2X1 NAND2X1_2538 ( .gnd(gnd), .vdd(vdd), .A(_9104_), .B(_204__12_), .Y(_13704_) );
NAND2X1 NAND2X1_2539 ( .gnd(gnd), .vdd(vdd), .A(_9099_), .B(_39__12_), .Y(_13705_) );
NAND3X1 NAND3X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_13705_), .B(_13704_), .C(_13703_), .Y(_13706_) );
NOR2X1 NOR2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_13702_), .B(_13706_), .Y(_13707_) );
NAND3X1 NAND3X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_13686_), .B(_13707_), .C(_13698_), .Y(_13708_) );
AOI22X1 AOI22X1_486 ( .gnd(gnd), .vdd(vdd), .A(_30__12_), .B(_9167_), .C(_227__12_), .D(_9170_), .Y(_13709_) );
AOI22X1 AOI22X1_487 ( .gnd(gnd), .vdd(vdd), .A(_209__12_), .B(_8957_), .C(_33__12_), .D(_8991_), .Y(_13710_) );
NAND2X1 NAND2X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_13709_), .B(_13710_), .Y(_13711_) );
AOI22X1 AOI22X1_488 ( .gnd(gnd), .vdd(vdd), .A(_44__12_), .B(_8968_), .C(_42__12_), .D(_8963_), .Y(_13712_) );
AOI22X1 AOI22X1_489 ( .gnd(gnd), .vdd(vdd), .A(_236__12_), .B(_8955_), .C(_208__12_), .D(_8950_), .Y(_13713_) );
NAND2X1 NAND2X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_13712_), .B(_13713_), .Y(_13714_) );
NOR2X1 NOR2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_13711_), .B(_13714_), .Y(_13715_) );
AOI22X1 AOI22X1_490 ( .gnd(gnd), .vdd(vdd), .A(_22__12_), .B(_9382_), .C(_3__12_), .D(_9383_), .Y(_13716_) );
AOI22X1 AOI22X1_491 ( .gnd(gnd), .vdd(vdd), .A(_232__12_), .B(_9354_), .C(_219__12_), .D(_9353_), .Y(_13717_) );
NAND2X1 NAND2X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_13716_), .B(_13717_), .Y(_13718_) );
AOI22X1 AOI22X1_492 ( .gnd(gnd), .vdd(vdd), .A(_255__12_), .B(_8986_), .C(_254__12_), .D(_8984_), .Y(_13719_) );
AOI22X1 AOI22X1_493 ( .gnd(gnd), .vdd(vdd), .A(_203__12_), .B(_9018_), .C(_156__12_), .D(_8973_), .Y(_13720_) );
NAND2X1 NAND2X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_13720_), .B(_13719_), .Y(_13721_) );
NOR2X1 NOR2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_13718_), .B(_13721_), .Y(_13722_) );
NAND2X1 NAND2X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_13715_), .B(_13722_), .Y(_13723_) );
AOI22X1 AOI22X1_494 ( .gnd(gnd), .vdd(vdd), .A(_234__12_), .B(_9182_), .C(_34__12_), .D(_9183_), .Y(_13724_) );
NAND2X1 NAND2X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_9185_), .B(_45__12_), .Y(_13725_) );
NAND2X1 NAND2X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_9188_), .B(_23__12_), .Y(_13726_) );
NAND3X1 NAND3X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_13725_), .B(_13726_), .C(_13724_), .Y(_13727_) );
NAND3X1 NAND3X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_15671_), .B(_9192_), .C(_15672_), .Y(_13728_) );
OAI21X1 OAI21X1_2540 ( .gnd(gnd), .vdd(vdd), .A(_15619_), .B(_9195_), .C(_13728_), .Y(_13729_) );
NAND2X1 NAND2X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_9197_), .B(_164__12_), .Y(_13730_) );
NAND3X1 NAND3X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_15727_), .B(_9199_), .C(_15728_), .Y(_13731_) );
NAND2X1 NAND2X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_13730_), .B(_13731_), .Y(_13732_) );
NOR2X1 NOR2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_13732_), .B(_13729_), .Y(_13733_) );
NAND2X1 NAND2X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_9203_), .B(_165__12_), .Y(_13734_) );
OAI21X1 OAI21X1_2541 ( .gnd(gnd), .vdd(vdd), .A(_15322_), .B(_9206_), .C(_13734_), .Y(_13735_) );
NAND2X1 NAND2X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_9208_), .B(_170__12_), .Y(_13736_) );
OAI21X1 OAI21X1_2542 ( .gnd(gnd), .vdd(vdd), .A(_15112_), .B(_9211_), .C(_13736_), .Y(_13737_) );
NOR2X1 NOR2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_13735_), .B(_13737_), .Y(_13738_) );
NOR3X1 NOR3X1_413 ( .gnd(gnd), .vdd(vdd), .A(_15987_), .B(_9215_), .C(_15988_), .Y(_13739_) );
NAND3X1 NAND3X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_15273_), .B(_9217_), .C(_15274_), .Y(_13740_) );
NAND3X1 NAND3X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_15221_), .B(_9219_), .C(_15220_), .Y(_13741_) );
NAND2X1 NAND2X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_13741_), .B(_13740_), .Y(_13742_) );
NAND3X1 NAND3X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_15495_), .B(_9222_), .C(_15496_), .Y(_13743_) );
NAND3X1 NAND3X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_15442_), .B(_9224_), .C(_15441_), .Y(_13744_) );
NAND2X1 NAND2X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_13743_), .B(_13744_), .Y(_13745_) );
NOR3X1 NOR3X1_414 ( .gnd(gnd), .vdd(vdd), .A(_13739_), .B(_13745_), .C(_13742_), .Y(_13746_) );
NAND3X1 NAND3X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_13738_), .B(_13746_), .C(_13733_), .Y(_13747_) );
NAND2X1 NAND2X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__12_), .Y(_13748_) );
NAND3X1 NAND3X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_15553_), .B(_9233_), .C(_15554_), .Y(_13749_) );
NOR2X1 NOR2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_8178_), .Y(_13750_) );
NOR2X1 NOR2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_9259_), .B(_6474_), .Y(_13751_) );
NOR2X1 NOR2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_13751_), .B(_13750_), .Y(_13752_) );
OAI21X1 OAI21X1_2543 ( .gnd(gnd), .vdd(vdd), .A(_3615_), .B(_9295_), .C(_13752_), .Y(_13753_) );
NAND3X1 NAND3X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_8208_), .B(_9286_), .C(_8209_), .Y(_13754_) );
OAI21X1 OAI21X1_2544 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_9263_), .C(_13754_), .Y(_13755_) );
NOR3X1 NOR3X1_415 ( .gnd(gnd), .vdd(vdd), .A(_7476_), .B(_10471_), .C(_7477_), .Y(_13756_) );
NOR2X1 NOR2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_9254_), .B(_4196_), .Y(_13757_) );
NOR3X1 NOR3X1_416 ( .gnd(gnd), .vdd(vdd), .A(_13755_), .B(_13757_), .C(_13756_), .Y(_13758_) );
NAND3X1 NAND3X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_8246_), .B(_9250_), .C(_8247_), .Y(_13759_) );
OAI21X1 OAI21X1_2545 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_10468_), .C(_13759_), .Y(_13760_) );
NAND3X1 NAND3X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_9268_), .C(_1182_), .Y(_13761_) );
OAI21X1 OAI21X1_2546 ( .gnd(gnd), .vdd(vdd), .A(_7646_), .B(_9301_), .C(_13761_), .Y(_13762_) );
NOR2X1 NOR2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_13760_), .B(_13762_), .Y(_13763_) );
NAND2X1 NAND2X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_13758_), .B(_13763_), .Y(_13764_) );
NOR2X1 NOR2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_13764_), .B(_13753_), .Y(_13765_) );
NAND3X1 NAND3X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_6441_), .B(_9281_), .C(_6442_), .Y(_13766_) );
NAND2X1 NAND2X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__12_), .Y(_13767_) );
NAND3X1 NAND3X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_7104_), .B(_9244_), .C(_7105_), .Y(_13768_) );
NAND3X1 NAND3X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_13766_), .B(_13767_), .C(_13768_), .Y(_13769_) );
NAND3X1 NAND3X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_2366_), .B(_9315_), .C(_2367_), .Y(_13770_) );
OAI21X1 OAI21X1_2547 ( .gnd(gnd), .vdd(vdd), .A(_5378_), .B(_9325_), .C(_13770_), .Y(_13771_) );
NOR2X1 NOR2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_13771_), .B(_13769_), .Y(_13772_) );
AOI22X1 AOI22X1_495 ( .gnd(gnd), .vdd(vdd), .A(_154__12_), .B(_9292_), .C(_180__12_), .D(_9248_), .Y(_13773_) );
AOI22X1 AOI22X1_496 ( .gnd(gnd), .vdd(vdd), .A(_186__12_), .B(_9298_), .C(_198__12_), .D(_9266_), .Y(_13774_) );
AND2X2 AND2X2_1606 ( .gnd(gnd), .vdd(vdd), .A(_13773_), .B(_13774_), .Y(_13775_) );
NAND2X1 NAND2X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_1__12_), .B(_9242_), .Y(_13776_) );
NAND2X1 NAND2X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_9255_), .B(_101__12_), .Y(_13777_) );
NAND2X1 NAND2X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_13776_), .B(_13777_), .Y(_13778_) );
NAND2X1 NAND2X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_9275_), .B(_173__12_), .Y(_13779_) );
OAI21X1 OAI21X1_2548 ( .gnd(gnd), .vdd(vdd), .A(_3568_), .B(_9306_), .C(_13779_), .Y(_13780_) );
NOR2X1 NOR2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_13778_), .B(_13780_), .Y(_13781_) );
NAND3X1 NAND3X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_13772_), .B(_13775_), .C(_13781_), .Y(_13782_) );
NAND3X1 NAND3X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_5971_), .B(_9310_), .C(_5972_), .Y(_13783_) );
OAI21X1 OAI21X1_2549 ( .gnd(gnd), .vdd(vdd), .A(_4828_), .B(_9273_), .C(_13783_), .Y(_13784_) );
AOI21X1 AOI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_235__12_), .B(_9324_), .C(_13784_), .Y(_13785_) );
AOI22X1 AOI22X1_497 ( .gnd(gnd), .vdd(vdd), .A(_181__12_), .B(_9321_), .C(_15__12_), .D(_9313_), .Y(_13786_) );
AOI22X1 AOI22X1_498 ( .gnd(gnd), .vdd(vdd), .A(_31__12_), .B(_9283_), .C(_251__12_), .D(_9320_), .Y(_13787_) );
NAND3X1 NAND3X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_13786_), .B(_13787_), .C(_13785_), .Y(_13788_) );
NOR2X1 NOR2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_13788_), .B(_13782_), .Y(_13789_) );
NAND3X1 NAND3X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_13749_), .B(_13765_), .C(_13789_), .Y(_13790_) );
AOI21X1 AOI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_157__12_), .B(_9232_), .C(_13790_), .Y(_13791_) );
AOI22X1 AOI22X1_499 ( .gnd(gnd), .vdd(vdd), .A(_155__12_), .B(_9333_), .C(_172__12_), .D(_9332_), .Y(_13792_) );
NAND3X1 NAND3X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_13792_), .B(_13791_), .C(_13748_), .Y(_13793_) );
NOR3X1 NOR3X1_417 ( .gnd(gnd), .vdd(vdd), .A(_13727_), .B(_13793_), .C(_13747_), .Y(_13794_) );
NAND2X1 NAND2X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__12_), .Y(_13795_) );
NAND3X1 NAND3X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_9339_), .C(_464_), .Y(_13796_) );
AOI22X1 AOI22X1_500 ( .gnd(gnd), .vdd(vdd), .A(_111__12_), .B(_9342_), .C(_12__12_), .D(_9341_), .Y(_13797_) );
NAND3X1 NAND3X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_13797_), .B(_13795_), .C(_13796_), .Y(_13798_) );
AOI22X1 AOI22X1_501 ( .gnd(gnd), .vdd(vdd), .A(_100__12_), .B(_9346_), .C(_212__12_), .D(_9345_), .Y(_13799_) );
AOI22X1 AOI22X1_502 ( .gnd(gnd), .vdd(vdd), .A(_245__12_), .B(_9348_), .C(_140__12_), .D(_9349_), .Y(_13800_) );
NAND2X1 NAND2X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_13800_), .B(_13799_), .Y(_13801_) );
NOR2X1 NOR2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_13798_), .B(_13801_), .Y(_13802_) );
AOI22X1 AOI22X1_503 ( .gnd(gnd), .vdd(vdd), .A(_40__12_), .B(_8952_), .C(_29__12_), .D(_9176_), .Y(_13803_) );
AOI22X1 AOI22X1_504 ( .gnd(gnd), .vdd(vdd), .A(_218__12_), .B(_9169_), .C(_247__12_), .D(_9165_), .Y(_13804_) );
NAND2X1 NAND2X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_13804_), .B(_13803_), .Y(_13805_) );
NAND3X1 NAND3X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_9362_), .B(_16196_), .C(_16197_), .Y(_13806_) );
OAI21X1 OAI21X1_2550 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_9361_), .C(_13806_), .Y(_13807_) );
NAND3X1 NAND3X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16098_), .C(_16099_), .Y(_13808_) );
NAND3X1 NAND3X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16043_), .C(_16044_), .Y(_13809_) );
NAND2X1 NAND2X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_13808_), .B(_13809_), .Y(_13810_) );
NOR2X1 NOR2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_13810_), .B(_13807_), .Y(_13811_) );
NAND3X1 NAND3X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_8685_), .B(_9371_), .C(_8684_), .Y(_13812_) );
NAND3X1 NAND3X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8577_), .C(_8576_), .Y(_13813_) );
NAND2X1 NAND2X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_13813_), .B(_13812_), .Y(_13814_) );
NAND3X1 NAND3X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8630_), .C(_8631_), .Y(_13815_) );
NAND3X1 NAND3X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_327_), .C(_328_), .Y(_13816_) );
NAND2X1 NAND2X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_13815_), .B(_13816_), .Y(_13817_) );
NOR2X1 NOR2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_13817_), .B(_13814_), .Y(_13818_) );
AOI22X1 AOI22X1_505 ( .gnd(gnd), .vdd(vdd), .A(_237__12_), .B(_8966_), .C(_177__12_), .D(_8961_), .Y(_13819_) );
NAND3X1 NAND3X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_13811_), .B(_13818_), .C(_13819_), .Y(_13820_) );
NOR2X1 NOR2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_13820_), .B(_13805_), .Y(_13821_) );
NAND3X1 NAND3X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_13802_), .B(_13794_), .C(_13821_), .Y(_13822_) );
NOR3X1 NOR3X1_418 ( .gnd(gnd), .vdd(vdd), .A(_13708_), .B(_13723_), .C(_13822_), .Y(_13823_) );
NAND3X1 NAND3X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_13552_), .B(_13823_), .C(_13679_), .Y(_13824_) );
NAND2X1 NAND2X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__12_), .Y(_13825_) );
NAND2X1 NAND2X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__12_), .Y(_13826_) );
NAND2X1 NAND2X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_13825_), .B(_13826_), .Y(_13827_) );
NOR3X1 NOR3X1_419 ( .gnd(gnd), .vdd(vdd), .A(_13544_), .B(_13827_), .C(_13824_), .Y(_13828_) );
NOR3X1 NOR3X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_9397_), .C(_1861_), .Y(_13829_) );
NAND3X1 NAND3X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_9399_), .B(_1330_), .C(_1329_), .Y(_13830_) );
NAND3X1 NAND3X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_1300_), .C(_1299_), .Y(_13831_) );
NAND2X1 NAND2X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_13830_), .B(_13831_), .Y(_13832_) );
NAND3X1 NAND3X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_1517_), .C(_1516_), .Y(_13833_) );
NAND3X1 NAND3X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_9406_), .B(_1473_), .C(_1472_), .Y(_13834_) );
NAND2X1 NAND2X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_13833_), .B(_13834_), .Y(_13835_) );
NOR2X1 NOR2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_13835_), .B(_13832_), .Y(_13836_) );
AOI22X1 AOI22X1_506 ( .gnd(gnd), .vdd(vdd), .A(_125__12_), .B(_9411_), .C(_122__12_), .D(_9444_), .Y(_13837_) );
NAND3X1 NAND3X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_1119_), .B(_9413_), .C(_1118_), .Y(_13838_) );
NAND2X1 NAND2X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_9415_), .B(_120__12_), .Y(_13839_) );
NAND3X1 NAND3X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_13838_), .B(_13839_), .C(_13837_), .Y(_13840_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_9421_), .C(_823_), .D(_9419_), .Y(_13841_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_9426_), .C(_708_), .D(_9424_), .Y(_13842_) );
NOR2X1 NOR2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_13841_), .B(_13842_), .Y(_13843_) );
NAND3X1 NAND3X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_7423_), .C(_7424_), .Y(_13844_) );
NAND2X1 NAND2X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__12_), .Y(_13845_) );
AOI22X1 AOI22X1_507 ( .gnd(gnd), .vdd(vdd), .A(_229__12_), .B(_9433_), .C(_139__12_), .D(_9431_), .Y(_13846_) );
NAND3X1 NAND3X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_13845_), .B(_13844_), .C(_13846_), .Y(_13847_) );
NAND3X1 NAND3X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_670_), .C(_671_), .Y(_13848_) );
OAI21X1 OAI21X1_2551 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_9440_), .C(_13848_), .Y(_13849_) );
NOR2X1 NOR2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_13849_), .B(_13847_), .Y(_13850_) );
NAND2X1 NAND2X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_13850_), .B(_13843_), .Y(_13851_) );
NAND3X1 NAND3X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_1024_), .B(_9410_), .C(_1023_), .Y(_13852_) );
NAND2X1 NAND2X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__12_), .Y(_13853_) );
AOI22X1 AOI22X1_508 ( .gnd(gnd), .vdd(vdd), .A(_130__12_), .B(_9449_), .C(_127__12_), .D(_9448_), .Y(_13854_) );
NAND3X1 NAND3X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_13852_), .B(_13853_), .C(_13854_), .Y(_13855_) );
NOR3X1 NOR3X1_421 ( .gnd(gnd), .vdd(vdd), .A(_13855_), .B(_13840_), .C(_13851_), .Y(_13856_) );
AOI22X1 AOI22X1_509 ( .gnd(gnd), .vdd(vdd), .A(_114__12_), .B(_9454_), .C(_110__12_), .D(_9453_), .Y(_13857_) );
NAND3X1 NAND3X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_13836_), .B(_13857_), .C(_13856_), .Y(_13858_) );
NAND3X1 NAND3X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_1720_), .B(_9457_), .C(_1721_), .Y(_13859_) );
NAND2X1 NAND2X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_9459_), .B(_102__12_), .Y(_13860_) );
NAND2X1 NAND2X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_13860_), .B(_13859_), .Y(_13861_) );
NOR3X1 NOR3X1_422 ( .gnd(gnd), .vdd(vdd), .A(_13861_), .B(_13829_), .C(_13858_), .Y(_13862_) );
NAND3X1 NAND3X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_13537_), .B(_13862_), .C(_13828_), .Y(_13863_) );
NOR2X1 NOR2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_13536_), .B(_13863_), .Y(_13864_) );
NAND3X1 NAND3X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_13525_), .B(_13532_), .C(_13864_), .Y(_13865_) );
NAND2X1 NAND2X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__12_), .Y(_13866_) );
NAND3X1 NAND3X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_2448_), .B(_9468_), .C(_2449_), .Y(_13867_) );
NAND2X1 NAND2X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_13867_), .B(_13866_), .Y(_13868_) );
NOR3X1 NOR3X1_423 ( .gnd(gnd), .vdd(vdd), .A(_13517_), .B(_13868_), .C(_13865_), .Y(_13869_) );
NAND3X1 NAND3X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_13509_), .B(_13514_), .C(_13869_), .Y(_13870_) );
NAND3X1 NAND3X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_3076_), .B(_9473_), .C(_3077_), .Y(_13871_) );
NAND2X1 NAND2X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__12_), .Y(_13872_) );
NAND2X1 NAND2X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__12_), .Y(_13873_) );
NAND2X1 NAND2X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__12_), .Y(_13874_) );
NAND2X1 NAND2X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_9482_), .B(_76__12_), .Y(_13875_) );
NAND3X1 NAND3X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_13875_), .B(_13873_), .C(_13874_), .Y(_13876_) );
AOI21X1 AOI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_68__12_), .B(_9477_), .C(_13876_), .Y(_13877_) );
NAND3X1 NAND3X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_13871_), .B(_13877_), .C(_13872_), .Y(_13878_) );
NOR3X1 NOR3X1_424 ( .gnd(gnd), .vdd(vdd), .A(_13508_), .B(_13878_), .C(_13870_), .Y(_13879_) );
AOI21X1 AOI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_13503_), .B(_13879_), .C(rst), .Y(_0__12_) );
NAND2X1 NAND2X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__13_), .Y(_13880_) );
NAND2X1 NAND2X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__13_), .Y(_13881_) );
NAND2X1 NAND2X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_13880_), .B(_13881_), .Y(_13882_) );
NAND2X1 NAND2X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__13_), .Y(_13883_) );
NAND2X1 NAND2X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__13_), .Y(_13884_) );
NAND2X1 NAND2X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_13883_), .B(_13884_), .Y(_13885_) );
NOR2X1 NOR2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_13882_), .B(_13885_), .Y(_13886_) );
NAND3X1 NAND3X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_3296_), .B(_8762_), .C(_3295_), .Y(_13887_) );
NAND3X1 NAND3X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_3246_), .B(_8765_), .C(_3245_), .Y(_13888_) );
AND2X2 AND2X2_1607 ( .gnd(gnd), .vdd(vdd), .A(_13888_), .B(_13887_), .Y(_13889_) );
AOI22X1 AOI22X1_510 ( .gnd(gnd), .vdd(vdd), .A(_62__13_), .B(_8774_), .C(_57__13_), .D(_8771_), .Y(_13890_) );
NAND2X1 NAND2X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_13889_), .B(_13890_), .Y(_13891_) );
NAND2X1 NAND2X1_2590 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__13_), .Y(_13892_) );
NAND3X1 NAND3X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_2833_), .B(_8786_), .C(_2834_), .Y(_13893_) );
OAI21X1 OAI21X1_2552 ( .gnd(gnd), .vdd(vdd), .A(_2780_), .B(_8799_), .C(_13893_), .Y(_13894_) );
NAND3X1 NAND3X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_2662_), .B(_8794_), .C(_2663_), .Y(_13895_) );
OAI21X1 OAI21X1_2553 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .B(_8792_), .C(_13895_), .Y(_13896_) );
NOR2X1 NOR2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_13896_), .B(_13894_), .Y(_13897_) );
AOI22X1 AOI22X1_511 ( .gnd(gnd), .vdd(vdd), .A(_76__13_), .B(_9482_), .C(_75__13_), .D(_8802_), .Y(_13898_) );
NAND2X1 NAND2X1_2591 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__13_), .Y(_13899_) );
NAND2X1 NAND2X1_2592 ( .gnd(gnd), .vdd(vdd), .A(_9468_), .B(_81__13_), .Y(_13900_) );
NAND3X1 NAND3X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_13900_), .B(_13899_), .C(_13898_), .Y(_13901_) );
INVX1 INVX1_3882 ( .gnd(gnd), .vdd(vdd), .A(_84__13_), .Y(_13902_) );
NOR2X1 NOR2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_13902_), .Y(_13903_) );
NOR2X1 NOR2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2308_), .Y(_13904_) );
NAND2X1 NAND2X1_2593 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__13_), .Y(_13905_) );
NAND3X1 NAND3X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(_8843_), .C(_2023_), .Y(_13906_) );
NAND3X1 NAND3X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1931_), .C(_1932_), .Y(_13907_) );
NAND3X1 NAND3X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_13907_), .B(_13906_), .C(_13905_), .Y(_13908_) );
NOR3X1 NOR3X1_425 ( .gnd(gnd), .vdd(vdd), .A(_13903_), .B(_13908_), .C(_13904_), .Y(_13909_) );
NAND3X1 NAND3X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_8829_), .C(_2270_), .Y(_13910_) );
NAND3X1 NAND3X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_8831_), .C(_2164_), .Y(_13911_) );
NAND2X1 NAND2X1_2594 ( .gnd(gnd), .vdd(vdd), .A(_13910_), .B(_13911_), .Y(_13912_) );
NAND3X1 NAND3X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_2104_), .B(_8834_), .C(_2105_), .Y(_13913_) );
NAND3X1 NAND3X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .B(_8836_), .C(_2216_), .Y(_13914_) );
NAND2X1 NAND2X1_2595 ( .gnd(gnd), .vdd(vdd), .A(_13913_), .B(_13914_), .Y(_13915_) );
NOR2X1 NOR2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_13915_), .B(_13912_), .Y(_13916_) );
AOI22X1 AOI22X1_512 ( .gnd(gnd), .vdd(vdd), .A(_98__13_), .B(_8845_), .C(_93__13_), .D(_8840_), .Y(_13917_) );
AOI22X1 AOI22X1_513 ( .gnd(gnd), .vdd(vdd), .A(_94__13_), .B(_8841_), .C(_91__13_), .D(_8823_), .Y(_13918_) );
NAND2X1 NAND2X1_2596 ( .gnd(gnd), .vdd(vdd), .A(_13917_), .B(_13918_), .Y(_13919_) );
NAND2X1 NAND2X1_2597 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__13_), .Y(_13920_) );
NAND2X1 NAND2X1_2598 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__13_), .Y(_13921_) );
NAND2X1 NAND2X1_2599 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__13_), .Y(_13922_) );
NAND2X1 NAND2X1_2600 ( .gnd(gnd), .vdd(vdd), .A(_13921_), .B(_13922_), .Y(_13923_) );
NAND2X1 NAND2X1_2601 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__13_), .Y(_13924_) );
NAND2X1 NAND2X1_2602 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__13_), .Y(_13925_) );
NAND2X1 NAND2X1_2603 ( .gnd(gnd), .vdd(vdd), .A(_13924_), .B(_13925_), .Y(_13926_) );
NOR2X1 NOR2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_13923_), .B(_13926_), .Y(_13927_) );
NAND2X1 NAND2X1_2604 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__13_), .Y(_13928_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_7157_), .B(_9930_), .C(_7201_), .D(_9929_), .Y(_13929_) );
NOR2X1 NOR2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7336_), .Y(_13930_) );
NOR2X1 NOR2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7293_), .Y(_13931_) );
NOR3X1 NOR3X1_426 ( .gnd(gnd), .vdd(vdd), .A(_13930_), .B(_13931_), .C(_13929_), .Y(_13932_) );
NAND2X1 NAND2X1_2605 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__13_), .Y(_13933_) );
NAND2X1 NAND2X1_2606 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__13_), .Y(_13934_) );
NAND2X1 NAND2X1_2607 ( .gnd(gnd), .vdd(vdd), .A(_13933_), .B(_13934_), .Y(_13935_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_7379_), .B(_9940_), .C(_7247_), .D(_9941_), .Y(_13936_) );
NOR2X1 NOR2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_13936_), .B(_13935_), .Y(_13937_) );
NAND3X1 NAND3X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_13928_), .B(_13932_), .C(_13937_), .Y(_13938_) );
AOI22X1 AOI22X1_514 ( .gnd(gnd), .vdd(vdd), .A(_20__13_), .B(_8898_), .C(_250__13_), .D(_9082_), .Y(_13939_) );
AOI22X1 AOI22X1_515 ( .gnd(gnd), .vdd(vdd), .A(_243__13_), .B(_9153_), .C(_175__13_), .D(_8904_), .Y(_13940_) );
NAND2X1 NAND2X1_2608 ( .gnd(gnd), .vdd(vdd), .A(_13939_), .B(_13940_), .Y(_13941_) );
NAND2X1 NAND2X1_2609 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__13_), .Y(_13942_) );
NAND2X1 NAND2X1_2610 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__13_), .Y(_13943_) );
AOI22X1 AOI22X1_516 ( .gnd(gnd), .vdd(vdd), .A(_19__13_), .B(_8914_), .C(_210__13_), .D(_8918_), .Y(_13944_) );
NAND3X1 NAND3X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_13942_), .B(_13943_), .C(_13944_), .Y(_13945_) );
NOR2X1 NOR2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_13941_), .B(_13945_), .Y(_13946_) );
AOI22X1 AOI22X1_517 ( .gnd(gnd), .vdd(vdd), .A(_134__13_), .B(_8933_), .C(_9__13_), .D(_8926_), .Y(_13947_) );
NAND2X1 NAND2X1_2611 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__13_), .Y(_13948_) );
NAND2X1 NAND2X1_2612 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_145__13_), .Y(_13949_) );
NAND3X1 NAND3X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_13948_), .B(_13949_), .C(_13947_), .Y(_13950_) );
AOI22X1 AOI22X1_518 ( .gnd(gnd), .vdd(vdd), .A(_4__13_), .B(_8937_), .C(_176__13_), .D(_8939_), .Y(_13951_) );
NAND2X1 NAND2X1_2613 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__13_), .Y(_13952_) );
NAND2X1 NAND2X1_2614 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__13_), .Y(_13953_) );
NAND3X1 NAND3X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_13952_), .B(_13953_), .C(_13951_), .Y(_13954_) );
NOR2X1 NOR2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_13954_), .B(_13950_), .Y(_13955_) );
NAND2X1 NAND2X1_2615 ( .gnd(gnd), .vdd(vdd), .A(_13946_), .B(_13955_), .Y(_13956_) );
NAND2X1 NAND2X1_2616 ( .gnd(gnd), .vdd(vdd), .A(_8950_), .B(_208__13_), .Y(_13957_) );
NAND2X1 NAND2X1_2617 ( .gnd(gnd), .vdd(vdd), .A(_8952_), .B(_40__13_), .Y(_13958_) );
AOI22X1 AOI22X1_519 ( .gnd(gnd), .vdd(vdd), .A(_249__13_), .B(_9053_), .C(_209__13_), .D(_8957_), .Y(_13959_) );
NAND3X1 NAND3X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_13957_), .B(_13958_), .C(_13959_), .Y(_13960_) );
AOI22X1 AOI22X1_520 ( .gnd(gnd), .vdd(vdd), .A(_42__13_), .B(_8963_), .C(_177__13_), .D(_8961_), .Y(_13961_) );
NAND2X1 NAND2X1_2618 ( .gnd(gnd), .vdd(vdd), .A(_9160_), .B(_244__13_), .Y(_13962_) );
NAND2X1 NAND2X1_2619 ( .gnd(gnd), .vdd(vdd), .A(_8968_), .B(_44__13_), .Y(_13963_) );
NAND3X1 NAND3X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_13962_), .B(_13963_), .C(_13961_), .Y(_13964_) );
NOR2X1 NOR2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_13960_), .B(_13964_), .Y(_13965_) );
NAND2X1 NAND2X1_2620 ( .gnd(gnd), .vdd(vdd), .A(_8986_), .B(_255__13_), .Y(_13966_) );
NAND2X1 NAND2X1_2621 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__13_), .Y(_13967_) );
AOI22X1 AOI22X1_521 ( .gnd(gnd), .vdd(vdd), .A(_37__13_), .B(_8978_), .C(_35__13_), .D(_8980_), .Y(_13968_) );
NAND3X1 NAND3X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_13966_), .B(_13967_), .C(_13968_), .Y(_13969_) );
NAND2X1 NAND2X1_2622 ( .gnd(gnd), .vdd(vdd), .A(_8984_), .B(_254__13_), .Y(_13970_) );
NAND2X1 NAND2X1_2623 ( .gnd(gnd), .vdd(vdd), .A(_8991_), .B(_33__13_), .Y(_13971_) );
AOI22X1 AOI22X1_522 ( .gnd(gnd), .vdd(vdd), .A(_203__13_), .B(_9018_), .C(_156__13_), .D(_8973_), .Y(_13972_) );
NAND3X1 NAND3X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_13970_), .B(_13971_), .C(_13972_), .Y(_13973_) );
NOR2X1 NOR2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_13973_), .B(_13969_), .Y(_13974_) );
NAND2X1 NAND2X1_2624 ( .gnd(gnd), .vdd(vdd), .A(_13965_), .B(_13974_), .Y(_13975_) );
NOR2X1 NOR2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_13956_), .B(_13975_), .Y(_13976_) );
NAND2X1 NAND2X1_2625 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__13_), .Y(_13977_) );
NAND2X1 NAND2X1_2626 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__13_), .Y(_13978_) );
AOI22X1 AOI22X1_523 ( .gnd(gnd), .vdd(vdd), .A(_13__13_), .B(_9007_), .C(_239__13_), .D(_9076_), .Y(_13979_) );
NAND3X1 NAND3X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_13977_), .B(_13978_), .C(_13979_), .Y(_13980_) );
AOI22X1 AOI22X1_524 ( .gnd(gnd), .vdd(vdd), .A(_206__13_), .B(_9013_), .C(_242__13_), .D(_9035_), .Y(_13981_) );
NAND2X1 NAND2X1_2627 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__13_), .Y(_13982_) );
NAND2X1 NAND2X1_2628 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__13_), .Y(_13983_) );
NAND3X1 NAND3X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_13982_), .B(_13983_), .C(_13981_), .Y(_13984_) );
NOR2X1 NOR2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_13980_), .B(_13984_), .Y(_13985_) );
AOI22X1 AOI22X1_525 ( .gnd(gnd), .vdd(vdd), .A(_222__13_), .B(_9024_), .C(_220__13_), .D(_9026_), .Y(_13986_) );
NAND2X1 NAND2X1_2629 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__13_), .Y(_13987_) );
NAND2X1 NAND2X1_2630 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__13_), .Y(_13988_) );
NAND3X1 NAND3X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_13987_), .B(_13988_), .C(_13986_), .Y(_13989_) );
AOI22X1 AOI22X1_526 ( .gnd(gnd), .vdd(vdd), .A(_18__13_), .B(_9037_), .C(_240__13_), .D(_9011_), .Y(_13990_) );
NAND2X1 NAND2X1_2631 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__13_), .Y(_13991_) );
NAND2X1 NAND2X1_2632 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__13_), .Y(_13992_) );
NAND3X1 NAND3X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_13991_), .B(_13992_), .C(_13990_), .Y(_13993_) );
NOR2X1 NOR2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_13989_), .B(_13993_), .Y(_13994_) );
NAND2X1 NAND2X1_2633 ( .gnd(gnd), .vdd(vdd), .A(_13985_), .B(_13994_), .Y(_13995_) );
AOI22X1 AOI22X1_527 ( .gnd(gnd), .vdd(vdd), .A(_225__13_), .B(_9048_), .C(_167__13_), .D(_9050_), .Y(_13996_) );
NAND2X1 NAND2X1_2634 ( .gnd(gnd), .vdd(vdd), .A(_8955_), .B(_236__13_), .Y(_13997_) );
NAND2X1 NAND2X1_2635 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__13_), .Y(_13998_) );
NAND3X1 NAND3X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_13997_), .B(_13998_), .C(_13996_), .Y(_13999_) );
NAND2X1 NAND2X1_2636 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__13_), .Y(_14000_) );
NAND2X1 NAND2X1_2637 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__13_), .Y(_14001_) );
AOI22X1 AOI22X1_528 ( .gnd(gnd), .vdd(vdd), .A(_224__13_), .B(_9064_), .C(_27__13_), .D(_9066_), .Y(_14002_) );
NAND3X1 NAND3X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_14000_), .B(_14001_), .C(_14002_), .Y(_14003_) );
NOR2X1 NOR2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_13999_), .B(_14003_), .Y(_14004_) );
AOI22X1 AOI22X1_529 ( .gnd(gnd), .vdd(vdd), .A(_184__13_), .B(_9073_), .C(_183__13_), .D(_9071_), .Y(_14005_) );
NAND2X1 NAND2X1_2638 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__13_), .Y(_14006_) );
NAND2X1 NAND2X1_2639 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__13_), .Y(_14007_) );
NAND3X1 NAND3X1_2895 ( .gnd(gnd), .vdd(vdd), .A(_14006_), .B(_14007_), .C(_14005_), .Y(_14008_) );
AOI22X1 AOI22X1_530 ( .gnd(gnd), .vdd(vdd), .A(_43__13_), .B(_9084_), .C(_248__13_), .D(_8901_), .Y(_14009_) );
NAND2X1 NAND2X1_2640 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__13_), .Y(_14010_) );
NAND2X1 NAND2X1_2641 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__13_), .Y(_14011_) );
NAND3X1 NAND3X1_2896 ( .gnd(gnd), .vdd(vdd), .A(_14010_), .B(_14011_), .C(_14009_), .Y(_14012_) );
NOR2X1 NOR2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(_14008_), .B(_14012_), .Y(_14013_) );
NAND2X1 NAND2X1_2642 ( .gnd(gnd), .vdd(vdd), .A(_14004_), .B(_14013_), .Y(_14014_) );
NOR2X1 NOR2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_13995_), .B(_14014_), .Y(_14015_) );
NAND3X1 NAND3X1_2897 ( .gnd(gnd), .vdd(vdd), .A(_6869_), .B(_9104_), .C(_6870_), .Y(_14016_) );
NAND3X1 NAND3X1_2898 ( .gnd(gnd), .vdd(vdd), .A(_3977_), .B(_9099_), .C(_3978_), .Y(_14017_) );
NAND2X1 NAND2X1_2643 ( .gnd(gnd), .vdd(vdd), .A(_14016_), .B(_14017_), .Y(_14018_) );
NAND2X1 NAND2X1_2644 ( .gnd(gnd), .vdd(vdd), .A(_9097_), .B(_10__13_), .Y(_14019_) );
NAND3X1 NAND3X1_2899 ( .gnd(gnd), .vdd(vdd), .A(_5112_), .B(_9102_), .C(_5113_), .Y(_14020_) );
NAND2X1 NAND2X1_2645 ( .gnd(gnd), .vdd(vdd), .A(_14020_), .B(_14019_), .Y(_14021_) );
NOR2X1 NOR2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_14018_), .B(_14021_), .Y(_14022_) );
NAND3X1 NAND3X1_2900 ( .gnd(gnd), .vdd(vdd), .A(_8330_), .B(_9188_), .C(_8331_), .Y(_14023_) );
NAND3X1 NAND3X1_2901 ( .gnd(gnd), .vdd(vdd), .A(_15941_), .B(_9109_), .C(_15942_), .Y(_14024_) );
NAND3X1 NAND3X1_2902 ( .gnd(gnd), .vdd(vdd), .A(_16146_), .B(_9115_), .C(_16147_), .Y(_14025_) );
NAND3X1 NAND3X1_2903 ( .gnd(gnd), .vdd(vdd), .A(_14024_), .B(_14025_), .C(_14023_), .Y(_14026_) );
AOI22X1 AOI22X1_531 ( .gnd(gnd), .vdd(vdd), .A(_234__13_), .B(_9182_), .C(_34__13_), .D(_9183_), .Y(_14027_) );
AOI22X1 AOI22X1_532 ( .gnd(gnd), .vdd(vdd), .A(_100__13_), .B(_9346_), .C(_45__13_), .D(_9185_), .Y(_14028_) );
NAND2X1 NAND2X1_2646 ( .gnd(gnd), .vdd(vdd), .A(_14028_), .B(_14027_), .Y(_14029_) );
NAND3X1 NAND3X1_2904 ( .gnd(gnd), .vdd(vdd), .A(_4757_), .B(_9127_), .C(_4756_), .Y(_14030_) );
NAND3X1 NAND3X1_2905 ( .gnd(gnd), .vdd(vdd), .A(_4021_), .B(_9129_), .C(_4022_), .Y(_14031_) );
NAND2X1 NAND2X1_2647 ( .gnd(gnd), .vdd(vdd), .A(_14030_), .B(_14031_), .Y(_14032_) );
NOR3X1 NOR3X1_427 ( .gnd(gnd), .vdd(vdd), .A(_14026_), .B(_14032_), .C(_14029_), .Y(_14033_) );
NAND3X1 NAND3X1_2906 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_9133_), .C(_3441_), .Y(_14034_) );
NAND3X1 NAND3X1_2907 ( .gnd(gnd), .vdd(vdd), .A(_5066_), .B(_9135_), .C(_5067_), .Y(_14035_) );
NAND3X1 NAND3X1_2908 ( .gnd(gnd), .vdd(vdd), .A(_6948_), .B(_9137_), .C(_6949_), .Y(_14036_) );
NAND3X1 NAND3X1_2909 ( .gnd(gnd), .vdd(vdd), .A(_14035_), .B(_14036_), .C(_14034_), .Y(_14037_) );
AOI22X1 AOI22X1_533 ( .gnd(gnd), .vdd(vdd), .A(_17__13_), .B(_9140_), .C(_2__13_), .D(_9141_), .Y(_14038_) );
AOI22X1 AOI22X1_534 ( .gnd(gnd), .vdd(vdd), .A(_205__13_), .B(_9143_), .C(_200__13_), .D(_9145_), .Y(_14039_) );
NAND2X1 NAND2X1_2648 ( .gnd(gnd), .vdd(vdd), .A(_14038_), .B(_14039_), .Y(_14040_) );
NOR2X1 NOR2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_14037_), .B(_14040_), .Y(_14041_) );
NAND3X1 NAND3X1_2910 ( .gnd(gnd), .vdd(vdd), .A(_14022_), .B(_14033_), .C(_14041_), .Y(_14042_) );
AOI22X1 AOI22X1_535 ( .gnd(gnd), .vdd(vdd), .A(_21__13_), .B(_9150_), .C(_185__13_), .D(_9151_), .Y(_14043_) );
AOI22X1 AOI22X1_536 ( .gnd(gnd), .vdd(vdd), .A(_237__13_), .B(_8966_), .C(_253__13_), .D(_9154_), .Y(_14044_) );
NAND2X1 NAND2X1_2649 ( .gnd(gnd), .vdd(vdd), .A(_14043_), .B(_14044_), .Y(_14045_) );
AOI22X1 AOI22X1_537 ( .gnd(gnd), .vdd(vdd), .A(_46__13_), .B(_9158_), .C(_231__13_), .D(_9157_), .Y(_14046_) );
AOI22X1 AOI22X1_538 ( .gnd(gnd), .vdd(vdd), .A(_47__13_), .B(_9161_), .C(_238__13_), .D(_8893_), .Y(_14047_) );
NAND2X1 NAND2X1_2650 ( .gnd(gnd), .vdd(vdd), .A(_14047_), .B(_14046_), .Y(_14048_) );
NOR2X1 NOR2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_14045_), .B(_14048_), .Y(_14049_) );
AOI22X1 AOI22X1_539 ( .gnd(gnd), .vdd(vdd), .A(_247__13_), .B(_9165_), .C(_30__13_), .D(_9167_), .Y(_14050_) );
AOI22X1 AOI22X1_540 ( .gnd(gnd), .vdd(vdd), .A(_227__13_), .B(_9170_), .C(_218__13_), .D(_9169_), .Y(_14051_) );
NAND2X1 NAND2X1_2651 ( .gnd(gnd), .vdd(vdd), .A(_14050_), .B(_14051_), .Y(_14052_) );
AOI22X1 AOI22X1_541 ( .gnd(gnd), .vdd(vdd), .A(_123__13_), .B(_8928_), .C(_213__13_), .D(_8989_), .Y(_14053_) );
AOI22X1 AOI22X1_542 ( .gnd(gnd), .vdd(vdd), .A(_29__13_), .B(_9176_), .C(_178__13_), .D(_9173_), .Y(_14054_) );
NAND2X1 NAND2X1_2652 ( .gnd(gnd), .vdd(vdd), .A(_14053_), .B(_14054_), .Y(_14055_) );
NOR2X1 NOR2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_14052_), .B(_14055_), .Y(_14056_) );
NAND2X1 NAND2X1_2653 ( .gnd(gnd), .vdd(vdd), .A(_14049_), .B(_14056_), .Y(_14057_) );
AOI22X1 AOI22X1_543 ( .gnd(gnd), .vdd(vdd), .A(_201__13_), .B(_9124_), .C(_212__13_), .D(_9345_), .Y(_14058_) );
NAND3X1 NAND3X1_2911 ( .gnd(gnd), .vdd(vdd), .A(_8444_), .B(_9348_), .C(_8443_), .Y(_14059_) );
NAND3X1 NAND3X1_2912 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_504_), .C(_505_), .Y(_14060_) );
AND2X2 AND2X2_1608 ( .gnd(gnd), .vdd(vdd), .A(_14060_), .B(_14059_), .Y(_14061_) );
NAND2X1 NAND2X1_2654 ( .gnd(gnd), .vdd(vdd), .A(_14058_), .B(_14061_), .Y(_14062_) );
NAND3X1 NAND3X1_2913 ( .gnd(gnd), .vdd(vdd), .A(_15150_), .B(_9208_), .C(_15151_), .Y(_14063_) );
OAI21X1 OAI21X1_2554 ( .gnd(gnd), .vdd(vdd), .A(_15114_), .B(_9211_), .C(_14063_), .Y(_14064_) );
NAND3X1 NAND3X1_2914 ( .gnd(gnd), .vdd(vdd), .A(_15498_), .B(_9222_), .C(_15499_), .Y(_14065_) );
NAND3X1 NAND3X1_2915 ( .gnd(gnd), .vdd(vdd), .A(_15445_), .B(_9224_), .C(_15444_), .Y(_14066_) );
NAND2X1 NAND2X1_2655 ( .gnd(gnd), .vdd(vdd), .A(_14065_), .B(_14066_), .Y(_14067_) );
NOR2X1 NOR2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_14067_), .B(_14064_), .Y(_14068_) );
NAND3X1 NAND3X1_2916 ( .gnd(gnd), .vdd(vdd), .A(_15276_), .B(_9217_), .C(_15277_), .Y(_14069_) );
NAND3X1 NAND3X1_2917 ( .gnd(gnd), .vdd(vdd), .A(_15224_), .B(_9219_), .C(_15223_), .Y(_14070_) );
NAND2X1 NAND2X1_2656 ( .gnd(gnd), .vdd(vdd), .A(_14070_), .B(_14069_), .Y(_14071_) );
NAND3X1 NAND3X1_2918 ( .gnd(gnd), .vdd(vdd), .A(_15674_), .B(_9192_), .C(_15675_), .Y(_14072_) );
NAND3X1 NAND3X1_2919 ( .gnd(gnd), .vdd(vdd), .A(_15731_), .B(_9199_), .C(_15730_), .Y(_14073_) );
NAND2X1 NAND2X1_2657 ( .gnd(gnd), .vdd(vdd), .A(_14073_), .B(_14072_), .Y(_14074_) );
NOR2X1 NOR2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_14074_), .B(_14071_), .Y(_14075_) );
NOR3X1 NOR3X1_428 ( .gnd(gnd), .vdd(vdd), .A(_16198_), .B(_10083_), .C(_16199_), .Y(_14076_) );
NAND3X1 NAND3X1_2920 ( .gnd(gnd), .vdd(vdd), .A(_15324_), .B(_9205_), .C(_15325_), .Y(_14077_) );
OAI21X1 OAI21X1_2555 ( .gnd(gnd), .vdd(vdd), .A(_15354_), .B(_10085_), .C(_14077_), .Y(_14078_) );
NAND3X1 NAND3X1_2921 ( .gnd(gnd), .vdd(vdd), .A(_15556_), .B(_9233_), .C(_15557_), .Y(_14079_) );
NAND3X1 NAND3X1_2922 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15622_), .C(_15621_), .Y(_14080_) );
NAND2X1 NAND2X1_2658 ( .gnd(gnd), .vdd(vdd), .A(_14079_), .B(_14080_), .Y(_14081_) );
NOR3X1 NOR3X1_429 ( .gnd(gnd), .vdd(vdd), .A(_14078_), .B(_14081_), .C(_14076_), .Y(_14082_) );
NAND3X1 NAND3X1_2923 ( .gnd(gnd), .vdd(vdd), .A(_14068_), .B(_14075_), .C(_14082_), .Y(_14083_) );
NAND3X1 NAND3X1_2924 ( .gnd(gnd), .vdd(vdd), .A(_15884_), .B(_9120_), .C(_15885_), .Y(_14084_) );
NAND3X1 NAND3X1_2925 ( .gnd(gnd), .vdd(vdd), .A(_15391_), .B(_9197_), .C(_15392_), .Y(_14085_) );
NOR3X1 NOR3X1_430 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_8180_), .C(_8179_), .Y(_14086_) );
AND2X2 AND2X2_1609 ( .gnd(gnd), .vdd(vdd), .A(_186__13_), .B(_9298_), .Y(_14087_) );
NOR3X1 NOR3X1_431 ( .gnd(gnd), .vdd(vdd), .A(_15823_), .B(_11264_), .C(_15822_), .Y(_14088_) );
NOR3X1 NOR3X1_432 ( .gnd(gnd), .vdd(vdd), .A(_14086_), .B(_14087_), .C(_14088_), .Y(_14089_) );
NOR3X1 NOR3X1_433 ( .gnd(gnd), .vdd(vdd), .A(_7478_), .B(_10471_), .C(_7479_), .Y(_14090_) );
NOR2X1 NOR2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_9263_), .B(_624_), .Y(_14091_) );
NAND3X1 NAND3X1_2926 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_9268_), .C(_1184_), .Y(_14092_) );
OAI21X1 OAI21X1_2556 ( .gnd(gnd), .vdd(vdd), .A(_2927_), .B(_10468_), .C(_14092_), .Y(_14093_) );
NOR3X1 NOR3X1_434 ( .gnd(gnd), .vdd(vdd), .A(_14091_), .B(_14093_), .C(_14090_), .Y(_14094_) );
NAND3X1 NAND3X1_2927 ( .gnd(gnd), .vdd(vdd), .A(_14923_), .B(_9275_), .C(_14925_), .Y(_14095_) );
OAI21X1 OAI21X1_2557 ( .gnd(gnd), .vdd(vdd), .A(_7649_), .B(_9301_), .C(_14095_), .Y(_14096_) );
NAND3X1 NAND3X1_2928 ( .gnd(gnd), .vdd(vdd), .A(_8211_), .B(_9286_), .C(_8212_), .Y(_14097_) );
OAI21X1 OAI21X1_2558 ( .gnd(gnd), .vdd(vdd), .A(_7108_), .B(_9245_), .C(_14097_), .Y(_14098_) );
NOR2X1 NOR2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_14096_), .B(_14098_), .Y(_14099_) );
NAND3X1 NAND3X1_2929 ( .gnd(gnd), .vdd(vdd), .A(_14099_), .B(_14089_), .C(_14094_), .Y(_14100_) );
NOR3X1 NOR3X1_435 ( .gnd(gnd), .vdd(vdd), .A(_5935_), .B(_9323_), .C(_5936_), .Y(_14101_) );
NAND3X1 NAND3X1_2930 ( .gnd(gnd), .vdd(vdd), .A(_7734_), .B(_9248_), .C(_7733_), .Y(_14102_) );
OAI21X1 OAI21X1_2559 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(_12340_), .C(_14102_), .Y(_14103_) );
NAND3X1 NAND3X1_2931 ( .gnd(gnd), .vdd(vdd), .A(_2370_), .B(_9315_), .C(_2369_), .Y(_14104_) );
OAI21X1 OAI21X1_2560 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_9282_), .C(_14104_), .Y(_14105_) );
NOR3X1 NOR3X1_436 ( .gnd(gnd), .vdd(vdd), .A(_14103_), .B(_14105_), .C(_14101_), .Y(_14106_) );
NAND3X1 NAND3X1_2932 ( .gnd(gnd), .vdd(vdd), .A(_7062_), .B(_9266_), .C(_7063_), .Y(_14107_) );
OAI21X1 OAI21X1_2561 ( .gnd(gnd), .vdd(vdd), .A(_4198_), .B(_9254_), .C(_14107_), .Y(_14108_) );
NAND2X1 NAND2X1_2659 ( .gnd(gnd), .vdd(vdd), .A(_9289_), .B(_199__13_), .Y(_14109_) );
OAI21X1 OAI21X1_2562 ( .gnd(gnd), .vdd(vdd), .A(_8250_), .B(_10875_), .C(_14109_), .Y(_14110_) );
NOR2X1 NOR2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_14110_), .B(_14108_), .Y(_14111_) );
NAND2X1 NAND2X1_2660 ( .gnd(gnd), .vdd(vdd), .A(_1__13_), .B(_9242_), .Y(_14112_) );
OAI21X1 OAI21X1_2563 ( .gnd(gnd), .vdd(vdd), .A(_6477_), .B(_9259_), .C(_14112_), .Y(_14113_) );
NAND3X1 NAND3X1_2933 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_9294_), .C(_3618_), .Y(_14114_) );
OAI21X1 OAI21X1_2564 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_9306_), .C(_14114_), .Y(_14115_) );
NOR2X1 NOR2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_14115_), .B(_14113_), .Y(_14116_) );
NAND3X1 NAND3X1_2934 ( .gnd(gnd), .vdd(vdd), .A(_14106_), .B(_14111_), .C(_14116_), .Y(_14117_) );
NOR2X1 NOR2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_10121_), .B(_7689_), .Y(_14118_) );
NOR3X1 NOR3X1_437 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_9312_), .C(_4791_), .Y(_14119_) );
NOR2X1 NOR2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .B(_4831_), .Y(_14120_) );
NOR3X1 NOR3X1_438 ( .gnd(gnd), .vdd(vdd), .A(_14118_), .B(_14120_), .C(_14119_), .Y(_14121_) );
AOI22X1 AOI22X1_544 ( .gnd(gnd), .vdd(vdd), .A(_217__13_), .B(_9281_), .C(_251__13_), .D(_9320_), .Y(_14122_) );
AOI22X1 AOI22X1_545 ( .gnd(gnd), .vdd(vdd), .A(_252__13_), .B(_9326_), .C(_233__13_), .D(_9310_), .Y(_14123_) );
NAND3X1 NAND3X1_2935 ( .gnd(gnd), .vdd(vdd), .A(_14121_), .B(_14122_), .C(_14123_), .Y(_14124_) );
NOR3X1 NOR3X1_439 ( .gnd(gnd), .vdd(vdd), .A(_14100_), .B(_14124_), .C(_14117_), .Y(_14125_) );
NAND2X1 NAND2X1_2661 ( .gnd(gnd), .vdd(vdd), .A(_14085_), .B(_14125_), .Y(_14126_) );
AOI21X1 AOI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_157__13_), .B(_9232_), .C(_14126_), .Y(_14127_) );
AOI22X1 AOI22X1_546 ( .gnd(gnd), .vdd(vdd), .A(_155__13_), .B(_9333_), .C(_172__13_), .D(_9332_), .Y(_14128_) );
NAND3X1 NAND3X1_2936 ( .gnd(gnd), .vdd(vdd), .A(_14084_), .B(_14128_), .C(_14127_), .Y(_14129_) );
NOR3X1 NOR3X1_440 ( .gnd(gnd), .vdd(vdd), .A(_14083_), .B(_14129_), .C(_14062_), .Y(_14130_) );
AOI22X1 AOI22X1_547 ( .gnd(gnd), .vdd(vdd), .A(_256__13_), .B(_9113_), .C(_142__13_), .D(_9118_), .Y(_14131_) );
NAND2X1 NAND2X1_2662 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__13_), .Y(_14132_) );
NAND2X1 NAND2X1_2663 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__13_), .Y(_14133_) );
NAND3X1 NAND3X1_2937 ( .gnd(gnd), .vdd(vdd), .A(_14132_), .B(_14133_), .C(_14131_), .Y(_14134_) );
NAND2X1 NAND2X1_2664 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__13_), .Y(_14135_) );
NAND3X1 NAND3X1_2938 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_9339_), .C(_467_), .Y(_14136_) );
AOI22X1 AOI22X1_548 ( .gnd(gnd), .vdd(vdd), .A(_111__13_), .B(_9342_), .C(_12__13_), .D(_9341_), .Y(_14137_) );
NAND3X1 NAND3X1_2939 ( .gnd(gnd), .vdd(vdd), .A(_14137_), .B(_14135_), .C(_14136_), .Y(_14138_) );
NOR2X1 NOR2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_14134_), .B(_14138_), .Y(_14139_) );
AOI22X1 AOI22X1_549 ( .gnd(gnd), .vdd(vdd), .A(_232__13_), .B(_9354_), .C(_219__13_), .D(_9353_), .Y(_14140_) );
AOI22X1 AOI22X1_550 ( .gnd(gnd), .vdd(vdd), .A(_246__13_), .B(_9356_), .C(_226__13_), .D(_9357_), .Y(_14141_) );
NAND2X1 NAND2X1_2665 ( .gnd(gnd), .vdd(vdd), .A(_14140_), .B(_14141_), .Y(_14142_) );
NAND3X1 NAND3X1_2940 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16101_), .C(_16102_), .Y(_14143_) );
NAND3X1 NAND3X1_2941 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16046_), .C(_16047_), .Y(_14144_) );
NAND2X1 NAND2X1_2666 ( .gnd(gnd), .vdd(vdd), .A(_14143_), .B(_14144_), .Y(_14145_) );
NAND3X1 NAND3X1_2942 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8580_), .C(_8579_), .Y(_14146_) );
OAI21X1 OAI21X1_2565 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_9361_), .C(_14146_), .Y(_14147_) );
NOR2X1 NOR2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_14145_), .B(_14147_), .Y(_14148_) );
NAND2X1 NAND2X1_2667 ( .gnd(gnd), .vdd(vdd), .A(_15990_), .B(_15991_), .Y(_14149_) );
NAND3X1 NAND3X1_2943 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8633_), .C(_8634_), .Y(_14150_) );
OAI21X1 OAI21X1_2566 ( .gnd(gnd), .vdd(vdd), .A(_14149_), .B(_9215_), .C(_14150_), .Y(_14151_) );
NAND3X1 NAND3X1_2944 ( .gnd(gnd), .vdd(vdd), .A(_8688_), .B(_9371_), .C(_8687_), .Y(_14152_) );
NAND3X1 NAND3X1_2945 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_330_), .C(_331_), .Y(_14153_) );
NAND2X1 NAND2X1_2668 ( .gnd(gnd), .vdd(vdd), .A(_14153_), .B(_14152_), .Y(_14154_) );
NOR2X1 NOR2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_14151_), .B(_14154_), .Y(_14155_) );
AOI22X1 AOI22X1_551 ( .gnd(gnd), .vdd(vdd), .A(_22__13_), .B(_9382_), .C(_3__13_), .D(_9383_), .Y(_14156_) );
NAND3X1 NAND3X1_2946 ( .gnd(gnd), .vdd(vdd), .A(_14148_), .B(_14155_), .C(_14156_), .Y(_14157_) );
NOR2X1 NOR2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_14142_), .B(_14157_), .Y(_14158_) );
NAND3X1 NAND3X1_2947 ( .gnd(gnd), .vdd(vdd), .A(_14130_), .B(_14139_), .C(_14158_), .Y(_14159_) );
NOR3X1 NOR3X1_441 ( .gnd(gnd), .vdd(vdd), .A(_14042_), .B(_14057_), .C(_14159_), .Y(_14160_) );
NAND3X1 NAND3X1_2948 ( .gnd(gnd), .vdd(vdd), .A(_13976_), .B(_14015_), .C(_14160_), .Y(_14161_) );
NAND3X1 NAND3X1_2949 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1597_), .C(_1598_), .Y(_14162_) );
NAND3X1 NAND3X1_2950 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .B(_8862_), .C(_1259_), .Y(_14163_) );
NAND2X1 NAND2X1_2669 ( .gnd(gnd), .vdd(vdd), .A(_14162_), .B(_14163_), .Y(_14164_) );
NOR3X1 NOR3X1_442 ( .gnd(gnd), .vdd(vdd), .A(_13938_), .B(_14164_), .C(_14161_), .Y(_14165_) );
NAND3X1 NAND3X1_2951 ( .gnd(gnd), .vdd(vdd), .A(_13920_), .B(_13927_), .C(_14165_), .Y(_14166_) );
NAND2X1 NAND2X1_2670 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__13_), .Y(_14167_) );
NAND3X1 NAND3X1_2952 ( .gnd(gnd), .vdd(vdd), .A(_1475_), .B(_9406_), .C(_1476_), .Y(_14168_) );
NAND3X1 NAND3X1_2953 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_9453_), .C(_1428_), .Y(_14169_) );
AND2X2 AND2X2_1610 ( .gnd(gnd), .vdd(vdd), .A(_14168_), .B(_14169_), .Y(_14170_) );
NAND2X1 NAND2X1_2671 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_108__13_), .Y(_14171_) );
NAND2X1 NAND2X1_2672 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_116__13_), .Y(_14172_) );
NAND3X1 NAND3X1_2954 ( .gnd(gnd), .vdd(vdd), .A(_14171_), .B(_14172_), .C(_14170_), .Y(_14173_) );
AOI22X1 AOI22X1_552 ( .gnd(gnd), .vdd(vdd), .A(_125__13_), .B(_9411_), .C(_124__13_), .D(_9410_), .Y(_14174_) );
AOI22X1 AOI22X1_553 ( .gnd(gnd), .vdd(vdd), .A(_120__13_), .B(_9415_), .C(_121__13_), .D(_9413_), .Y(_14175_) );
AND2X2 AND2X2_1611 ( .gnd(gnd), .vdd(vdd), .A(_14175_), .B(_14174_), .Y(_14176_) );
AOI22X1 AOI22X1_554 ( .gnd(gnd), .vdd(vdd), .A(_132__13_), .B(_9420_), .C(_131__13_), .D(_9418_), .Y(_14177_) );
NAND2X1 NAND2X1_2673 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__13_), .Y(_14178_) );
NAND2X1 NAND2X1_2674 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__13_), .Y(_14179_) );
NAND3X1 NAND3X1_2955 ( .gnd(gnd), .vdd(vdd), .A(_14178_), .B(_14179_), .C(_14177_), .Y(_14180_) );
NAND3X1 NAND3X1_2956 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_9431_), .C(_562_), .Y(_14181_) );
NAND2X1 NAND2X1_2675 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__13_), .Y(_14182_) );
NAND2X1 NAND2X1_2676 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__13_), .Y(_14183_) );
NAND3X1 NAND3X1_2957 ( .gnd(gnd), .vdd(vdd), .A(_14183_), .B(_14181_), .C(_14182_), .Y(_14184_) );
AOI21X1 AOI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_136__13_), .B(_9429_), .C(_14184_), .Y(_14185_) );
NAND2X1 NAND2X1_2677 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__13_), .Y(_14186_) );
NAND2X1 NAND2X1_2678 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__13_), .Y(_14187_) );
NAND3X1 NAND3X1_2958 ( .gnd(gnd), .vdd(vdd), .A(_14186_), .B(_14187_), .C(_14185_), .Y(_14188_) );
NAND3X1 NAND3X1_2959 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_9444_), .C(_1067_), .Y(_14189_) );
NAND2X1 NAND2X1_2679 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__13_), .Y(_14190_) );
AOI22X1 AOI22X1_555 ( .gnd(gnd), .vdd(vdd), .A(_130__13_), .B(_9449_), .C(_127__13_), .D(_9448_), .Y(_14191_) );
NAND3X1 NAND3X1_2960 ( .gnd(gnd), .vdd(vdd), .A(_14189_), .B(_14191_), .C(_14190_), .Y(_14192_) );
NOR3X1 NOR3X1_443 ( .gnd(gnd), .vdd(vdd), .A(_14180_), .B(_14188_), .C(_14192_), .Y(_14193_) );
AOI22X1 AOI22X1_556 ( .gnd(gnd), .vdd(vdd), .A(_115__13_), .B(_9399_), .C(_114__13_), .D(_9454_), .Y(_14194_) );
NAND3X1 NAND3X1_2961 ( .gnd(gnd), .vdd(vdd), .A(_14194_), .B(_14176_), .C(_14193_), .Y(_14195_) );
NOR2X1 NOR2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_14173_), .B(_14195_), .Y(_14196_) );
AOI22X1 AOI22X1_557 ( .gnd(gnd), .vdd(vdd), .A(_102__13_), .B(_9459_), .C(_103__13_), .D(_9457_), .Y(_14197_) );
NAND3X1 NAND3X1_2962 ( .gnd(gnd), .vdd(vdd), .A(_14167_), .B(_14197_), .C(_14196_), .Y(_14198_) );
NOR3X1 NOR3X1_444 ( .gnd(gnd), .vdd(vdd), .A(_13919_), .B(_14198_), .C(_14166_), .Y(_14199_) );
NAND3X1 NAND3X1_2963 ( .gnd(gnd), .vdd(vdd), .A(_13909_), .B(_13916_), .C(_14199_), .Y(_14200_) );
NAND2X1 NAND2X1_2680 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__13_), .Y(_14201_) );
NAND2X1 NAND2X1_2681 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__13_), .Y(_14202_) );
NAND2X1 NAND2X1_2682 ( .gnd(gnd), .vdd(vdd), .A(_14201_), .B(_14202_), .Y(_14203_) );
NOR3X1 NOR3X1_445 ( .gnd(gnd), .vdd(vdd), .A(_13901_), .B(_14203_), .C(_14200_), .Y(_14204_) );
NAND3X1 NAND3X1_2964 ( .gnd(gnd), .vdd(vdd), .A(_13892_), .B(_13897_), .C(_14204_), .Y(_14205_) );
NAND3X1 NAND3X1_2965 ( .gnd(gnd), .vdd(vdd), .A(_3079_), .B(_9473_), .C(_3080_), .Y(_14206_) );
NAND2X1 NAND2X1_2683 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__13_), .Y(_14207_) );
NAND3X1 NAND3X1_2966 ( .gnd(gnd), .vdd(vdd), .A(_2594_), .B(_8803_), .C(_2593_), .Y(_14208_) );
NAND2X1 NAND2X1_2684 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__13_), .Y(_14209_) );
NAND3X1 NAND3X1_2967 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .B(_8806_), .C(_2411_), .Y(_14210_) );
NAND3X1 NAND3X1_2968 ( .gnd(gnd), .vdd(vdd), .A(_14208_), .B(_14210_), .C(_14209_), .Y(_14211_) );
AOI21X1 AOI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_68__13_), .B(_9477_), .C(_14211_), .Y(_14212_) );
NAND3X1 NAND3X1_2969 ( .gnd(gnd), .vdd(vdd), .A(_14206_), .B(_14212_), .C(_14207_), .Y(_14213_) );
NOR3X1 NOR3X1_446 ( .gnd(gnd), .vdd(vdd), .A(_13891_), .B(_14213_), .C(_14205_), .Y(_14214_) );
AOI21X1 AOI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_13886_), .B(_14214_), .C(rst), .Y(_0__13_) );
NAND2X1 NAND2X1_2685 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__14_), .Y(_14215_) );
NAND2X1 NAND2X1_2686 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__14_), .Y(_14216_) );
NAND2X1 NAND2X1_2687 ( .gnd(gnd), .vdd(vdd), .A(_14215_), .B(_14216_), .Y(_14217_) );
NAND2X1 NAND2X1_2688 ( .gnd(gnd), .vdd(vdd), .A(_8765_), .B(_55__14_), .Y(_14218_) );
NAND2X1 NAND2X1_2689 ( .gnd(gnd), .vdd(vdd), .A(_8771_), .B(_57__14_), .Y(_14219_) );
NAND2X1 NAND2X1_2690 ( .gnd(gnd), .vdd(vdd), .A(_14219_), .B(_14218_), .Y(_14220_) );
NOR2X1 NOR2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_14220_), .B(_14217_), .Y(_14221_) );
NAND3X1 NAND3X1_2970 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .B(_8750_), .C(_3170_), .Y(_14222_) );
NAND3X1 NAND3X1_2971 ( .gnd(gnd), .vdd(vdd), .A(_3119_), .B(_8757_), .C(_3118_), .Y(_14223_) );
NAND2X1 NAND2X1_2691 ( .gnd(gnd), .vdd(vdd), .A(_14222_), .B(_14223_), .Y(_14224_) );
NAND3X1 NAND3X1_2972 ( .gnd(gnd), .vdd(vdd), .A(_3299_), .B(_8762_), .C(_3298_), .Y(_14225_) );
NAND3X1 NAND3X1_2973 ( .gnd(gnd), .vdd(vdd), .A(_3028_), .B(_8774_), .C(_3027_), .Y(_14226_) );
NAND2X1 NAND2X1_2692 ( .gnd(gnd), .vdd(vdd), .A(_14225_), .B(_14226_), .Y(_14227_) );
OR2X2 OR2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_14224_), .B(_14227_), .Y(_14228_) );
NAND2X1 NAND2X1_2693 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__14_), .Y(_14229_) );
NAND3X1 NAND3X1_2974 ( .gnd(gnd), .vdd(vdd), .A(_2836_), .B(_8786_), .C(_2837_), .Y(_14230_) );
OAI21X1 OAI21X1_2567 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .B(_8792_), .C(_14230_), .Y(_14231_) );
NAND3X1 NAND3X1_2975 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_8794_), .C(_2666_), .Y(_14232_) );
OAI21X1 OAI21X1_2568 ( .gnd(gnd), .vdd(vdd), .A(_2783_), .B(_8799_), .C(_14232_), .Y(_14233_) );
NOR2X1 NOR2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_14233_), .B(_14231_), .Y(_14234_) );
AOI22X1 AOI22X1_558 ( .gnd(gnd), .vdd(vdd), .A(_76__14_), .B(_9482_), .C(_77__14_), .D(_9478_), .Y(_14235_) );
NAND2X1 NAND2X1_2694 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__14_), .Y(_14236_) );
NAND2X1 NAND2X1_2695 ( .gnd(gnd), .vdd(vdd), .A(_8806_), .B(_82__14_), .Y(_14237_) );
NAND3X1 NAND3X1_2976 ( .gnd(gnd), .vdd(vdd), .A(_14236_), .B(_14237_), .C(_14235_), .Y(_14238_) );
NAND2X1 NAND2X1_2696 ( .gnd(gnd), .vdd(vdd), .A(_9480_), .B(_73__14_), .Y(_14239_) );
NAND3X1 NAND3X1_2977 ( .gnd(gnd), .vdd(vdd), .A(_2596_), .B(_8803_), .C(_2595_), .Y(_14240_) );
NAND2X1 NAND2X1_2697 ( .gnd(gnd), .vdd(vdd), .A(_14240_), .B(_14239_), .Y(_14241_) );
INVX1 INVX1_3883 ( .gnd(gnd), .vdd(vdd), .A(_84__14_), .Y(_14242_) );
NOR2X1 NOR2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_14242_), .Y(_14243_) );
NOR2X1 NOR2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2310_), .Y(_14244_) );
NAND2X1 NAND2X1_2698 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__14_), .Y(_14245_) );
NAND3X1 NAND3X1_2978 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1934_), .C(_1935_), .Y(_14246_) );
NAND2X1 NAND2X1_2699 ( .gnd(gnd), .vdd(vdd), .A(_8845_), .B(_98__14_), .Y(_14247_) );
NAND3X1 NAND3X1_2979 ( .gnd(gnd), .vdd(vdd), .A(_14246_), .B(_14245_), .C(_14247_), .Y(_14248_) );
NOR3X1 NOR3X1_447 ( .gnd(gnd), .vdd(vdd), .A(_14243_), .B(_14248_), .C(_14244_), .Y(_14249_) );
NAND3X1 NAND3X1_2980 ( .gnd(gnd), .vdd(vdd), .A(_2272_), .B(_8829_), .C(_2273_), .Y(_14250_) );
NAND3X1 NAND3X1_2981 ( .gnd(gnd), .vdd(vdd), .A(_2166_), .B(_8831_), .C(_2167_), .Y(_14251_) );
NAND2X1 NAND2X1_2700 ( .gnd(gnd), .vdd(vdd), .A(_14250_), .B(_14251_), .Y(_14252_) );
NAND3X1 NAND3X1_2982 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_8834_), .C(_2108_), .Y(_14253_) );
NAND3X1 NAND3X1_2983 ( .gnd(gnd), .vdd(vdd), .A(_2218_), .B(_8836_), .C(_2219_), .Y(_14254_) );
NAND2X1 NAND2X1_2701 ( .gnd(gnd), .vdd(vdd), .A(_14253_), .B(_14254_), .Y(_14255_) );
NOR2X1 NOR2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_14255_), .B(_14252_), .Y(_14256_) );
AOI22X1 AOI22X1_559 ( .gnd(gnd), .vdd(vdd), .A(_92__14_), .B(_8843_), .C(_91__14_), .D(_8823_), .Y(_14257_) );
AOI22X1 AOI22X1_560 ( .gnd(gnd), .vdd(vdd), .A(_94__14_), .B(_8841_), .C(_93__14_), .D(_8840_), .Y(_14258_) );
NAND2X1 NAND2X1_2702 ( .gnd(gnd), .vdd(vdd), .A(_14258_), .B(_14257_), .Y(_14259_) );
NAND2X1 NAND2X1_2703 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__14_), .Y(_14260_) );
NAND2X1 NAND2X1_2704 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_106__14_), .Y(_14261_) );
NAND2X1 NAND2X1_2705 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__14_), .Y(_14262_) );
NAND2X1 NAND2X1_2706 ( .gnd(gnd), .vdd(vdd), .A(_14261_), .B(_14262_), .Y(_14263_) );
NAND2X1 NAND2X1_2707 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__14_), .Y(_14264_) );
NAND2X1 NAND2X1_2708 ( .gnd(gnd), .vdd(vdd), .A(_8862_), .B(_117__14_), .Y(_14265_) );
NAND2X1 NAND2X1_2709 ( .gnd(gnd), .vdd(vdd), .A(_14265_), .B(_14264_), .Y(_14266_) );
NOR2X1 NOR2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_14266_), .B(_14263_), .Y(_14267_) );
NAND2X1 NAND2X1_2710 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__14_), .Y(_14268_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_7160_), .B(_9930_), .C(_7204_), .D(_9929_), .Y(_14269_) );
NOR2X1 NOR2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7339_), .Y(_14270_) );
NOR2X1 NOR2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7296_), .Y(_14271_) );
NOR3X1 NOR3X1_448 ( .gnd(gnd), .vdd(vdd), .A(_14270_), .B(_14271_), .C(_14269_), .Y(_14272_) );
NAND2X1 NAND2X1_2711 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__14_), .Y(_14273_) );
NAND2X1 NAND2X1_2712 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__14_), .Y(_14274_) );
NAND2X1 NAND2X1_2713 ( .gnd(gnd), .vdd(vdd), .A(_14273_), .B(_14274_), .Y(_14275_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_7382_), .B(_9940_), .C(_7250_), .D(_9941_), .Y(_14276_) );
NOR2X1 NOR2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_14276_), .B(_14275_), .Y(_14277_) );
NAND3X1 NAND3X1_2984 ( .gnd(gnd), .vdd(vdd), .A(_14268_), .B(_14272_), .C(_14277_), .Y(_14278_) );
AOI22X1 AOI22X1_561 ( .gnd(gnd), .vdd(vdd), .A(_20__14_), .B(_8898_), .C(_249__14_), .D(_9053_), .Y(_14279_) );
AOI22X1 AOI22X1_562 ( .gnd(gnd), .vdd(vdd), .A(_250__14_), .B(_9082_), .C(_175__14_), .D(_8904_), .Y(_14280_) );
NAND2X1 NAND2X1_2714 ( .gnd(gnd), .vdd(vdd), .A(_14279_), .B(_14280_), .Y(_14281_) );
NAND2X1 NAND2X1_2715 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__14_), .Y(_14282_) );
NAND2X1 NAND2X1_2716 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__14_), .Y(_14283_) );
AOI22X1 AOI22X1_563 ( .gnd(gnd), .vdd(vdd), .A(_19__14_), .B(_8914_), .C(_210__14_), .D(_8918_), .Y(_14284_) );
NAND3X1 NAND3X1_2985 ( .gnd(gnd), .vdd(vdd), .A(_14282_), .B(_14283_), .C(_14284_), .Y(_14285_) );
NOR2X1 NOR2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_14281_), .B(_14285_), .Y(_14286_) );
AOI22X1 AOI22X1_564 ( .gnd(gnd), .vdd(vdd), .A(_123__14_), .B(_8928_), .C(_9__14_), .D(_8926_), .Y(_14287_) );
NAND2X1 NAND2X1_2717 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__14_), .Y(_14288_) );
NAND2X1 NAND2X1_2718 ( .gnd(gnd), .vdd(vdd), .A(_8933_), .B(_134__14_), .Y(_14289_) );
NAND3X1 NAND3X1_2986 ( .gnd(gnd), .vdd(vdd), .A(_14288_), .B(_14289_), .C(_14287_), .Y(_14290_) );
AOI22X1 AOI22X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4__14_), .B(_8937_), .C(_176__14_), .D(_8939_), .Y(_14291_) );
NAND2X1 NAND2X1_2719 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__14_), .Y(_14292_) );
NAND2X1 NAND2X1_2720 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__14_), .Y(_14293_) );
NAND3X1 NAND3X1_2987 ( .gnd(gnd), .vdd(vdd), .A(_14292_), .B(_14293_), .C(_14291_), .Y(_14294_) );
NOR2X1 NOR2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_14294_), .B(_14290_), .Y(_14295_) );
NAND2X1 NAND2X1_2721 ( .gnd(gnd), .vdd(vdd), .A(_14286_), .B(_14295_), .Y(_14296_) );
AOI22X1 AOI22X1_566 ( .gnd(gnd), .vdd(vdd), .A(_47__14_), .B(_9161_), .C(_238__14_), .D(_8893_), .Y(_14297_) );
NAND2X1 NAND2X1_2722 ( .gnd(gnd), .vdd(vdd), .A(_9150_), .B(_21__14_), .Y(_14298_) );
NAND2X1 NAND2X1_2723 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .B(_185__14_), .Y(_14299_) );
NAND3X1 NAND3X1_2988 ( .gnd(gnd), .vdd(vdd), .A(_14298_), .B(_14299_), .C(_14297_), .Y(_14300_) );
AOI22X1 AOI22X1_567 ( .gnd(gnd), .vdd(vdd), .A(_246__14_), .B(_9356_), .C(_226__14_), .D(_9357_), .Y(_14301_) );
NAND2X1 NAND2X1_2724 ( .gnd(gnd), .vdd(vdd), .A(_9157_), .B(_231__14_), .Y(_14302_) );
NAND2X1 NAND2X1_2725 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_46__14_), .Y(_14303_) );
NAND3X1 NAND3X1_2989 ( .gnd(gnd), .vdd(vdd), .A(_14302_), .B(_14303_), .C(_14301_), .Y(_14304_) );
NOR2X1 NOR2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_14300_), .B(_14304_), .Y(_14305_) );
NAND2X1 NAND2X1_2726 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_178__14_), .Y(_14306_) );
NAND2X1 NAND2X1_2727 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__14_), .Y(_14307_) );
AOI22X1 AOI22X1_568 ( .gnd(gnd), .vdd(vdd), .A(_37__14_), .B(_8978_), .C(_35__14_), .D(_8980_), .Y(_14308_) );
NAND3X1 NAND3X1_2990 ( .gnd(gnd), .vdd(vdd), .A(_14306_), .B(_14307_), .C(_14308_), .Y(_14309_) );
NAND2X1 NAND2X1_2728 ( .gnd(gnd), .vdd(vdd), .A(_8966_), .B(_237__14_), .Y(_14310_) );
NAND2X1 NAND2X1_2729 ( .gnd(gnd), .vdd(vdd), .A(_9154_), .B(_253__14_), .Y(_14311_) );
AOI22X1 AOI22X1_569 ( .gnd(gnd), .vdd(vdd), .A(_145__14_), .B(_9177_), .C(_213__14_), .D(_8989_), .Y(_14312_) );
NAND3X1 NAND3X1_2991 ( .gnd(gnd), .vdd(vdd), .A(_14310_), .B(_14311_), .C(_14312_), .Y(_14313_) );
NOR2X1 NOR2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_14313_), .B(_14309_), .Y(_14314_) );
NAND2X1 NAND2X1_2730 ( .gnd(gnd), .vdd(vdd), .A(_14305_), .B(_14314_), .Y(_14315_) );
NOR2X1 NOR2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_14296_), .B(_14315_), .Y(_14316_) );
NAND2X1 NAND2X1_2731 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__14_), .Y(_14317_) );
NAND2X1 NAND2X1_2732 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__14_), .Y(_14318_) );
AOI22X1 AOI22X1_570 ( .gnd(gnd), .vdd(vdd), .A(_13__14_), .B(_9007_), .C(_239__14_), .D(_9076_), .Y(_14319_) );
NAND3X1 NAND3X1_2992 ( .gnd(gnd), .vdd(vdd), .A(_14317_), .B(_14318_), .C(_14319_), .Y(_14320_) );
AOI22X1 AOI22X1_571 ( .gnd(gnd), .vdd(vdd), .A(_206__14_), .B(_9013_), .C(_242__14_), .D(_9035_), .Y(_14321_) );
NAND2X1 NAND2X1_2733 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__14_), .Y(_14322_) );
NAND2X1 NAND2X1_2734 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__14_), .Y(_14323_) );
NAND3X1 NAND3X1_2993 ( .gnd(gnd), .vdd(vdd), .A(_14322_), .B(_14323_), .C(_14321_), .Y(_14324_) );
NOR2X1 NOR2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(_14320_), .B(_14324_), .Y(_14325_) );
AOI22X1 AOI22X1_572 ( .gnd(gnd), .vdd(vdd), .A(_222__14_), .B(_9024_), .C(_220__14_), .D(_9026_), .Y(_14326_) );
NAND2X1 NAND2X1_2735 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__14_), .Y(_14327_) );
NAND2X1 NAND2X1_2736 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__14_), .Y(_14328_) );
NAND3X1 NAND3X1_2994 ( .gnd(gnd), .vdd(vdd), .A(_14327_), .B(_14328_), .C(_14326_), .Y(_14329_) );
AOI22X1 AOI22X1_573 ( .gnd(gnd), .vdd(vdd), .A(_18__14_), .B(_9037_), .C(_240__14_), .D(_9011_), .Y(_14330_) );
NAND2X1 NAND2X1_2737 ( .gnd(gnd), .vdd(vdd), .A(_9040_), .B(_221__14_), .Y(_14331_) );
NAND2X1 NAND2X1_2738 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__14_), .Y(_14332_) );
NAND3X1 NAND3X1_2995 ( .gnd(gnd), .vdd(vdd), .A(_14331_), .B(_14332_), .C(_14330_), .Y(_14333_) );
NOR2X1 NOR2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_14329_), .B(_14333_), .Y(_14334_) );
NAND2X1 NAND2X1_2739 ( .gnd(gnd), .vdd(vdd), .A(_14325_), .B(_14334_), .Y(_14335_) );
AOI22X1 AOI22X1_574 ( .gnd(gnd), .vdd(vdd), .A(_225__14_), .B(_9048_), .C(_167__14_), .D(_9050_), .Y(_14336_) );
NAND2X1 NAND2X1_2740 ( .gnd(gnd), .vdd(vdd), .A(_8955_), .B(_236__14_), .Y(_14337_) );
NAND2X1 NAND2X1_2741 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__14_), .Y(_14338_) );
NAND3X1 NAND3X1_2996 ( .gnd(gnd), .vdd(vdd), .A(_14337_), .B(_14338_), .C(_14336_), .Y(_14339_) );
NAND2X1 NAND2X1_2742 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__14_), .Y(_14340_) );
NAND2X1 NAND2X1_2743 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__14_), .Y(_14341_) );
AOI22X1 AOI22X1_575 ( .gnd(gnd), .vdd(vdd), .A(_224__14_), .B(_9064_), .C(_27__14_), .D(_9066_), .Y(_14342_) );
NAND3X1 NAND3X1_2997 ( .gnd(gnd), .vdd(vdd), .A(_14340_), .B(_14341_), .C(_14342_), .Y(_14343_) );
NOR2X1 NOR2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_14339_), .B(_14343_), .Y(_14344_) );
AOI22X1 AOI22X1_576 ( .gnd(gnd), .vdd(vdd), .A(_184__14_), .B(_9073_), .C(_183__14_), .D(_9071_), .Y(_14345_) );
NAND2X1 NAND2X1_2744 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__14_), .Y(_14346_) );
NAND2X1 NAND2X1_2745 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__14_), .Y(_14347_) );
NAND3X1 NAND3X1_2998 ( .gnd(gnd), .vdd(vdd), .A(_14346_), .B(_14347_), .C(_14345_), .Y(_14348_) );
AOI22X1 AOI22X1_577 ( .gnd(gnd), .vdd(vdd), .A(_43__14_), .B(_9084_), .C(_248__14_), .D(_8901_), .Y(_14349_) );
NAND2X1 NAND2X1_2746 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__14_), .Y(_14350_) );
NAND2X1 NAND2X1_2747 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__14_), .Y(_14351_) );
NAND3X1 NAND3X1_2999 ( .gnd(gnd), .vdd(vdd), .A(_14350_), .B(_14351_), .C(_14349_), .Y(_14352_) );
NOR2X1 NOR2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_14348_), .B(_14352_), .Y(_14353_) );
NAND2X1 NAND2X1_2748 ( .gnd(gnd), .vdd(vdd), .A(_14344_), .B(_14353_), .Y(_14354_) );
NOR2X1 NOR2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_14335_), .B(_14354_), .Y(_14355_) );
NAND3X1 NAND3X1_3000 ( .gnd(gnd), .vdd(vdd), .A(_6833_), .B(_9143_), .C(_6834_), .Y(_14356_) );
NAND3X1 NAND3X1_3001 ( .gnd(gnd), .vdd(vdd), .A(_6985_), .B(_9145_), .C(_6986_), .Y(_14357_) );
NAND2X1 NAND2X1_2749 ( .gnd(gnd), .vdd(vdd), .A(_14356_), .B(_14357_), .Y(_14358_) );
NAND3X1 NAND3X1_3002 ( .gnd(gnd), .vdd(vdd), .A(_5069_), .B(_9135_), .C(_5070_), .Y(_14359_) );
NAND3X1 NAND3X1_3003 ( .gnd(gnd), .vdd(vdd), .A(_6951_), .B(_9137_), .C(_6952_), .Y(_14360_) );
NAND2X1 NAND2X1_2750 ( .gnd(gnd), .vdd(vdd), .A(_14360_), .B(_14359_), .Y(_14361_) );
NOR2X1 NOR2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_14358_), .B(_14361_), .Y(_14362_) );
NAND3X1 NAND3X1_3004 ( .gnd(gnd), .vdd(vdd), .A(_8333_), .B(_9188_), .C(_8334_), .Y(_14363_) );
NAND3X1 NAND3X1_3005 ( .gnd(gnd), .vdd(vdd), .A(_15944_), .B(_9109_), .C(_15945_), .Y(_14364_) );
NAND3X1 NAND3X1_3006 ( .gnd(gnd), .vdd(vdd), .A(_16149_), .B(_9115_), .C(_16150_), .Y(_14365_) );
NAND3X1 NAND3X1_3007 ( .gnd(gnd), .vdd(vdd), .A(_14364_), .B(_14365_), .C(_14363_), .Y(_14366_) );
AOI22X1 AOI22X1_578 ( .gnd(gnd), .vdd(vdd), .A(_234__14_), .B(_9182_), .C(_34__14_), .D(_9183_), .Y(_14367_) );
AOI22X1 AOI22X1_579 ( .gnd(gnd), .vdd(vdd), .A(_100__14_), .B(_9346_), .C(_45__14_), .D(_9185_), .Y(_14368_) );
NAND2X1 NAND2X1_2751 ( .gnd(gnd), .vdd(vdd), .A(_14368_), .B(_14367_), .Y(_14369_) );
NAND3X1 NAND3X1_3008 ( .gnd(gnd), .vdd(vdd), .A(_4717_), .B(_9140_), .C(_4716_), .Y(_14370_) );
OAI21X1 OAI21X1_2569 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_10036_), .C(_14370_), .Y(_14371_) );
NOR3X1 NOR3X1_449 ( .gnd(gnd), .vdd(vdd), .A(_14371_), .B(_14366_), .C(_14369_), .Y(_14372_) );
NAND3X1 NAND3X1_3009 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_9133_), .C(_3444_), .Y(_14373_) );
NAND3X1 NAND3X1_3010 ( .gnd(gnd), .vdd(vdd), .A(_4941_), .B(_9097_), .C(_4942_), .Y(_14374_) );
NAND3X1 NAND3X1_3011 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .B(_9102_), .C(_5116_), .Y(_14375_) );
NAND3X1 NAND3X1_3012 ( .gnd(gnd), .vdd(vdd), .A(_14374_), .B(_14375_), .C(_14373_), .Y(_14376_) );
AOI22X1 AOI22X1_580 ( .gnd(gnd), .vdd(vdd), .A(_38__14_), .B(_9129_), .C(_16__14_), .D(_9127_), .Y(_14377_) );
AOI22X1 AOI22X1_581 ( .gnd(gnd), .vdd(vdd), .A(_39__14_), .B(_9099_), .C(_204__14_), .D(_9104_), .Y(_14378_) );
NAND2X1 NAND2X1_2752 ( .gnd(gnd), .vdd(vdd), .A(_14377_), .B(_14378_), .Y(_14379_) );
NOR2X1 NOR2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_14376_), .B(_14379_), .Y(_14380_) );
NAND3X1 NAND3X1_3013 ( .gnd(gnd), .vdd(vdd), .A(_14362_), .B(_14372_), .C(_14380_), .Y(_14381_) );
AOI22X1 AOI22X1_582 ( .gnd(gnd), .vdd(vdd), .A(_227__14_), .B(_9170_), .C(_30__14_), .D(_9167_), .Y(_14382_) );
AOI22X1 AOI22X1_583 ( .gnd(gnd), .vdd(vdd), .A(_209__14_), .B(_8957_), .C(_33__14_), .D(_8991_), .Y(_14383_) );
NAND2X1 NAND2X1_2753 ( .gnd(gnd), .vdd(vdd), .A(_14382_), .B(_14383_), .Y(_14384_) );
AOI22X1 AOI22X1_584 ( .gnd(gnd), .vdd(vdd), .A(_44__14_), .B(_8968_), .C(_42__14_), .D(_8963_), .Y(_14385_) );
AOI22X1 AOI22X1_585 ( .gnd(gnd), .vdd(vdd), .A(_208__14_), .B(_8950_), .C(_243__14_), .D(_9153_), .Y(_14386_) );
NAND2X1 NAND2X1_2754 ( .gnd(gnd), .vdd(vdd), .A(_14385_), .B(_14386_), .Y(_14387_) );
NOR2X1 NOR2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_14384_), .B(_14387_), .Y(_14388_) );
AOI22X1 AOI22X1_586 ( .gnd(gnd), .vdd(vdd), .A(_22__14_), .B(_9382_), .C(_3__14_), .D(_9383_), .Y(_14389_) );
NAND2X1 NAND2X1_2755 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_219__14_), .Y(_14390_) );
NAND2X1 NAND2X1_2756 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(_232__14_), .Y(_14391_) );
NAND3X1 NAND3X1_3014 ( .gnd(gnd), .vdd(vdd), .A(_14390_), .B(_14391_), .C(_14389_), .Y(_14392_) );
AOI22X1 AOI22X1_587 ( .gnd(gnd), .vdd(vdd), .A(_255__14_), .B(_8986_), .C(_254__14_), .D(_8984_), .Y(_14393_) );
AOI22X1 AOI22X1_588 ( .gnd(gnd), .vdd(vdd), .A(_203__14_), .B(_9018_), .C(_156__14_), .D(_8973_), .Y(_14394_) );
NAND2X1 NAND2X1_2757 ( .gnd(gnd), .vdd(vdd), .A(_14393_), .B(_14394_), .Y(_14395_) );
NOR2X1 NOR2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_14392_), .B(_14395_), .Y(_14396_) );
NAND2X1 NAND2X1_2758 ( .gnd(gnd), .vdd(vdd), .A(_14388_), .B(_14396_), .Y(_14397_) );
AOI22X1 AOI22X1_589 ( .gnd(gnd), .vdd(vdd), .A(_201__14_), .B(_9124_), .C(_212__14_), .D(_9345_), .Y(_14398_) );
NAND3X1 NAND3X1_3015 ( .gnd(gnd), .vdd(vdd), .A(_8447_), .B(_9348_), .C(_8446_), .Y(_14399_) );
NAND3X1 NAND3X1_3016 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_507_), .C(_508_), .Y(_14400_) );
AND2X2 AND2X2_1612 ( .gnd(gnd), .vdd(vdd), .A(_14400_), .B(_14399_), .Y(_14401_) );
NAND2X1 NAND2X1_2759 ( .gnd(gnd), .vdd(vdd), .A(_14398_), .B(_14401_), .Y(_14402_) );
NAND3X1 NAND3X1_3017 ( .gnd(gnd), .vdd(vdd), .A(_15153_), .B(_9208_), .C(_15154_), .Y(_14403_) );
OAI21X1 OAI21X1_2570 ( .gnd(gnd), .vdd(vdd), .A(_15116_), .B(_9211_), .C(_14403_), .Y(_14404_) );
NAND3X1 NAND3X1_3018 ( .gnd(gnd), .vdd(vdd), .A(_15501_), .B(_9222_), .C(_15502_), .Y(_14405_) );
NAND3X1 NAND3X1_3019 ( .gnd(gnd), .vdd(vdd), .A(_15448_), .B(_9224_), .C(_15447_), .Y(_14406_) );
NAND2X1 NAND2X1_2760 ( .gnd(gnd), .vdd(vdd), .A(_14405_), .B(_14406_), .Y(_14407_) );
NOR2X1 NOR2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_14407_), .B(_14404_), .Y(_14408_) );
NAND3X1 NAND3X1_3020 ( .gnd(gnd), .vdd(vdd), .A(_15279_), .B(_9217_), .C(_15280_), .Y(_14409_) );
NAND3X1 NAND3X1_3021 ( .gnd(gnd), .vdd(vdd), .A(_15227_), .B(_9219_), .C(_15226_), .Y(_14410_) );
NAND2X1 NAND2X1_2761 ( .gnd(gnd), .vdd(vdd), .A(_14410_), .B(_14409_), .Y(_14411_) );
NAND3X1 NAND3X1_3022 ( .gnd(gnd), .vdd(vdd), .A(_15677_), .B(_9192_), .C(_15678_), .Y(_14412_) );
NAND3X1 NAND3X1_3023 ( .gnd(gnd), .vdd(vdd), .A(_15734_), .B(_9199_), .C(_15733_), .Y(_14413_) );
NAND2X1 NAND2X1_2762 ( .gnd(gnd), .vdd(vdd), .A(_14413_), .B(_14412_), .Y(_14414_) );
NOR2X1 NOR2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_14414_), .B(_14411_), .Y(_14415_) );
NOR3X1 NOR3X1_450 ( .gnd(gnd), .vdd(vdd), .A(_16200_), .B(_10083_), .C(_16201_), .Y(_14416_) );
NAND3X1 NAND3X1_3024 ( .gnd(gnd), .vdd(vdd), .A(_15327_), .B(_9205_), .C(_15328_), .Y(_14417_) );
OAI21X1 OAI21X1_2571 ( .gnd(gnd), .vdd(vdd), .A(_15356_), .B(_10085_), .C(_14417_), .Y(_14418_) );
NAND3X1 NAND3X1_3025 ( .gnd(gnd), .vdd(vdd), .A(_15559_), .B(_9233_), .C(_15560_), .Y(_14419_) );
NAND3X1 NAND3X1_3026 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15625_), .C(_15624_), .Y(_14420_) );
NAND2X1 NAND2X1_2763 ( .gnd(gnd), .vdd(vdd), .A(_14419_), .B(_14420_), .Y(_14421_) );
NOR3X1 NOR3X1_451 ( .gnd(gnd), .vdd(vdd), .A(_14418_), .B(_14421_), .C(_14416_), .Y(_14422_) );
NAND3X1 NAND3X1_3027 ( .gnd(gnd), .vdd(vdd), .A(_14408_), .B(_14415_), .C(_14422_), .Y(_14423_) );
NAND3X1 NAND3X1_3028 ( .gnd(gnd), .vdd(vdd), .A(_15887_), .B(_9120_), .C(_15888_), .Y(_14424_) );
NAND3X1 NAND3X1_3029 ( .gnd(gnd), .vdd(vdd), .A(_15394_), .B(_9197_), .C(_15395_), .Y(_14425_) );
AOI22X1 AOI22X1_590 ( .gnd(gnd), .vdd(vdd), .A(_251__14_), .B(_9320_), .C(_235__14_), .D(_9324_), .Y(_14426_) );
AOI22X1 AOI22X1_591 ( .gnd(gnd), .vdd(vdd), .A(_14__14_), .B(_9274_), .C(_252__14_), .D(_9326_), .Y(_14427_) );
NAND2X1 NAND2X1_2764 ( .gnd(gnd), .vdd(vdd), .A(_14427_), .B(_14426_), .Y(_14428_) );
NAND2X1 NAND2X1_2765 ( .gnd(gnd), .vdd(vdd), .A(_9298_), .B(_186__14_), .Y(_14429_) );
AOI22X1 AOI22X1_592 ( .gnd(gnd), .vdd(vdd), .A(_67__14_), .B(_9286_), .C(_199__14_), .D(_9289_), .Y(_14430_) );
NAND2X1 NAND2X1_2766 ( .gnd(gnd), .vdd(vdd), .A(_14429_), .B(_14430_), .Y(_14431_) );
AOI21X1 AOI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_216__14_), .B(_9260_), .C(_14431_), .Y(_14432_) );
OAI21X1 OAI21X1_2572 ( .gnd(gnd), .vdd(vdd), .A(_7691_), .B(_10121_), .C(_14432_), .Y(_14433_) );
NOR2X1 NOR2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_14428_), .B(_14433_), .Y(_14434_) );
NAND2X1 NAND2X1_2767 ( .gnd(gnd), .vdd(vdd), .A(_10110_), .B(_32__14_), .Y(_14435_) );
AOI22X1 AOI22X1_593 ( .gnd(gnd), .vdd(vdd), .A(_50__14_), .B(_9778_), .C(_65__14_), .D(_9277_), .Y(_14436_) );
NAND3X1 NAND3X1_3030 ( .gnd(gnd), .vdd(vdd), .A(_1781_), .B(_9255_), .C(_1780_), .Y(_14437_) );
OAI21X1 OAI21X1_2573 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_8722_), .C(_14437_), .Y(_14438_) );
NOR2X1 NOR2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_9295_), .B(_3621_), .Y(_14439_) );
INVX1 INVX1_3884 ( .gnd(gnd), .vdd(vdd), .A(_9315_), .Y(_14440_) );
NOR3X1 NOR3X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_14440_), .C(_2371_), .Y(_14441_) );
NOR3X1 NOR3X1_453 ( .gnd(gnd), .vdd(vdd), .A(_14439_), .B(_14441_), .C(_14438_), .Y(_14442_) );
NAND3X1 NAND3X1_3031 ( .gnd(gnd), .vdd(vdd), .A(_14435_), .B(_14436_), .C(_14442_), .Y(_14443_) );
NAND2X1 NAND2X1_2768 ( .gnd(gnd), .vdd(vdd), .A(_9235_), .B(_187__14_), .Y(_14444_) );
NAND3X1 NAND3X1_3032 ( .gnd(gnd), .vdd(vdd), .A(_7066_), .B(_9266_), .C(_7065_), .Y(_14445_) );
OAI21X1 OAI21X1_2574 ( .gnd(gnd), .vdd(vdd), .A(_7111_), .B(_9245_), .C(_14445_), .Y(_14446_) );
AOI21X1 AOI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_182__14_), .B(_9300_), .C(_14446_), .Y(_14447_) );
NAND3X1 NAND3X1_3033 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_9268_), .C(_1187_), .Y(_14448_) );
OAI21X1 OAI21X1_2575 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_9263_), .C(_14448_), .Y(_14449_) );
NAND3X1 NAND3X1_3034 ( .gnd(gnd), .vdd(vdd), .A(_15826_), .B(_9292_), .C(_15825_), .Y(_14450_) );
OAI21X1 OAI21X1_2576 ( .gnd(gnd), .vdd(vdd), .A(_14928_), .B(_9276_), .C(_14450_), .Y(_14451_) );
NOR2X1 NOR2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_14451_), .B(_14449_), .Y(_14452_) );
NAND3X1 NAND3X1_3035 ( .gnd(gnd), .vdd(vdd), .A(_14444_), .B(_14452_), .C(_14447_), .Y(_14453_) );
NOR3X1 NOR3X1_454 ( .gnd(gnd), .vdd(vdd), .A(_9304_), .B(_8182_), .C(_8181_), .Y(_14454_) );
NOR2X1 NOR2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_10875_), .B(_8253_), .Y(_14455_) );
NOR3X1 NOR3X1_455 ( .gnd(gnd), .vdd(vdd), .A(_9249_), .B(_7735_), .C(_7736_), .Y(_14456_) );
NOR3X1 NOR3X1_456 ( .gnd(gnd), .vdd(vdd), .A(_14455_), .B(_14456_), .C(_14454_), .Y(_14457_) );
AOI22X1 AOI22X1_594 ( .gnd(gnd), .vdd(vdd), .A(_217__14_), .B(_9281_), .C(_233__14_), .D(_9310_), .Y(_14458_) );
AOI22X1 AOI22X1_595 ( .gnd(gnd), .vdd(vdd), .A(_31__14_), .B(_9283_), .C(_15__14_), .D(_9313_), .Y(_14459_) );
NAND3X1 NAND3X1_3036 ( .gnd(gnd), .vdd(vdd), .A(_14457_), .B(_14458_), .C(_14459_), .Y(_14460_) );
NOR3X1 NOR3X1_457 ( .gnd(gnd), .vdd(vdd), .A(_14460_), .B(_14453_), .C(_14443_), .Y(_14461_) );
NAND3X1 NAND3X1_3037 ( .gnd(gnd), .vdd(vdd), .A(_14434_), .B(_14425_), .C(_14461_), .Y(_14462_) );
AOI21X1 AOI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_157__14_), .B(_9232_), .C(_14462_), .Y(_14463_) );
AOI22X1 AOI22X1_596 ( .gnd(gnd), .vdd(vdd), .A(_155__14_), .B(_9333_), .C(_172__14_), .D(_9332_), .Y(_14464_) );
NAND3X1 NAND3X1_3038 ( .gnd(gnd), .vdd(vdd), .A(_14424_), .B(_14464_), .C(_14463_), .Y(_14465_) );
NOR3X1 NOR3X1_458 ( .gnd(gnd), .vdd(vdd), .A(_14423_), .B(_14465_), .C(_14402_), .Y(_14466_) );
AOI22X1 AOI22X1_597 ( .gnd(gnd), .vdd(vdd), .A(_256__14_), .B(_9113_), .C(_142__14_), .D(_9118_), .Y(_14467_) );
NAND2X1 NAND2X1_2769 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__14_), .Y(_14468_) );
NAND2X1 NAND2X1_2770 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__14_), .Y(_14469_) );
NAND3X1 NAND3X1_3039 ( .gnd(gnd), .vdd(vdd), .A(_14468_), .B(_14469_), .C(_14467_), .Y(_14470_) );
NAND2X1 NAND2X1_2771 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__14_), .Y(_14471_) );
NAND3X1 NAND3X1_3040 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_9339_), .C(_470_), .Y(_14472_) );
AOI22X1 AOI22X1_598 ( .gnd(gnd), .vdd(vdd), .A(_111__14_), .B(_9342_), .C(_12__14_), .D(_9341_), .Y(_14473_) );
NAND3X1 NAND3X1_3041 ( .gnd(gnd), .vdd(vdd), .A(_14473_), .B(_14471_), .C(_14472_), .Y(_14474_) );
NOR2X1 NOR2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_14470_), .B(_14474_), .Y(_14475_) );
AOI22X1 AOI22X1_599 ( .gnd(gnd), .vdd(vdd), .A(_40__14_), .B(_8952_), .C(_29__14_), .D(_9176_), .Y(_14476_) );
AOI22X1 AOI22X1_600 ( .gnd(gnd), .vdd(vdd), .A(_247__14_), .B(_9165_), .C(_218__14_), .D(_9169_), .Y(_14477_) );
NAND2X1 NAND2X1_2772 ( .gnd(gnd), .vdd(vdd), .A(_14477_), .B(_14476_), .Y(_14478_) );
NAND3X1 NAND3X1_3042 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16104_), .C(_16105_), .Y(_14479_) );
NAND3X1 NAND3X1_3043 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16049_), .C(_16050_), .Y(_14480_) );
NAND2X1 NAND2X1_2773 ( .gnd(gnd), .vdd(vdd), .A(_14479_), .B(_14480_), .Y(_14481_) );
NAND3X1 NAND3X1_3044 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8583_), .C(_8582_), .Y(_14482_) );
OAI21X1 OAI21X1_2577 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_9361_), .C(_14482_), .Y(_14483_) );
NOR2X1 NOR2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_14481_), .B(_14483_), .Y(_14484_) );
NAND2X1 NAND2X1_2774 ( .gnd(gnd), .vdd(vdd), .A(_15993_), .B(_15994_), .Y(_14485_) );
NAND3X1 NAND3X1_3045 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8636_), .C(_8637_), .Y(_14486_) );
OAI21X1 OAI21X1_2578 ( .gnd(gnd), .vdd(vdd), .A(_14485_), .B(_9215_), .C(_14486_), .Y(_14487_) );
NAND3X1 NAND3X1_3046 ( .gnd(gnd), .vdd(vdd), .A(_8691_), .B(_9371_), .C(_8690_), .Y(_14488_) );
NAND3X1 NAND3X1_3047 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_333_), .C(_334_), .Y(_14489_) );
NAND2X1 NAND2X1_2775 ( .gnd(gnd), .vdd(vdd), .A(_14489_), .B(_14488_), .Y(_14490_) );
NOR2X1 NOR2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_14487_), .B(_14490_), .Y(_14491_) );
AOI22X1 AOI22X1_601 ( .gnd(gnd), .vdd(vdd), .A(_244__14_), .B(_9160_), .C(_177__14_), .D(_8961_), .Y(_14492_) );
NAND3X1 NAND3X1_3048 ( .gnd(gnd), .vdd(vdd), .A(_14484_), .B(_14491_), .C(_14492_), .Y(_14493_) );
NOR2X1 NOR2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_14478_), .B(_14493_), .Y(_14494_) );
NAND3X1 NAND3X1_3049 ( .gnd(gnd), .vdd(vdd), .A(_14466_), .B(_14475_), .C(_14494_), .Y(_14495_) );
NOR3X1 NOR3X1_459 ( .gnd(gnd), .vdd(vdd), .A(_14381_), .B(_14397_), .C(_14495_), .Y(_14496_) );
NAND3X1 NAND3X1_3050 ( .gnd(gnd), .vdd(vdd), .A(_14316_), .B(_14355_), .C(_14496_), .Y(_14497_) );
NAND3X1 NAND3X1_3051 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_1557_), .C(_1558_), .Y(_14498_) );
NAND3X1 NAND3X1_3052 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_1642_), .C(_1643_), .Y(_14499_) );
NAND2X1 NAND2X1_2776 ( .gnd(gnd), .vdd(vdd), .A(_14498_), .B(_14499_), .Y(_14500_) );
NOR3X1 NOR3X1_460 ( .gnd(gnd), .vdd(vdd), .A(_14278_), .B(_14500_), .C(_14497_), .Y(_14501_) );
NAND3X1 NAND3X1_3053 ( .gnd(gnd), .vdd(vdd), .A(_14260_), .B(_14267_), .C(_14501_), .Y(_14502_) );
NAND2X1 NAND2X1_2777 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__14_), .Y(_14503_) );
AOI22X1 AOI22X1_602 ( .gnd(gnd), .vdd(vdd), .A(_115__14_), .B(_9399_), .C(_116__14_), .D(_9401_), .Y(_14504_) );
AOI22X1 AOI22X1_603 ( .gnd(gnd), .vdd(vdd), .A(_108__14_), .B(_9404_), .C(_109__14_), .D(_9406_), .Y(_14505_) );
NAND2X1 NAND2X1_2778 ( .gnd(gnd), .vdd(vdd), .A(_14504_), .B(_14505_), .Y(_14506_) );
NAND2X1 NAND2X1_2779 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_125__14_), .Y(_14507_) );
NAND2X1 NAND2X1_2780 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_122__14_), .Y(_14508_) );
NAND2X1 NAND2X1_2781 ( .gnd(gnd), .vdd(vdd), .A(_14507_), .B(_14508_), .Y(_14509_) );
NOR2X1 NOR2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_1125_), .Y(_14510_) );
AND2X2 AND2X2_1613 ( .gnd(gnd), .vdd(vdd), .A(_120__14_), .B(_9415_), .Y(_14511_) );
NOR3X1 NOR3X1_461 ( .gnd(gnd), .vdd(vdd), .A(_14510_), .B(_14511_), .C(_14509_), .Y(_14512_) );
AOI22X1 AOI22X1_604 ( .gnd(gnd), .vdd(vdd), .A(_132__14_), .B(_9420_), .C(_131__14_), .D(_9418_), .Y(_14513_) );
NAND2X1 NAND2X1_2782 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__14_), .Y(_14514_) );
NAND2X1 NAND2X1_2783 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__14_), .Y(_14515_) );
NAND3X1 NAND3X1_3054 ( .gnd(gnd), .vdd(vdd), .A(_14514_), .B(_14515_), .C(_14513_), .Y(_14516_) );
NAND3X1 NAND3X1_3055 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_9431_), .C(_565_), .Y(_14517_) );
NAND2X1 NAND2X1_2784 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__14_), .Y(_14518_) );
NAND2X1 NAND2X1_2785 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__14_), .Y(_14519_) );
NAND3X1 NAND3X1_3056 ( .gnd(gnd), .vdd(vdd), .A(_14519_), .B(_14517_), .C(_14518_), .Y(_14520_) );
AOI21X1 AOI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__14_), .C(_14520_), .Y(_14521_) );
NAND2X1 NAND2X1_2786 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__14_), .Y(_14522_) );
NAND2X1 NAND2X1_2787 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_136__14_), .Y(_14523_) );
NAND3X1 NAND3X1_3057 ( .gnd(gnd), .vdd(vdd), .A(_14522_), .B(_14523_), .C(_14521_), .Y(_14524_) );
NAND3X1 NAND3X1_3058 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_9410_), .C(_1028_), .Y(_14525_) );
NAND2X1 NAND2X1_2788 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__14_), .Y(_14526_) );
AOI22X1 AOI22X1_605 ( .gnd(gnd), .vdd(vdd), .A(_130__14_), .B(_9449_), .C(_127__14_), .D(_9448_), .Y(_14527_) );
NAND3X1 NAND3X1_3059 ( .gnd(gnd), .vdd(vdd), .A(_14525_), .B(_14527_), .C(_14526_), .Y(_14528_) );
NOR3X1 NOR3X1_462 ( .gnd(gnd), .vdd(vdd), .A(_14516_), .B(_14524_), .C(_14528_), .Y(_14529_) );
AOI22X1 AOI22X1_606 ( .gnd(gnd), .vdd(vdd), .A(_110__14_), .B(_9453_), .C(_114__14_), .D(_9454_), .Y(_14530_) );
NAND3X1 NAND3X1_3060 ( .gnd(gnd), .vdd(vdd), .A(_14512_), .B(_14530_), .C(_14529_), .Y(_14531_) );
NOR2X1 NOR2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_14506_), .B(_14531_), .Y(_14532_) );
AOI22X1 AOI22X1_607 ( .gnd(gnd), .vdd(vdd), .A(_102__14_), .B(_9459_), .C(_103__14_), .D(_9457_), .Y(_14533_) );
NAND3X1 NAND3X1_3061 ( .gnd(gnd), .vdd(vdd), .A(_14503_), .B(_14533_), .C(_14532_), .Y(_14534_) );
NOR3X1 NOR3X1_463 ( .gnd(gnd), .vdd(vdd), .A(_14259_), .B(_14534_), .C(_14502_), .Y(_14535_) );
NAND3X1 NAND3X1_3062 ( .gnd(gnd), .vdd(vdd), .A(_14249_), .B(_14256_), .C(_14535_), .Y(_14536_) );
NOR3X1 NOR3X1_464 ( .gnd(gnd), .vdd(vdd), .A(_14238_), .B(_14241_), .C(_14536_), .Y(_14537_) );
NAND3X1 NAND3X1_3063 ( .gnd(gnd), .vdd(vdd), .A(_14229_), .B(_14234_), .C(_14537_), .Y(_14538_) );
NAND3X1 NAND3X1_3064 ( .gnd(gnd), .vdd(vdd), .A(_3082_), .B(_9473_), .C(_3083_), .Y(_14539_) );
NAND2X1 NAND2X1_2789 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__14_), .Y(_14540_) );
NAND2X1 NAND2X1_2790 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__14_), .Y(_14541_) );
NAND2X1 NAND2X1_2791 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__14_), .Y(_14542_) );
NAND3X1 NAND3X1_3065 ( .gnd(gnd), .vdd(vdd), .A(_2452_), .B(_9468_), .C(_2453_), .Y(_14543_) );
NAND3X1 NAND3X1_3066 ( .gnd(gnd), .vdd(vdd), .A(_14543_), .B(_14541_), .C(_14542_), .Y(_14544_) );
AOI21X1 AOI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_68__14_), .B(_9477_), .C(_14544_), .Y(_14545_) );
NAND3X1 NAND3X1_3067 ( .gnd(gnd), .vdd(vdd), .A(_14545_), .B(_14539_), .C(_14540_), .Y(_14546_) );
NOR3X1 NOR3X1_465 ( .gnd(gnd), .vdd(vdd), .A(_14228_), .B(_14546_), .C(_14538_), .Y(_14547_) );
AOI21X1 AOI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_14221_), .B(_14547_), .C(rst), .Y(_0__14_) );
NAND2X1 NAND2X1_2792 ( .gnd(gnd), .vdd(vdd), .A(_8736_), .B(_63__15_), .Y(_14548_) );
NAND2X1 NAND2X1_2793 ( .gnd(gnd), .vdd(vdd), .A(_8742_), .B(_59__15_), .Y(_14549_) );
NAND2X1 NAND2X1_2794 ( .gnd(gnd), .vdd(vdd), .A(_14548_), .B(_14549_), .Y(_14550_) );
NAND2X1 NAND2X1_2795 ( .gnd(gnd), .vdd(vdd), .A(_8750_), .B(_58__15_), .Y(_14551_) );
NAND2X1 NAND2X1_2796 ( .gnd(gnd), .vdd(vdd), .A(_8757_), .B(_60__15_), .Y(_14552_) );
NAND2X1 NAND2X1_2797 ( .gnd(gnd), .vdd(vdd), .A(_14551_), .B(_14552_), .Y(_14553_) );
NOR2X1 NOR2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_14550_), .B(_14553_), .Y(_14554_) );
NAND3X1 NAND3X1_3068 ( .gnd(gnd), .vdd(vdd), .A(_3302_), .B(_8762_), .C(_3301_), .Y(_14555_) );
NAND3X1 NAND3X1_3069 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_8765_), .C(_3249_), .Y(_14556_) );
AND2X2 AND2X2_1614 ( .gnd(gnd), .vdd(vdd), .A(_14556_), .B(_14555_), .Y(_14557_) );
AOI22X1 AOI22X1_608 ( .gnd(gnd), .vdd(vdd), .A(_62__15_), .B(_8774_), .C(_57__15_), .D(_8771_), .Y(_14558_) );
NAND2X1 NAND2X1_2798 ( .gnd(gnd), .vdd(vdd), .A(_14557_), .B(_14558_), .Y(_14559_) );
NAND2X1 NAND2X1_2799 ( .gnd(gnd), .vdd(vdd), .A(_8779_), .B(_64__15_), .Y(_14560_) );
NAND3X1 NAND3X1_3070 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .B(_8794_), .C(_2669_), .Y(_14561_) );
OAI21X1 OAI21X1_2579 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .B(_8792_), .C(_14561_), .Y(_14562_) );
NAND3X1 NAND3X1_3071 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(_8786_), .C(_2840_), .Y(_14563_) );
OAI21X1 OAI21X1_2580 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_8799_), .C(_14563_), .Y(_14564_) );
NOR2X1 NOR2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_14562_), .B(_14564_), .Y(_14565_) );
AOI22X1 AOI22X1_609 ( .gnd(gnd), .vdd(vdd), .A(_73__15_), .B(_9480_), .C(_74__15_), .D(_8803_), .Y(_14566_) );
AOI22X1 AOI22X1_610 ( .gnd(gnd), .vdd(vdd), .A(_76__15_), .B(_9482_), .C(_81__15_), .D(_9468_), .Y(_14567_) );
NAND2X1 NAND2X1_2800 ( .gnd(gnd), .vdd(vdd), .A(_14567_), .B(_14566_), .Y(_14568_) );
NOR2X1 NOR2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_8812_), .B(_2336_), .Y(_14569_) );
NOR2X1 NOR2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_8818_), .B(_2312_), .Y(_14570_) );
NAND2X1 NAND2X1_2801 ( .gnd(gnd), .vdd(vdd), .A(_8821_), .B(_96__15_), .Y(_14571_) );
NAND3X1 NAND3X1_3072 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .B(_8843_), .C(_2028_), .Y(_14572_) );
NAND3X1 NAND3X1_3073 ( .gnd(gnd), .vdd(vdd), .A(_8825_), .B(_1937_), .C(_1938_), .Y(_14573_) );
NAND3X1 NAND3X1_3074 ( .gnd(gnd), .vdd(vdd), .A(_14573_), .B(_14572_), .C(_14571_), .Y(_14574_) );
NOR3X1 NOR3X1_466 ( .gnd(gnd), .vdd(vdd), .A(_14569_), .B(_14574_), .C(_14570_), .Y(_14575_) );
NAND3X1 NAND3X1_3075 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_8829_), .C(_2276_), .Y(_14576_) );
NAND3X1 NAND3X1_3076 ( .gnd(gnd), .vdd(vdd), .A(_2169_), .B(_8831_), .C(_2170_), .Y(_14577_) );
NAND2X1 NAND2X1_2802 ( .gnd(gnd), .vdd(vdd), .A(_14576_), .B(_14577_), .Y(_14578_) );
NAND3X1 NAND3X1_3077 ( .gnd(gnd), .vdd(vdd), .A(_2110_), .B(_8834_), .C(_2109_), .Y(_14579_) );
NAND3X1 NAND3X1_3078 ( .gnd(gnd), .vdd(vdd), .A(_2221_), .B(_8836_), .C(_2222_), .Y(_14580_) );
NAND2X1 NAND2X1_2803 ( .gnd(gnd), .vdd(vdd), .A(_14580_), .B(_14579_), .Y(_14581_) );
NOR2X1 NOR2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_14578_), .B(_14581_), .Y(_14582_) );
AOI22X1 AOI22X1_611 ( .gnd(gnd), .vdd(vdd), .A(_98__15_), .B(_8845_), .C(_93__15_), .D(_8840_), .Y(_14583_) );
AOI22X1 AOI22X1_612 ( .gnd(gnd), .vdd(vdd), .A(_94__15_), .B(_8841_), .C(_91__15_), .D(_8823_), .Y(_14584_) );
NAND2X1 NAND2X1_2804 ( .gnd(gnd), .vdd(vdd), .A(_14583_), .B(_14584_), .Y(_14585_) );
NAND2X1 NAND2X1_2805 ( .gnd(gnd), .vdd(vdd), .A(_8848_), .B(_99__15_), .Y(_14586_) );
NAND2X1 NAND2X1_2806 ( .gnd(gnd), .vdd(vdd), .A(_9390_), .B(_107__15_), .Y(_14587_) );
NAND2X1 NAND2X1_2807 ( .gnd(gnd), .vdd(vdd), .A(_9392_), .B(_105__15_), .Y(_14588_) );
NAND2X1 NAND2X1_2808 ( .gnd(gnd), .vdd(vdd), .A(_14587_), .B(_14588_), .Y(_14589_) );
NAND2X1 NAND2X1_2809 ( .gnd(gnd), .vdd(vdd), .A(_8860_), .B(_104__15_), .Y(_14590_) );
NAND2X1 NAND2X1_2810 ( .gnd(gnd), .vdd(vdd), .A(_8857_), .B(_113__15_), .Y(_14591_) );
NAND2X1 NAND2X1_2811 ( .gnd(gnd), .vdd(vdd), .A(_14590_), .B(_14591_), .Y(_14592_) );
NOR2X1 NOR2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_14589_), .B(_14592_), .Y(_14593_) );
NAND2X1 NAND2X1_2812 ( .gnd(gnd), .vdd(vdd), .A(_8866_), .B(_118__15_), .Y(_14594_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_7163_), .B(_9930_), .C(_7207_), .D(_9929_), .Y(_14595_) );
NOR2X1 NOR2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_9932_), .B(_7342_), .Y(_14596_) );
NOR2X1 NOR2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_9934_), .B(_7299_), .Y(_14597_) );
NOR3X1 NOR3X1_467 ( .gnd(gnd), .vdd(vdd), .A(_14596_), .B(_14597_), .C(_14595_), .Y(_14598_) );
NAND2X1 NAND2X1_2813 ( .gnd(gnd), .vdd(vdd), .A(_8879_), .B(_188__15_), .Y(_14599_) );
NAND2X1 NAND2X1_2814 ( .gnd(gnd), .vdd(vdd), .A(_8881_), .B(_126__15_), .Y(_14600_) );
NAND2X1 NAND2X1_2815 ( .gnd(gnd), .vdd(vdd), .A(_14599_), .B(_14600_), .Y(_14601_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_7385_), .B(_9940_), .C(_7253_), .D(_9941_), .Y(_14602_) );
NOR2X1 NOR2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_14602_), .B(_14601_), .Y(_14603_) );
NAND3X1 NAND3X1_3079 ( .gnd(gnd), .vdd(vdd), .A(_14594_), .B(_14598_), .C(_14603_), .Y(_14604_) );
AOI22X1 AOI22X1_613 ( .gnd(gnd), .vdd(vdd), .A(_20__15_), .B(_8898_), .C(_250__15_), .D(_9082_), .Y(_14605_) );
AOI22X1 AOI22X1_614 ( .gnd(gnd), .vdd(vdd), .A(_243__15_), .B(_9153_), .C(_175__15_), .D(_8904_), .Y(_14606_) );
NAND2X1 NAND2X1_2816 ( .gnd(gnd), .vdd(vdd), .A(_14605_), .B(_14606_), .Y(_14607_) );
NAND2X1 NAND2X1_2817 ( .gnd(gnd), .vdd(vdd), .A(_8909_), .B(_36__15_), .Y(_14608_) );
NAND2X1 NAND2X1_2818 ( .gnd(gnd), .vdd(vdd), .A(_8911_), .B(_41__15_), .Y(_14609_) );
AOI22X1 AOI22X1_615 ( .gnd(gnd), .vdd(vdd), .A(_19__15_), .B(_8914_), .C(_210__15_), .D(_8918_), .Y(_14610_) );
NAND3X1 NAND3X1_3080 ( .gnd(gnd), .vdd(vdd), .A(_14608_), .B(_14609_), .C(_14610_), .Y(_14611_) );
NOR2X1 NOR2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_14607_), .B(_14611_), .Y(_14612_) );
AOI22X1 AOI22X1_616 ( .gnd(gnd), .vdd(vdd), .A(_134__15_), .B(_8933_), .C(_9__15_), .D(_8926_), .Y(_14613_) );
NAND2X1 NAND2X1_2819 ( .gnd(gnd), .vdd(vdd), .A(_8931_), .B(_24__15_), .Y(_14614_) );
NAND2X1 NAND2X1_2820 ( .gnd(gnd), .vdd(vdd), .A(_9177_), .B(_145__15_), .Y(_14615_) );
NAND3X1 NAND3X1_3081 ( .gnd(gnd), .vdd(vdd), .A(_14614_), .B(_14615_), .C(_14613_), .Y(_14616_) );
AOI22X1 AOI22X1_617 ( .gnd(gnd), .vdd(vdd), .A(_4__15_), .B(_8937_), .C(_176__15_), .D(_8939_), .Y(_14617_) );
NAND2X1 NAND2X1_2821 ( .gnd(gnd), .vdd(vdd), .A(_8942_), .B(_5__15_), .Y(_14618_) );
NAND2X1 NAND2X1_2822 ( .gnd(gnd), .vdd(vdd), .A(_8944_), .B(_8__15_), .Y(_14619_) );
NAND3X1 NAND3X1_3082 ( .gnd(gnd), .vdd(vdd), .A(_14618_), .B(_14619_), .C(_14617_), .Y(_14620_) );
NOR2X1 NOR2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_14620_), .B(_14616_), .Y(_14621_) );
NAND2X1 NAND2X1_2823 ( .gnd(gnd), .vdd(vdd), .A(_14612_), .B(_14621_), .Y(_14622_) );
AOI22X1 AOI22X1_618 ( .gnd(gnd), .vdd(vdd), .A(_47__15_), .B(_9161_), .C(_238__15_), .D(_8893_), .Y(_14623_) );
NAND2X1 NAND2X1_2824 ( .gnd(gnd), .vdd(vdd), .A(_9150_), .B(_21__15_), .Y(_14624_) );
NAND2X1 NAND2X1_2825 ( .gnd(gnd), .vdd(vdd), .A(_9151_), .B(_185__15_), .Y(_14625_) );
NAND3X1 NAND3X1_3083 ( .gnd(gnd), .vdd(vdd), .A(_14624_), .B(_14625_), .C(_14623_), .Y(_14626_) );
AOI22X1 AOI22X1_619 ( .gnd(gnd), .vdd(vdd), .A(_246__15_), .B(_9356_), .C(_226__15_), .D(_9357_), .Y(_14627_) );
NAND2X1 NAND2X1_2826 ( .gnd(gnd), .vdd(vdd), .A(_9157_), .B(_231__15_), .Y(_14628_) );
NAND2X1 NAND2X1_2827 ( .gnd(gnd), .vdd(vdd), .A(_9158_), .B(_46__15_), .Y(_14629_) );
NAND3X1 NAND3X1_3084 ( .gnd(gnd), .vdd(vdd), .A(_14628_), .B(_14629_), .C(_14627_), .Y(_14630_) );
NOR2X1 NOR2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_14626_), .B(_14630_), .Y(_14631_) );
NAND2X1 NAND2X1_2828 ( .gnd(gnd), .vdd(vdd), .A(_9173_), .B(_178__15_), .Y(_14632_) );
NAND2X1 NAND2X1_2829 ( .gnd(gnd), .vdd(vdd), .A(_8975_), .B(_52__15_), .Y(_14633_) );
AOI22X1 AOI22X1_620 ( .gnd(gnd), .vdd(vdd), .A(_37__15_), .B(_8978_), .C(_35__15_), .D(_8980_), .Y(_14634_) );
NAND3X1 NAND3X1_3085 ( .gnd(gnd), .vdd(vdd), .A(_14632_), .B(_14633_), .C(_14634_), .Y(_14635_) );
AOI22X1 AOI22X1_621 ( .gnd(gnd), .vdd(vdd), .A(_237__15_), .B(_8966_), .C(_253__15_), .D(_9154_), .Y(_14636_) );
NAND2X1 NAND2X1_2830 ( .gnd(gnd), .vdd(vdd), .A(_8928_), .B(_123__15_), .Y(_14637_) );
NAND2X1 NAND2X1_2831 ( .gnd(gnd), .vdd(vdd), .A(_8989_), .B(_213__15_), .Y(_14638_) );
NAND3X1 NAND3X1_3086 ( .gnd(gnd), .vdd(vdd), .A(_14637_), .B(_14638_), .C(_14636_), .Y(_14639_) );
NOR2X1 NOR2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_14635_), .B(_14639_), .Y(_14640_) );
NAND2X1 NAND2X1_2832 ( .gnd(gnd), .vdd(vdd), .A(_14631_), .B(_14640_), .Y(_14641_) );
NOR2X1 NOR2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_14622_), .B(_14641_), .Y(_14642_) );
NAND2X1 NAND2X1_2833 ( .gnd(gnd), .vdd(vdd), .A(_8998_), .B(_11__15_), .Y(_14643_) );
NAND2X1 NAND2X1_2834 ( .gnd(gnd), .vdd(vdd), .A(_9002_), .B(_215__15_), .Y(_14644_) );
AOI22X1 AOI22X1_622 ( .gnd(gnd), .vdd(vdd), .A(_13__15_), .B(_9007_), .C(_239__15_), .D(_9076_), .Y(_14645_) );
NAND3X1 NAND3X1_3087 ( .gnd(gnd), .vdd(vdd), .A(_14643_), .B(_14644_), .C(_14645_), .Y(_14646_) );
AOI22X1 AOI22X1_623 ( .gnd(gnd), .vdd(vdd), .A(_206__15_), .B(_9013_), .C(_242__15_), .D(_9035_), .Y(_14647_) );
NAND2X1 NAND2X1_2835 ( .gnd(gnd), .vdd(vdd), .A(_9016_), .B(_207__15_), .Y(_14648_) );
NAND2X1 NAND2X1_2836 ( .gnd(gnd), .vdd(vdd), .A(_9174_), .B(_214__15_), .Y(_14649_) );
NAND3X1 NAND3X1_3088 ( .gnd(gnd), .vdd(vdd), .A(_14648_), .B(_14649_), .C(_14647_), .Y(_14650_) );
NOR2X1 NOR2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_14646_), .B(_14650_), .Y(_14651_) );
AOI22X1 AOI22X1_624 ( .gnd(gnd), .vdd(vdd), .A(_222__15_), .B(_9024_), .C(_220__15_), .D(_9026_), .Y(_14652_) );
NAND2X1 NAND2X1_2837 ( .gnd(gnd), .vdd(vdd), .A(_9029_), .B(_230__15_), .Y(_14653_) );
NAND2X1 NAND2X1_2838 ( .gnd(gnd), .vdd(vdd), .A(_9031_), .B(_228__15_), .Y(_14654_) );
NAND3X1 NAND3X1_3089 ( .gnd(gnd), .vdd(vdd), .A(_14653_), .B(_14654_), .C(_14652_), .Y(_14655_) );
AOI22X1 AOI22X1_625 ( .gnd(gnd), .vdd(vdd), .A(_18__15_), .B(_9037_), .C(_240__15_), .D(_9011_), .Y(_14656_) );
NAND2X1 NAND2X1_2839 ( .gnd(gnd), .vdd(vdd), .A(_9061_), .B(_26__15_), .Y(_14657_) );
NAND2X1 NAND2X1_2840 ( .gnd(gnd), .vdd(vdd), .A(_9042_), .B(_28__15_), .Y(_14658_) );
NAND3X1 NAND3X1_3090 ( .gnd(gnd), .vdd(vdd), .A(_14657_), .B(_14658_), .C(_14656_), .Y(_14659_) );
NOR2X1 NOR2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_14655_), .B(_14659_), .Y(_14660_) );
NAND2X1 NAND2X1_2841 ( .gnd(gnd), .vdd(vdd), .A(_14651_), .B(_14660_), .Y(_14661_) );
AOI22X1 AOI22X1_626 ( .gnd(gnd), .vdd(vdd), .A(_225__15_), .B(_9048_), .C(_167__15_), .D(_9050_), .Y(_14662_) );
NAND2X1 NAND2X1_2842 ( .gnd(gnd), .vdd(vdd), .A(_8955_), .B(_236__15_), .Y(_14663_) );
NAND2X1 NAND2X1_2843 ( .gnd(gnd), .vdd(vdd), .A(_9055_), .B(_174__15_), .Y(_14664_) );
NAND3X1 NAND3X1_3091 ( .gnd(gnd), .vdd(vdd), .A(_14663_), .B(_14664_), .C(_14662_), .Y(_14665_) );
NAND2X1 NAND2X1_2844 ( .gnd(gnd), .vdd(vdd), .A(_9059_), .B(_25__15_), .Y(_14666_) );
NAND2X1 NAND2X1_2845 ( .gnd(gnd), .vdd(vdd), .A(_9066_), .B(_27__15_), .Y(_14667_) );
AOI22X1 AOI22X1_627 ( .gnd(gnd), .vdd(vdd), .A(_224__15_), .B(_9064_), .C(_221__15_), .D(_9040_), .Y(_14668_) );
NAND3X1 NAND3X1_3092 ( .gnd(gnd), .vdd(vdd), .A(_14666_), .B(_14667_), .C(_14668_), .Y(_14669_) );
NOR2X1 NOR2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_14665_), .B(_14669_), .Y(_14670_) );
AOI22X1 AOI22X1_628 ( .gnd(gnd), .vdd(vdd), .A(_184__15_), .B(_9073_), .C(_183__15_), .D(_9071_), .Y(_14671_) );
NAND2X1 NAND2X1_2846 ( .gnd(gnd), .vdd(vdd), .A(_9005_), .B(_241__15_), .Y(_14672_) );
NAND2X1 NAND2X1_2847 ( .gnd(gnd), .vdd(vdd), .A(_9078_), .B(_51__15_), .Y(_14673_) );
NAND3X1 NAND3X1_3093 ( .gnd(gnd), .vdd(vdd), .A(_14672_), .B(_14673_), .C(_14671_), .Y(_14674_) );
AOI22X1 AOI22X1_629 ( .gnd(gnd), .vdd(vdd), .A(_43__15_), .B(_9084_), .C(_248__15_), .D(_8901_), .Y(_14675_) );
NAND2X1 NAND2X1_2848 ( .gnd(gnd), .vdd(vdd), .A(_9087_), .B(_211__15_), .Y(_14676_) );
NAND2X1 NAND2X1_2849 ( .gnd(gnd), .vdd(vdd), .A(_9089_), .B(_48__15_), .Y(_14677_) );
NAND3X1 NAND3X1_3094 ( .gnd(gnd), .vdd(vdd), .A(_14676_), .B(_14677_), .C(_14675_), .Y(_14678_) );
NOR2X1 NOR2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_14674_), .B(_14678_), .Y(_14679_) );
NAND2X1 NAND2X1_2850 ( .gnd(gnd), .vdd(vdd), .A(_14670_), .B(_14679_), .Y(_14680_) );
NOR2X1 NOR2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_14661_), .B(_14680_), .Y(_14681_) );
NAND3X1 NAND3X1_3095 ( .gnd(gnd), .vdd(vdd), .A(_6836_), .B(_9143_), .C(_6837_), .Y(_14682_) );
NAND3X1 NAND3X1_3096 ( .gnd(gnd), .vdd(vdd), .A(_6988_), .B(_9145_), .C(_6989_), .Y(_14683_) );
NAND2X1 NAND2X1_2851 ( .gnd(gnd), .vdd(vdd), .A(_14682_), .B(_14683_), .Y(_14684_) );
NAND3X1 NAND3X1_3097 ( .gnd(gnd), .vdd(vdd), .A(_5072_), .B(_9135_), .C(_5073_), .Y(_14685_) );
NAND3X1 NAND3X1_3098 ( .gnd(gnd), .vdd(vdd), .A(_6954_), .B(_9137_), .C(_6955_), .Y(_14686_) );
NAND2X1 NAND2X1_2852 ( .gnd(gnd), .vdd(vdd), .A(_14686_), .B(_14685_), .Y(_14687_) );
NOR2X1 NOR2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_14684_), .B(_14687_), .Y(_14688_) );
NAND3X1 NAND3X1_3099 ( .gnd(gnd), .vdd(vdd), .A(_8336_), .B(_9188_), .C(_8337_), .Y(_14689_) );
NAND3X1 NAND3X1_3100 ( .gnd(gnd), .vdd(vdd), .A(_15947_), .B(_9109_), .C(_15948_), .Y(_14690_) );
NAND3X1 NAND3X1_3101 ( .gnd(gnd), .vdd(vdd), .A(_16152_), .B(_9115_), .C(_16153_), .Y(_14691_) );
NAND3X1 NAND3X1_3102 ( .gnd(gnd), .vdd(vdd), .A(_14690_), .B(_14691_), .C(_14689_), .Y(_14692_) );
AOI22X1 AOI22X1_630 ( .gnd(gnd), .vdd(vdd), .A(_234__15_), .B(_9182_), .C(_34__15_), .D(_9183_), .Y(_14693_) );
AOI22X1 AOI22X1_631 ( .gnd(gnd), .vdd(vdd), .A(_100__15_), .B(_9346_), .C(_45__15_), .D(_9185_), .Y(_14694_) );
NAND2X1 NAND2X1_2853 ( .gnd(gnd), .vdd(vdd), .A(_14694_), .B(_14693_), .Y(_14695_) );
NAND3X1 NAND3X1_3103 ( .gnd(gnd), .vdd(vdd), .A(_4720_), .B(_9140_), .C(_4719_), .Y(_14696_) );
OAI21X1 OAI21X1_2581 ( .gnd(gnd), .vdd(vdd), .A(_5258_), .B(_10036_), .C(_14696_), .Y(_14697_) );
NOR3X1 NOR3X1_468 ( .gnd(gnd), .vdd(vdd), .A(_14697_), .B(_14692_), .C(_14695_), .Y(_14698_) );
NAND3X1 NAND3X1_3104 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_9133_), .C(_3447_), .Y(_14699_) );
NAND3X1 NAND3X1_3105 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(_9097_), .C(_4945_), .Y(_14700_) );
NAND3X1 NAND3X1_3106 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .B(_9102_), .C(_5119_), .Y(_14701_) );
NAND3X1 NAND3X1_3107 ( .gnd(gnd), .vdd(vdd), .A(_14700_), .B(_14701_), .C(_14699_), .Y(_14702_) );
AOI22X1 AOI22X1_632 ( .gnd(gnd), .vdd(vdd), .A(_38__15_), .B(_9129_), .C(_16__15_), .D(_9127_), .Y(_14703_) );
AOI22X1 AOI22X1_633 ( .gnd(gnd), .vdd(vdd), .A(_39__15_), .B(_9099_), .C(_204__15_), .D(_9104_), .Y(_14704_) );
NAND2X1 NAND2X1_2854 ( .gnd(gnd), .vdd(vdd), .A(_14703_), .B(_14704_), .Y(_14705_) );
NOR2X1 NOR2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_14702_), .B(_14705_), .Y(_14706_) );
NAND3X1 NAND3X1_3108 ( .gnd(gnd), .vdd(vdd), .A(_14688_), .B(_14698_), .C(_14706_), .Y(_14707_) );
AOI22X1 AOI22X1_634 ( .gnd(gnd), .vdd(vdd), .A(_227__15_), .B(_9170_), .C(_30__15_), .D(_9167_), .Y(_14708_) );
AOI22X1 AOI22X1_635 ( .gnd(gnd), .vdd(vdd), .A(_209__15_), .B(_8957_), .C(_33__15_), .D(_8991_), .Y(_14709_) );
NAND2X1 NAND2X1_2855 ( .gnd(gnd), .vdd(vdd), .A(_14708_), .B(_14709_), .Y(_14710_) );
AOI22X1 AOI22X1_636 ( .gnd(gnd), .vdd(vdd), .A(_44__15_), .B(_8968_), .C(_42__15_), .D(_8963_), .Y(_14711_) );
AOI22X1 AOI22X1_637 ( .gnd(gnd), .vdd(vdd), .A(_249__15_), .B(_9053_), .C(_208__15_), .D(_8950_), .Y(_14712_) );
NAND2X1 NAND2X1_2856 ( .gnd(gnd), .vdd(vdd), .A(_14711_), .B(_14712_), .Y(_14713_) );
NOR2X1 NOR2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_14710_), .B(_14713_), .Y(_14714_) );
AOI22X1 AOI22X1_638 ( .gnd(gnd), .vdd(vdd), .A(_22__15_), .B(_9382_), .C(_3__15_), .D(_9383_), .Y(_14715_) );
NAND2X1 NAND2X1_2857 ( .gnd(gnd), .vdd(vdd), .A(_9353_), .B(_219__15_), .Y(_14716_) );
NAND2X1 NAND2X1_2858 ( .gnd(gnd), .vdd(vdd), .A(_9354_), .B(_232__15_), .Y(_14717_) );
NAND3X1 NAND3X1_3109 ( .gnd(gnd), .vdd(vdd), .A(_14716_), .B(_14717_), .C(_14715_), .Y(_14718_) );
AOI22X1 AOI22X1_639 ( .gnd(gnd), .vdd(vdd), .A(_255__15_), .B(_8986_), .C(_254__15_), .D(_8984_), .Y(_14719_) );
AOI22X1 AOI22X1_640 ( .gnd(gnd), .vdd(vdd), .A(_203__15_), .B(_9018_), .C(_156__15_), .D(_8973_), .Y(_14720_) );
NAND2X1 NAND2X1_2859 ( .gnd(gnd), .vdd(vdd), .A(_14719_), .B(_14720_), .Y(_14721_) );
NOR2X1 NOR2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_14718_), .B(_14721_), .Y(_14722_) );
NAND2X1 NAND2X1_2860 ( .gnd(gnd), .vdd(vdd), .A(_14714_), .B(_14722_), .Y(_14723_) );
AOI22X1 AOI22X1_641 ( .gnd(gnd), .vdd(vdd), .A(_201__15_), .B(_9124_), .C(_212__15_), .D(_9345_), .Y(_14724_) );
NAND3X1 NAND3X1_3110 ( .gnd(gnd), .vdd(vdd), .A(_8450_), .B(_9348_), .C(_8449_), .Y(_14725_) );
NAND3X1 NAND3X1_3111 ( .gnd(gnd), .vdd(vdd), .A(_9349_), .B(_510_), .C(_511_), .Y(_14726_) );
AND2X2 AND2X2_1615 ( .gnd(gnd), .vdd(vdd), .A(_14726_), .B(_14725_), .Y(_14727_) );
NAND2X1 NAND2X1_2861 ( .gnd(gnd), .vdd(vdd), .A(_14724_), .B(_14727_), .Y(_14728_) );
NAND3X1 NAND3X1_3112 ( .gnd(gnd), .vdd(vdd), .A(_15156_), .B(_9208_), .C(_15157_), .Y(_14729_) );
OAI21X1 OAI21X1_2582 ( .gnd(gnd), .vdd(vdd), .A(_15118_), .B(_9211_), .C(_14729_), .Y(_14730_) );
NAND3X1 NAND3X1_3113 ( .gnd(gnd), .vdd(vdd), .A(_15504_), .B(_9222_), .C(_15505_), .Y(_14731_) );
NAND3X1 NAND3X1_3114 ( .gnd(gnd), .vdd(vdd), .A(_15451_), .B(_9224_), .C(_15450_), .Y(_14732_) );
NAND2X1 NAND2X1_2862 ( .gnd(gnd), .vdd(vdd), .A(_14731_), .B(_14732_), .Y(_14733_) );
NOR2X1 NOR2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_14733_), .B(_14730_), .Y(_14734_) );
NAND3X1 NAND3X1_3115 ( .gnd(gnd), .vdd(vdd), .A(_15282_), .B(_9217_), .C(_15283_), .Y(_14735_) );
NAND3X1 NAND3X1_3116 ( .gnd(gnd), .vdd(vdd), .A(_15230_), .B(_9219_), .C(_15229_), .Y(_14736_) );
NAND2X1 NAND2X1_2863 ( .gnd(gnd), .vdd(vdd), .A(_14736_), .B(_14735_), .Y(_14737_) );
NAND3X1 NAND3X1_3117 ( .gnd(gnd), .vdd(vdd), .A(_15680_), .B(_9192_), .C(_15681_), .Y(_14738_) );
NAND3X1 NAND3X1_3118 ( .gnd(gnd), .vdd(vdd), .A(_15737_), .B(_9199_), .C(_15736_), .Y(_14739_) );
NAND2X1 NAND2X1_2864 ( .gnd(gnd), .vdd(vdd), .A(_14739_), .B(_14738_), .Y(_14740_) );
NOR2X1 NOR2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_14740_), .B(_14737_), .Y(_14741_) );
NOR3X1 NOR3X1_469 ( .gnd(gnd), .vdd(vdd), .A(_16202_), .B(_10083_), .C(_16203_), .Y(_14742_) );
NAND3X1 NAND3X1_3119 ( .gnd(gnd), .vdd(vdd), .A(_15330_), .B(_9205_), .C(_15331_), .Y(_14743_) );
OAI21X1 OAI21X1_2583 ( .gnd(gnd), .vdd(vdd), .A(_15358_), .B(_10085_), .C(_14743_), .Y(_14744_) );
NAND3X1 NAND3X1_3120 ( .gnd(gnd), .vdd(vdd), .A(_15562_), .B(_9233_), .C(_15563_), .Y(_14745_) );
NAND3X1 NAND3X1_3121 ( .gnd(gnd), .vdd(vdd), .A(_9194_), .B(_15628_), .C(_15627_), .Y(_14746_) );
NAND2X1 NAND2X1_2865 ( .gnd(gnd), .vdd(vdd), .A(_14745_), .B(_14746_), .Y(_14747_) );
NOR3X1 NOR3X1_470 ( .gnd(gnd), .vdd(vdd), .A(_14744_), .B(_14747_), .C(_14742_), .Y(_14748_) );
NAND3X1 NAND3X1_3122 ( .gnd(gnd), .vdd(vdd), .A(_14734_), .B(_14741_), .C(_14748_), .Y(_14749_) );
NAND3X1 NAND3X1_3123 ( .gnd(gnd), .vdd(vdd), .A(_15890_), .B(_9120_), .C(_15891_), .Y(_14750_) );
NAND3X1 NAND3X1_3124 ( .gnd(gnd), .vdd(vdd), .A(_15397_), .B(_9197_), .C(_15396_), .Y(_14751_) );
NOR2X1 NOR2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_9288_), .B(_7021_), .Y(_14752_) );
NOR2X1 NOR2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_9301_), .B(_7653_), .Y(_14753_) );
NOR3X1 NOR3X1_471 ( .gnd(gnd), .vdd(vdd), .A(_15828_), .B(_11264_), .C(_15827_), .Y(_14754_) );
NOR3X1 NOR3X1_472 ( .gnd(gnd), .vdd(vdd), .A(_14752_), .B(_14753_), .C(_14754_), .Y(_14755_) );
NAND3X1 NAND3X1_3125 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_9255_), .C(_1783_), .Y(_14756_) );
OAI21X1 OAI21X1_2584 ( .gnd(gnd), .vdd(vdd), .A(_9765_), .B(_8725_), .C(_14756_), .Y(_14757_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_8185_), .B(_9304_), .C(_4201_), .D(_9254_), .Y(_14758_) );
NOR2X1 NOR2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_14758_), .B(_14757_), .Y(_14759_) );
NAND3X1 NAND3X1_3126 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_9262_), .C(_629_), .Y(_14760_) );
OAI21X1 OAI21X1_2585 ( .gnd(gnd), .vdd(vdd), .A(_2932_), .B(_10468_), .C(_14760_), .Y(_14761_) );
NOR3X1 NOR3X1_473 ( .gnd(gnd), .vdd(vdd), .A(_7481_), .B(_10471_), .C(_7482_), .Y(_14762_) );
NOR3X1 NOR3X1_474 ( .gnd(gnd), .vdd(vdd), .A(_7113_), .B(_9245_), .C(_7112_), .Y(_14763_) );
NOR3X1 NOR3X1_475 ( .gnd(gnd), .vdd(vdd), .A(_14761_), .B(_14763_), .C(_14762_), .Y(_14764_) );
NAND3X1 NAND3X1_3127 ( .gnd(gnd), .vdd(vdd), .A(_14755_), .B(_14759_), .C(_14764_), .Y(_14765_) );
NAND3X1 NAND3X1_3128 ( .gnd(gnd), .vdd(vdd), .A(_6448_), .B(_9281_), .C(_6449_), .Y(_14766_) );
NAND3X1 NAND3X1_3129 ( .gnd(gnd), .vdd(vdd), .A(_7739_), .B(_9248_), .C(_7738_), .Y(_14767_) );
NAND3X1 NAND3X1_3130 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(_9268_), .C(_1190_), .Y(_14768_) );
NAND3X1 NAND3X1_3131 ( .gnd(gnd), .vdd(vdd), .A(_14767_), .B(_14768_), .C(_14766_), .Y(_14769_) );
NOR2X1 NOR2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_9323_), .B(_5940_), .Y(_14770_) );
NOR2X1 NOR2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_9273_), .B(_4835_), .Y(_14771_) );
NOR3X1 NOR3X1_476 ( .gnd(gnd), .vdd(vdd), .A(_14770_), .B(_14771_), .C(_14769_), .Y(_14772_) );
NAND3X1 NAND3X1_3132 ( .gnd(gnd), .vdd(vdd), .A(_7068_), .B(_9266_), .C(_7069_), .Y(_14773_) );
OAI21X1 OAI21X1_2586 ( .gnd(gnd), .vdd(vdd), .A(_8256_), .B(_10875_), .C(_14773_), .Y(_14774_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_7505_), .B(_11613_), .C(_3577_), .D(_9306_), .Y(_14775_) );
NOR2X1 NOR2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_14775_), .B(_14774_), .Y(_14776_) );
NAND2X1 NAND2X1_2866 ( .gnd(gnd), .vdd(vdd), .A(_9286_), .B(_67__15_), .Y(_14777_) );
OAI21X1 OAI21X1_2587 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .B(_9295_), .C(_14777_), .Y(_14778_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_6481_), .B(_9259_), .C(_14931_), .D(_9276_), .Y(_14779_) );
NOR2X1 NOR2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_14779_), .B(_14778_), .Y(_14780_) );
NAND3X1 NAND3X1_3133 ( .gnd(gnd), .vdd(vdd), .A(_14772_), .B(_14780_), .C(_14776_), .Y(_14781_) );
NOR3X1 NOR3X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2374_), .B(_14440_), .C(_2373_), .Y(_14782_) );
NOR3X1 NOR3X1_478 ( .gnd(gnd), .vdd(vdd), .A(_4796_), .B(_9312_), .C(_4795_), .Y(_14783_) );
NOR2X1 NOR2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_9282_), .B(_4241_), .Y(_14784_) );
NOR3X1 NOR3X1_479 ( .gnd(gnd), .vdd(vdd), .A(_14783_), .B(_14784_), .C(_14782_), .Y(_14785_) );
AOI22X1 AOI22X1_642 ( .gnd(gnd), .vdd(vdd), .A(_181__15_), .B(_9321_), .C(_252__15_), .D(_9326_), .Y(_14786_) );
AOI22X1 AOI22X1_643 ( .gnd(gnd), .vdd(vdd), .A(_251__15_), .B(_9320_), .C(_233__15_), .D(_9310_), .Y(_14787_) );
NAND3X1 NAND3X1_3134 ( .gnd(gnd), .vdd(vdd), .A(_14786_), .B(_14787_), .C(_14785_), .Y(_14788_) );
NOR3X1 NOR3X1_480 ( .gnd(gnd), .vdd(vdd), .A(_14765_), .B(_14788_), .C(_14781_), .Y(_14789_) );
NAND2X1 NAND2X1_2867 ( .gnd(gnd), .vdd(vdd), .A(_14751_), .B(_14789_), .Y(_14790_) );
AOI21X1 AOI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_157__15_), .B(_9232_), .C(_14790_), .Y(_14791_) );
AOI22X1 AOI22X1_644 ( .gnd(gnd), .vdd(vdd), .A(_155__15_), .B(_9333_), .C(_172__15_), .D(_9332_), .Y(_14792_) );
NAND3X1 NAND3X1_3135 ( .gnd(gnd), .vdd(vdd), .A(_14750_), .B(_14792_), .C(_14791_), .Y(_14793_) );
NOR3X1 NOR3X1_481 ( .gnd(gnd), .vdd(vdd), .A(_14749_), .B(_14793_), .C(_14728_), .Y(_14794_) );
AOI22X1 AOI22X1_645 ( .gnd(gnd), .vdd(vdd), .A(_256__15_), .B(_9113_), .C(_142__15_), .D(_9118_), .Y(_14795_) );
NAND2X1 NAND2X1_2868 ( .gnd(gnd), .vdd(vdd), .A(_9123_), .B(_89__15_), .Y(_14796_) );
NAND2X1 NAND2X1_2869 ( .gnd(gnd), .vdd(vdd), .A(_9229_), .B(_223__15_), .Y(_14797_) );
NAND3X1 NAND3X1_3136 ( .gnd(gnd), .vdd(vdd), .A(_14796_), .B(_14797_), .C(_14795_), .Y(_14798_) );
NAND2X1 NAND2X1_2870 ( .gnd(gnd), .vdd(vdd), .A(_9337_), .B(_143__15_), .Y(_14799_) );
NAND3X1 NAND3X1_3137 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_9339_), .C(_473_), .Y(_14800_) );
AOI22X1 AOI22X1_646 ( .gnd(gnd), .vdd(vdd), .A(_111__15_), .B(_9342_), .C(_12__15_), .D(_9341_), .Y(_14801_) );
NAND3X1 NAND3X1_3138 ( .gnd(gnd), .vdd(vdd), .A(_14801_), .B(_14799_), .C(_14800_), .Y(_14802_) );
NOR2X1 NOR2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_14798_), .B(_14802_), .Y(_14803_) );
AOI22X1 AOI22X1_647 ( .gnd(gnd), .vdd(vdd), .A(_40__15_), .B(_8952_), .C(_29__15_), .D(_9176_), .Y(_14804_) );
AOI22X1 AOI22X1_648 ( .gnd(gnd), .vdd(vdd), .A(_247__15_), .B(_9165_), .C(_218__15_), .D(_9169_), .Y(_14805_) );
NAND2X1 NAND2X1_2871 ( .gnd(gnd), .vdd(vdd), .A(_14805_), .B(_14804_), .Y(_14806_) );
NAND3X1 NAND3X1_3139 ( .gnd(gnd), .vdd(vdd), .A(_9365_), .B(_16107_), .C(_16108_), .Y(_14807_) );
NAND3X1 NAND3X1_3140 ( .gnd(gnd), .vdd(vdd), .A(_9367_), .B(_16052_), .C(_16053_), .Y(_14808_) );
NAND2X1 NAND2X1_2872 ( .gnd(gnd), .vdd(vdd), .A(_14807_), .B(_14808_), .Y(_14809_) );
NAND3X1 NAND3X1_3141 ( .gnd(gnd), .vdd(vdd), .A(_9373_), .B(_8586_), .C(_8585_), .Y(_14810_) );
OAI21X1 OAI21X1_2588 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_9361_), .C(_14810_), .Y(_14811_) );
NOR2X1 NOR2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_14809_), .B(_14811_), .Y(_14812_) );
NAND2X1 NAND2X1_2873 ( .gnd(gnd), .vdd(vdd), .A(_15996_), .B(_15997_), .Y(_14813_) );
NAND3X1 NAND3X1_3142 ( .gnd(gnd), .vdd(vdd), .A(_9376_), .B(_8639_), .C(_8640_), .Y(_14814_) );
OAI21X1 OAI21X1_2589 ( .gnd(gnd), .vdd(vdd), .A(_14813_), .B(_9215_), .C(_14814_), .Y(_14815_) );
NAND3X1 NAND3X1_3143 ( .gnd(gnd), .vdd(vdd), .A(_8694_), .B(_9371_), .C(_8693_), .Y(_14816_) );
NAND3X1 NAND3X1_3144 ( .gnd(gnd), .vdd(vdd), .A(_9378_), .B(_336_), .C(_337_), .Y(_14817_) );
NAND2X1 NAND2X1_2874 ( .gnd(gnd), .vdd(vdd), .A(_14817_), .B(_14816_), .Y(_14818_) );
NOR2X1 NOR2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_14815_), .B(_14818_), .Y(_14819_) );
AOI22X1 AOI22X1_649 ( .gnd(gnd), .vdd(vdd), .A(_244__15_), .B(_9160_), .C(_177__15_), .D(_8961_), .Y(_14820_) );
NAND3X1 NAND3X1_3145 ( .gnd(gnd), .vdd(vdd), .A(_14812_), .B(_14819_), .C(_14820_), .Y(_14821_) );
NOR2X1 NOR2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_14806_), .B(_14821_), .Y(_14822_) );
NAND3X1 NAND3X1_3146 ( .gnd(gnd), .vdd(vdd), .A(_14794_), .B(_14803_), .C(_14822_), .Y(_14823_) );
NOR3X1 NOR3X1_482 ( .gnd(gnd), .vdd(vdd), .A(_14707_), .B(_14723_), .C(_14823_), .Y(_14824_) );
NAND3X1 NAND3X1_3147 ( .gnd(gnd), .vdd(vdd), .A(_14642_), .B(_14681_), .C(_14824_), .Y(_14825_) );
NAND3X1 NAND3X1_3148 ( .gnd(gnd), .vdd(vdd), .A(_8855_), .B(_1601_), .C(_1602_), .Y(_14826_) );
NAND3X1 NAND3X1_3149 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_8862_), .C(_1263_), .Y(_14827_) );
NAND2X1 NAND2X1_2875 ( .gnd(gnd), .vdd(vdd), .A(_14826_), .B(_14827_), .Y(_14828_) );
NOR3X1 NOR3X1_483 ( .gnd(gnd), .vdd(vdd), .A(_14604_), .B(_14828_), .C(_14825_), .Y(_14829_) );
NAND3X1 NAND3X1_3150 ( .gnd(gnd), .vdd(vdd), .A(_14586_), .B(_14593_), .C(_14829_), .Y(_14830_) );
NAND2X1 NAND2X1_2876 ( .gnd(gnd), .vdd(vdd), .A(_9396_), .B(_97__15_), .Y(_14831_) );
NAND3X1 NAND3X1_3151 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_9406_), .C(_1480_), .Y(_14832_) );
NAND3X1 NAND3X1_3152 ( .gnd(gnd), .vdd(vdd), .A(_1431_), .B(_9453_), .C(_1432_), .Y(_14833_) );
AND2X2 AND2X2_1616 ( .gnd(gnd), .vdd(vdd), .A(_14832_), .B(_14833_), .Y(_14834_) );
NAND2X1 NAND2X1_2877 ( .gnd(gnd), .vdd(vdd), .A(_9404_), .B(_108__15_), .Y(_14835_) );
NAND2X1 NAND2X1_2878 ( .gnd(gnd), .vdd(vdd), .A(_9401_), .B(_116__15_), .Y(_14836_) );
NAND3X1 NAND3X1_3153 ( .gnd(gnd), .vdd(vdd), .A(_14835_), .B(_14836_), .C(_14834_), .Y(_14837_) );
NAND2X1 NAND2X1_2879 ( .gnd(gnd), .vdd(vdd), .A(_9411_), .B(_125__15_), .Y(_14838_) );
NAND2X1 NAND2X1_2880 ( .gnd(gnd), .vdd(vdd), .A(_9444_), .B(_122__15_), .Y(_14839_) );
NAND2X1 NAND2X1_2881 ( .gnd(gnd), .vdd(vdd), .A(_14838_), .B(_14839_), .Y(_14840_) );
NOR2X1 NOR2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_10176_), .B(_1128_), .Y(_14841_) );
AND2X2 AND2X2_1617 ( .gnd(gnd), .vdd(vdd), .A(_120__15_), .B(_9415_), .Y(_14842_) );
NOR3X1 NOR3X1_484 ( .gnd(gnd), .vdd(vdd), .A(_14841_), .B(_14842_), .C(_14840_), .Y(_14843_) );
AOI22X1 AOI22X1_650 ( .gnd(gnd), .vdd(vdd), .A(_132__15_), .B(_9420_), .C(_131__15_), .D(_9418_), .Y(_14844_) );
NAND2X1 NAND2X1_2882 ( .gnd(gnd), .vdd(vdd), .A(_9423_), .B(_135__15_), .Y(_14845_) );
NAND2X1 NAND2X1_2883 ( .gnd(gnd), .vdd(vdd), .A(_9425_), .B(_133__15_), .Y(_14846_) );
NAND3X1 NAND3X1_3154 ( .gnd(gnd), .vdd(vdd), .A(_14845_), .B(_14846_), .C(_14844_), .Y(_14847_) );
NAND3X1 NAND3X1_3155 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_9431_), .C(_568_), .Y(_14848_) );
NAND2X1 NAND2X1_2884 ( .gnd(gnd), .vdd(vdd), .A(_9433_), .B(_229__15_), .Y(_14849_) );
NAND2X1 NAND2X1_2885 ( .gnd(gnd), .vdd(vdd), .A(_9434_), .B(_138__15_), .Y(_14850_) );
NAND3X1 NAND3X1_3156 ( .gnd(gnd), .vdd(vdd), .A(_14850_), .B(_14848_), .C(_14849_), .Y(_14851_) );
AOI21X1 AOI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_9437_), .B(_189__15_), .C(_14851_), .Y(_14852_) );
NAND2X1 NAND2X1_2886 ( .gnd(gnd), .vdd(vdd), .A(_9439_), .B(_129__15_), .Y(_14853_) );
NAND2X1 NAND2X1_2887 ( .gnd(gnd), .vdd(vdd), .A(_9429_), .B(_136__15_), .Y(_14854_) );
NAND3X1 NAND3X1_3157 ( .gnd(gnd), .vdd(vdd), .A(_14853_), .B(_14854_), .C(_14852_), .Y(_14855_) );
NAND3X1 NAND3X1_3158 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_9410_), .C(_1031_), .Y(_14856_) );
NAND2X1 NAND2X1_2888 ( .gnd(gnd), .vdd(vdd), .A(_9446_), .B(_128__15_), .Y(_14857_) );
AOI22X1 AOI22X1_651 ( .gnd(gnd), .vdd(vdd), .A(_130__15_), .B(_9449_), .C(_127__15_), .D(_9448_), .Y(_14858_) );
NAND3X1 NAND3X1_3159 ( .gnd(gnd), .vdd(vdd), .A(_14856_), .B(_14858_), .C(_14857_), .Y(_14859_) );
NOR3X1 NOR3X1_485 ( .gnd(gnd), .vdd(vdd), .A(_14847_), .B(_14855_), .C(_14859_), .Y(_14860_) );
AOI22X1 AOI22X1_652 ( .gnd(gnd), .vdd(vdd), .A(_115__15_), .B(_9399_), .C(_114__15_), .D(_9454_), .Y(_14861_) );
NAND3X1 NAND3X1_3160 ( .gnd(gnd), .vdd(vdd), .A(_14843_), .B(_14861_), .C(_14860_), .Y(_14862_) );
NOR2X1 NOR2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_14837_), .B(_14862_), .Y(_14863_) );
AOI22X1 AOI22X1_653 ( .gnd(gnd), .vdd(vdd), .A(_102__15_), .B(_9459_), .C(_103__15_), .D(_9457_), .Y(_14864_) );
NAND3X1 NAND3X1_3161 ( .gnd(gnd), .vdd(vdd), .A(_14831_), .B(_14864_), .C(_14863_), .Y(_14865_) );
NOR3X1 NOR3X1_486 ( .gnd(gnd), .vdd(vdd), .A(_14585_), .B(_14865_), .C(_14830_), .Y(_14866_) );
NAND3X1 NAND3X1_3162 ( .gnd(gnd), .vdd(vdd), .A(_14575_), .B(_14582_), .C(_14866_), .Y(_14867_) );
NAND2X1 NAND2X1_2889 ( .gnd(gnd), .vdd(vdd), .A(_8802_), .B(_75__15_), .Y(_14868_) );
NAND3X1 NAND3X1_3163 ( .gnd(gnd), .vdd(vdd), .A(_2414_), .B(_8806_), .C(_2415_), .Y(_14869_) );
NAND2X1 NAND2X1_2890 ( .gnd(gnd), .vdd(vdd), .A(_14869_), .B(_14868_), .Y(_14870_) );
NOR3X1 NOR3X1_487 ( .gnd(gnd), .vdd(vdd), .A(_14568_), .B(_14870_), .C(_14867_), .Y(_14871_) );
NAND3X1 NAND3X1_3164 ( .gnd(gnd), .vdd(vdd), .A(_14560_), .B(_14565_), .C(_14871_), .Y(_14872_) );
NAND3X1 NAND3X1_3165 ( .gnd(gnd), .vdd(vdd), .A(_3085_), .B(_9473_), .C(_3086_), .Y(_14873_) );
NAND2X1 NAND2X1_2891 ( .gnd(gnd), .vdd(vdd), .A(_9475_), .B(_66__15_), .Y(_14874_) );
NAND2X1 NAND2X1_2892 ( .gnd(gnd), .vdd(vdd), .A(_9466_), .B(_79__15_), .Y(_14875_) );
NAND2X1 NAND2X1_2893 ( .gnd(gnd), .vdd(vdd), .A(_8805_), .B(_80__15_), .Y(_14876_) );
NAND2X1 NAND2X1_2894 ( .gnd(gnd), .vdd(vdd), .A(_9478_), .B(_77__15_), .Y(_14877_) );
NAND3X1 NAND3X1_3166 ( .gnd(gnd), .vdd(vdd), .A(_14875_), .B(_14876_), .C(_14877_), .Y(_14878_) );
AOI21X1 AOI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_68__15_), .B(_9477_), .C(_14878_), .Y(_14879_) );
NAND3X1 NAND3X1_3167 ( .gnd(gnd), .vdd(vdd), .A(_14873_), .B(_14879_), .C(_14874_), .Y(_14880_) );
NOR3X1 NOR3X1_488 ( .gnd(gnd), .vdd(vdd), .A(_14559_), .B(_14880_), .C(_14872_), .Y(_14881_) );
AOI21X1 AOI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_14554_), .B(_14881_), .C(rst), .Y(_0__15_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_16233__0_), .Y(IDATA_CORE_out[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_16233__1_), .Y(IDATA_CORE_out[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_16233__2_), .Y(IDATA_CORE_out[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_16233__3_), .Y(IDATA_CORE_out[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_16233__4_), .Y(IDATA_CORE_out[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_16233__5_), .Y(IDATA_CORE_out[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_16233__6_), .Y(IDATA_CORE_out[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_16233__7_), .Y(IDATA_CORE_out[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_16233__8_), .Y(IDATA_CORE_out[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_16233__9_), .Y(IDATA_CORE_out[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_16233__10_), .Y(IDATA_CORE_out[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_16233__11_), .Y(IDATA_CORE_out[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_16233__12_), .Y(IDATA_CORE_out[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_16233__13_), .Y(IDATA_CORE_out[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_16233__14_), .Y(IDATA_CORE_out[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_16233__15_), .Y(IDATA_CORE_out[15]) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf3), .D(_0__0_), .Q(_16233__0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf3), .D(_0__1_), .Q(_16233__1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf3), .D(_0__2_), .Q(_16233__2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf3), .D(_0__3_), .Q(_16233__3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf3), .D(_0__4_), .Q(_16233__4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf3), .D(_0__5_), .Q(_16233__5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf3), .D(_0__6_), .Q(_16233__6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf3), .D(_0__7_), .Q(_16233__7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf3), .D(_0__8_), .Q(_16233__8_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf3), .D(_0__9_), .Q(_16233__9_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf3), .D(_0__10_), .Q(_16233__10_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf3), .D(_0__11_), .Q(_16233__11_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf3), .D(_0__12_), .Q(_16233__12_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf3), .D(_0__13_), .Q(_16233__13_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf3), .D(_0__14_), .Q(_16233__14_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf3), .D(_0__15_), .Q(_16233__15_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_1__0_), .Q(data_0__0_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_1__1_), .Q(data_0__1_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_1__2_), .Q(data_0__2_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_1__3_), .Q(data_0__3_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_1__4_), .Q(data_0__4_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_1__5_), .Q(data_0__5_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_1__6_), .Q(data_0__6_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_1__7_), .Q(data_0__7_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_1__8_), .Q(data_0__8_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_1__9_), .Q(data_0__9_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_1__10_), .Q(data_0__10_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_1__11_), .Q(data_0__11_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_1__12_), .Q(data_0__12_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_1__13_), .Q(data_0__13_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_1__14_), .Q(data_0__14_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_1__15_), .Q(data_0__15_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_112__0_), .Q(data_1__0_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_112__1_), .Q(data_1__1_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_112__2_), .Q(data_1__2_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_112__3_), .Q(data_1__3_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_112__4_), .Q(data_1__4_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_112__5_), .Q(data_1__5_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_112__6_), .Q(data_1__6_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_112__7_), .Q(data_1__7_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_112__8_), .Q(data_1__8_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_112__9_), .Q(data_1__9_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_112__10_), .Q(data_1__10_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_112__11_), .Q(data_1__11_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_112__12_), .Q(data_1__12_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_112__13_), .Q(data_1__13_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_112__14_), .Q(data_1__14_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_112__15_), .Q(data_1__15_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_179__0_), .Q(data_2__0_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_179__1_), .Q(data_2__1_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_179__2_), .Q(data_2__2_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_179__3_), .Q(data_2__3_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_179__4_), .Q(data_2__4_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_179__5_), .Q(data_2__5_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_179__6_), .Q(data_2__6_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_179__7_), .Q(data_2__7_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_179__8_), .Q(data_2__8_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_179__9_), .Q(data_2__9_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_179__10_), .Q(data_2__10_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_179__11_), .Q(data_2__11_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_179__12_), .Q(data_2__12_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_179__13_), .Q(data_2__13_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_179__14_), .Q(data_2__14_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_179__15_), .Q(data_2__15_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_190__0_), .Q(data_3__0_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_190__1_), .Q(data_3__1_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_190__2_), .Q(data_3__2_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_190__3_), .Q(data_3__3_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_190__4_), .Q(data_3__4_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_190__5_), .Q(data_3__5_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_190__6_), .Q(data_3__6_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_190__7_), .Q(data_3__7_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_190__8_), .Q(data_3__8_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_190__9_), .Q(data_3__9_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_190__10_), .Q(data_3__10_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_190__11_), .Q(data_3__11_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_190__12_), .Q(data_3__12_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_190__13_), .Q(data_3__13_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_190__14_), .Q(data_3__14_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_190__15_), .Q(data_3__15_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_201__0_), .Q(data_4__0_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_201__1_), .Q(data_4__1_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_201__2_), .Q(data_4__2_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_201__3_), .Q(data_4__3_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_201__4_), .Q(data_4__4_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_201__5_), .Q(data_4__5_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_201__6_), .Q(data_4__6_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_201__7_), .Q(data_4__7_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_201__8_), .Q(data_4__8_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_201__9_), .Q(data_4__9_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_201__10_), .Q(data_4__10_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_201__11_), .Q(data_4__11_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_201__12_), .Q(data_4__12_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_201__13_), .Q(data_4__13_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_201__14_), .Q(data_4__14_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_201__15_), .Q(data_4__15_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_212__0_), .Q(data_5__0_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_212__1_), .Q(data_5__1_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_212__2_), .Q(data_5__2_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_212__3_), .Q(data_5__3_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_212__4_), .Q(data_5__4_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_212__5_), .Q(data_5__5_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_212__6_), .Q(data_5__6_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_212__7_), .Q(data_5__7_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_212__8_), .Q(data_5__8_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_212__9_), .Q(data_5__9_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_212__10_), .Q(data_5__10_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_212__11_), .Q(data_5__11_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_212__12_), .Q(data_5__12_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_212__13_), .Q(data_5__13_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_212__14_), .Q(data_5__14_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_212__15_), .Q(data_5__15_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_223__0_), .Q(data_6__0_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_223__1_), .Q(data_6__1_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_223__2_), .Q(data_6__2_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_223__3_), .Q(data_6__3_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_223__4_), .Q(data_6__4_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_223__5_), .Q(data_6__5_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_223__6_), .Q(data_6__6_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_223__7_), .Q(data_6__7_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_223__8_), .Q(data_6__8_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_223__9_), .Q(data_6__9_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_223__10_), .Q(data_6__10_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_223__11_), .Q(data_6__11_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_223__12_), .Q(data_6__12_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_223__13_), .Q(data_6__13_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_223__14_), .Q(data_6__14_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_223__15_), .Q(data_6__15_) );
DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_234__0_), .Q(data_7__0_) );
DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_234__1_), .Q(data_7__1_) );
DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_234__2_), .Q(data_7__2_) );
DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_234__3_), .Q(data_7__3_) );
DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_234__4_), .Q(data_7__4_) );
DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_234__5_), .Q(data_7__5_) );
DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_234__6_), .Q(data_7__6_) );
DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_234__7_), .Q(data_7__7_) );
DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_234__8_), .Q(data_7__8_) );
DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_234__9_), .Q(data_7__9_) );
DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_234__10_), .Q(data_7__10_) );
DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_234__11_), .Q(data_7__11_) );
DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_234__12_), .Q(data_7__12_) );
DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_234__13_), .Q(data_7__13_) );
DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_234__14_), .Q(data_7__14_) );
DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_234__15_), .Q(data_7__15_) );
DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_245__0_), .Q(data_8__0_) );
DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_245__1_), .Q(data_8__1_) );
DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_245__2_), .Q(data_8__2_) );
DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_245__3_), .Q(data_8__3_) );
DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_245__4_), .Q(data_8__4_) );
DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_245__5_), .Q(data_8__5_) );
DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_245__6_), .Q(data_8__6_) );
DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_245__7_), .Q(data_8__7_) );
DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_245__8_), .Q(data_8__8_) );
DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_245__9_), .Q(data_8__9_) );
DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_245__10_), .Q(data_8__10_) );
DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_245__11_), .Q(data_8__11_) );
DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_245__12_), .Q(data_8__12_) );
DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_245__13_), .Q(data_8__13_) );
DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_245__14_), .Q(data_8__14_) );
DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_245__15_), .Q(data_8__15_) );
DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_256__0_), .Q(data_9__0_) );
DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_256__1_), .Q(data_9__1_) );
DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_256__2_), .Q(data_9__2_) );
DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_256__3_), .Q(data_9__3_) );
DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_256__4_), .Q(data_9__4_) );
DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_256__5_), .Q(data_9__5_) );
DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_256__6_), .Q(data_9__6_) );
DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_256__7_), .Q(data_9__7_) );
DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_256__8_), .Q(data_9__8_) );
DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_256__9_), .Q(data_9__9_) );
DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_256__10_), .Q(data_9__10_) );
DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_256__11_), .Q(data_9__11_) );
DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_256__12_), .Q(data_9__12_) );
DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_256__13_), .Q(data_9__13_) );
DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_256__14_), .Q(data_9__14_) );
DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_256__15_), .Q(data_9__15_) );
DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_12__0_), .Q(data_10__0_) );
DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_12__1_), .Q(data_10__1_) );
DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_12__2_), .Q(data_10__2_) );
DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_12__3_), .Q(data_10__3_) );
DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_12__4_), .Q(data_10__4_) );
DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_12__5_), .Q(data_10__5_) );
DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_12__6_), .Q(data_10__6_) );
DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_12__7_), .Q(data_10__7_) );
DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_12__8_), .Q(data_10__8_) );
DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_12__9_), .Q(data_10__9_) );
DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_12__10_), .Q(data_10__10_) );
DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_12__11_), .Q(data_10__11_) );
DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_12__12_), .Q(data_10__12_) );
DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_12__13_), .Q(data_10__13_) );
DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_12__14_), .Q(data_10__14_) );
DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_12__15_), .Q(data_10__15_) );
DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_23__0_), .Q(data_11__0_) );
DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_23__1_), .Q(data_11__1_) );
DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_23__2_), .Q(data_11__2_) );
DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_23__3_), .Q(data_11__3_) );
DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_23__4_), .Q(data_11__4_) );
DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_23__5_), .Q(data_11__5_) );
DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_23__6_), .Q(data_11__6_) );
DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_23__7_), .Q(data_11__7_) );
DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_23__8_), .Q(data_11__8_) );
DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_23__9_), .Q(data_11__9_) );
DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_23__10_), .Q(data_11__10_) );
DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_23__11_), .Q(data_11__11_) );
DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_23__12_), .Q(data_11__12_) );
DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_23__13_), .Q(data_11__13_) );
DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_23__14_), .Q(data_11__14_) );
DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_23__15_), .Q(data_11__15_) );
DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_34__0_), .Q(data_12__0_) );
DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_34__1_), .Q(data_12__1_) );
DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_34__2_), .Q(data_12__2_) );
DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_34__3_), .Q(data_12__3_) );
DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_34__4_), .Q(data_12__4_) );
DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_34__5_), .Q(data_12__5_) );
DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_34__6_), .Q(data_12__6_) );
DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_34__7_), .Q(data_12__7_) );
DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_34__8_), .Q(data_12__8_) );
DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_34__9_), .Q(data_12__9_) );
DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_34__10_), .Q(data_12__10_) );
DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_34__11_), .Q(data_12__11_) );
DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_34__12_), .Q(data_12__12_) );
DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_34__13_), .Q(data_12__13_) );
DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_34__14_), .Q(data_12__14_) );
DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_34__15_), .Q(data_12__15_) );
DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_45__0_), .Q(data_13__0_) );
DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_45__1_), .Q(data_13__1_) );
DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_45__2_), .Q(data_13__2_) );
DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_45__3_), .Q(data_13__3_) );
DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_45__4_), .Q(data_13__4_) );
DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_45__5_), .Q(data_13__5_) );
DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_45__6_), .Q(data_13__6_) );
DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_45__7_), .Q(data_13__7_) );
DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_45__8_), .Q(data_13__8_) );
DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_45__9_), .Q(data_13__9_) );
DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_45__10_), .Q(data_13__10_) );
DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_45__11_), .Q(data_13__11_) );
DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_45__12_), .Q(data_13__12_) );
DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_45__13_), .Q(data_13__13_) );
DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_45__14_), .Q(data_13__14_) );
DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_45__15_), .Q(data_13__15_) );
DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_56__0_), .Q(data_14__0_) );
DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_56__1_), .Q(data_14__1_) );
DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_56__2_), .Q(data_14__2_) );
DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_56__3_), .Q(data_14__3_) );
DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_56__4_), .Q(data_14__4_) );
DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_56__5_), .Q(data_14__5_) );
DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_56__6_), .Q(data_14__6_) );
DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_56__7_), .Q(data_14__7_) );
DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_56__8_), .Q(data_14__8_) );
DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_56__9_), .Q(data_14__9_) );
DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_56__10_), .Q(data_14__10_) );
DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_56__11_), .Q(data_14__11_) );
DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_56__12_), .Q(data_14__12_) );
DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_56__13_), .Q(data_14__13_) );
DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_56__14_), .Q(data_14__14_) );
DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_56__15_), .Q(data_14__15_) );
DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf2), .D(_67__0_), .Q(data_15__0_) );
DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf2), .D(_67__1_), .Q(data_15__1_) );
DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf2), .D(_67__2_), .Q(data_15__2_) );
DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf2), .D(_67__3_), .Q(data_15__3_) );
DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf2), .D(_67__4_), .Q(data_15__4_) );
DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf2), .D(_67__5_), .Q(data_15__5_) );
DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf2), .D(_67__6_), .Q(data_15__6_) );
DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf2), .D(_67__7_), .Q(data_15__7_) );
DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf2), .D(_67__8_), .Q(data_15__8_) );
DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf2), .D(_67__9_), .Q(data_15__9_) );
DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf2), .D(_67__10_), .Q(data_15__10_) );
DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf2), .D(_67__11_), .Q(data_15__11_) );
DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf2), .D(_67__12_), .Q(data_15__12_) );
DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf2), .D(_67__13_), .Q(data_15__13_) );
DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf2), .D(_67__14_), .Q(data_15__14_) );
DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf2), .D(_67__15_), .Q(data_15__15_) );
DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_78__0_), .Q(data_16__0_) );
DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_78__1_), .Q(data_16__1_) );
DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_78__2_), .Q(data_16__2_) );
DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_78__3_), .Q(data_16__3_) );
DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_78__4_), .Q(data_16__4_) );
DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_78__5_), .Q(data_16__5_) );
DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_78__6_), .Q(data_16__6_) );
DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_78__7_), .Q(data_16__7_) );
DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_78__8_), .Q(data_16__8_) );
DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_78__9_), .Q(data_16__9_) );
DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_78__10_), .Q(data_16__10_) );
DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_78__11_), .Q(data_16__11_) );
DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_78__12_), .Q(data_16__12_) );
DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_78__13_), .Q(data_16__13_) );
DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_78__14_), .Q(data_16__14_) );
DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_78__15_), .Q(data_16__15_) );
DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_89__0_), .Q(data_17__0_) );
DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_89__1_), .Q(data_17__1_) );
DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_89__2_), .Q(data_17__2_) );
DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_89__3_), .Q(data_17__3_) );
DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_89__4_), .Q(data_17__4_) );
DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_89__5_), .Q(data_17__5_) );
DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_89__6_), .Q(data_17__6_) );
DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_89__7_), .Q(data_17__7_) );
DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_89__8_), .Q(data_17__8_) );
DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_89__9_), .Q(data_17__9_) );
DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_89__10_), .Q(data_17__10_) );
DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_89__11_), .Q(data_17__11_) );
DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_89__12_), .Q(data_17__12_) );
DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_89__13_), .Q(data_17__13_) );
DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_89__14_), .Q(data_17__14_) );
DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_89__15_), .Q(data_17__15_) );
DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_100__0_), .Q(data_18__0_) );
DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_100__1_), .Q(data_18__1_) );
DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_100__2_), .Q(data_18__2_) );
DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_100__3_), .Q(data_18__3_) );
DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_100__4_), .Q(data_18__4_) );
DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_100__5_), .Q(data_18__5_) );
DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_100__6_), .Q(data_18__6_) );
DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_100__7_), .Q(data_18__7_) );
DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_100__8_), .Q(data_18__8_) );
DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_100__9_), .Q(data_18__9_) );
DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_100__10_), .Q(data_18__10_) );
DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_100__11_), .Q(data_18__11_) );
DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_100__12_), .Q(data_18__12_) );
DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_100__13_), .Q(data_18__13_) );
DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_100__14_), .Q(data_18__14_) );
DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_100__15_), .Q(data_18__15_) );
DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_111__0_), .Q(data_19__0_) );
DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_111__1_), .Q(data_19__1_) );
DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_111__2_), .Q(data_19__2_) );
DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_111__3_), .Q(data_19__3_) );
DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_111__4_), .Q(data_19__4_) );
DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_111__5_), .Q(data_19__5_) );
DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_111__6_), .Q(data_19__6_) );
DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_111__7_), .Q(data_19__7_) );
DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_111__8_), .Q(data_19__8_) );
DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_111__9_), .Q(data_19__9_) );
DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_111__10_), .Q(data_19__10_) );
DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_111__11_), .Q(data_19__11_) );
DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_111__12_), .Q(data_19__12_) );
DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_111__13_), .Q(data_19__13_) );
DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_111__14_), .Q(data_19__14_) );
DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_111__15_), .Q(data_19__15_) );
DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_123__0_), .Q(data_20__0_) );
DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_123__1_), .Q(data_20__1_) );
DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_123__2_), .Q(data_20__2_) );
DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_123__3_), .Q(data_20__3_) );
DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_123__4_), .Q(data_20__4_) );
DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_123__5_), .Q(data_20__5_) );
DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_123__6_), .Q(data_20__6_) );
DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_123__7_), .Q(data_20__7_) );
DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_123__8_), .Q(data_20__8_) );
DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_123__9_), .Q(data_20__9_) );
DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_123__10_), .Q(data_20__10_) );
DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_123__11_), .Q(data_20__11_) );
DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_123__12_), .Q(data_20__12_) );
DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_123__13_), .Q(data_20__13_) );
DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_123__14_), .Q(data_20__14_) );
DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_123__15_), .Q(data_20__15_) );
DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_134__0_), .Q(data_21__0_) );
DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_134__1_), .Q(data_21__1_) );
DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_134__2_), .Q(data_21__2_) );
DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_134__3_), .Q(data_21__3_) );
DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_134__4_), .Q(data_21__4_) );
DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_134__5_), .Q(data_21__5_) );
DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_134__6_), .Q(data_21__6_) );
DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_134__7_), .Q(data_21__7_) );
DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_134__8_), .Q(data_21__8_) );
DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_134__9_), .Q(data_21__9_) );
DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_134__10_), .Q(data_21__10_) );
DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_134__11_), .Q(data_21__11_) );
DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_134__12_), .Q(data_21__12_) );
DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_134__13_), .Q(data_21__13_) );
DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_134__14_), .Q(data_21__14_) );
DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_134__15_), .Q(data_21__15_) );
DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_145__0_), .Q(data_22__0_) );
DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_145__1_), .Q(data_22__1_) );
DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_145__2_), .Q(data_22__2_) );
DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_145__3_), .Q(data_22__3_) );
DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_145__4_), .Q(data_22__4_) );
DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_145__5_), .Q(data_22__5_) );
DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_145__6_), .Q(data_22__6_) );
DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_145__7_), .Q(data_22__7_) );
DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_145__8_), .Q(data_22__8_) );
DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_145__9_), .Q(data_22__9_) );
DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_145__10_), .Q(data_22__10_) );
DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_145__11_), .Q(data_22__11_) );
DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_145__12_), .Q(data_22__12_) );
DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_145__13_), .Q(data_22__13_) );
DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_145__14_), .Q(data_22__14_) );
DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_145__15_), .Q(data_22__15_) );
DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_156__0_), .Q(data_23__0_) );
DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_156__1_), .Q(data_23__1_) );
DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_156__2_), .Q(data_23__2_) );
DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_156__3_), .Q(data_23__3_) );
DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_156__4_), .Q(data_23__4_) );
DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_156__5_), .Q(data_23__5_) );
DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_156__6_), .Q(data_23__6_) );
DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_156__7_), .Q(data_23__7_) );
DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_156__8_), .Q(data_23__8_) );
DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_156__9_), .Q(data_23__9_) );
DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_156__10_), .Q(data_23__10_) );
DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_156__11_), .Q(data_23__11_) );
DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_156__12_), .Q(data_23__12_) );
DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_156__13_), .Q(data_23__13_) );
DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_156__14_), .Q(data_23__14_) );
DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_156__15_), .Q(data_23__15_) );
DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_167__0_), .Q(data_24__0_) );
DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_167__1_), .Q(data_24__1_) );
DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_167__2_), .Q(data_24__2_) );
DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_167__3_), .Q(data_24__3_) );
DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_167__4_), .Q(data_24__4_) );
DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_167__5_), .Q(data_24__5_) );
DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_167__6_), .Q(data_24__6_) );
DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_167__7_), .Q(data_24__7_) );
DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_167__8_), .Q(data_24__8_) );
DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_167__9_), .Q(data_24__9_) );
DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_167__10_), .Q(data_24__10_) );
DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_167__11_), .Q(data_24__11_) );
DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_167__12_), .Q(data_24__12_) );
DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_167__13_), .Q(data_24__13_) );
DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_167__14_), .Q(data_24__14_) );
DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_167__15_), .Q(data_24__15_) );
DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_174__0_), .Q(data_25__0_) );
DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_174__1_), .Q(data_25__1_) );
DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_174__2_), .Q(data_25__2_) );
DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_174__3_), .Q(data_25__3_) );
DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_174__4_), .Q(data_25__4_) );
DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_174__5_), .Q(data_25__5_) );
DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_174__6_), .Q(data_25__6_) );
DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_174__7_), .Q(data_25__7_) );
DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_174__8_), .Q(data_25__8_) );
DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_174__9_), .Q(data_25__9_) );
DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_174__10_), .Q(data_25__10_) );
DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_174__11_), .Q(data_25__11_) );
DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_174__12_), .Q(data_25__12_) );
DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_174__13_), .Q(data_25__13_) );
DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_174__14_), .Q(data_25__14_) );
DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_174__15_), .Q(data_25__15_) );
DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_175__0_), .Q(data_26__0_) );
DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_175__1_), .Q(data_26__1_) );
DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_175__2_), .Q(data_26__2_) );
DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_175__3_), .Q(data_26__3_) );
DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_175__4_), .Q(data_26__4_) );
DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_175__5_), .Q(data_26__5_) );
DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_175__6_), .Q(data_26__6_) );
DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_175__7_), .Q(data_26__7_) );
DFFPOSX1 DFFPOSX1_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_175__8_), .Q(data_26__8_) );
DFFPOSX1 DFFPOSX1_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_175__9_), .Q(data_26__9_) );
DFFPOSX1 DFFPOSX1_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_175__10_), .Q(data_26__10_) );
DFFPOSX1 DFFPOSX1_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_175__11_), .Q(data_26__11_) );
DFFPOSX1 DFFPOSX1_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_175__12_), .Q(data_26__12_) );
DFFPOSX1 DFFPOSX1_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_175__13_), .Q(data_26__13_) );
DFFPOSX1 DFFPOSX1_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_175__14_), .Q(data_26__14_) );
DFFPOSX1 DFFPOSX1_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_175__15_), .Q(data_26__15_) );
DFFPOSX1 DFFPOSX1_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_176__0_), .Q(data_27__0_) );
DFFPOSX1 DFFPOSX1_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_176__1_), .Q(data_27__1_) );
DFFPOSX1 DFFPOSX1_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_176__2_), .Q(data_27__2_) );
DFFPOSX1 DFFPOSX1_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_176__3_), .Q(data_27__3_) );
DFFPOSX1 DFFPOSX1_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_176__4_), .Q(data_27__4_) );
DFFPOSX1 DFFPOSX1_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_176__5_), .Q(data_27__5_) );
DFFPOSX1 DFFPOSX1_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_176__6_), .Q(data_27__6_) );
DFFPOSX1 DFFPOSX1_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_176__7_), .Q(data_27__7_) );
DFFPOSX1 DFFPOSX1_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_176__8_), .Q(data_27__8_) );
DFFPOSX1 DFFPOSX1_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_176__9_), .Q(data_27__9_) );
DFFPOSX1 DFFPOSX1_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_176__10_), .Q(data_27__10_) );
DFFPOSX1 DFFPOSX1_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_176__11_), .Q(data_27__11_) );
DFFPOSX1 DFFPOSX1_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_176__12_), .Q(data_27__12_) );
DFFPOSX1 DFFPOSX1_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_176__13_), .Q(data_27__13_) );
DFFPOSX1 DFFPOSX1_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_176__14_), .Q(data_27__14_) );
DFFPOSX1 DFFPOSX1_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_176__15_), .Q(data_27__15_) );
DFFPOSX1 DFFPOSX1_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_177__0_), .Q(data_28__0_) );
DFFPOSX1 DFFPOSX1_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_177__1_), .Q(data_28__1_) );
DFFPOSX1 DFFPOSX1_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_177__2_), .Q(data_28__2_) );
DFFPOSX1 DFFPOSX1_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_177__3_), .Q(data_28__3_) );
DFFPOSX1 DFFPOSX1_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_177__4_), .Q(data_28__4_) );
DFFPOSX1 DFFPOSX1_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_177__5_), .Q(data_28__5_) );
DFFPOSX1 DFFPOSX1_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_177__6_), .Q(data_28__6_) );
DFFPOSX1 DFFPOSX1_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_177__7_), .Q(data_28__7_) );
DFFPOSX1 DFFPOSX1_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_177__8_), .Q(data_28__8_) );
DFFPOSX1 DFFPOSX1_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_177__9_), .Q(data_28__9_) );
DFFPOSX1 DFFPOSX1_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_177__10_), .Q(data_28__10_) );
DFFPOSX1 DFFPOSX1_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_177__11_), .Q(data_28__11_) );
DFFPOSX1 DFFPOSX1_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_177__12_), .Q(data_28__12_) );
DFFPOSX1 DFFPOSX1_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_177__13_), .Q(data_28__13_) );
DFFPOSX1 DFFPOSX1_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_177__14_), .Q(data_28__14_) );
DFFPOSX1 DFFPOSX1_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_177__15_), .Q(data_28__15_) );
DFFPOSX1 DFFPOSX1_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_178__0_), .Q(data_29__0_) );
DFFPOSX1 DFFPOSX1_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_178__1_), .Q(data_29__1_) );
DFFPOSX1 DFFPOSX1_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_178__2_), .Q(data_29__2_) );
DFFPOSX1 DFFPOSX1_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_178__3_), .Q(data_29__3_) );
DFFPOSX1 DFFPOSX1_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_178__4_), .Q(data_29__4_) );
DFFPOSX1 DFFPOSX1_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_178__5_), .Q(data_29__5_) );
DFFPOSX1 DFFPOSX1_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_178__6_), .Q(data_29__6_) );
DFFPOSX1 DFFPOSX1_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_178__7_), .Q(data_29__7_) );
DFFPOSX1 DFFPOSX1_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_178__8_), .Q(data_29__8_) );
DFFPOSX1 DFFPOSX1_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_178__9_), .Q(data_29__9_) );
DFFPOSX1 DFFPOSX1_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_178__10_), .Q(data_29__10_) );
DFFPOSX1 DFFPOSX1_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_178__11_), .Q(data_29__11_) );
DFFPOSX1 DFFPOSX1_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_178__12_), .Q(data_29__12_) );
DFFPOSX1 DFFPOSX1_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_178__13_), .Q(data_29__13_) );
DFFPOSX1 DFFPOSX1_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_178__14_), .Q(data_29__14_) );
DFFPOSX1 DFFPOSX1_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_178__15_), .Q(data_29__15_) );
DFFPOSX1 DFFPOSX1_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_180__0_), .Q(data_30__0_) );
DFFPOSX1 DFFPOSX1_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_180__1_), .Q(data_30__1_) );
DFFPOSX1 DFFPOSX1_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_180__2_), .Q(data_30__2_) );
DFFPOSX1 DFFPOSX1_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_180__3_), .Q(data_30__3_) );
DFFPOSX1 DFFPOSX1_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_180__4_), .Q(data_30__4_) );
DFFPOSX1 DFFPOSX1_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_180__5_), .Q(data_30__5_) );
DFFPOSX1 DFFPOSX1_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_180__6_), .Q(data_30__6_) );
DFFPOSX1 DFFPOSX1_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_180__7_), .Q(data_30__7_) );
DFFPOSX1 DFFPOSX1_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_180__8_), .Q(data_30__8_) );
DFFPOSX1 DFFPOSX1_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_180__9_), .Q(data_30__9_) );
DFFPOSX1 DFFPOSX1_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_180__10_), .Q(data_30__10_) );
DFFPOSX1 DFFPOSX1_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_180__11_), .Q(data_30__11_) );
DFFPOSX1 DFFPOSX1_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_180__12_), .Q(data_30__12_) );
DFFPOSX1 DFFPOSX1_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_180__13_), .Q(data_30__13_) );
DFFPOSX1 DFFPOSX1_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_180__14_), .Q(data_30__14_) );
DFFPOSX1 DFFPOSX1_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_180__15_), .Q(data_30__15_) );
DFFPOSX1 DFFPOSX1_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf1), .D(_181__0_), .Q(data_31__0_) );
DFFPOSX1 DFFPOSX1_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf1), .D(_181__1_), .Q(data_31__1_) );
DFFPOSX1 DFFPOSX1_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf1), .D(_181__2_), .Q(data_31__2_) );
DFFPOSX1 DFFPOSX1_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf1), .D(_181__3_), .Q(data_31__3_) );
DFFPOSX1 DFFPOSX1_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf1), .D(_181__4_), .Q(data_31__4_) );
DFFPOSX1 DFFPOSX1_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf1), .D(_181__5_), .Q(data_31__5_) );
DFFPOSX1 DFFPOSX1_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf1), .D(_181__6_), .Q(data_31__6_) );
DFFPOSX1 DFFPOSX1_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf1), .D(_181__7_), .Q(data_31__7_) );
DFFPOSX1 DFFPOSX1_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf1), .D(_181__8_), .Q(data_31__8_) );
DFFPOSX1 DFFPOSX1_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf1), .D(_181__9_), .Q(data_31__9_) );
DFFPOSX1 DFFPOSX1_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf1), .D(_181__10_), .Q(data_31__10_) );
DFFPOSX1 DFFPOSX1_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf1), .D(_181__11_), .Q(data_31__11_) );
DFFPOSX1 DFFPOSX1_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf1), .D(_181__12_), .Q(data_31__12_) );
DFFPOSX1 DFFPOSX1_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf1), .D(_181__13_), .Q(data_31__13_) );
DFFPOSX1 DFFPOSX1_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf1), .D(_181__14_), .Q(data_31__14_) );
DFFPOSX1 DFFPOSX1_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf1), .D(_181__15_), .Q(data_31__15_) );
DFFPOSX1 DFFPOSX1_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_182__0_), .Q(data_32__0_) );
DFFPOSX1 DFFPOSX1_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_182__1_), .Q(data_32__1_) );
DFFPOSX1 DFFPOSX1_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_182__2_), .Q(data_32__2_) );
DFFPOSX1 DFFPOSX1_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_182__3_), .Q(data_32__3_) );
DFFPOSX1 DFFPOSX1_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_182__4_), .Q(data_32__4_) );
DFFPOSX1 DFFPOSX1_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_182__5_), .Q(data_32__5_) );
DFFPOSX1 DFFPOSX1_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_182__6_), .Q(data_32__6_) );
DFFPOSX1 DFFPOSX1_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_182__7_), .Q(data_32__7_) );
DFFPOSX1 DFFPOSX1_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_182__8_), .Q(data_32__8_) );
DFFPOSX1 DFFPOSX1_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_182__9_), .Q(data_32__9_) );
DFFPOSX1 DFFPOSX1_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_182__10_), .Q(data_32__10_) );
DFFPOSX1 DFFPOSX1_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_182__11_), .Q(data_32__11_) );
DFFPOSX1 DFFPOSX1_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_182__12_), .Q(data_32__12_) );
DFFPOSX1 DFFPOSX1_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_182__13_), .Q(data_32__13_) );
DFFPOSX1 DFFPOSX1_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_182__14_), .Q(data_32__14_) );
DFFPOSX1 DFFPOSX1_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_182__15_), .Q(data_32__15_) );
DFFPOSX1 DFFPOSX1_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_183__0_), .Q(data_33__0_) );
DFFPOSX1 DFFPOSX1_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_183__1_), .Q(data_33__1_) );
DFFPOSX1 DFFPOSX1_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_183__2_), .Q(data_33__2_) );
DFFPOSX1 DFFPOSX1_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_183__3_), .Q(data_33__3_) );
DFFPOSX1 DFFPOSX1_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_183__4_), .Q(data_33__4_) );
DFFPOSX1 DFFPOSX1_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_183__5_), .Q(data_33__5_) );
DFFPOSX1 DFFPOSX1_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_183__6_), .Q(data_33__6_) );
DFFPOSX1 DFFPOSX1_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_183__7_), .Q(data_33__7_) );
DFFPOSX1 DFFPOSX1_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_183__8_), .Q(data_33__8_) );
DFFPOSX1 DFFPOSX1_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_183__9_), .Q(data_33__9_) );
DFFPOSX1 DFFPOSX1_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_183__10_), .Q(data_33__10_) );
DFFPOSX1 DFFPOSX1_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_183__11_), .Q(data_33__11_) );
DFFPOSX1 DFFPOSX1_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_183__12_), .Q(data_33__12_) );
DFFPOSX1 DFFPOSX1_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_183__13_), .Q(data_33__13_) );
DFFPOSX1 DFFPOSX1_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_183__14_), .Q(data_33__14_) );
DFFPOSX1 DFFPOSX1_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_183__15_), .Q(data_33__15_) );
DFFPOSX1 DFFPOSX1_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_184__0_), .Q(data_34__0_) );
DFFPOSX1 DFFPOSX1_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_184__1_), .Q(data_34__1_) );
DFFPOSX1 DFFPOSX1_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_184__2_), .Q(data_34__2_) );
DFFPOSX1 DFFPOSX1_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_184__3_), .Q(data_34__3_) );
DFFPOSX1 DFFPOSX1_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_184__4_), .Q(data_34__4_) );
DFFPOSX1 DFFPOSX1_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_184__5_), .Q(data_34__5_) );
DFFPOSX1 DFFPOSX1_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_184__6_), .Q(data_34__6_) );
DFFPOSX1 DFFPOSX1_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_184__7_), .Q(data_34__7_) );
DFFPOSX1 DFFPOSX1_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_184__8_), .Q(data_34__8_) );
DFFPOSX1 DFFPOSX1_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_184__9_), .Q(data_34__9_) );
DFFPOSX1 DFFPOSX1_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_184__10_), .Q(data_34__10_) );
DFFPOSX1 DFFPOSX1_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_184__11_), .Q(data_34__11_) );
DFFPOSX1 DFFPOSX1_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_184__12_), .Q(data_34__12_) );
DFFPOSX1 DFFPOSX1_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_184__13_), .Q(data_34__13_) );
DFFPOSX1 DFFPOSX1_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_184__14_), .Q(data_34__14_) );
DFFPOSX1 DFFPOSX1_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_184__15_), .Q(data_34__15_) );
DFFPOSX1 DFFPOSX1_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_185__0_), .Q(data_35__0_) );
DFFPOSX1 DFFPOSX1_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_185__1_), .Q(data_35__1_) );
DFFPOSX1 DFFPOSX1_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_185__2_), .Q(data_35__2_) );
DFFPOSX1 DFFPOSX1_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_185__3_), .Q(data_35__3_) );
DFFPOSX1 DFFPOSX1_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_185__4_), .Q(data_35__4_) );
DFFPOSX1 DFFPOSX1_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_185__5_), .Q(data_35__5_) );
DFFPOSX1 DFFPOSX1_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_185__6_), .Q(data_35__6_) );
DFFPOSX1 DFFPOSX1_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_185__7_), .Q(data_35__7_) );
DFFPOSX1 DFFPOSX1_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_185__8_), .Q(data_35__8_) );
DFFPOSX1 DFFPOSX1_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_185__9_), .Q(data_35__9_) );
DFFPOSX1 DFFPOSX1_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_185__10_), .Q(data_35__10_) );
DFFPOSX1 DFFPOSX1_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_185__11_), .Q(data_35__11_) );
DFFPOSX1 DFFPOSX1_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_185__12_), .Q(data_35__12_) );
DFFPOSX1 DFFPOSX1_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_185__13_), .Q(data_35__13_) );
DFFPOSX1 DFFPOSX1_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_185__14_), .Q(data_35__14_) );
DFFPOSX1 DFFPOSX1_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_185__15_), .Q(data_35__15_) );
DFFPOSX1 DFFPOSX1_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_186__0_), .Q(data_36__0_) );
DFFPOSX1 DFFPOSX1_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_186__1_), .Q(data_36__1_) );
DFFPOSX1 DFFPOSX1_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_186__2_), .Q(data_36__2_) );
DFFPOSX1 DFFPOSX1_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_186__3_), .Q(data_36__3_) );
DFFPOSX1 DFFPOSX1_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_186__4_), .Q(data_36__4_) );
DFFPOSX1 DFFPOSX1_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_186__5_), .Q(data_36__5_) );
DFFPOSX1 DFFPOSX1_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_186__6_), .Q(data_36__6_) );
DFFPOSX1 DFFPOSX1_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_186__7_), .Q(data_36__7_) );
DFFPOSX1 DFFPOSX1_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_186__8_), .Q(data_36__8_) );
DFFPOSX1 DFFPOSX1_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_186__9_), .Q(data_36__9_) );
DFFPOSX1 DFFPOSX1_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_186__10_), .Q(data_36__10_) );
DFFPOSX1 DFFPOSX1_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_186__11_), .Q(data_36__11_) );
DFFPOSX1 DFFPOSX1_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_186__12_), .Q(data_36__12_) );
DFFPOSX1 DFFPOSX1_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_186__13_), .Q(data_36__13_) );
DFFPOSX1 DFFPOSX1_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_186__14_), .Q(data_36__14_) );
DFFPOSX1 DFFPOSX1_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_186__15_), .Q(data_36__15_) );
DFFPOSX1 DFFPOSX1_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_187__0_), .Q(data_37__0_) );
DFFPOSX1 DFFPOSX1_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_187__1_), .Q(data_37__1_) );
DFFPOSX1 DFFPOSX1_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_187__2_), .Q(data_37__2_) );
DFFPOSX1 DFFPOSX1_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_187__3_), .Q(data_37__3_) );
DFFPOSX1 DFFPOSX1_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_187__4_), .Q(data_37__4_) );
DFFPOSX1 DFFPOSX1_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_187__5_), .Q(data_37__5_) );
DFFPOSX1 DFFPOSX1_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_187__6_), .Q(data_37__6_) );
DFFPOSX1 DFFPOSX1_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_187__7_), .Q(data_37__7_) );
DFFPOSX1 DFFPOSX1_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_187__8_), .Q(data_37__8_) );
DFFPOSX1 DFFPOSX1_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_187__9_), .Q(data_37__9_) );
DFFPOSX1 DFFPOSX1_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_187__10_), .Q(data_37__10_) );
DFFPOSX1 DFFPOSX1_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_187__11_), .Q(data_37__11_) );
DFFPOSX1 DFFPOSX1_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_187__12_), .Q(data_37__12_) );
DFFPOSX1 DFFPOSX1_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_187__13_), .Q(data_37__13_) );
DFFPOSX1 DFFPOSX1_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_187__14_), .Q(data_37__14_) );
DFFPOSX1 DFFPOSX1_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_187__15_), .Q(data_37__15_) );
DFFPOSX1 DFFPOSX1_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_188__0_), .Q(data_38__0_) );
DFFPOSX1 DFFPOSX1_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_188__1_), .Q(data_38__1_) );
DFFPOSX1 DFFPOSX1_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_188__2_), .Q(data_38__2_) );
DFFPOSX1 DFFPOSX1_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_188__3_), .Q(data_38__3_) );
DFFPOSX1 DFFPOSX1_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_188__4_), .Q(data_38__4_) );
DFFPOSX1 DFFPOSX1_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_188__5_), .Q(data_38__5_) );
DFFPOSX1 DFFPOSX1_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_188__6_), .Q(data_38__6_) );
DFFPOSX1 DFFPOSX1_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_188__7_), .Q(data_38__7_) );
DFFPOSX1 DFFPOSX1_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_188__8_), .Q(data_38__8_) );
DFFPOSX1 DFFPOSX1_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_188__9_), .Q(data_38__9_) );
DFFPOSX1 DFFPOSX1_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_188__10_), .Q(data_38__10_) );
DFFPOSX1 DFFPOSX1_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_188__11_), .Q(data_38__11_) );
DFFPOSX1 DFFPOSX1_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_188__12_), .Q(data_38__12_) );
DFFPOSX1 DFFPOSX1_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_188__13_), .Q(data_38__13_) );
DFFPOSX1 DFFPOSX1_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_188__14_), .Q(data_38__14_) );
DFFPOSX1 DFFPOSX1_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_188__15_), .Q(data_38__15_) );
DFFPOSX1 DFFPOSX1_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_189__0_), .Q(data_39__0_) );
DFFPOSX1 DFFPOSX1_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_189__1_), .Q(data_39__1_) );
DFFPOSX1 DFFPOSX1_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_189__2_), .Q(data_39__2_) );
DFFPOSX1 DFFPOSX1_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_189__3_), .Q(data_39__3_) );
DFFPOSX1 DFFPOSX1_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_189__4_), .Q(data_39__4_) );
DFFPOSX1 DFFPOSX1_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_189__5_), .Q(data_39__5_) );
DFFPOSX1 DFFPOSX1_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_189__6_), .Q(data_39__6_) );
DFFPOSX1 DFFPOSX1_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_189__7_), .Q(data_39__7_) );
DFFPOSX1 DFFPOSX1_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_189__8_), .Q(data_39__8_) );
DFFPOSX1 DFFPOSX1_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_189__9_), .Q(data_39__9_) );
DFFPOSX1 DFFPOSX1_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_189__10_), .Q(data_39__10_) );
DFFPOSX1 DFFPOSX1_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_189__11_), .Q(data_39__11_) );
DFFPOSX1 DFFPOSX1_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_189__12_), .Q(data_39__12_) );
DFFPOSX1 DFFPOSX1_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_189__13_), .Q(data_39__13_) );
DFFPOSX1 DFFPOSX1_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_189__14_), .Q(data_39__14_) );
DFFPOSX1 DFFPOSX1_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_189__15_), .Q(data_39__15_) );
DFFPOSX1 DFFPOSX1_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_191__0_), .Q(data_40__0_) );
DFFPOSX1 DFFPOSX1_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_191__1_), .Q(data_40__1_) );
DFFPOSX1 DFFPOSX1_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_191__2_), .Q(data_40__2_) );
DFFPOSX1 DFFPOSX1_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_191__3_), .Q(data_40__3_) );
DFFPOSX1 DFFPOSX1_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_191__4_), .Q(data_40__4_) );
DFFPOSX1 DFFPOSX1_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_191__5_), .Q(data_40__5_) );
DFFPOSX1 DFFPOSX1_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_191__6_), .Q(data_40__6_) );
DFFPOSX1 DFFPOSX1_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_191__7_), .Q(data_40__7_) );
DFFPOSX1 DFFPOSX1_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_191__8_), .Q(data_40__8_) );
DFFPOSX1 DFFPOSX1_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_191__9_), .Q(data_40__9_) );
DFFPOSX1 DFFPOSX1_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_191__10_), .Q(data_40__10_) );
DFFPOSX1 DFFPOSX1_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_191__11_), .Q(data_40__11_) );
DFFPOSX1 DFFPOSX1_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_191__12_), .Q(data_40__12_) );
DFFPOSX1 DFFPOSX1_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_191__13_), .Q(data_40__13_) );
DFFPOSX1 DFFPOSX1_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_191__14_), .Q(data_40__14_) );
DFFPOSX1 DFFPOSX1_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_191__15_), .Q(data_40__15_) );
DFFPOSX1 DFFPOSX1_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_192__0_), .Q(data_41__0_) );
DFFPOSX1 DFFPOSX1_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_192__1_), .Q(data_41__1_) );
DFFPOSX1 DFFPOSX1_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_192__2_), .Q(data_41__2_) );
DFFPOSX1 DFFPOSX1_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_192__3_), .Q(data_41__3_) );
DFFPOSX1 DFFPOSX1_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_192__4_), .Q(data_41__4_) );
DFFPOSX1 DFFPOSX1_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_192__5_), .Q(data_41__5_) );
DFFPOSX1 DFFPOSX1_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_192__6_), .Q(data_41__6_) );
DFFPOSX1 DFFPOSX1_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_192__7_), .Q(data_41__7_) );
DFFPOSX1 DFFPOSX1_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_192__8_), .Q(data_41__8_) );
DFFPOSX1 DFFPOSX1_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_192__9_), .Q(data_41__9_) );
DFFPOSX1 DFFPOSX1_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_192__10_), .Q(data_41__10_) );
DFFPOSX1 DFFPOSX1_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_192__11_), .Q(data_41__11_) );
DFFPOSX1 DFFPOSX1_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_192__12_), .Q(data_41__12_) );
DFFPOSX1 DFFPOSX1_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_192__13_), .Q(data_41__13_) );
DFFPOSX1 DFFPOSX1_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_192__14_), .Q(data_41__14_) );
DFFPOSX1 DFFPOSX1_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_192__15_), .Q(data_41__15_) );
DFFPOSX1 DFFPOSX1_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_193__0_), .Q(data_42__0_) );
DFFPOSX1 DFFPOSX1_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_193__1_), .Q(data_42__1_) );
DFFPOSX1 DFFPOSX1_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_193__2_), .Q(data_42__2_) );
DFFPOSX1 DFFPOSX1_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_193__3_), .Q(data_42__3_) );
DFFPOSX1 DFFPOSX1_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_193__4_), .Q(data_42__4_) );
DFFPOSX1 DFFPOSX1_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_193__5_), .Q(data_42__5_) );
DFFPOSX1 DFFPOSX1_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_193__6_), .Q(data_42__6_) );
DFFPOSX1 DFFPOSX1_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_193__7_), .Q(data_42__7_) );
DFFPOSX1 DFFPOSX1_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_193__8_), .Q(data_42__8_) );
DFFPOSX1 DFFPOSX1_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_193__9_), .Q(data_42__9_) );
DFFPOSX1 DFFPOSX1_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_193__10_), .Q(data_42__10_) );
DFFPOSX1 DFFPOSX1_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_193__11_), .Q(data_42__11_) );
DFFPOSX1 DFFPOSX1_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_193__12_), .Q(data_42__12_) );
DFFPOSX1 DFFPOSX1_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_193__13_), .Q(data_42__13_) );
DFFPOSX1 DFFPOSX1_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_193__14_), .Q(data_42__14_) );
DFFPOSX1 DFFPOSX1_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_193__15_), .Q(data_42__15_) );
DFFPOSX1 DFFPOSX1_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_194__0_), .Q(data_43__0_) );
DFFPOSX1 DFFPOSX1_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_194__1_), .Q(data_43__1_) );
DFFPOSX1 DFFPOSX1_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_194__2_), .Q(data_43__2_) );
DFFPOSX1 DFFPOSX1_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_194__3_), .Q(data_43__3_) );
DFFPOSX1 DFFPOSX1_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_194__4_), .Q(data_43__4_) );
DFFPOSX1 DFFPOSX1_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_194__5_), .Q(data_43__5_) );
DFFPOSX1 DFFPOSX1_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_194__6_), .Q(data_43__6_) );
DFFPOSX1 DFFPOSX1_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_194__7_), .Q(data_43__7_) );
DFFPOSX1 DFFPOSX1_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_194__8_), .Q(data_43__8_) );
DFFPOSX1 DFFPOSX1_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_194__9_), .Q(data_43__9_) );
DFFPOSX1 DFFPOSX1_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_194__10_), .Q(data_43__10_) );
DFFPOSX1 DFFPOSX1_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_194__11_), .Q(data_43__11_) );
DFFPOSX1 DFFPOSX1_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_194__12_), .Q(data_43__12_) );
DFFPOSX1 DFFPOSX1_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_194__13_), .Q(data_43__13_) );
DFFPOSX1 DFFPOSX1_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_194__14_), .Q(data_43__14_) );
DFFPOSX1 DFFPOSX1_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_194__15_), .Q(data_43__15_) );
DFFPOSX1 DFFPOSX1_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_195__0_), .Q(data_44__0_) );
DFFPOSX1 DFFPOSX1_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_195__1_), .Q(data_44__1_) );
DFFPOSX1 DFFPOSX1_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_195__2_), .Q(data_44__2_) );
DFFPOSX1 DFFPOSX1_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_195__3_), .Q(data_44__3_) );
DFFPOSX1 DFFPOSX1_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_195__4_), .Q(data_44__4_) );
DFFPOSX1 DFFPOSX1_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_195__5_), .Q(data_44__5_) );
DFFPOSX1 DFFPOSX1_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_195__6_), .Q(data_44__6_) );
DFFPOSX1 DFFPOSX1_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_195__7_), .Q(data_44__7_) );
DFFPOSX1 DFFPOSX1_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_195__8_), .Q(data_44__8_) );
DFFPOSX1 DFFPOSX1_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_195__9_), .Q(data_44__9_) );
DFFPOSX1 DFFPOSX1_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_195__10_), .Q(data_44__10_) );
DFFPOSX1 DFFPOSX1_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_195__11_), .Q(data_44__11_) );
DFFPOSX1 DFFPOSX1_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_195__12_), .Q(data_44__12_) );
DFFPOSX1 DFFPOSX1_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_195__13_), .Q(data_44__13_) );
DFFPOSX1 DFFPOSX1_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_195__14_), .Q(data_44__14_) );
DFFPOSX1 DFFPOSX1_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_195__15_), .Q(data_44__15_) );
DFFPOSX1 DFFPOSX1_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_196__0_), .Q(data_45__0_) );
DFFPOSX1 DFFPOSX1_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_196__1_), .Q(data_45__1_) );
DFFPOSX1 DFFPOSX1_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_196__2_), .Q(data_45__2_) );
DFFPOSX1 DFFPOSX1_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_196__3_), .Q(data_45__3_) );
DFFPOSX1 DFFPOSX1_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_196__4_), .Q(data_45__4_) );
DFFPOSX1 DFFPOSX1_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_196__5_), .Q(data_45__5_) );
DFFPOSX1 DFFPOSX1_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_196__6_), .Q(data_45__6_) );
DFFPOSX1 DFFPOSX1_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_196__7_), .Q(data_45__7_) );
DFFPOSX1 DFFPOSX1_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_196__8_), .Q(data_45__8_) );
DFFPOSX1 DFFPOSX1_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_196__9_), .Q(data_45__9_) );
DFFPOSX1 DFFPOSX1_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_196__10_), .Q(data_45__10_) );
DFFPOSX1 DFFPOSX1_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_196__11_), .Q(data_45__11_) );
DFFPOSX1 DFFPOSX1_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_196__12_), .Q(data_45__12_) );
DFFPOSX1 DFFPOSX1_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_196__13_), .Q(data_45__13_) );
DFFPOSX1 DFFPOSX1_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_196__14_), .Q(data_45__14_) );
DFFPOSX1 DFFPOSX1_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_196__15_), .Q(data_45__15_) );
DFFPOSX1 DFFPOSX1_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_197__0_), .Q(data_46__0_) );
DFFPOSX1 DFFPOSX1_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_197__1_), .Q(data_46__1_) );
DFFPOSX1 DFFPOSX1_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_197__2_), .Q(data_46__2_) );
DFFPOSX1 DFFPOSX1_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_197__3_), .Q(data_46__3_) );
DFFPOSX1 DFFPOSX1_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_197__4_), .Q(data_46__4_) );
DFFPOSX1 DFFPOSX1_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_197__5_), .Q(data_46__5_) );
DFFPOSX1 DFFPOSX1_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_197__6_), .Q(data_46__6_) );
DFFPOSX1 DFFPOSX1_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_197__7_), .Q(data_46__7_) );
DFFPOSX1 DFFPOSX1_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_197__8_), .Q(data_46__8_) );
DFFPOSX1 DFFPOSX1_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_197__9_), .Q(data_46__9_) );
DFFPOSX1 DFFPOSX1_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_197__10_), .Q(data_46__10_) );
DFFPOSX1 DFFPOSX1_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_197__11_), .Q(data_46__11_) );
DFFPOSX1 DFFPOSX1_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_197__12_), .Q(data_46__12_) );
DFFPOSX1 DFFPOSX1_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_197__13_), .Q(data_46__13_) );
DFFPOSX1 DFFPOSX1_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_197__14_), .Q(data_46__14_) );
DFFPOSX1 DFFPOSX1_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_197__15_), .Q(data_46__15_) );
DFFPOSX1 DFFPOSX1_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf0), .D(_198__0_), .Q(data_47__0_) );
DFFPOSX1 DFFPOSX1_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf0), .D(_198__1_), .Q(data_47__1_) );
DFFPOSX1 DFFPOSX1_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf0), .D(_198__2_), .Q(data_47__2_) );
DFFPOSX1 DFFPOSX1_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf0), .D(_198__3_), .Q(data_47__3_) );
DFFPOSX1 DFFPOSX1_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf0), .D(_198__4_), .Q(data_47__4_) );
DFFPOSX1 DFFPOSX1_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf0), .D(_198__5_), .Q(data_47__5_) );
DFFPOSX1 DFFPOSX1_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf0), .D(_198__6_), .Q(data_47__6_) );
DFFPOSX1 DFFPOSX1_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf0), .D(_198__7_), .Q(data_47__7_) );
DFFPOSX1 DFFPOSX1_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf0), .D(_198__8_), .Q(data_47__8_) );
DFFPOSX1 DFFPOSX1_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf0), .D(_198__9_), .Q(data_47__9_) );
DFFPOSX1 DFFPOSX1_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf0), .D(_198__10_), .Q(data_47__10_) );
DFFPOSX1 DFFPOSX1_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf0), .D(_198__11_), .Q(data_47__11_) );
DFFPOSX1 DFFPOSX1_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf0), .D(_198__12_), .Q(data_47__12_) );
DFFPOSX1 DFFPOSX1_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf0), .D(_198__13_), .Q(data_47__13_) );
DFFPOSX1 DFFPOSX1_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf0), .D(_198__14_), .Q(data_47__14_) );
DFFPOSX1 DFFPOSX1_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf0), .D(_198__15_), .Q(data_47__15_) );
DFFPOSX1 DFFPOSX1_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_199__0_), .Q(data_48__0_) );
DFFPOSX1 DFFPOSX1_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_199__1_), .Q(data_48__1_) );
DFFPOSX1 DFFPOSX1_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_199__2_), .Q(data_48__2_) );
DFFPOSX1 DFFPOSX1_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_199__3_), .Q(data_48__3_) );
DFFPOSX1 DFFPOSX1_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_199__4_), .Q(data_48__4_) );
DFFPOSX1 DFFPOSX1_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_199__5_), .Q(data_48__5_) );
DFFPOSX1 DFFPOSX1_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_199__6_), .Q(data_48__6_) );
DFFPOSX1 DFFPOSX1_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_199__7_), .Q(data_48__7_) );
DFFPOSX1 DFFPOSX1_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_199__8_), .Q(data_48__8_) );
DFFPOSX1 DFFPOSX1_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_199__9_), .Q(data_48__9_) );
DFFPOSX1 DFFPOSX1_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_199__10_), .Q(data_48__10_) );
DFFPOSX1 DFFPOSX1_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_199__11_), .Q(data_48__11_) );
DFFPOSX1 DFFPOSX1_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_199__12_), .Q(data_48__12_) );
DFFPOSX1 DFFPOSX1_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_199__13_), .Q(data_48__13_) );
DFFPOSX1 DFFPOSX1_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_199__14_), .Q(data_48__14_) );
DFFPOSX1 DFFPOSX1_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_199__15_), .Q(data_48__15_) );
DFFPOSX1 DFFPOSX1_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_200__0_), .Q(data_49__0_) );
DFFPOSX1 DFFPOSX1_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_200__1_), .Q(data_49__1_) );
DFFPOSX1 DFFPOSX1_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_200__2_), .Q(data_49__2_) );
DFFPOSX1 DFFPOSX1_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_200__3_), .Q(data_49__3_) );
DFFPOSX1 DFFPOSX1_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_200__4_), .Q(data_49__4_) );
DFFPOSX1 DFFPOSX1_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_200__5_), .Q(data_49__5_) );
DFFPOSX1 DFFPOSX1_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_200__6_), .Q(data_49__6_) );
DFFPOSX1 DFFPOSX1_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_200__7_), .Q(data_49__7_) );
DFFPOSX1 DFFPOSX1_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_200__8_), .Q(data_49__8_) );
DFFPOSX1 DFFPOSX1_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_200__9_), .Q(data_49__9_) );
DFFPOSX1 DFFPOSX1_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_200__10_), .Q(data_49__10_) );
DFFPOSX1 DFFPOSX1_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_200__11_), .Q(data_49__11_) );
DFFPOSX1 DFFPOSX1_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_200__12_), .Q(data_49__12_) );
DFFPOSX1 DFFPOSX1_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_200__13_), .Q(data_49__13_) );
DFFPOSX1 DFFPOSX1_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_200__14_), .Q(data_49__14_) );
DFFPOSX1 DFFPOSX1_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_200__15_), .Q(data_49__15_) );
DFFPOSX1 DFFPOSX1_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_202__0_), .Q(data_50__0_) );
DFFPOSX1 DFFPOSX1_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_202__1_), .Q(data_50__1_) );
DFFPOSX1 DFFPOSX1_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_202__2_), .Q(data_50__2_) );
DFFPOSX1 DFFPOSX1_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_202__3_), .Q(data_50__3_) );
DFFPOSX1 DFFPOSX1_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_202__4_), .Q(data_50__4_) );
DFFPOSX1 DFFPOSX1_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_202__5_), .Q(data_50__5_) );
DFFPOSX1 DFFPOSX1_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_202__6_), .Q(data_50__6_) );
DFFPOSX1 DFFPOSX1_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_202__7_), .Q(data_50__7_) );
DFFPOSX1 DFFPOSX1_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_202__8_), .Q(data_50__8_) );
DFFPOSX1 DFFPOSX1_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_202__9_), .Q(data_50__9_) );
DFFPOSX1 DFFPOSX1_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_202__10_), .Q(data_50__10_) );
DFFPOSX1 DFFPOSX1_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_202__11_), .Q(data_50__11_) );
DFFPOSX1 DFFPOSX1_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_202__12_), .Q(data_50__12_) );
DFFPOSX1 DFFPOSX1_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_202__13_), .Q(data_50__13_) );
DFFPOSX1 DFFPOSX1_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_202__14_), .Q(data_50__14_) );
DFFPOSX1 DFFPOSX1_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_202__15_), .Q(data_50__15_) );
DFFPOSX1 DFFPOSX1_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_203__0_), .Q(data_51__0_) );
DFFPOSX1 DFFPOSX1_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_203__1_), .Q(data_51__1_) );
DFFPOSX1 DFFPOSX1_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_203__2_), .Q(data_51__2_) );
DFFPOSX1 DFFPOSX1_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_203__3_), .Q(data_51__3_) );
DFFPOSX1 DFFPOSX1_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_203__4_), .Q(data_51__4_) );
DFFPOSX1 DFFPOSX1_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_203__5_), .Q(data_51__5_) );
DFFPOSX1 DFFPOSX1_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_203__6_), .Q(data_51__6_) );
DFFPOSX1 DFFPOSX1_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_203__7_), .Q(data_51__7_) );
DFFPOSX1 DFFPOSX1_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_203__8_), .Q(data_51__8_) );
DFFPOSX1 DFFPOSX1_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_203__9_), .Q(data_51__9_) );
DFFPOSX1 DFFPOSX1_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_203__10_), .Q(data_51__10_) );
DFFPOSX1 DFFPOSX1_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_203__11_), .Q(data_51__11_) );
DFFPOSX1 DFFPOSX1_845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_203__12_), .Q(data_51__12_) );
DFFPOSX1 DFFPOSX1_846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_203__13_), .Q(data_51__13_) );
DFFPOSX1 DFFPOSX1_847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_203__14_), .Q(data_51__14_) );
DFFPOSX1 DFFPOSX1_848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_203__15_), .Q(data_51__15_) );
DFFPOSX1 DFFPOSX1_849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_204__0_), .Q(data_52__0_) );
DFFPOSX1 DFFPOSX1_850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_204__1_), .Q(data_52__1_) );
DFFPOSX1 DFFPOSX1_851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_204__2_), .Q(data_52__2_) );
DFFPOSX1 DFFPOSX1_852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_204__3_), .Q(data_52__3_) );
DFFPOSX1 DFFPOSX1_853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_204__4_), .Q(data_52__4_) );
DFFPOSX1 DFFPOSX1_854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_204__5_), .Q(data_52__5_) );
DFFPOSX1 DFFPOSX1_855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_204__6_), .Q(data_52__6_) );
DFFPOSX1 DFFPOSX1_856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_204__7_), .Q(data_52__7_) );
DFFPOSX1 DFFPOSX1_857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_204__8_), .Q(data_52__8_) );
DFFPOSX1 DFFPOSX1_858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_204__9_), .Q(data_52__9_) );
DFFPOSX1 DFFPOSX1_859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_204__10_), .Q(data_52__10_) );
DFFPOSX1 DFFPOSX1_860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_204__11_), .Q(data_52__11_) );
DFFPOSX1 DFFPOSX1_861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_204__12_), .Q(data_52__12_) );
DFFPOSX1 DFFPOSX1_862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_204__13_), .Q(data_52__13_) );
DFFPOSX1 DFFPOSX1_863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_204__14_), .Q(data_52__14_) );
DFFPOSX1 DFFPOSX1_864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_204__15_), .Q(data_52__15_) );
DFFPOSX1 DFFPOSX1_865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_205__0_), .Q(data_53__0_) );
DFFPOSX1 DFFPOSX1_866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_205__1_), .Q(data_53__1_) );
DFFPOSX1 DFFPOSX1_867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_205__2_), .Q(data_53__2_) );
DFFPOSX1 DFFPOSX1_868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_205__3_), .Q(data_53__3_) );
DFFPOSX1 DFFPOSX1_869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_205__4_), .Q(data_53__4_) );
DFFPOSX1 DFFPOSX1_870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_205__5_), .Q(data_53__5_) );
DFFPOSX1 DFFPOSX1_871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_205__6_), .Q(data_53__6_) );
DFFPOSX1 DFFPOSX1_872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_205__7_), .Q(data_53__7_) );
DFFPOSX1 DFFPOSX1_873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_205__8_), .Q(data_53__8_) );
DFFPOSX1 DFFPOSX1_874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_205__9_), .Q(data_53__9_) );
DFFPOSX1 DFFPOSX1_875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_205__10_), .Q(data_53__10_) );
DFFPOSX1 DFFPOSX1_876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_205__11_), .Q(data_53__11_) );
DFFPOSX1 DFFPOSX1_877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_205__12_), .Q(data_53__12_) );
DFFPOSX1 DFFPOSX1_878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_205__13_), .Q(data_53__13_) );
DFFPOSX1 DFFPOSX1_879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_205__14_), .Q(data_53__14_) );
DFFPOSX1 DFFPOSX1_880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_205__15_), .Q(data_53__15_) );
DFFPOSX1 DFFPOSX1_881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_206__0_), .Q(data_54__0_) );
DFFPOSX1 DFFPOSX1_882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_206__1_), .Q(data_54__1_) );
DFFPOSX1 DFFPOSX1_883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_206__2_), .Q(data_54__2_) );
DFFPOSX1 DFFPOSX1_884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_206__3_), .Q(data_54__3_) );
DFFPOSX1 DFFPOSX1_885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_206__4_), .Q(data_54__4_) );
DFFPOSX1 DFFPOSX1_886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_206__5_), .Q(data_54__5_) );
DFFPOSX1 DFFPOSX1_887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_206__6_), .Q(data_54__6_) );
DFFPOSX1 DFFPOSX1_888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_206__7_), .Q(data_54__7_) );
DFFPOSX1 DFFPOSX1_889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_206__8_), .Q(data_54__8_) );
DFFPOSX1 DFFPOSX1_890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_206__9_), .Q(data_54__9_) );
DFFPOSX1 DFFPOSX1_891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_206__10_), .Q(data_54__10_) );
DFFPOSX1 DFFPOSX1_892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_206__11_), .Q(data_54__11_) );
DFFPOSX1 DFFPOSX1_893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_206__12_), .Q(data_54__12_) );
DFFPOSX1 DFFPOSX1_894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_206__13_), .Q(data_54__13_) );
DFFPOSX1 DFFPOSX1_895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_206__14_), .Q(data_54__14_) );
DFFPOSX1 DFFPOSX1_896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_206__15_), .Q(data_54__15_) );
DFFPOSX1 DFFPOSX1_897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_207__0_), .Q(data_55__0_) );
DFFPOSX1 DFFPOSX1_898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_207__1_), .Q(data_55__1_) );
DFFPOSX1 DFFPOSX1_899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_207__2_), .Q(data_55__2_) );
DFFPOSX1 DFFPOSX1_900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_207__3_), .Q(data_55__3_) );
DFFPOSX1 DFFPOSX1_901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_207__4_), .Q(data_55__4_) );
DFFPOSX1 DFFPOSX1_902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_207__5_), .Q(data_55__5_) );
DFFPOSX1 DFFPOSX1_903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_207__6_), .Q(data_55__6_) );
DFFPOSX1 DFFPOSX1_904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_207__7_), .Q(data_55__7_) );
DFFPOSX1 DFFPOSX1_905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_207__8_), .Q(data_55__8_) );
DFFPOSX1 DFFPOSX1_906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_207__9_), .Q(data_55__9_) );
DFFPOSX1 DFFPOSX1_907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_207__10_), .Q(data_55__10_) );
DFFPOSX1 DFFPOSX1_908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_207__11_), .Q(data_55__11_) );
DFFPOSX1 DFFPOSX1_909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_207__12_), .Q(data_55__12_) );
DFFPOSX1 DFFPOSX1_910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_207__13_), .Q(data_55__13_) );
DFFPOSX1 DFFPOSX1_911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_207__14_), .Q(data_55__14_) );
DFFPOSX1 DFFPOSX1_912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_207__15_), .Q(data_55__15_) );
DFFPOSX1 DFFPOSX1_913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_208__0_), .Q(data_56__0_) );
DFFPOSX1 DFFPOSX1_914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_208__1_), .Q(data_56__1_) );
DFFPOSX1 DFFPOSX1_915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_208__2_), .Q(data_56__2_) );
DFFPOSX1 DFFPOSX1_916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_208__3_), .Q(data_56__3_) );
DFFPOSX1 DFFPOSX1_917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_208__4_), .Q(data_56__4_) );
DFFPOSX1 DFFPOSX1_918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_208__5_), .Q(data_56__5_) );
DFFPOSX1 DFFPOSX1_919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_208__6_), .Q(data_56__6_) );
DFFPOSX1 DFFPOSX1_920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_208__7_), .Q(data_56__7_) );
DFFPOSX1 DFFPOSX1_921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_208__8_), .Q(data_56__8_) );
DFFPOSX1 DFFPOSX1_922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_208__9_), .Q(data_56__9_) );
DFFPOSX1 DFFPOSX1_923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_208__10_), .Q(data_56__10_) );
DFFPOSX1 DFFPOSX1_924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_208__11_), .Q(data_56__11_) );
DFFPOSX1 DFFPOSX1_925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_208__12_), .Q(data_56__12_) );
DFFPOSX1 DFFPOSX1_926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_208__13_), .Q(data_56__13_) );
DFFPOSX1 DFFPOSX1_927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_208__14_), .Q(data_56__14_) );
DFFPOSX1 DFFPOSX1_928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_208__15_), .Q(data_56__15_) );
DFFPOSX1 DFFPOSX1_929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_209__0_), .Q(data_57__0_) );
DFFPOSX1 DFFPOSX1_930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_209__1_), .Q(data_57__1_) );
DFFPOSX1 DFFPOSX1_931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_209__2_), .Q(data_57__2_) );
DFFPOSX1 DFFPOSX1_932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_209__3_), .Q(data_57__3_) );
DFFPOSX1 DFFPOSX1_933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_209__4_), .Q(data_57__4_) );
DFFPOSX1 DFFPOSX1_934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_209__5_), .Q(data_57__5_) );
DFFPOSX1 DFFPOSX1_935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_209__6_), .Q(data_57__6_) );
DFFPOSX1 DFFPOSX1_936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_209__7_), .Q(data_57__7_) );
DFFPOSX1 DFFPOSX1_937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_209__8_), .Q(data_57__8_) );
DFFPOSX1 DFFPOSX1_938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_209__9_), .Q(data_57__9_) );
DFFPOSX1 DFFPOSX1_939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_209__10_), .Q(data_57__10_) );
DFFPOSX1 DFFPOSX1_940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_209__11_), .Q(data_57__11_) );
DFFPOSX1 DFFPOSX1_941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_209__12_), .Q(data_57__12_) );
DFFPOSX1 DFFPOSX1_942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_209__13_), .Q(data_57__13_) );
DFFPOSX1 DFFPOSX1_943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_209__14_), .Q(data_57__14_) );
DFFPOSX1 DFFPOSX1_944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_209__15_), .Q(data_57__15_) );
DFFPOSX1 DFFPOSX1_945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_210__0_), .Q(data_58__0_) );
DFFPOSX1 DFFPOSX1_946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_210__1_), .Q(data_58__1_) );
DFFPOSX1 DFFPOSX1_947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_210__2_), .Q(data_58__2_) );
DFFPOSX1 DFFPOSX1_948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_210__3_), .Q(data_58__3_) );
DFFPOSX1 DFFPOSX1_949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_210__4_), .Q(data_58__4_) );
DFFPOSX1 DFFPOSX1_950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_210__5_), .Q(data_58__5_) );
DFFPOSX1 DFFPOSX1_951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_210__6_), .Q(data_58__6_) );
DFFPOSX1 DFFPOSX1_952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_210__7_), .Q(data_58__7_) );
DFFPOSX1 DFFPOSX1_953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_210__8_), .Q(data_58__8_) );
DFFPOSX1 DFFPOSX1_954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_210__9_), .Q(data_58__9_) );
DFFPOSX1 DFFPOSX1_955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_210__10_), .Q(data_58__10_) );
DFFPOSX1 DFFPOSX1_956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_210__11_), .Q(data_58__11_) );
DFFPOSX1 DFFPOSX1_957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_210__12_), .Q(data_58__12_) );
DFFPOSX1 DFFPOSX1_958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_210__13_), .Q(data_58__13_) );
DFFPOSX1 DFFPOSX1_959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_210__14_), .Q(data_58__14_) );
DFFPOSX1 DFFPOSX1_960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_210__15_), .Q(data_58__15_) );
DFFPOSX1 DFFPOSX1_961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_211__0_), .Q(data_59__0_) );
DFFPOSX1 DFFPOSX1_962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_211__1_), .Q(data_59__1_) );
DFFPOSX1 DFFPOSX1_963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_211__2_), .Q(data_59__2_) );
DFFPOSX1 DFFPOSX1_964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_211__3_), .Q(data_59__3_) );
DFFPOSX1 DFFPOSX1_965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_211__4_), .Q(data_59__4_) );
DFFPOSX1 DFFPOSX1_966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_211__5_), .Q(data_59__5_) );
DFFPOSX1 DFFPOSX1_967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_211__6_), .Q(data_59__6_) );
DFFPOSX1 DFFPOSX1_968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_211__7_), .Q(data_59__7_) );
DFFPOSX1 DFFPOSX1_969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_211__8_), .Q(data_59__8_) );
DFFPOSX1 DFFPOSX1_970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_211__9_), .Q(data_59__9_) );
DFFPOSX1 DFFPOSX1_971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_211__10_), .Q(data_59__10_) );
DFFPOSX1 DFFPOSX1_972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_211__11_), .Q(data_59__11_) );
DFFPOSX1 DFFPOSX1_973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_211__12_), .Q(data_59__12_) );
DFFPOSX1 DFFPOSX1_974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_211__13_), .Q(data_59__13_) );
DFFPOSX1 DFFPOSX1_975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_211__14_), .Q(data_59__14_) );
DFFPOSX1 DFFPOSX1_976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_211__15_), .Q(data_59__15_) );
DFFPOSX1 DFFPOSX1_977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_213__0_), .Q(data_60__0_) );
DFFPOSX1 DFFPOSX1_978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_213__1_), .Q(data_60__1_) );
DFFPOSX1 DFFPOSX1_979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_213__2_), .Q(data_60__2_) );
DFFPOSX1 DFFPOSX1_980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_213__3_), .Q(data_60__3_) );
DFFPOSX1 DFFPOSX1_981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_213__4_), .Q(data_60__4_) );
DFFPOSX1 DFFPOSX1_982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_213__5_), .Q(data_60__5_) );
DFFPOSX1 DFFPOSX1_983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_213__6_), .Q(data_60__6_) );
DFFPOSX1 DFFPOSX1_984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_213__7_), .Q(data_60__7_) );
DFFPOSX1 DFFPOSX1_985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_213__8_), .Q(data_60__8_) );
DFFPOSX1 DFFPOSX1_986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_213__9_), .Q(data_60__9_) );
DFFPOSX1 DFFPOSX1_987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_213__10_), .Q(data_60__10_) );
DFFPOSX1 DFFPOSX1_988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_213__11_), .Q(data_60__11_) );
DFFPOSX1 DFFPOSX1_989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_213__12_), .Q(data_60__12_) );
DFFPOSX1 DFFPOSX1_990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_213__13_), .Q(data_60__13_) );
DFFPOSX1 DFFPOSX1_991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_213__14_), .Q(data_60__14_) );
DFFPOSX1 DFFPOSX1_992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_213__15_), .Q(data_60__15_) );
DFFPOSX1 DFFPOSX1_993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_214__0_), .Q(data_61__0_) );
DFFPOSX1 DFFPOSX1_994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_214__1_), .Q(data_61__1_) );
DFFPOSX1 DFFPOSX1_995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_214__2_), .Q(data_61__2_) );
DFFPOSX1 DFFPOSX1_996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_214__3_), .Q(data_61__3_) );
DFFPOSX1 DFFPOSX1_997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_214__4_), .Q(data_61__4_) );
DFFPOSX1 DFFPOSX1_998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_214__5_), .Q(data_61__5_) );
DFFPOSX1 DFFPOSX1_999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_214__6_), .Q(data_61__6_) );
DFFPOSX1 DFFPOSX1_1000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_214__7_), .Q(data_61__7_) );
DFFPOSX1 DFFPOSX1_1001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_214__8_), .Q(data_61__8_) );
DFFPOSX1 DFFPOSX1_1002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_214__9_), .Q(data_61__9_) );
DFFPOSX1 DFFPOSX1_1003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_214__10_), .Q(data_61__10_) );
DFFPOSX1 DFFPOSX1_1004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_214__11_), .Q(data_61__11_) );
DFFPOSX1 DFFPOSX1_1005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_214__12_), .Q(data_61__12_) );
DFFPOSX1 DFFPOSX1_1006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_214__13_), .Q(data_61__13_) );
DFFPOSX1 DFFPOSX1_1007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_214__14_), .Q(data_61__14_) );
DFFPOSX1 DFFPOSX1_1008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_214__15_), .Q(data_61__15_) );
DFFPOSX1 DFFPOSX1_1009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_215__0_), .Q(data_62__0_) );
DFFPOSX1 DFFPOSX1_1010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_215__1_), .Q(data_62__1_) );
DFFPOSX1 DFFPOSX1_1011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_215__2_), .Q(data_62__2_) );
DFFPOSX1 DFFPOSX1_1012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_215__3_), .Q(data_62__3_) );
DFFPOSX1 DFFPOSX1_1013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_215__4_), .Q(data_62__4_) );
DFFPOSX1 DFFPOSX1_1014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_215__5_), .Q(data_62__5_) );
DFFPOSX1 DFFPOSX1_1015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_215__6_), .Q(data_62__6_) );
DFFPOSX1 DFFPOSX1_1016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_215__7_), .Q(data_62__7_) );
DFFPOSX1 DFFPOSX1_1017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_215__8_), .Q(data_62__8_) );
DFFPOSX1 DFFPOSX1_1018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_215__9_), .Q(data_62__9_) );
DFFPOSX1 DFFPOSX1_1019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_215__10_), .Q(data_62__10_) );
DFFPOSX1 DFFPOSX1_1020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_215__11_), .Q(data_62__11_) );
DFFPOSX1 DFFPOSX1_1021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_215__12_), .Q(data_62__12_) );
DFFPOSX1 DFFPOSX1_1022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_215__13_), .Q(data_62__13_) );
DFFPOSX1 DFFPOSX1_1023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_215__14_), .Q(data_62__14_) );
DFFPOSX1 DFFPOSX1_1024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_215__15_), .Q(data_62__15_) );
DFFPOSX1 DFFPOSX1_1025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf3), .D(_216__0_), .Q(data_63__0_) );
DFFPOSX1 DFFPOSX1_1026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf3), .D(_216__1_), .Q(data_63__1_) );
DFFPOSX1 DFFPOSX1_1027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf3), .D(_216__2_), .Q(data_63__2_) );
DFFPOSX1 DFFPOSX1_1028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf3), .D(_216__3_), .Q(data_63__3_) );
DFFPOSX1 DFFPOSX1_1029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf3), .D(_216__4_), .Q(data_63__4_) );
DFFPOSX1 DFFPOSX1_1030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf3), .D(_216__5_), .Q(data_63__5_) );
DFFPOSX1 DFFPOSX1_1031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf3), .D(_216__6_), .Q(data_63__6_) );
DFFPOSX1 DFFPOSX1_1032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf3), .D(_216__7_), .Q(data_63__7_) );
DFFPOSX1 DFFPOSX1_1033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf3), .D(_216__8_), .Q(data_63__8_) );
DFFPOSX1 DFFPOSX1_1034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf3), .D(_216__9_), .Q(data_63__9_) );
DFFPOSX1 DFFPOSX1_1035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf3), .D(_216__10_), .Q(data_63__10_) );
DFFPOSX1 DFFPOSX1_1036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf3), .D(_216__11_), .Q(data_63__11_) );
DFFPOSX1 DFFPOSX1_1037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf3), .D(_216__12_), .Q(data_63__12_) );
DFFPOSX1 DFFPOSX1_1038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf3), .D(_216__13_), .Q(data_63__13_) );
DFFPOSX1 DFFPOSX1_1039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf3), .D(_216__14_), .Q(data_63__14_) );
DFFPOSX1 DFFPOSX1_1040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf3), .D(_216__15_), .Q(data_63__15_) );
DFFPOSX1 DFFPOSX1_1041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_217__0_), .Q(data_64__0_) );
DFFPOSX1 DFFPOSX1_1042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_217__1_), .Q(data_64__1_) );
DFFPOSX1 DFFPOSX1_1043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_217__2_), .Q(data_64__2_) );
DFFPOSX1 DFFPOSX1_1044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_217__3_), .Q(data_64__3_) );
DFFPOSX1 DFFPOSX1_1045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_217__4_), .Q(data_64__4_) );
DFFPOSX1 DFFPOSX1_1046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_217__5_), .Q(data_64__5_) );
DFFPOSX1 DFFPOSX1_1047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_217__6_), .Q(data_64__6_) );
DFFPOSX1 DFFPOSX1_1048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_217__7_), .Q(data_64__7_) );
DFFPOSX1 DFFPOSX1_1049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_217__8_), .Q(data_64__8_) );
DFFPOSX1 DFFPOSX1_1050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_217__9_), .Q(data_64__9_) );
DFFPOSX1 DFFPOSX1_1051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_217__10_), .Q(data_64__10_) );
DFFPOSX1 DFFPOSX1_1052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_217__11_), .Q(data_64__11_) );
DFFPOSX1 DFFPOSX1_1053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_217__12_), .Q(data_64__12_) );
DFFPOSX1 DFFPOSX1_1054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_217__13_), .Q(data_64__13_) );
DFFPOSX1 DFFPOSX1_1055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_217__14_), .Q(data_64__14_) );
DFFPOSX1 DFFPOSX1_1056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_217__15_), .Q(data_64__15_) );
DFFPOSX1 DFFPOSX1_1057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_218__0_), .Q(data_65__0_) );
DFFPOSX1 DFFPOSX1_1058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_218__1_), .Q(data_65__1_) );
DFFPOSX1 DFFPOSX1_1059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_218__2_), .Q(data_65__2_) );
DFFPOSX1 DFFPOSX1_1060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_218__3_), .Q(data_65__3_) );
DFFPOSX1 DFFPOSX1_1061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_218__4_), .Q(data_65__4_) );
DFFPOSX1 DFFPOSX1_1062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_218__5_), .Q(data_65__5_) );
DFFPOSX1 DFFPOSX1_1063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_218__6_), .Q(data_65__6_) );
DFFPOSX1 DFFPOSX1_1064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_218__7_), .Q(data_65__7_) );
DFFPOSX1 DFFPOSX1_1065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_218__8_), .Q(data_65__8_) );
DFFPOSX1 DFFPOSX1_1066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_218__9_), .Q(data_65__9_) );
DFFPOSX1 DFFPOSX1_1067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_218__10_), .Q(data_65__10_) );
DFFPOSX1 DFFPOSX1_1068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_218__11_), .Q(data_65__11_) );
DFFPOSX1 DFFPOSX1_1069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_218__12_), .Q(data_65__12_) );
DFFPOSX1 DFFPOSX1_1070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_218__13_), .Q(data_65__13_) );
DFFPOSX1 DFFPOSX1_1071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_218__14_), .Q(data_65__14_) );
DFFPOSX1 DFFPOSX1_1072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_218__15_), .Q(data_65__15_) );
DFFPOSX1 DFFPOSX1_1073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_219__0_), .Q(data_66__0_) );
DFFPOSX1 DFFPOSX1_1074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_219__1_), .Q(data_66__1_) );
DFFPOSX1 DFFPOSX1_1075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_219__2_), .Q(data_66__2_) );
DFFPOSX1 DFFPOSX1_1076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_219__3_), .Q(data_66__3_) );
DFFPOSX1 DFFPOSX1_1077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_219__4_), .Q(data_66__4_) );
DFFPOSX1 DFFPOSX1_1078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_219__5_), .Q(data_66__5_) );
DFFPOSX1 DFFPOSX1_1079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_219__6_), .Q(data_66__6_) );
DFFPOSX1 DFFPOSX1_1080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_219__7_), .Q(data_66__7_) );
DFFPOSX1 DFFPOSX1_1081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_219__8_), .Q(data_66__8_) );
DFFPOSX1 DFFPOSX1_1082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_219__9_), .Q(data_66__9_) );
DFFPOSX1 DFFPOSX1_1083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_219__10_), .Q(data_66__10_) );
DFFPOSX1 DFFPOSX1_1084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_219__11_), .Q(data_66__11_) );
DFFPOSX1 DFFPOSX1_1085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_219__12_), .Q(data_66__12_) );
DFFPOSX1 DFFPOSX1_1086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_219__13_), .Q(data_66__13_) );
DFFPOSX1 DFFPOSX1_1087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_219__14_), .Q(data_66__14_) );
DFFPOSX1 DFFPOSX1_1088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_219__15_), .Q(data_66__15_) );
DFFPOSX1 DFFPOSX1_1089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_220__0_), .Q(data_67__0_) );
DFFPOSX1 DFFPOSX1_1090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_220__1_), .Q(data_67__1_) );
DFFPOSX1 DFFPOSX1_1091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_220__2_), .Q(data_67__2_) );
DFFPOSX1 DFFPOSX1_1092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_220__3_), .Q(data_67__3_) );
DFFPOSX1 DFFPOSX1_1093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_220__4_), .Q(data_67__4_) );
DFFPOSX1 DFFPOSX1_1094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_220__5_), .Q(data_67__5_) );
DFFPOSX1 DFFPOSX1_1095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_220__6_), .Q(data_67__6_) );
DFFPOSX1 DFFPOSX1_1096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_220__7_), .Q(data_67__7_) );
DFFPOSX1 DFFPOSX1_1097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_220__8_), .Q(data_67__8_) );
DFFPOSX1 DFFPOSX1_1098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_220__9_), .Q(data_67__9_) );
DFFPOSX1 DFFPOSX1_1099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_220__10_), .Q(data_67__10_) );
DFFPOSX1 DFFPOSX1_1100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_220__11_), .Q(data_67__11_) );
DFFPOSX1 DFFPOSX1_1101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_220__12_), .Q(data_67__12_) );
DFFPOSX1 DFFPOSX1_1102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_220__13_), .Q(data_67__13_) );
DFFPOSX1 DFFPOSX1_1103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_220__14_), .Q(data_67__14_) );
DFFPOSX1 DFFPOSX1_1104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_220__15_), .Q(data_67__15_) );
DFFPOSX1 DFFPOSX1_1105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_221__0_), .Q(data_68__0_) );
DFFPOSX1 DFFPOSX1_1106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_221__1_), .Q(data_68__1_) );
DFFPOSX1 DFFPOSX1_1107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_221__2_), .Q(data_68__2_) );
DFFPOSX1 DFFPOSX1_1108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_221__3_), .Q(data_68__3_) );
DFFPOSX1 DFFPOSX1_1109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_221__4_), .Q(data_68__4_) );
DFFPOSX1 DFFPOSX1_1110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_221__5_), .Q(data_68__5_) );
DFFPOSX1 DFFPOSX1_1111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_221__6_), .Q(data_68__6_) );
DFFPOSX1 DFFPOSX1_1112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_221__7_), .Q(data_68__7_) );
DFFPOSX1 DFFPOSX1_1113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_221__8_), .Q(data_68__8_) );
DFFPOSX1 DFFPOSX1_1114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_221__9_), .Q(data_68__9_) );
DFFPOSX1 DFFPOSX1_1115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_221__10_), .Q(data_68__10_) );
DFFPOSX1 DFFPOSX1_1116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_221__11_), .Q(data_68__11_) );
DFFPOSX1 DFFPOSX1_1117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_221__12_), .Q(data_68__12_) );
DFFPOSX1 DFFPOSX1_1118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_221__13_), .Q(data_68__13_) );
DFFPOSX1 DFFPOSX1_1119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_221__14_), .Q(data_68__14_) );
DFFPOSX1 DFFPOSX1_1120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_221__15_), .Q(data_68__15_) );
DFFPOSX1 DFFPOSX1_1121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_222__0_), .Q(data_69__0_) );
DFFPOSX1 DFFPOSX1_1122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_222__1_), .Q(data_69__1_) );
DFFPOSX1 DFFPOSX1_1123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_222__2_), .Q(data_69__2_) );
DFFPOSX1 DFFPOSX1_1124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_222__3_), .Q(data_69__3_) );
DFFPOSX1 DFFPOSX1_1125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_222__4_), .Q(data_69__4_) );
DFFPOSX1 DFFPOSX1_1126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_222__5_), .Q(data_69__5_) );
DFFPOSX1 DFFPOSX1_1127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_222__6_), .Q(data_69__6_) );
DFFPOSX1 DFFPOSX1_1128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_222__7_), .Q(data_69__7_) );
DFFPOSX1 DFFPOSX1_1129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_222__8_), .Q(data_69__8_) );
DFFPOSX1 DFFPOSX1_1130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_222__9_), .Q(data_69__9_) );
DFFPOSX1 DFFPOSX1_1131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_222__10_), .Q(data_69__10_) );
DFFPOSX1 DFFPOSX1_1132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_222__11_), .Q(data_69__11_) );
DFFPOSX1 DFFPOSX1_1133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_222__12_), .Q(data_69__12_) );
DFFPOSX1 DFFPOSX1_1134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_222__13_), .Q(data_69__13_) );
DFFPOSX1 DFFPOSX1_1135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_222__14_), .Q(data_69__14_) );
DFFPOSX1 DFFPOSX1_1136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_222__15_), .Q(data_69__15_) );
DFFPOSX1 DFFPOSX1_1137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_224__0_), .Q(data_70__0_) );
DFFPOSX1 DFFPOSX1_1138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_224__1_), .Q(data_70__1_) );
DFFPOSX1 DFFPOSX1_1139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_224__2_), .Q(data_70__2_) );
DFFPOSX1 DFFPOSX1_1140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_224__3_), .Q(data_70__3_) );
DFFPOSX1 DFFPOSX1_1141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_224__4_), .Q(data_70__4_) );
DFFPOSX1 DFFPOSX1_1142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_224__5_), .Q(data_70__5_) );
DFFPOSX1 DFFPOSX1_1143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_224__6_), .Q(data_70__6_) );
DFFPOSX1 DFFPOSX1_1144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_224__7_), .Q(data_70__7_) );
DFFPOSX1 DFFPOSX1_1145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_224__8_), .Q(data_70__8_) );
DFFPOSX1 DFFPOSX1_1146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_224__9_), .Q(data_70__9_) );
DFFPOSX1 DFFPOSX1_1147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_224__10_), .Q(data_70__10_) );
DFFPOSX1 DFFPOSX1_1148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_224__11_), .Q(data_70__11_) );
DFFPOSX1 DFFPOSX1_1149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_224__12_), .Q(data_70__12_) );
DFFPOSX1 DFFPOSX1_1150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_224__13_), .Q(data_70__13_) );
DFFPOSX1 DFFPOSX1_1151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_224__14_), .Q(data_70__14_) );
DFFPOSX1 DFFPOSX1_1152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_224__15_), .Q(data_70__15_) );
DFFPOSX1 DFFPOSX1_1153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_225__0_), .Q(data_71__0_) );
DFFPOSX1 DFFPOSX1_1154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_225__1_), .Q(data_71__1_) );
DFFPOSX1 DFFPOSX1_1155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_225__2_), .Q(data_71__2_) );
DFFPOSX1 DFFPOSX1_1156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_225__3_), .Q(data_71__3_) );
DFFPOSX1 DFFPOSX1_1157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_225__4_), .Q(data_71__4_) );
DFFPOSX1 DFFPOSX1_1158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_225__5_), .Q(data_71__5_) );
DFFPOSX1 DFFPOSX1_1159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_225__6_), .Q(data_71__6_) );
DFFPOSX1 DFFPOSX1_1160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_225__7_), .Q(data_71__7_) );
DFFPOSX1 DFFPOSX1_1161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_225__8_), .Q(data_71__8_) );
DFFPOSX1 DFFPOSX1_1162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_225__9_), .Q(data_71__9_) );
DFFPOSX1 DFFPOSX1_1163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_225__10_), .Q(data_71__10_) );
DFFPOSX1 DFFPOSX1_1164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_225__11_), .Q(data_71__11_) );
DFFPOSX1 DFFPOSX1_1165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_225__12_), .Q(data_71__12_) );
DFFPOSX1 DFFPOSX1_1166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_225__13_), .Q(data_71__13_) );
DFFPOSX1 DFFPOSX1_1167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_225__14_), .Q(data_71__14_) );
DFFPOSX1 DFFPOSX1_1168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_225__15_), .Q(data_71__15_) );
DFFPOSX1 DFFPOSX1_1169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_226__0_), .Q(data_72__0_) );
DFFPOSX1 DFFPOSX1_1170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_226__1_), .Q(data_72__1_) );
DFFPOSX1 DFFPOSX1_1171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_226__2_), .Q(data_72__2_) );
DFFPOSX1 DFFPOSX1_1172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_226__3_), .Q(data_72__3_) );
DFFPOSX1 DFFPOSX1_1173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_226__4_), .Q(data_72__4_) );
DFFPOSX1 DFFPOSX1_1174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_226__5_), .Q(data_72__5_) );
DFFPOSX1 DFFPOSX1_1175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_226__6_), .Q(data_72__6_) );
DFFPOSX1 DFFPOSX1_1176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_226__7_), .Q(data_72__7_) );
DFFPOSX1 DFFPOSX1_1177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_226__8_), .Q(data_72__8_) );
DFFPOSX1 DFFPOSX1_1178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_226__9_), .Q(data_72__9_) );
DFFPOSX1 DFFPOSX1_1179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_226__10_), .Q(data_72__10_) );
DFFPOSX1 DFFPOSX1_1180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_226__11_), .Q(data_72__11_) );
DFFPOSX1 DFFPOSX1_1181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_226__12_), .Q(data_72__12_) );
DFFPOSX1 DFFPOSX1_1182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_226__13_), .Q(data_72__13_) );
DFFPOSX1 DFFPOSX1_1183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_226__14_), .Q(data_72__14_) );
DFFPOSX1 DFFPOSX1_1184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_226__15_), .Q(data_72__15_) );
DFFPOSX1 DFFPOSX1_1185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_227__0_), .Q(data_73__0_) );
DFFPOSX1 DFFPOSX1_1186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_227__1_), .Q(data_73__1_) );
DFFPOSX1 DFFPOSX1_1187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_227__2_), .Q(data_73__2_) );
DFFPOSX1 DFFPOSX1_1188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_227__3_), .Q(data_73__3_) );
DFFPOSX1 DFFPOSX1_1189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_227__4_), .Q(data_73__4_) );
DFFPOSX1 DFFPOSX1_1190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_227__5_), .Q(data_73__5_) );
DFFPOSX1 DFFPOSX1_1191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_227__6_), .Q(data_73__6_) );
DFFPOSX1 DFFPOSX1_1192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_227__7_), .Q(data_73__7_) );
DFFPOSX1 DFFPOSX1_1193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_227__8_), .Q(data_73__8_) );
DFFPOSX1 DFFPOSX1_1194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_227__9_), .Q(data_73__9_) );
DFFPOSX1 DFFPOSX1_1195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_227__10_), .Q(data_73__10_) );
DFFPOSX1 DFFPOSX1_1196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_227__11_), .Q(data_73__11_) );
DFFPOSX1 DFFPOSX1_1197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_227__12_), .Q(data_73__12_) );
DFFPOSX1 DFFPOSX1_1198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_227__13_), .Q(data_73__13_) );
DFFPOSX1 DFFPOSX1_1199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_227__14_), .Q(data_73__14_) );
DFFPOSX1 DFFPOSX1_1200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_227__15_), .Q(data_73__15_) );
DFFPOSX1 DFFPOSX1_1201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_228__0_), .Q(data_74__0_) );
DFFPOSX1 DFFPOSX1_1202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_228__1_), .Q(data_74__1_) );
DFFPOSX1 DFFPOSX1_1203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_228__2_), .Q(data_74__2_) );
DFFPOSX1 DFFPOSX1_1204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_228__3_), .Q(data_74__3_) );
DFFPOSX1 DFFPOSX1_1205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_228__4_), .Q(data_74__4_) );
DFFPOSX1 DFFPOSX1_1206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_228__5_), .Q(data_74__5_) );
DFFPOSX1 DFFPOSX1_1207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_228__6_), .Q(data_74__6_) );
DFFPOSX1 DFFPOSX1_1208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_228__7_), .Q(data_74__7_) );
DFFPOSX1 DFFPOSX1_1209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_228__8_), .Q(data_74__8_) );
DFFPOSX1 DFFPOSX1_1210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_228__9_), .Q(data_74__9_) );
DFFPOSX1 DFFPOSX1_1211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_228__10_), .Q(data_74__10_) );
DFFPOSX1 DFFPOSX1_1212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_228__11_), .Q(data_74__11_) );
DFFPOSX1 DFFPOSX1_1213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_228__12_), .Q(data_74__12_) );
DFFPOSX1 DFFPOSX1_1214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_228__13_), .Q(data_74__13_) );
DFFPOSX1 DFFPOSX1_1215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_228__14_), .Q(data_74__14_) );
DFFPOSX1 DFFPOSX1_1216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_228__15_), .Q(data_74__15_) );
DFFPOSX1 DFFPOSX1_1217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_229__0_), .Q(data_75__0_) );
DFFPOSX1 DFFPOSX1_1218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_229__1_), .Q(data_75__1_) );
DFFPOSX1 DFFPOSX1_1219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_229__2_), .Q(data_75__2_) );
DFFPOSX1 DFFPOSX1_1220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_229__3_), .Q(data_75__3_) );
DFFPOSX1 DFFPOSX1_1221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_229__4_), .Q(data_75__4_) );
DFFPOSX1 DFFPOSX1_1222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_229__5_), .Q(data_75__5_) );
DFFPOSX1 DFFPOSX1_1223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_229__6_), .Q(data_75__6_) );
DFFPOSX1 DFFPOSX1_1224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_229__7_), .Q(data_75__7_) );
DFFPOSX1 DFFPOSX1_1225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_229__8_), .Q(data_75__8_) );
DFFPOSX1 DFFPOSX1_1226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_229__9_), .Q(data_75__9_) );
DFFPOSX1 DFFPOSX1_1227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_229__10_), .Q(data_75__10_) );
DFFPOSX1 DFFPOSX1_1228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_229__11_), .Q(data_75__11_) );
DFFPOSX1 DFFPOSX1_1229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_229__12_), .Q(data_75__12_) );
DFFPOSX1 DFFPOSX1_1230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_229__13_), .Q(data_75__13_) );
DFFPOSX1 DFFPOSX1_1231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_229__14_), .Q(data_75__14_) );
DFFPOSX1 DFFPOSX1_1232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_229__15_), .Q(data_75__15_) );
DFFPOSX1 DFFPOSX1_1233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_230__0_), .Q(data_76__0_) );
DFFPOSX1 DFFPOSX1_1234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_230__1_), .Q(data_76__1_) );
DFFPOSX1 DFFPOSX1_1235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_230__2_), .Q(data_76__2_) );
DFFPOSX1 DFFPOSX1_1236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_230__3_), .Q(data_76__3_) );
DFFPOSX1 DFFPOSX1_1237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_230__4_), .Q(data_76__4_) );
DFFPOSX1 DFFPOSX1_1238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_230__5_), .Q(data_76__5_) );
DFFPOSX1 DFFPOSX1_1239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_230__6_), .Q(data_76__6_) );
DFFPOSX1 DFFPOSX1_1240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_230__7_), .Q(data_76__7_) );
DFFPOSX1 DFFPOSX1_1241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_230__8_), .Q(data_76__8_) );
DFFPOSX1 DFFPOSX1_1242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_230__9_), .Q(data_76__9_) );
DFFPOSX1 DFFPOSX1_1243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_230__10_), .Q(data_76__10_) );
DFFPOSX1 DFFPOSX1_1244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_230__11_), .Q(data_76__11_) );
DFFPOSX1 DFFPOSX1_1245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_230__12_), .Q(data_76__12_) );
DFFPOSX1 DFFPOSX1_1246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_230__13_), .Q(data_76__13_) );
DFFPOSX1 DFFPOSX1_1247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_230__14_), .Q(data_76__14_) );
DFFPOSX1 DFFPOSX1_1248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_230__15_), .Q(data_76__15_) );
DFFPOSX1 DFFPOSX1_1249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_231__0_), .Q(data_77__0_) );
DFFPOSX1 DFFPOSX1_1250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_231__1_), .Q(data_77__1_) );
DFFPOSX1 DFFPOSX1_1251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_231__2_), .Q(data_77__2_) );
DFFPOSX1 DFFPOSX1_1252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_231__3_), .Q(data_77__3_) );
DFFPOSX1 DFFPOSX1_1253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_231__4_), .Q(data_77__4_) );
DFFPOSX1 DFFPOSX1_1254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_231__5_), .Q(data_77__5_) );
DFFPOSX1 DFFPOSX1_1255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_231__6_), .Q(data_77__6_) );
DFFPOSX1 DFFPOSX1_1256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_231__7_), .Q(data_77__7_) );
DFFPOSX1 DFFPOSX1_1257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_231__8_), .Q(data_77__8_) );
DFFPOSX1 DFFPOSX1_1258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_231__9_), .Q(data_77__9_) );
DFFPOSX1 DFFPOSX1_1259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_231__10_), .Q(data_77__10_) );
DFFPOSX1 DFFPOSX1_1260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_231__11_), .Q(data_77__11_) );
DFFPOSX1 DFFPOSX1_1261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_231__12_), .Q(data_77__12_) );
DFFPOSX1 DFFPOSX1_1262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_231__13_), .Q(data_77__13_) );
DFFPOSX1 DFFPOSX1_1263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_231__14_), .Q(data_77__14_) );
DFFPOSX1 DFFPOSX1_1264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_231__15_), .Q(data_77__15_) );
DFFPOSX1 DFFPOSX1_1265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_232__0_), .Q(data_78__0_) );
DFFPOSX1 DFFPOSX1_1266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_232__1_), .Q(data_78__1_) );
DFFPOSX1 DFFPOSX1_1267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_232__2_), .Q(data_78__2_) );
DFFPOSX1 DFFPOSX1_1268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_232__3_), .Q(data_78__3_) );
DFFPOSX1 DFFPOSX1_1269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_232__4_), .Q(data_78__4_) );
DFFPOSX1 DFFPOSX1_1270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_232__5_), .Q(data_78__5_) );
DFFPOSX1 DFFPOSX1_1271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_232__6_), .Q(data_78__6_) );
DFFPOSX1 DFFPOSX1_1272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_232__7_), .Q(data_78__7_) );
DFFPOSX1 DFFPOSX1_1273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_232__8_), .Q(data_78__8_) );
DFFPOSX1 DFFPOSX1_1274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_232__9_), .Q(data_78__9_) );
DFFPOSX1 DFFPOSX1_1275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_232__10_), .Q(data_78__10_) );
DFFPOSX1 DFFPOSX1_1276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_232__11_), .Q(data_78__11_) );
DFFPOSX1 DFFPOSX1_1277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_232__12_), .Q(data_78__12_) );
DFFPOSX1 DFFPOSX1_1278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_232__13_), .Q(data_78__13_) );
DFFPOSX1 DFFPOSX1_1279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_232__14_), .Q(data_78__14_) );
DFFPOSX1 DFFPOSX1_1280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_232__15_), .Q(data_78__15_) );
DFFPOSX1 DFFPOSX1_1281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf2), .D(_233__0_), .Q(data_79__0_) );
DFFPOSX1 DFFPOSX1_1282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf2), .D(_233__1_), .Q(data_79__1_) );
DFFPOSX1 DFFPOSX1_1283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf2), .D(_233__2_), .Q(data_79__2_) );
DFFPOSX1 DFFPOSX1_1284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf2), .D(_233__3_), .Q(data_79__3_) );
DFFPOSX1 DFFPOSX1_1285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf2), .D(_233__4_), .Q(data_79__4_) );
DFFPOSX1 DFFPOSX1_1286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf2), .D(_233__5_), .Q(data_79__5_) );
DFFPOSX1 DFFPOSX1_1287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf2), .D(_233__6_), .Q(data_79__6_) );
DFFPOSX1 DFFPOSX1_1288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf2), .D(_233__7_), .Q(data_79__7_) );
DFFPOSX1 DFFPOSX1_1289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf2), .D(_233__8_), .Q(data_79__8_) );
DFFPOSX1 DFFPOSX1_1290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf2), .D(_233__9_), .Q(data_79__9_) );
DFFPOSX1 DFFPOSX1_1291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf2), .D(_233__10_), .Q(data_79__10_) );
DFFPOSX1 DFFPOSX1_1292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf2), .D(_233__11_), .Q(data_79__11_) );
DFFPOSX1 DFFPOSX1_1293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf2), .D(_233__12_), .Q(data_79__12_) );
DFFPOSX1 DFFPOSX1_1294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf2), .D(_233__13_), .Q(data_79__13_) );
DFFPOSX1 DFFPOSX1_1295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf2), .D(_233__14_), .Q(data_79__14_) );
DFFPOSX1 DFFPOSX1_1296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf2), .D(_233__15_), .Q(data_79__15_) );
DFFPOSX1 DFFPOSX1_1297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_235__0_), .Q(data_80__0_) );
DFFPOSX1 DFFPOSX1_1298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_235__1_), .Q(data_80__1_) );
DFFPOSX1 DFFPOSX1_1299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_235__2_), .Q(data_80__2_) );
DFFPOSX1 DFFPOSX1_1300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_235__3_), .Q(data_80__3_) );
DFFPOSX1 DFFPOSX1_1301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_235__4_), .Q(data_80__4_) );
DFFPOSX1 DFFPOSX1_1302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_235__5_), .Q(data_80__5_) );
DFFPOSX1 DFFPOSX1_1303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_235__6_), .Q(data_80__6_) );
DFFPOSX1 DFFPOSX1_1304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_235__7_), .Q(data_80__7_) );
DFFPOSX1 DFFPOSX1_1305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_235__8_), .Q(data_80__8_) );
DFFPOSX1 DFFPOSX1_1306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_235__9_), .Q(data_80__9_) );
DFFPOSX1 DFFPOSX1_1307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_235__10_), .Q(data_80__10_) );
DFFPOSX1 DFFPOSX1_1308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_235__11_), .Q(data_80__11_) );
DFFPOSX1 DFFPOSX1_1309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_235__12_), .Q(data_80__12_) );
DFFPOSX1 DFFPOSX1_1310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_235__13_), .Q(data_80__13_) );
DFFPOSX1 DFFPOSX1_1311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_235__14_), .Q(data_80__14_) );
DFFPOSX1 DFFPOSX1_1312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_235__15_), .Q(data_80__15_) );
DFFPOSX1 DFFPOSX1_1313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_236__0_), .Q(data_81__0_) );
DFFPOSX1 DFFPOSX1_1314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_236__1_), .Q(data_81__1_) );
DFFPOSX1 DFFPOSX1_1315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_236__2_), .Q(data_81__2_) );
DFFPOSX1 DFFPOSX1_1316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_236__3_), .Q(data_81__3_) );
DFFPOSX1 DFFPOSX1_1317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_236__4_), .Q(data_81__4_) );
DFFPOSX1 DFFPOSX1_1318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_236__5_), .Q(data_81__5_) );
DFFPOSX1 DFFPOSX1_1319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_236__6_), .Q(data_81__6_) );
DFFPOSX1 DFFPOSX1_1320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_236__7_), .Q(data_81__7_) );
DFFPOSX1 DFFPOSX1_1321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_236__8_), .Q(data_81__8_) );
DFFPOSX1 DFFPOSX1_1322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_236__9_), .Q(data_81__9_) );
DFFPOSX1 DFFPOSX1_1323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_236__10_), .Q(data_81__10_) );
DFFPOSX1 DFFPOSX1_1324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_236__11_), .Q(data_81__11_) );
DFFPOSX1 DFFPOSX1_1325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_236__12_), .Q(data_81__12_) );
DFFPOSX1 DFFPOSX1_1326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_236__13_), .Q(data_81__13_) );
DFFPOSX1 DFFPOSX1_1327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_236__14_), .Q(data_81__14_) );
DFFPOSX1 DFFPOSX1_1328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_236__15_), .Q(data_81__15_) );
DFFPOSX1 DFFPOSX1_1329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_237__0_), .Q(data_82__0_) );
DFFPOSX1 DFFPOSX1_1330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_237__1_), .Q(data_82__1_) );
DFFPOSX1 DFFPOSX1_1331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_237__2_), .Q(data_82__2_) );
DFFPOSX1 DFFPOSX1_1332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_237__3_), .Q(data_82__3_) );
DFFPOSX1 DFFPOSX1_1333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_237__4_), .Q(data_82__4_) );
DFFPOSX1 DFFPOSX1_1334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_237__5_), .Q(data_82__5_) );
DFFPOSX1 DFFPOSX1_1335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_237__6_), .Q(data_82__6_) );
DFFPOSX1 DFFPOSX1_1336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_237__7_), .Q(data_82__7_) );
DFFPOSX1 DFFPOSX1_1337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_237__8_), .Q(data_82__8_) );
DFFPOSX1 DFFPOSX1_1338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_237__9_), .Q(data_82__9_) );
DFFPOSX1 DFFPOSX1_1339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_237__10_), .Q(data_82__10_) );
DFFPOSX1 DFFPOSX1_1340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_237__11_), .Q(data_82__11_) );
DFFPOSX1 DFFPOSX1_1341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_237__12_), .Q(data_82__12_) );
DFFPOSX1 DFFPOSX1_1342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_237__13_), .Q(data_82__13_) );
DFFPOSX1 DFFPOSX1_1343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_237__14_), .Q(data_82__14_) );
DFFPOSX1 DFFPOSX1_1344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_237__15_), .Q(data_82__15_) );
DFFPOSX1 DFFPOSX1_1345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_238__0_), .Q(data_83__0_) );
DFFPOSX1 DFFPOSX1_1346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_238__1_), .Q(data_83__1_) );
DFFPOSX1 DFFPOSX1_1347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_238__2_), .Q(data_83__2_) );
DFFPOSX1 DFFPOSX1_1348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_238__3_), .Q(data_83__3_) );
DFFPOSX1 DFFPOSX1_1349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_238__4_), .Q(data_83__4_) );
DFFPOSX1 DFFPOSX1_1350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_238__5_), .Q(data_83__5_) );
DFFPOSX1 DFFPOSX1_1351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_238__6_), .Q(data_83__6_) );
DFFPOSX1 DFFPOSX1_1352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_238__7_), .Q(data_83__7_) );
DFFPOSX1 DFFPOSX1_1353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_238__8_), .Q(data_83__8_) );
DFFPOSX1 DFFPOSX1_1354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_238__9_), .Q(data_83__9_) );
DFFPOSX1 DFFPOSX1_1355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_238__10_), .Q(data_83__10_) );
DFFPOSX1 DFFPOSX1_1356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_238__11_), .Q(data_83__11_) );
DFFPOSX1 DFFPOSX1_1357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_238__12_), .Q(data_83__12_) );
DFFPOSX1 DFFPOSX1_1358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_238__13_), .Q(data_83__13_) );
DFFPOSX1 DFFPOSX1_1359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_238__14_), .Q(data_83__14_) );
DFFPOSX1 DFFPOSX1_1360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_238__15_), .Q(data_83__15_) );
DFFPOSX1 DFFPOSX1_1361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_239__0_), .Q(data_84__0_) );
DFFPOSX1 DFFPOSX1_1362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_239__1_), .Q(data_84__1_) );
DFFPOSX1 DFFPOSX1_1363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_239__2_), .Q(data_84__2_) );
DFFPOSX1 DFFPOSX1_1364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_239__3_), .Q(data_84__3_) );
DFFPOSX1 DFFPOSX1_1365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_239__4_), .Q(data_84__4_) );
DFFPOSX1 DFFPOSX1_1366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_239__5_), .Q(data_84__5_) );
DFFPOSX1 DFFPOSX1_1367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_239__6_), .Q(data_84__6_) );
DFFPOSX1 DFFPOSX1_1368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_239__7_), .Q(data_84__7_) );
DFFPOSX1 DFFPOSX1_1369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_239__8_), .Q(data_84__8_) );
DFFPOSX1 DFFPOSX1_1370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_239__9_), .Q(data_84__9_) );
DFFPOSX1 DFFPOSX1_1371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_239__10_), .Q(data_84__10_) );
DFFPOSX1 DFFPOSX1_1372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_239__11_), .Q(data_84__11_) );
DFFPOSX1 DFFPOSX1_1373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_239__12_), .Q(data_84__12_) );
DFFPOSX1 DFFPOSX1_1374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_239__13_), .Q(data_84__13_) );
DFFPOSX1 DFFPOSX1_1375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_239__14_), .Q(data_84__14_) );
DFFPOSX1 DFFPOSX1_1376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_239__15_), .Q(data_84__15_) );
DFFPOSX1 DFFPOSX1_1377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_240__0_), .Q(data_85__0_) );
DFFPOSX1 DFFPOSX1_1378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_240__1_), .Q(data_85__1_) );
DFFPOSX1 DFFPOSX1_1379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_240__2_), .Q(data_85__2_) );
DFFPOSX1 DFFPOSX1_1380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_240__3_), .Q(data_85__3_) );
DFFPOSX1 DFFPOSX1_1381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_240__4_), .Q(data_85__4_) );
DFFPOSX1 DFFPOSX1_1382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_240__5_), .Q(data_85__5_) );
DFFPOSX1 DFFPOSX1_1383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_240__6_), .Q(data_85__6_) );
DFFPOSX1 DFFPOSX1_1384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_240__7_), .Q(data_85__7_) );
DFFPOSX1 DFFPOSX1_1385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_240__8_), .Q(data_85__8_) );
DFFPOSX1 DFFPOSX1_1386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_240__9_), .Q(data_85__9_) );
DFFPOSX1 DFFPOSX1_1387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_240__10_), .Q(data_85__10_) );
DFFPOSX1 DFFPOSX1_1388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_240__11_), .Q(data_85__11_) );
DFFPOSX1 DFFPOSX1_1389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_240__12_), .Q(data_85__12_) );
DFFPOSX1 DFFPOSX1_1390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_240__13_), .Q(data_85__13_) );
DFFPOSX1 DFFPOSX1_1391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_240__14_), .Q(data_85__14_) );
DFFPOSX1 DFFPOSX1_1392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_240__15_), .Q(data_85__15_) );
DFFPOSX1 DFFPOSX1_1393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_241__0_), .Q(data_86__0_) );
DFFPOSX1 DFFPOSX1_1394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_241__1_), .Q(data_86__1_) );
DFFPOSX1 DFFPOSX1_1395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_241__2_), .Q(data_86__2_) );
DFFPOSX1 DFFPOSX1_1396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_241__3_), .Q(data_86__3_) );
DFFPOSX1 DFFPOSX1_1397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_241__4_), .Q(data_86__4_) );
DFFPOSX1 DFFPOSX1_1398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_241__5_), .Q(data_86__5_) );
DFFPOSX1 DFFPOSX1_1399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_241__6_), .Q(data_86__6_) );
DFFPOSX1 DFFPOSX1_1400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_241__7_), .Q(data_86__7_) );
DFFPOSX1 DFFPOSX1_1401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_241__8_), .Q(data_86__8_) );
DFFPOSX1 DFFPOSX1_1402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_241__9_), .Q(data_86__9_) );
DFFPOSX1 DFFPOSX1_1403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_241__10_), .Q(data_86__10_) );
DFFPOSX1 DFFPOSX1_1404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_241__11_), .Q(data_86__11_) );
DFFPOSX1 DFFPOSX1_1405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_241__12_), .Q(data_86__12_) );
DFFPOSX1 DFFPOSX1_1406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_241__13_), .Q(data_86__13_) );
DFFPOSX1 DFFPOSX1_1407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_241__14_), .Q(data_86__14_) );
DFFPOSX1 DFFPOSX1_1408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_241__15_), .Q(data_86__15_) );
DFFPOSX1 DFFPOSX1_1409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_242__0_), .Q(data_87__0_) );
DFFPOSX1 DFFPOSX1_1410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_242__1_), .Q(data_87__1_) );
DFFPOSX1 DFFPOSX1_1411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_242__2_), .Q(data_87__2_) );
DFFPOSX1 DFFPOSX1_1412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_242__3_), .Q(data_87__3_) );
DFFPOSX1 DFFPOSX1_1413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_242__4_), .Q(data_87__4_) );
DFFPOSX1 DFFPOSX1_1414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_242__5_), .Q(data_87__5_) );
DFFPOSX1 DFFPOSX1_1415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_242__6_), .Q(data_87__6_) );
DFFPOSX1 DFFPOSX1_1416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_242__7_), .Q(data_87__7_) );
DFFPOSX1 DFFPOSX1_1417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_242__8_), .Q(data_87__8_) );
DFFPOSX1 DFFPOSX1_1418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_242__9_), .Q(data_87__9_) );
DFFPOSX1 DFFPOSX1_1419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_242__10_), .Q(data_87__10_) );
DFFPOSX1 DFFPOSX1_1420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_242__11_), .Q(data_87__11_) );
DFFPOSX1 DFFPOSX1_1421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_242__12_), .Q(data_87__12_) );
DFFPOSX1 DFFPOSX1_1422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_242__13_), .Q(data_87__13_) );
DFFPOSX1 DFFPOSX1_1423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_242__14_), .Q(data_87__14_) );
DFFPOSX1 DFFPOSX1_1424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_242__15_), .Q(data_87__15_) );
DFFPOSX1 DFFPOSX1_1425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_243__0_), .Q(data_88__0_) );
DFFPOSX1 DFFPOSX1_1426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_243__1_), .Q(data_88__1_) );
DFFPOSX1 DFFPOSX1_1427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_243__2_), .Q(data_88__2_) );
DFFPOSX1 DFFPOSX1_1428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_243__3_), .Q(data_88__3_) );
DFFPOSX1 DFFPOSX1_1429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_243__4_), .Q(data_88__4_) );
DFFPOSX1 DFFPOSX1_1430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_243__5_), .Q(data_88__5_) );
DFFPOSX1 DFFPOSX1_1431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_243__6_), .Q(data_88__6_) );
DFFPOSX1 DFFPOSX1_1432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_243__7_), .Q(data_88__7_) );
DFFPOSX1 DFFPOSX1_1433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_243__8_), .Q(data_88__8_) );
DFFPOSX1 DFFPOSX1_1434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_243__9_), .Q(data_88__9_) );
DFFPOSX1 DFFPOSX1_1435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_243__10_), .Q(data_88__10_) );
DFFPOSX1 DFFPOSX1_1436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_243__11_), .Q(data_88__11_) );
DFFPOSX1 DFFPOSX1_1437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_243__12_), .Q(data_88__12_) );
DFFPOSX1 DFFPOSX1_1438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_243__13_), .Q(data_88__13_) );
DFFPOSX1 DFFPOSX1_1439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_243__14_), .Q(data_88__14_) );
DFFPOSX1 DFFPOSX1_1440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_243__15_), .Q(data_88__15_) );
DFFPOSX1 DFFPOSX1_1441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_244__0_), .Q(data_89__0_) );
DFFPOSX1 DFFPOSX1_1442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_244__1_), .Q(data_89__1_) );
DFFPOSX1 DFFPOSX1_1443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_244__2_), .Q(data_89__2_) );
DFFPOSX1 DFFPOSX1_1444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_244__3_), .Q(data_89__3_) );
DFFPOSX1 DFFPOSX1_1445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_244__4_), .Q(data_89__4_) );
DFFPOSX1 DFFPOSX1_1446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_244__5_), .Q(data_89__5_) );
DFFPOSX1 DFFPOSX1_1447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_244__6_), .Q(data_89__6_) );
DFFPOSX1 DFFPOSX1_1448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_244__7_), .Q(data_89__7_) );
DFFPOSX1 DFFPOSX1_1449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_244__8_), .Q(data_89__8_) );
DFFPOSX1 DFFPOSX1_1450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_244__9_), .Q(data_89__9_) );
DFFPOSX1 DFFPOSX1_1451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_244__10_), .Q(data_89__10_) );
DFFPOSX1 DFFPOSX1_1452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_244__11_), .Q(data_89__11_) );
DFFPOSX1 DFFPOSX1_1453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_244__12_), .Q(data_89__12_) );
DFFPOSX1 DFFPOSX1_1454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_244__13_), .Q(data_89__13_) );
DFFPOSX1 DFFPOSX1_1455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_244__14_), .Q(data_89__14_) );
DFFPOSX1 DFFPOSX1_1456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_244__15_), .Q(data_89__15_) );
DFFPOSX1 DFFPOSX1_1457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_246__0_), .Q(data_90__0_) );
DFFPOSX1 DFFPOSX1_1458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_246__1_), .Q(data_90__1_) );
DFFPOSX1 DFFPOSX1_1459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_246__2_), .Q(data_90__2_) );
DFFPOSX1 DFFPOSX1_1460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_246__3_), .Q(data_90__3_) );
DFFPOSX1 DFFPOSX1_1461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_246__4_), .Q(data_90__4_) );
DFFPOSX1 DFFPOSX1_1462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_246__5_), .Q(data_90__5_) );
DFFPOSX1 DFFPOSX1_1463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_246__6_), .Q(data_90__6_) );
DFFPOSX1 DFFPOSX1_1464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_246__7_), .Q(data_90__7_) );
DFFPOSX1 DFFPOSX1_1465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_246__8_), .Q(data_90__8_) );
DFFPOSX1 DFFPOSX1_1466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_246__9_), .Q(data_90__9_) );
DFFPOSX1 DFFPOSX1_1467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_246__10_), .Q(data_90__10_) );
DFFPOSX1 DFFPOSX1_1468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_246__11_), .Q(data_90__11_) );
DFFPOSX1 DFFPOSX1_1469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_246__12_), .Q(data_90__12_) );
DFFPOSX1 DFFPOSX1_1470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_246__13_), .Q(data_90__13_) );
DFFPOSX1 DFFPOSX1_1471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_246__14_), .Q(data_90__14_) );
DFFPOSX1 DFFPOSX1_1472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_246__15_), .Q(data_90__15_) );
DFFPOSX1 DFFPOSX1_1473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_247__0_), .Q(data_91__0_) );
DFFPOSX1 DFFPOSX1_1474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_247__1_), .Q(data_91__1_) );
DFFPOSX1 DFFPOSX1_1475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_247__2_), .Q(data_91__2_) );
DFFPOSX1 DFFPOSX1_1476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_247__3_), .Q(data_91__3_) );
DFFPOSX1 DFFPOSX1_1477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_247__4_), .Q(data_91__4_) );
DFFPOSX1 DFFPOSX1_1478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_247__5_), .Q(data_91__5_) );
DFFPOSX1 DFFPOSX1_1479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_247__6_), .Q(data_91__6_) );
DFFPOSX1 DFFPOSX1_1480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_247__7_), .Q(data_91__7_) );
DFFPOSX1 DFFPOSX1_1481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_247__8_), .Q(data_91__8_) );
DFFPOSX1 DFFPOSX1_1482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_247__9_), .Q(data_91__9_) );
DFFPOSX1 DFFPOSX1_1483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_247__10_), .Q(data_91__10_) );
DFFPOSX1 DFFPOSX1_1484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_247__11_), .Q(data_91__11_) );
DFFPOSX1 DFFPOSX1_1485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_247__12_), .Q(data_91__12_) );
DFFPOSX1 DFFPOSX1_1486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_247__13_), .Q(data_91__13_) );
DFFPOSX1 DFFPOSX1_1487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_247__14_), .Q(data_91__14_) );
DFFPOSX1 DFFPOSX1_1488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_247__15_), .Q(data_91__15_) );
DFFPOSX1 DFFPOSX1_1489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_248__0_), .Q(data_92__0_) );
DFFPOSX1 DFFPOSX1_1490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_248__1_), .Q(data_92__1_) );
DFFPOSX1 DFFPOSX1_1491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_248__2_), .Q(data_92__2_) );
DFFPOSX1 DFFPOSX1_1492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_248__3_), .Q(data_92__3_) );
DFFPOSX1 DFFPOSX1_1493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_248__4_), .Q(data_92__4_) );
DFFPOSX1 DFFPOSX1_1494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_248__5_), .Q(data_92__5_) );
DFFPOSX1 DFFPOSX1_1495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_248__6_), .Q(data_92__6_) );
DFFPOSX1 DFFPOSX1_1496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_248__7_), .Q(data_92__7_) );
DFFPOSX1 DFFPOSX1_1497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_248__8_), .Q(data_92__8_) );
DFFPOSX1 DFFPOSX1_1498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_248__9_), .Q(data_92__9_) );
DFFPOSX1 DFFPOSX1_1499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_248__10_), .Q(data_92__10_) );
DFFPOSX1 DFFPOSX1_1500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_248__11_), .Q(data_92__11_) );
DFFPOSX1 DFFPOSX1_1501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_248__12_), .Q(data_92__12_) );
DFFPOSX1 DFFPOSX1_1502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_248__13_), .Q(data_92__13_) );
DFFPOSX1 DFFPOSX1_1503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_248__14_), .Q(data_92__14_) );
DFFPOSX1 DFFPOSX1_1504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_248__15_), .Q(data_92__15_) );
DFFPOSX1 DFFPOSX1_1505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_249__0_), .Q(data_93__0_) );
DFFPOSX1 DFFPOSX1_1506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_249__1_), .Q(data_93__1_) );
DFFPOSX1 DFFPOSX1_1507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_249__2_), .Q(data_93__2_) );
DFFPOSX1 DFFPOSX1_1508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_249__3_), .Q(data_93__3_) );
DFFPOSX1 DFFPOSX1_1509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_249__4_), .Q(data_93__4_) );
DFFPOSX1 DFFPOSX1_1510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_249__5_), .Q(data_93__5_) );
DFFPOSX1 DFFPOSX1_1511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_249__6_), .Q(data_93__6_) );
DFFPOSX1 DFFPOSX1_1512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_249__7_), .Q(data_93__7_) );
DFFPOSX1 DFFPOSX1_1513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_249__8_), .Q(data_93__8_) );
DFFPOSX1 DFFPOSX1_1514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_249__9_), .Q(data_93__9_) );
DFFPOSX1 DFFPOSX1_1515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_249__10_), .Q(data_93__10_) );
DFFPOSX1 DFFPOSX1_1516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_249__11_), .Q(data_93__11_) );
DFFPOSX1 DFFPOSX1_1517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_249__12_), .Q(data_93__12_) );
DFFPOSX1 DFFPOSX1_1518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_249__13_), .Q(data_93__13_) );
DFFPOSX1 DFFPOSX1_1519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_249__14_), .Q(data_93__14_) );
DFFPOSX1 DFFPOSX1_1520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_249__15_), .Q(data_93__15_) );
DFFPOSX1 DFFPOSX1_1521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_250__0_), .Q(data_94__0_) );
DFFPOSX1 DFFPOSX1_1522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_250__1_), .Q(data_94__1_) );
DFFPOSX1 DFFPOSX1_1523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_250__2_), .Q(data_94__2_) );
DFFPOSX1 DFFPOSX1_1524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_250__3_), .Q(data_94__3_) );
DFFPOSX1 DFFPOSX1_1525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_250__4_), .Q(data_94__4_) );
DFFPOSX1 DFFPOSX1_1526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_250__5_), .Q(data_94__5_) );
DFFPOSX1 DFFPOSX1_1527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_250__6_), .Q(data_94__6_) );
DFFPOSX1 DFFPOSX1_1528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_250__7_), .Q(data_94__7_) );
DFFPOSX1 DFFPOSX1_1529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_250__8_), .Q(data_94__8_) );
DFFPOSX1 DFFPOSX1_1530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_250__9_), .Q(data_94__9_) );
DFFPOSX1 DFFPOSX1_1531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_250__10_), .Q(data_94__10_) );
DFFPOSX1 DFFPOSX1_1532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_250__11_), .Q(data_94__11_) );
DFFPOSX1 DFFPOSX1_1533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_250__12_), .Q(data_94__12_) );
DFFPOSX1 DFFPOSX1_1534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_250__13_), .Q(data_94__13_) );
DFFPOSX1 DFFPOSX1_1535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_250__14_), .Q(data_94__14_) );
DFFPOSX1 DFFPOSX1_1536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_250__15_), .Q(data_94__15_) );
DFFPOSX1 DFFPOSX1_1537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf1), .D(_251__0_), .Q(data_95__0_) );
DFFPOSX1 DFFPOSX1_1538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf1), .D(_251__1_), .Q(data_95__1_) );
DFFPOSX1 DFFPOSX1_1539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf1), .D(_251__2_), .Q(data_95__2_) );
DFFPOSX1 DFFPOSX1_1540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf1), .D(_251__3_), .Q(data_95__3_) );
DFFPOSX1 DFFPOSX1_1541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf1), .D(_251__4_), .Q(data_95__4_) );
DFFPOSX1 DFFPOSX1_1542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf1), .D(_251__5_), .Q(data_95__5_) );
DFFPOSX1 DFFPOSX1_1543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf1), .D(_251__6_), .Q(data_95__6_) );
DFFPOSX1 DFFPOSX1_1544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf1), .D(_251__7_), .Q(data_95__7_) );
DFFPOSX1 DFFPOSX1_1545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf1), .D(_251__8_), .Q(data_95__8_) );
DFFPOSX1 DFFPOSX1_1546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf1), .D(_251__9_), .Q(data_95__9_) );
DFFPOSX1 DFFPOSX1_1547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf1), .D(_251__10_), .Q(data_95__10_) );
DFFPOSX1 DFFPOSX1_1548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf1), .D(_251__11_), .Q(data_95__11_) );
DFFPOSX1 DFFPOSX1_1549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf1), .D(_251__12_), .Q(data_95__12_) );
DFFPOSX1 DFFPOSX1_1550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf1), .D(_251__13_), .Q(data_95__13_) );
DFFPOSX1 DFFPOSX1_1551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf1), .D(_251__14_), .Q(data_95__14_) );
DFFPOSX1 DFFPOSX1_1552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf1), .D(_251__15_), .Q(data_95__15_) );
DFFPOSX1 DFFPOSX1_1553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_252__0_), .Q(data_96__0_) );
DFFPOSX1 DFFPOSX1_1554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_252__1_), .Q(data_96__1_) );
DFFPOSX1 DFFPOSX1_1555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_252__2_), .Q(data_96__2_) );
DFFPOSX1 DFFPOSX1_1556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_252__3_), .Q(data_96__3_) );
DFFPOSX1 DFFPOSX1_1557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_252__4_), .Q(data_96__4_) );
DFFPOSX1 DFFPOSX1_1558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_252__5_), .Q(data_96__5_) );
DFFPOSX1 DFFPOSX1_1559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_252__6_), .Q(data_96__6_) );
DFFPOSX1 DFFPOSX1_1560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_252__7_), .Q(data_96__7_) );
DFFPOSX1 DFFPOSX1_1561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_252__8_), .Q(data_96__8_) );
DFFPOSX1 DFFPOSX1_1562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_252__9_), .Q(data_96__9_) );
DFFPOSX1 DFFPOSX1_1563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_252__10_), .Q(data_96__10_) );
DFFPOSX1 DFFPOSX1_1564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_252__11_), .Q(data_96__11_) );
DFFPOSX1 DFFPOSX1_1565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_252__12_), .Q(data_96__12_) );
DFFPOSX1 DFFPOSX1_1566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_252__13_), .Q(data_96__13_) );
DFFPOSX1 DFFPOSX1_1567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_252__14_), .Q(data_96__14_) );
DFFPOSX1 DFFPOSX1_1568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_252__15_), .Q(data_96__15_) );
DFFPOSX1 DFFPOSX1_1569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_253__0_), .Q(data_97__0_) );
DFFPOSX1 DFFPOSX1_1570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_253__1_), .Q(data_97__1_) );
DFFPOSX1 DFFPOSX1_1571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_253__2_), .Q(data_97__2_) );
DFFPOSX1 DFFPOSX1_1572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_253__3_), .Q(data_97__3_) );
DFFPOSX1 DFFPOSX1_1573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_253__4_), .Q(data_97__4_) );
DFFPOSX1 DFFPOSX1_1574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_253__5_), .Q(data_97__5_) );
DFFPOSX1 DFFPOSX1_1575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_253__6_), .Q(data_97__6_) );
DFFPOSX1 DFFPOSX1_1576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_253__7_), .Q(data_97__7_) );
DFFPOSX1 DFFPOSX1_1577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_253__8_), .Q(data_97__8_) );
DFFPOSX1 DFFPOSX1_1578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_253__9_), .Q(data_97__9_) );
DFFPOSX1 DFFPOSX1_1579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_253__10_), .Q(data_97__10_) );
DFFPOSX1 DFFPOSX1_1580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_253__11_), .Q(data_97__11_) );
DFFPOSX1 DFFPOSX1_1581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_253__12_), .Q(data_97__12_) );
DFFPOSX1 DFFPOSX1_1582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_253__13_), .Q(data_97__13_) );
DFFPOSX1 DFFPOSX1_1583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_253__14_), .Q(data_97__14_) );
DFFPOSX1 DFFPOSX1_1584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_253__15_), .Q(data_97__15_) );
DFFPOSX1 DFFPOSX1_1585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_254__0_), .Q(data_98__0_) );
DFFPOSX1 DFFPOSX1_1586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_254__1_), .Q(data_98__1_) );
DFFPOSX1 DFFPOSX1_1587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_254__2_), .Q(data_98__2_) );
DFFPOSX1 DFFPOSX1_1588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_254__3_), .Q(data_98__3_) );
DFFPOSX1 DFFPOSX1_1589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_254__4_), .Q(data_98__4_) );
DFFPOSX1 DFFPOSX1_1590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_254__5_), .Q(data_98__5_) );
DFFPOSX1 DFFPOSX1_1591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_254__6_), .Q(data_98__6_) );
DFFPOSX1 DFFPOSX1_1592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_254__7_), .Q(data_98__7_) );
DFFPOSX1 DFFPOSX1_1593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_254__8_), .Q(data_98__8_) );
DFFPOSX1 DFFPOSX1_1594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_254__9_), .Q(data_98__9_) );
DFFPOSX1 DFFPOSX1_1595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_254__10_), .Q(data_98__10_) );
DFFPOSX1 DFFPOSX1_1596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_254__11_), .Q(data_98__11_) );
DFFPOSX1 DFFPOSX1_1597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_254__12_), .Q(data_98__12_) );
DFFPOSX1 DFFPOSX1_1598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_254__13_), .Q(data_98__13_) );
DFFPOSX1 DFFPOSX1_1599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_254__14_), .Q(data_98__14_) );
DFFPOSX1 DFFPOSX1_1600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_254__15_), .Q(data_98__15_) );
DFFPOSX1 DFFPOSX1_1601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_255__0_), .Q(data_99__0_) );
DFFPOSX1 DFFPOSX1_1602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_255__1_), .Q(data_99__1_) );
DFFPOSX1 DFFPOSX1_1603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_255__2_), .Q(data_99__2_) );
DFFPOSX1 DFFPOSX1_1604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_255__3_), .Q(data_99__3_) );
DFFPOSX1 DFFPOSX1_1605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_255__4_), .Q(data_99__4_) );
DFFPOSX1 DFFPOSX1_1606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_255__5_), .Q(data_99__5_) );
DFFPOSX1 DFFPOSX1_1607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_255__6_), .Q(data_99__6_) );
DFFPOSX1 DFFPOSX1_1608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_255__7_), .Q(data_99__7_) );
DFFPOSX1 DFFPOSX1_1609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_255__8_), .Q(data_99__8_) );
DFFPOSX1 DFFPOSX1_1610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_255__9_), .Q(data_99__9_) );
DFFPOSX1 DFFPOSX1_1611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_255__10_), .Q(data_99__10_) );
DFFPOSX1 DFFPOSX1_1612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_255__11_), .Q(data_99__11_) );
DFFPOSX1 DFFPOSX1_1613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_255__12_), .Q(data_99__12_) );
DFFPOSX1 DFFPOSX1_1614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_255__13_), .Q(data_99__13_) );
DFFPOSX1 DFFPOSX1_1615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_255__14_), .Q(data_99__14_) );
DFFPOSX1 DFFPOSX1_1616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_255__15_), .Q(data_99__15_) );
DFFPOSX1 DFFPOSX1_1617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_2__0_), .Q(data_100__0_) );
DFFPOSX1 DFFPOSX1_1618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_2__1_), .Q(data_100__1_) );
DFFPOSX1 DFFPOSX1_1619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_2__2_), .Q(data_100__2_) );
DFFPOSX1 DFFPOSX1_1620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_2__3_), .Q(data_100__3_) );
DFFPOSX1 DFFPOSX1_1621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_2__4_), .Q(data_100__4_) );
DFFPOSX1 DFFPOSX1_1622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_2__5_), .Q(data_100__5_) );
DFFPOSX1 DFFPOSX1_1623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_2__6_), .Q(data_100__6_) );
DFFPOSX1 DFFPOSX1_1624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_2__7_), .Q(data_100__7_) );
DFFPOSX1 DFFPOSX1_1625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_2__8_), .Q(data_100__8_) );
DFFPOSX1 DFFPOSX1_1626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_2__9_), .Q(data_100__9_) );
DFFPOSX1 DFFPOSX1_1627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_2__10_), .Q(data_100__10_) );
DFFPOSX1 DFFPOSX1_1628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_2__11_), .Q(data_100__11_) );
DFFPOSX1 DFFPOSX1_1629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_2__12_), .Q(data_100__12_) );
DFFPOSX1 DFFPOSX1_1630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_2__13_), .Q(data_100__13_) );
DFFPOSX1 DFFPOSX1_1631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_2__14_), .Q(data_100__14_) );
DFFPOSX1 DFFPOSX1_1632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_2__15_), .Q(data_100__15_) );
DFFPOSX1 DFFPOSX1_1633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_3__0_), .Q(data_101__0_) );
DFFPOSX1 DFFPOSX1_1634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_3__1_), .Q(data_101__1_) );
DFFPOSX1 DFFPOSX1_1635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_3__2_), .Q(data_101__2_) );
DFFPOSX1 DFFPOSX1_1636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_3__3_), .Q(data_101__3_) );
DFFPOSX1 DFFPOSX1_1637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_3__4_), .Q(data_101__4_) );
DFFPOSX1 DFFPOSX1_1638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_3__5_), .Q(data_101__5_) );
DFFPOSX1 DFFPOSX1_1639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_3__6_), .Q(data_101__6_) );
DFFPOSX1 DFFPOSX1_1640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_3__7_), .Q(data_101__7_) );
DFFPOSX1 DFFPOSX1_1641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_3__8_), .Q(data_101__8_) );
DFFPOSX1 DFFPOSX1_1642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_3__9_), .Q(data_101__9_) );
DFFPOSX1 DFFPOSX1_1643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_3__10_), .Q(data_101__10_) );
DFFPOSX1 DFFPOSX1_1644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_3__11_), .Q(data_101__11_) );
DFFPOSX1 DFFPOSX1_1645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_3__12_), .Q(data_101__12_) );
DFFPOSX1 DFFPOSX1_1646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_3__13_), .Q(data_101__13_) );
DFFPOSX1 DFFPOSX1_1647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_3__14_), .Q(data_101__14_) );
DFFPOSX1 DFFPOSX1_1648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_3__15_), .Q(data_101__15_) );
DFFPOSX1 DFFPOSX1_1649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_4__0_), .Q(data_102__0_) );
DFFPOSX1 DFFPOSX1_1650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_4__1_), .Q(data_102__1_) );
DFFPOSX1 DFFPOSX1_1651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_4__2_), .Q(data_102__2_) );
DFFPOSX1 DFFPOSX1_1652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_4__3_), .Q(data_102__3_) );
DFFPOSX1 DFFPOSX1_1653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_4__4_), .Q(data_102__4_) );
DFFPOSX1 DFFPOSX1_1654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_4__5_), .Q(data_102__5_) );
DFFPOSX1 DFFPOSX1_1655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_4__6_), .Q(data_102__6_) );
DFFPOSX1 DFFPOSX1_1656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_4__7_), .Q(data_102__7_) );
DFFPOSX1 DFFPOSX1_1657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_4__8_), .Q(data_102__8_) );
DFFPOSX1 DFFPOSX1_1658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_4__9_), .Q(data_102__9_) );
DFFPOSX1 DFFPOSX1_1659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_4__10_), .Q(data_102__10_) );
DFFPOSX1 DFFPOSX1_1660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_4__11_), .Q(data_102__11_) );
DFFPOSX1 DFFPOSX1_1661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_4__12_), .Q(data_102__12_) );
DFFPOSX1 DFFPOSX1_1662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_4__13_), .Q(data_102__13_) );
DFFPOSX1 DFFPOSX1_1663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_4__14_), .Q(data_102__14_) );
DFFPOSX1 DFFPOSX1_1664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_4__15_), .Q(data_102__15_) );
DFFPOSX1 DFFPOSX1_1665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_5__0_), .Q(data_103__0_) );
DFFPOSX1 DFFPOSX1_1666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_5__1_), .Q(data_103__1_) );
DFFPOSX1 DFFPOSX1_1667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_5__2_), .Q(data_103__2_) );
DFFPOSX1 DFFPOSX1_1668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_5__3_), .Q(data_103__3_) );
DFFPOSX1 DFFPOSX1_1669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_5__4_), .Q(data_103__4_) );
DFFPOSX1 DFFPOSX1_1670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_5__5_), .Q(data_103__5_) );
DFFPOSX1 DFFPOSX1_1671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_5__6_), .Q(data_103__6_) );
DFFPOSX1 DFFPOSX1_1672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_5__7_), .Q(data_103__7_) );
DFFPOSX1 DFFPOSX1_1673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_5__8_), .Q(data_103__8_) );
DFFPOSX1 DFFPOSX1_1674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_5__9_), .Q(data_103__9_) );
DFFPOSX1 DFFPOSX1_1675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_5__10_), .Q(data_103__10_) );
DFFPOSX1 DFFPOSX1_1676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_5__11_), .Q(data_103__11_) );
DFFPOSX1 DFFPOSX1_1677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_5__12_), .Q(data_103__12_) );
DFFPOSX1 DFFPOSX1_1678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_5__13_), .Q(data_103__13_) );
DFFPOSX1 DFFPOSX1_1679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_5__14_), .Q(data_103__14_) );
DFFPOSX1 DFFPOSX1_1680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_5__15_), .Q(data_103__15_) );
DFFPOSX1 DFFPOSX1_1681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_6__0_), .Q(data_104__0_) );
DFFPOSX1 DFFPOSX1_1682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_6__1_), .Q(data_104__1_) );
DFFPOSX1 DFFPOSX1_1683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_6__2_), .Q(data_104__2_) );
DFFPOSX1 DFFPOSX1_1684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_6__3_), .Q(data_104__3_) );
DFFPOSX1 DFFPOSX1_1685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_6__4_), .Q(data_104__4_) );
DFFPOSX1 DFFPOSX1_1686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_6__5_), .Q(data_104__5_) );
DFFPOSX1 DFFPOSX1_1687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_6__6_), .Q(data_104__6_) );
DFFPOSX1 DFFPOSX1_1688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_6__7_), .Q(data_104__7_) );
DFFPOSX1 DFFPOSX1_1689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_6__8_), .Q(data_104__8_) );
DFFPOSX1 DFFPOSX1_1690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_6__9_), .Q(data_104__9_) );
DFFPOSX1 DFFPOSX1_1691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_6__10_), .Q(data_104__10_) );
DFFPOSX1 DFFPOSX1_1692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_6__11_), .Q(data_104__11_) );
DFFPOSX1 DFFPOSX1_1693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_6__12_), .Q(data_104__12_) );
DFFPOSX1 DFFPOSX1_1694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_6__13_), .Q(data_104__13_) );
DFFPOSX1 DFFPOSX1_1695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_6__14_), .Q(data_104__14_) );
DFFPOSX1 DFFPOSX1_1696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_6__15_), .Q(data_104__15_) );
DFFPOSX1 DFFPOSX1_1697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_7__0_), .Q(data_105__0_) );
DFFPOSX1 DFFPOSX1_1698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_7__1_), .Q(data_105__1_) );
DFFPOSX1 DFFPOSX1_1699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_7__2_), .Q(data_105__2_) );
DFFPOSX1 DFFPOSX1_1700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_7__3_), .Q(data_105__3_) );
DFFPOSX1 DFFPOSX1_1701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_7__4_), .Q(data_105__4_) );
DFFPOSX1 DFFPOSX1_1702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_7__5_), .Q(data_105__5_) );
DFFPOSX1 DFFPOSX1_1703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_7__6_), .Q(data_105__6_) );
DFFPOSX1 DFFPOSX1_1704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_7__7_), .Q(data_105__7_) );
DFFPOSX1 DFFPOSX1_1705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_7__8_), .Q(data_105__8_) );
DFFPOSX1 DFFPOSX1_1706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_7__9_), .Q(data_105__9_) );
DFFPOSX1 DFFPOSX1_1707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_7__10_), .Q(data_105__10_) );
DFFPOSX1 DFFPOSX1_1708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_7__11_), .Q(data_105__11_) );
DFFPOSX1 DFFPOSX1_1709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_7__12_), .Q(data_105__12_) );
DFFPOSX1 DFFPOSX1_1710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_7__13_), .Q(data_105__13_) );
DFFPOSX1 DFFPOSX1_1711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_7__14_), .Q(data_105__14_) );
DFFPOSX1 DFFPOSX1_1712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_7__15_), .Q(data_105__15_) );
DFFPOSX1 DFFPOSX1_1713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_8__0_), .Q(data_106__0_) );
DFFPOSX1 DFFPOSX1_1714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_8__1_), .Q(data_106__1_) );
DFFPOSX1 DFFPOSX1_1715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_8__2_), .Q(data_106__2_) );
DFFPOSX1 DFFPOSX1_1716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_8__3_), .Q(data_106__3_) );
DFFPOSX1 DFFPOSX1_1717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_8__4_), .Q(data_106__4_) );
DFFPOSX1 DFFPOSX1_1718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_8__5_), .Q(data_106__5_) );
DFFPOSX1 DFFPOSX1_1719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_8__6_), .Q(data_106__6_) );
DFFPOSX1 DFFPOSX1_1720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_8__7_), .Q(data_106__7_) );
DFFPOSX1 DFFPOSX1_1721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_8__8_), .Q(data_106__8_) );
DFFPOSX1 DFFPOSX1_1722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_8__9_), .Q(data_106__9_) );
DFFPOSX1 DFFPOSX1_1723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_8__10_), .Q(data_106__10_) );
DFFPOSX1 DFFPOSX1_1724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_8__11_), .Q(data_106__11_) );
DFFPOSX1 DFFPOSX1_1725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_8__12_), .Q(data_106__12_) );
DFFPOSX1 DFFPOSX1_1726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_8__13_), .Q(data_106__13_) );
DFFPOSX1 DFFPOSX1_1727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_8__14_), .Q(data_106__14_) );
DFFPOSX1 DFFPOSX1_1728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_8__15_), .Q(data_106__15_) );
DFFPOSX1 DFFPOSX1_1729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_9__0_), .Q(data_107__0_) );
DFFPOSX1 DFFPOSX1_1730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_9__1_), .Q(data_107__1_) );
DFFPOSX1 DFFPOSX1_1731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_9__2_), .Q(data_107__2_) );
DFFPOSX1 DFFPOSX1_1732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_9__3_), .Q(data_107__3_) );
DFFPOSX1 DFFPOSX1_1733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_9__4_), .Q(data_107__4_) );
DFFPOSX1 DFFPOSX1_1734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_9__5_), .Q(data_107__5_) );
DFFPOSX1 DFFPOSX1_1735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_9__6_), .Q(data_107__6_) );
DFFPOSX1 DFFPOSX1_1736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_9__7_), .Q(data_107__7_) );
DFFPOSX1 DFFPOSX1_1737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_9__8_), .Q(data_107__8_) );
DFFPOSX1 DFFPOSX1_1738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_9__9_), .Q(data_107__9_) );
DFFPOSX1 DFFPOSX1_1739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_9__10_), .Q(data_107__10_) );
DFFPOSX1 DFFPOSX1_1740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_9__11_), .Q(data_107__11_) );
DFFPOSX1 DFFPOSX1_1741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_9__12_), .Q(data_107__12_) );
DFFPOSX1 DFFPOSX1_1742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_9__13_), .Q(data_107__13_) );
DFFPOSX1 DFFPOSX1_1743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_9__14_), .Q(data_107__14_) );
DFFPOSX1 DFFPOSX1_1744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_9__15_), .Q(data_107__15_) );
DFFPOSX1 DFFPOSX1_1745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_10__0_), .Q(data_108__0_) );
DFFPOSX1 DFFPOSX1_1746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_10__1_), .Q(data_108__1_) );
DFFPOSX1 DFFPOSX1_1747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_10__2_), .Q(data_108__2_) );
DFFPOSX1 DFFPOSX1_1748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_10__3_), .Q(data_108__3_) );
DFFPOSX1 DFFPOSX1_1749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_10__4_), .Q(data_108__4_) );
DFFPOSX1 DFFPOSX1_1750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_10__5_), .Q(data_108__5_) );
DFFPOSX1 DFFPOSX1_1751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_10__6_), .Q(data_108__6_) );
DFFPOSX1 DFFPOSX1_1752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_10__7_), .Q(data_108__7_) );
DFFPOSX1 DFFPOSX1_1753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_10__8_), .Q(data_108__8_) );
DFFPOSX1 DFFPOSX1_1754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_10__9_), .Q(data_108__9_) );
DFFPOSX1 DFFPOSX1_1755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_10__10_), .Q(data_108__10_) );
DFFPOSX1 DFFPOSX1_1756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_10__11_), .Q(data_108__11_) );
DFFPOSX1 DFFPOSX1_1757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10__12_), .Q(data_108__12_) );
DFFPOSX1 DFFPOSX1_1758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_10__13_), .Q(data_108__13_) );
DFFPOSX1 DFFPOSX1_1759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__14_), .Q(data_108__14_) );
DFFPOSX1 DFFPOSX1_1760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_10__15_), .Q(data_108__15_) );
DFFPOSX1 DFFPOSX1_1761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_11__0_), .Q(data_109__0_) );
DFFPOSX1 DFFPOSX1_1762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_11__1_), .Q(data_109__1_) );
DFFPOSX1 DFFPOSX1_1763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_11__2_), .Q(data_109__2_) );
DFFPOSX1 DFFPOSX1_1764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_11__3_), .Q(data_109__3_) );
DFFPOSX1 DFFPOSX1_1765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_11__4_), .Q(data_109__4_) );
DFFPOSX1 DFFPOSX1_1766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_11__5_), .Q(data_109__5_) );
DFFPOSX1 DFFPOSX1_1767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_11__6_), .Q(data_109__6_) );
DFFPOSX1 DFFPOSX1_1768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_11__7_), .Q(data_109__7_) );
DFFPOSX1 DFFPOSX1_1769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_11__8_), .Q(data_109__8_) );
DFFPOSX1 DFFPOSX1_1770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_11__9_), .Q(data_109__9_) );
DFFPOSX1 DFFPOSX1_1771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_11__10_), .Q(data_109__10_) );
DFFPOSX1 DFFPOSX1_1772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_11__11_), .Q(data_109__11_) );
DFFPOSX1 DFFPOSX1_1773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_11__12_), .Q(data_109__12_) );
DFFPOSX1 DFFPOSX1_1774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_11__13_), .Q(data_109__13_) );
DFFPOSX1 DFFPOSX1_1775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_11__14_), .Q(data_109__14_) );
DFFPOSX1 DFFPOSX1_1776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_11__15_), .Q(data_109__15_) );
DFFPOSX1 DFFPOSX1_1777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_13__0_), .Q(data_110__0_) );
DFFPOSX1 DFFPOSX1_1778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_13__1_), .Q(data_110__1_) );
DFFPOSX1 DFFPOSX1_1779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_13__2_), .Q(data_110__2_) );
DFFPOSX1 DFFPOSX1_1780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_13__3_), .Q(data_110__3_) );
DFFPOSX1 DFFPOSX1_1781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_13__4_), .Q(data_110__4_) );
DFFPOSX1 DFFPOSX1_1782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_13__5_), .Q(data_110__5_) );
DFFPOSX1 DFFPOSX1_1783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_13__6_), .Q(data_110__6_) );
DFFPOSX1 DFFPOSX1_1784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_13__7_), .Q(data_110__7_) );
DFFPOSX1 DFFPOSX1_1785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_13__8_), .Q(data_110__8_) );
DFFPOSX1 DFFPOSX1_1786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_13__9_), .Q(data_110__9_) );
DFFPOSX1 DFFPOSX1_1787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_13__10_), .Q(data_110__10_) );
DFFPOSX1 DFFPOSX1_1788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_13__11_), .Q(data_110__11_) );
DFFPOSX1 DFFPOSX1_1789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_13__12_), .Q(data_110__12_) );
DFFPOSX1 DFFPOSX1_1790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_13__13_), .Q(data_110__13_) );
DFFPOSX1 DFFPOSX1_1791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_13__14_), .Q(data_110__14_) );
DFFPOSX1 DFFPOSX1_1792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_13__15_), .Q(data_110__15_) );
DFFPOSX1 DFFPOSX1_1793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf0), .D(_14__0_), .Q(data_111__0_) );
DFFPOSX1 DFFPOSX1_1794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf0), .D(_14__1_), .Q(data_111__1_) );
DFFPOSX1 DFFPOSX1_1795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf0), .D(_14__2_), .Q(data_111__2_) );
DFFPOSX1 DFFPOSX1_1796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf0), .D(_14__3_), .Q(data_111__3_) );
DFFPOSX1 DFFPOSX1_1797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf0), .D(_14__4_), .Q(data_111__4_) );
DFFPOSX1 DFFPOSX1_1798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf0), .D(_14__5_), .Q(data_111__5_) );
DFFPOSX1 DFFPOSX1_1799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf0), .D(_14__6_), .Q(data_111__6_) );
DFFPOSX1 DFFPOSX1_1800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf0), .D(_14__7_), .Q(data_111__7_) );
DFFPOSX1 DFFPOSX1_1801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf0), .D(_14__8_), .Q(data_111__8_) );
DFFPOSX1 DFFPOSX1_1802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf0), .D(_14__9_), .Q(data_111__9_) );
DFFPOSX1 DFFPOSX1_1803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf0), .D(_14__10_), .Q(data_111__10_) );
DFFPOSX1 DFFPOSX1_1804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf0), .D(_14__11_), .Q(data_111__11_) );
DFFPOSX1 DFFPOSX1_1805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf0), .D(_14__12_), .Q(data_111__12_) );
DFFPOSX1 DFFPOSX1_1806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf0), .D(_14__13_), .Q(data_111__13_) );
DFFPOSX1 DFFPOSX1_1807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf0), .D(_14__14_), .Q(data_111__14_) );
DFFPOSX1 DFFPOSX1_1808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf0), .D(_14__15_), .Q(data_111__15_) );
DFFPOSX1 DFFPOSX1_1809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_15__0_), .Q(data_112__0_) );
DFFPOSX1 DFFPOSX1_1810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_15__1_), .Q(data_112__1_) );
DFFPOSX1 DFFPOSX1_1811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_15__2_), .Q(data_112__2_) );
DFFPOSX1 DFFPOSX1_1812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_15__3_), .Q(data_112__3_) );
DFFPOSX1 DFFPOSX1_1813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_15__4_), .Q(data_112__4_) );
DFFPOSX1 DFFPOSX1_1814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_15__5_), .Q(data_112__5_) );
DFFPOSX1 DFFPOSX1_1815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_15__6_), .Q(data_112__6_) );
DFFPOSX1 DFFPOSX1_1816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_15__7_), .Q(data_112__7_) );
DFFPOSX1 DFFPOSX1_1817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_15__8_), .Q(data_112__8_) );
DFFPOSX1 DFFPOSX1_1818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_15__9_), .Q(data_112__9_) );
DFFPOSX1 DFFPOSX1_1819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_15__10_), .Q(data_112__10_) );
DFFPOSX1 DFFPOSX1_1820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_15__11_), .Q(data_112__11_) );
DFFPOSX1 DFFPOSX1_1821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_15__12_), .Q(data_112__12_) );
DFFPOSX1 DFFPOSX1_1822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_15__13_), .Q(data_112__13_) );
DFFPOSX1 DFFPOSX1_1823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_15__14_), .Q(data_112__14_) );
DFFPOSX1 DFFPOSX1_1824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_15__15_), .Q(data_112__15_) );
DFFPOSX1 DFFPOSX1_1825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_16__0_), .Q(data_113__0_) );
DFFPOSX1 DFFPOSX1_1826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_16__1_), .Q(data_113__1_) );
DFFPOSX1 DFFPOSX1_1827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_16__2_), .Q(data_113__2_) );
DFFPOSX1 DFFPOSX1_1828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_16__3_), .Q(data_113__3_) );
DFFPOSX1 DFFPOSX1_1829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_16__4_), .Q(data_113__4_) );
DFFPOSX1 DFFPOSX1_1830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_16__5_), .Q(data_113__5_) );
DFFPOSX1 DFFPOSX1_1831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_16__6_), .Q(data_113__6_) );
DFFPOSX1 DFFPOSX1_1832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_16__7_), .Q(data_113__7_) );
DFFPOSX1 DFFPOSX1_1833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_16__8_), .Q(data_113__8_) );
DFFPOSX1 DFFPOSX1_1834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_16__9_), .Q(data_113__9_) );
DFFPOSX1 DFFPOSX1_1835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_16__10_), .Q(data_113__10_) );
DFFPOSX1 DFFPOSX1_1836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_16__11_), .Q(data_113__11_) );
DFFPOSX1 DFFPOSX1_1837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_16__12_), .Q(data_113__12_) );
DFFPOSX1 DFFPOSX1_1838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_16__13_), .Q(data_113__13_) );
DFFPOSX1 DFFPOSX1_1839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_16__14_), .Q(data_113__14_) );
DFFPOSX1 DFFPOSX1_1840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_16__15_), .Q(data_113__15_) );
DFFPOSX1 DFFPOSX1_1841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_17__0_), .Q(data_114__0_) );
DFFPOSX1 DFFPOSX1_1842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_17__1_), .Q(data_114__1_) );
DFFPOSX1 DFFPOSX1_1843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_17__2_), .Q(data_114__2_) );
DFFPOSX1 DFFPOSX1_1844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_17__3_), .Q(data_114__3_) );
DFFPOSX1 DFFPOSX1_1845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_17__4_), .Q(data_114__4_) );
DFFPOSX1 DFFPOSX1_1846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_17__5_), .Q(data_114__5_) );
DFFPOSX1 DFFPOSX1_1847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_17__6_), .Q(data_114__6_) );
DFFPOSX1 DFFPOSX1_1848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_17__7_), .Q(data_114__7_) );
DFFPOSX1 DFFPOSX1_1849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_17__8_), .Q(data_114__8_) );
DFFPOSX1 DFFPOSX1_1850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_17__9_), .Q(data_114__9_) );
DFFPOSX1 DFFPOSX1_1851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_17__10_), .Q(data_114__10_) );
DFFPOSX1 DFFPOSX1_1852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_17__11_), .Q(data_114__11_) );
DFFPOSX1 DFFPOSX1_1853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_17__12_), .Q(data_114__12_) );
DFFPOSX1 DFFPOSX1_1854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_17__13_), .Q(data_114__13_) );
DFFPOSX1 DFFPOSX1_1855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_17__14_), .Q(data_114__14_) );
DFFPOSX1 DFFPOSX1_1856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_17__15_), .Q(data_114__15_) );
DFFPOSX1 DFFPOSX1_1857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_18__0_), .Q(data_115__0_) );
DFFPOSX1 DFFPOSX1_1858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_18__1_), .Q(data_115__1_) );
DFFPOSX1 DFFPOSX1_1859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_18__2_), .Q(data_115__2_) );
DFFPOSX1 DFFPOSX1_1860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_18__3_), .Q(data_115__3_) );
DFFPOSX1 DFFPOSX1_1861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_18__4_), .Q(data_115__4_) );
DFFPOSX1 DFFPOSX1_1862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_18__5_), .Q(data_115__5_) );
DFFPOSX1 DFFPOSX1_1863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_18__6_), .Q(data_115__6_) );
DFFPOSX1 DFFPOSX1_1864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_18__7_), .Q(data_115__7_) );
DFFPOSX1 DFFPOSX1_1865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_18__8_), .Q(data_115__8_) );
DFFPOSX1 DFFPOSX1_1866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_18__9_), .Q(data_115__9_) );
DFFPOSX1 DFFPOSX1_1867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_18__10_), .Q(data_115__10_) );
DFFPOSX1 DFFPOSX1_1868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_18__11_), .Q(data_115__11_) );
DFFPOSX1 DFFPOSX1_1869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_18__12_), .Q(data_115__12_) );
DFFPOSX1 DFFPOSX1_1870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_18__13_), .Q(data_115__13_) );
DFFPOSX1 DFFPOSX1_1871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_18__14_), .Q(data_115__14_) );
DFFPOSX1 DFFPOSX1_1872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_18__15_), .Q(data_115__15_) );
DFFPOSX1 DFFPOSX1_1873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_19__0_), .Q(data_116__0_) );
DFFPOSX1 DFFPOSX1_1874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_19__1_), .Q(data_116__1_) );
DFFPOSX1 DFFPOSX1_1875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_19__2_), .Q(data_116__2_) );
DFFPOSX1 DFFPOSX1_1876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_19__3_), .Q(data_116__3_) );
DFFPOSX1 DFFPOSX1_1877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_19__4_), .Q(data_116__4_) );
DFFPOSX1 DFFPOSX1_1878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_19__5_), .Q(data_116__5_) );
DFFPOSX1 DFFPOSX1_1879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_19__6_), .Q(data_116__6_) );
DFFPOSX1 DFFPOSX1_1880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_19__7_), .Q(data_116__7_) );
DFFPOSX1 DFFPOSX1_1881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_19__8_), .Q(data_116__8_) );
DFFPOSX1 DFFPOSX1_1882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_19__9_), .Q(data_116__9_) );
DFFPOSX1 DFFPOSX1_1883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_19__10_), .Q(data_116__10_) );
DFFPOSX1 DFFPOSX1_1884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_19__11_), .Q(data_116__11_) );
DFFPOSX1 DFFPOSX1_1885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_19__12_), .Q(data_116__12_) );
DFFPOSX1 DFFPOSX1_1886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_19__13_), .Q(data_116__13_) );
DFFPOSX1 DFFPOSX1_1887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_19__14_), .Q(data_116__14_) );
DFFPOSX1 DFFPOSX1_1888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_19__15_), .Q(data_116__15_) );
DFFPOSX1 DFFPOSX1_1889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_20__0_), .Q(data_117__0_) );
DFFPOSX1 DFFPOSX1_1890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_20__1_), .Q(data_117__1_) );
DFFPOSX1 DFFPOSX1_1891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_20__2_), .Q(data_117__2_) );
DFFPOSX1 DFFPOSX1_1892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_20__3_), .Q(data_117__3_) );
DFFPOSX1 DFFPOSX1_1893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_20__4_), .Q(data_117__4_) );
DFFPOSX1 DFFPOSX1_1894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_20__5_), .Q(data_117__5_) );
DFFPOSX1 DFFPOSX1_1895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_20__6_), .Q(data_117__6_) );
DFFPOSX1 DFFPOSX1_1896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_20__7_), .Q(data_117__7_) );
DFFPOSX1 DFFPOSX1_1897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_20__8_), .Q(data_117__8_) );
DFFPOSX1 DFFPOSX1_1898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_20__9_), .Q(data_117__9_) );
DFFPOSX1 DFFPOSX1_1899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_20__10_), .Q(data_117__10_) );
DFFPOSX1 DFFPOSX1_1900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_20__11_), .Q(data_117__11_) );
DFFPOSX1 DFFPOSX1_1901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_20__12_), .Q(data_117__12_) );
DFFPOSX1 DFFPOSX1_1902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_20__13_), .Q(data_117__13_) );
DFFPOSX1 DFFPOSX1_1903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_20__14_), .Q(data_117__14_) );
DFFPOSX1 DFFPOSX1_1904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_20__15_), .Q(data_117__15_) );
DFFPOSX1 DFFPOSX1_1905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_21__0_), .Q(data_118__0_) );
DFFPOSX1 DFFPOSX1_1906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_21__1_), .Q(data_118__1_) );
DFFPOSX1 DFFPOSX1_1907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_21__2_), .Q(data_118__2_) );
DFFPOSX1 DFFPOSX1_1908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_21__3_), .Q(data_118__3_) );
DFFPOSX1 DFFPOSX1_1909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_21__4_), .Q(data_118__4_) );
DFFPOSX1 DFFPOSX1_1910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_21__5_), .Q(data_118__5_) );
DFFPOSX1 DFFPOSX1_1911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_21__6_), .Q(data_118__6_) );
DFFPOSX1 DFFPOSX1_1912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_21__7_), .Q(data_118__7_) );
DFFPOSX1 DFFPOSX1_1913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_21__8_), .Q(data_118__8_) );
DFFPOSX1 DFFPOSX1_1914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_21__9_), .Q(data_118__9_) );
DFFPOSX1 DFFPOSX1_1915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_21__10_), .Q(data_118__10_) );
DFFPOSX1 DFFPOSX1_1916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_21__11_), .Q(data_118__11_) );
DFFPOSX1 DFFPOSX1_1917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_21__12_), .Q(data_118__12_) );
DFFPOSX1 DFFPOSX1_1918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_21__13_), .Q(data_118__13_) );
DFFPOSX1 DFFPOSX1_1919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_21__14_), .Q(data_118__14_) );
DFFPOSX1 DFFPOSX1_1920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_21__15_), .Q(data_118__15_) );
DFFPOSX1 DFFPOSX1_1921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_22__0_), .Q(data_119__0_) );
DFFPOSX1 DFFPOSX1_1922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_22__1_), .Q(data_119__1_) );
DFFPOSX1 DFFPOSX1_1923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_22__2_), .Q(data_119__2_) );
DFFPOSX1 DFFPOSX1_1924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_22__3_), .Q(data_119__3_) );
DFFPOSX1 DFFPOSX1_1925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_22__4_), .Q(data_119__4_) );
DFFPOSX1 DFFPOSX1_1926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_22__5_), .Q(data_119__5_) );
DFFPOSX1 DFFPOSX1_1927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_22__6_), .Q(data_119__6_) );
DFFPOSX1 DFFPOSX1_1928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_22__7_), .Q(data_119__7_) );
DFFPOSX1 DFFPOSX1_1929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_22__8_), .Q(data_119__8_) );
DFFPOSX1 DFFPOSX1_1930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_22__9_), .Q(data_119__9_) );
DFFPOSX1 DFFPOSX1_1931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_22__10_), .Q(data_119__10_) );
DFFPOSX1 DFFPOSX1_1932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_22__11_), .Q(data_119__11_) );
DFFPOSX1 DFFPOSX1_1933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_22__12_), .Q(data_119__12_) );
DFFPOSX1 DFFPOSX1_1934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_22__13_), .Q(data_119__13_) );
DFFPOSX1 DFFPOSX1_1935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_22__14_), .Q(data_119__14_) );
DFFPOSX1 DFFPOSX1_1936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_22__15_), .Q(data_119__15_) );
DFFPOSX1 DFFPOSX1_1937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_24__0_), .Q(data_120__0_) );
DFFPOSX1 DFFPOSX1_1938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_24__1_), .Q(data_120__1_) );
DFFPOSX1 DFFPOSX1_1939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_24__2_), .Q(data_120__2_) );
DFFPOSX1 DFFPOSX1_1940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_24__3_), .Q(data_120__3_) );
DFFPOSX1 DFFPOSX1_1941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_24__4_), .Q(data_120__4_) );
DFFPOSX1 DFFPOSX1_1942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_24__5_), .Q(data_120__5_) );
DFFPOSX1 DFFPOSX1_1943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_24__6_), .Q(data_120__6_) );
DFFPOSX1 DFFPOSX1_1944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_24__7_), .Q(data_120__7_) );
DFFPOSX1 DFFPOSX1_1945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_24__8_), .Q(data_120__8_) );
DFFPOSX1 DFFPOSX1_1946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_24__9_), .Q(data_120__9_) );
DFFPOSX1 DFFPOSX1_1947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_24__10_), .Q(data_120__10_) );
DFFPOSX1 DFFPOSX1_1948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_24__11_), .Q(data_120__11_) );
DFFPOSX1 DFFPOSX1_1949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_24__12_), .Q(data_120__12_) );
DFFPOSX1 DFFPOSX1_1950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_24__13_), .Q(data_120__13_) );
DFFPOSX1 DFFPOSX1_1951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_24__14_), .Q(data_120__14_) );
DFFPOSX1 DFFPOSX1_1952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_24__15_), .Q(data_120__15_) );
DFFPOSX1 DFFPOSX1_1953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_25__0_), .Q(data_121__0_) );
DFFPOSX1 DFFPOSX1_1954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_25__1_), .Q(data_121__1_) );
DFFPOSX1 DFFPOSX1_1955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_25__2_), .Q(data_121__2_) );
DFFPOSX1 DFFPOSX1_1956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_25__3_), .Q(data_121__3_) );
DFFPOSX1 DFFPOSX1_1957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_25__4_), .Q(data_121__4_) );
DFFPOSX1 DFFPOSX1_1958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_25__5_), .Q(data_121__5_) );
DFFPOSX1 DFFPOSX1_1959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_25__6_), .Q(data_121__6_) );
DFFPOSX1 DFFPOSX1_1960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_25__7_), .Q(data_121__7_) );
DFFPOSX1 DFFPOSX1_1961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_25__8_), .Q(data_121__8_) );
DFFPOSX1 DFFPOSX1_1962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_25__9_), .Q(data_121__9_) );
DFFPOSX1 DFFPOSX1_1963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_25__10_), .Q(data_121__10_) );
DFFPOSX1 DFFPOSX1_1964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_25__11_), .Q(data_121__11_) );
DFFPOSX1 DFFPOSX1_1965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_25__12_), .Q(data_121__12_) );
DFFPOSX1 DFFPOSX1_1966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_25__13_), .Q(data_121__13_) );
DFFPOSX1 DFFPOSX1_1967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_25__14_), .Q(data_121__14_) );
DFFPOSX1 DFFPOSX1_1968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_25__15_), .Q(data_121__15_) );
DFFPOSX1 DFFPOSX1_1969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_26__0_), .Q(data_122__0_) );
DFFPOSX1 DFFPOSX1_1970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_26__1_), .Q(data_122__1_) );
DFFPOSX1 DFFPOSX1_1971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_26__2_), .Q(data_122__2_) );
DFFPOSX1 DFFPOSX1_1972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_26__3_), .Q(data_122__3_) );
DFFPOSX1 DFFPOSX1_1973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_26__4_), .Q(data_122__4_) );
DFFPOSX1 DFFPOSX1_1974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_26__5_), .Q(data_122__5_) );
DFFPOSX1 DFFPOSX1_1975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_26__6_), .Q(data_122__6_) );
DFFPOSX1 DFFPOSX1_1976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_26__7_), .Q(data_122__7_) );
DFFPOSX1 DFFPOSX1_1977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_26__8_), .Q(data_122__8_) );
DFFPOSX1 DFFPOSX1_1978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_26__9_), .Q(data_122__9_) );
DFFPOSX1 DFFPOSX1_1979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_26__10_), .Q(data_122__10_) );
DFFPOSX1 DFFPOSX1_1980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_26__11_), .Q(data_122__11_) );
DFFPOSX1 DFFPOSX1_1981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_26__12_), .Q(data_122__12_) );
DFFPOSX1 DFFPOSX1_1982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_26__13_), .Q(data_122__13_) );
DFFPOSX1 DFFPOSX1_1983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_26__14_), .Q(data_122__14_) );
DFFPOSX1 DFFPOSX1_1984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_26__15_), .Q(data_122__15_) );
DFFPOSX1 DFFPOSX1_1985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_27__0_), .Q(data_123__0_) );
DFFPOSX1 DFFPOSX1_1986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_27__1_), .Q(data_123__1_) );
DFFPOSX1 DFFPOSX1_1987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_27__2_), .Q(data_123__2_) );
DFFPOSX1 DFFPOSX1_1988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_27__3_), .Q(data_123__3_) );
DFFPOSX1 DFFPOSX1_1989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_27__4_), .Q(data_123__4_) );
DFFPOSX1 DFFPOSX1_1990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_27__5_), .Q(data_123__5_) );
DFFPOSX1 DFFPOSX1_1991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_27__6_), .Q(data_123__6_) );
DFFPOSX1 DFFPOSX1_1992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_27__7_), .Q(data_123__7_) );
DFFPOSX1 DFFPOSX1_1993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_27__8_), .Q(data_123__8_) );
DFFPOSX1 DFFPOSX1_1994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_27__9_), .Q(data_123__9_) );
DFFPOSX1 DFFPOSX1_1995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_27__10_), .Q(data_123__10_) );
DFFPOSX1 DFFPOSX1_1996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_27__11_), .Q(data_123__11_) );
DFFPOSX1 DFFPOSX1_1997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_27__12_), .Q(data_123__12_) );
DFFPOSX1 DFFPOSX1_1998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_27__13_), .Q(data_123__13_) );
DFFPOSX1 DFFPOSX1_1999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_27__14_), .Q(data_123__14_) );
DFFPOSX1 DFFPOSX1_2000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_27__15_), .Q(data_123__15_) );
DFFPOSX1 DFFPOSX1_2001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_28__0_), .Q(data_124__0_) );
DFFPOSX1 DFFPOSX1_2002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_28__1_), .Q(data_124__1_) );
DFFPOSX1 DFFPOSX1_2003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_28__2_), .Q(data_124__2_) );
DFFPOSX1 DFFPOSX1_2004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_28__3_), .Q(data_124__3_) );
DFFPOSX1 DFFPOSX1_2005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_28__4_), .Q(data_124__4_) );
DFFPOSX1 DFFPOSX1_2006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_28__5_), .Q(data_124__5_) );
DFFPOSX1 DFFPOSX1_2007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_28__6_), .Q(data_124__6_) );
DFFPOSX1 DFFPOSX1_2008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_28__7_), .Q(data_124__7_) );
DFFPOSX1 DFFPOSX1_2009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_28__8_), .Q(data_124__8_) );
DFFPOSX1 DFFPOSX1_2010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_28__9_), .Q(data_124__9_) );
DFFPOSX1 DFFPOSX1_2011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_28__10_), .Q(data_124__10_) );
DFFPOSX1 DFFPOSX1_2012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_28__11_), .Q(data_124__11_) );
DFFPOSX1 DFFPOSX1_2013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_28__12_), .Q(data_124__12_) );
DFFPOSX1 DFFPOSX1_2014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_28__13_), .Q(data_124__13_) );
DFFPOSX1 DFFPOSX1_2015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_28__14_), .Q(data_124__14_) );
DFFPOSX1 DFFPOSX1_2016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_28__15_), .Q(data_124__15_) );
DFFPOSX1 DFFPOSX1_2017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_29__0_), .Q(data_125__0_) );
DFFPOSX1 DFFPOSX1_2018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_29__1_), .Q(data_125__1_) );
DFFPOSX1 DFFPOSX1_2019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_29__2_), .Q(data_125__2_) );
DFFPOSX1 DFFPOSX1_2020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_29__3_), .Q(data_125__3_) );
DFFPOSX1 DFFPOSX1_2021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_29__4_), .Q(data_125__4_) );
DFFPOSX1 DFFPOSX1_2022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_29__5_), .Q(data_125__5_) );
DFFPOSX1 DFFPOSX1_2023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_29__6_), .Q(data_125__6_) );
DFFPOSX1 DFFPOSX1_2024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_29__7_), .Q(data_125__7_) );
DFFPOSX1 DFFPOSX1_2025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_29__8_), .Q(data_125__8_) );
DFFPOSX1 DFFPOSX1_2026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_29__9_), .Q(data_125__9_) );
DFFPOSX1 DFFPOSX1_2027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_29__10_), .Q(data_125__10_) );
DFFPOSX1 DFFPOSX1_2028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_29__11_), .Q(data_125__11_) );
DFFPOSX1 DFFPOSX1_2029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_29__12_), .Q(data_125__12_) );
DFFPOSX1 DFFPOSX1_2030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_29__13_), .Q(data_125__13_) );
DFFPOSX1 DFFPOSX1_2031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_29__14_), .Q(data_125__14_) );
DFFPOSX1 DFFPOSX1_2032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_29__15_), .Q(data_125__15_) );
DFFPOSX1 DFFPOSX1_2033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_30__0_), .Q(data_126__0_) );
DFFPOSX1 DFFPOSX1_2034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_30__1_), .Q(data_126__1_) );
DFFPOSX1 DFFPOSX1_2035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_30__2_), .Q(data_126__2_) );
DFFPOSX1 DFFPOSX1_2036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_30__3_), .Q(data_126__3_) );
DFFPOSX1 DFFPOSX1_2037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_30__4_), .Q(data_126__4_) );
DFFPOSX1 DFFPOSX1_2038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_30__5_), .Q(data_126__5_) );
DFFPOSX1 DFFPOSX1_2039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_30__6_), .Q(data_126__6_) );
DFFPOSX1 DFFPOSX1_2040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_30__7_), .Q(data_126__7_) );
DFFPOSX1 DFFPOSX1_2041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_30__8_), .Q(data_126__8_) );
DFFPOSX1 DFFPOSX1_2042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_30__9_), .Q(data_126__9_) );
DFFPOSX1 DFFPOSX1_2043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_30__10_), .Q(data_126__10_) );
DFFPOSX1 DFFPOSX1_2044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_30__11_), .Q(data_126__11_) );
DFFPOSX1 DFFPOSX1_2045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_30__12_), .Q(data_126__12_) );
DFFPOSX1 DFFPOSX1_2046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_30__13_), .Q(data_126__13_) );
DFFPOSX1 DFFPOSX1_2047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_30__14_), .Q(data_126__14_) );
DFFPOSX1 DFFPOSX1_2048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_30__15_), .Q(data_126__15_) );
DFFPOSX1 DFFPOSX1_2049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf3), .D(_31__0_), .Q(data_127__0_) );
DFFPOSX1 DFFPOSX1_2050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf3), .D(_31__1_), .Q(data_127__1_) );
DFFPOSX1 DFFPOSX1_2051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf3), .D(_31__2_), .Q(data_127__2_) );
DFFPOSX1 DFFPOSX1_2052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf3), .D(_31__3_), .Q(data_127__3_) );
DFFPOSX1 DFFPOSX1_2053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf3), .D(_31__4_), .Q(data_127__4_) );
DFFPOSX1 DFFPOSX1_2054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf3), .D(_31__5_), .Q(data_127__5_) );
DFFPOSX1 DFFPOSX1_2055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf3), .D(_31__6_), .Q(data_127__6_) );
DFFPOSX1 DFFPOSX1_2056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf3), .D(_31__7_), .Q(data_127__7_) );
DFFPOSX1 DFFPOSX1_2057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf3), .D(_31__8_), .Q(data_127__8_) );
DFFPOSX1 DFFPOSX1_2058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf3), .D(_31__9_), .Q(data_127__9_) );
DFFPOSX1 DFFPOSX1_2059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf3), .D(_31__10_), .Q(data_127__10_) );
DFFPOSX1 DFFPOSX1_2060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf3), .D(_31__11_), .Q(data_127__11_) );
DFFPOSX1 DFFPOSX1_2061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf3), .D(_31__12_), .Q(data_127__12_) );
DFFPOSX1 DFFPOSX1_2062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf3), .D(_31__13_), .Q(data_127__13_) );
DFFPOSX1 DFFPOSX1_2063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf3), .D(_31__14_), .Q(data_127__14_) );
DFFPOSX1 DFFPOSX1_2064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf3), .D(_31__15_), .Q(data_127__15_) );
DFFPOSX1 DFFPOSX1_2065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_32__0_), .Q(data_128__0_) );
DFFPOSX1 DFFPOSX1_2066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_32__1_), .Q(data_128__1_) );
DFFPOSX1 DFFPOSX1_2067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_32__2_), .Q(data_128__2_) );
DFFPOSX1 DFFPOSX1_2068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_32__3_), .Q(data_128__3_) );
DFFPOSX1 DFFPOSX1_2069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_32__4_), .Q(data_128__4_) );
DFFPOSX1 DFFPOSX1_2070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_32__5_), .Q(data_128__5_) );
DFFPOSX1 DFFPOSX1_2071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_32__6_), .Q(data_128__6_) );
DFFPOSX1 DFFPOSX1_2072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_32__7_), .Q(data_128__7_) );
DFFPOSX1 DFFPOSX1_2073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_32__8_), .Q(data_128__8_) );
DFFPOSX1 DFFPOSX1_2074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_32__9_), .Q(data_128__9_) );
DFFPOSX1 DFFPOSX1_2075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_32__10_), .Q(data_128__10_) );
DFFPOSX1 DFFPOSX1_2076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_32__11_), .Q(data_128__11_) );
DFFPOSX1 DFFPOSX1_2077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_32__12_), .Q(data_128__12_) );
DFFPOSX1 DFFPOSX1_2078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_32__13_), .Q(data_128__13_) );
DFFPOSX1 DFFPOSX1_2079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_32__14_), .Q(data_128__14_) );
DFFPOSX1 DFFPOSX1_2080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_32__15_), .Q(data_128__15_) );
DFFPOSX1 DFFPOSX1_2081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_33__0_), .Q(data_129__0_) );
DFFPOSX1 DFFPOSX1_2082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_33__1_), .Q(data_129__1_) );
DFFPOSX1 DFFPOSX1_2083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_33__2_), .Q(data_129__2_) );
DFFPOSX1 DFFPOSX1_2084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_33__3_), .Q(data_129__3_) );
DFFPOSX1 DFFPOSX1_2085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_33__4_), .Q(data_129__4_) );
DFFPOSX1 DFFPOSX1_2086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_33__5_), .Q(data_129__5_) );
DFFPOSX1 DFFPOSX1_2087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_33__6_), .Q(data_129__6_) );
DFFPOSX1 DFFPOSX1_2088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_33__7_), .Q(data_129__7_) );
DFFPOSX1 DFFPOSX1_2089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_33__8_), .Q(data_129__8_) );
DFFPOSX1 DFFPOSX1_2090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_33__9_), .Q(data_129__9_) );
DFFPOSX1 DFFPOSX1_2091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_33__10_), .Q(data_129__10_) );
DFFPOSX1 DFFPOSX1_2092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_33__11_), .Q(data_129__11_) );
DFFPOSX1 DFFPOSX1_2093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_33__12_), .Q(data_129__12_) );
DFFPOSX1 DFFPOSX1_2094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_33__13_), .Q(data_129__13_) );
DFFPOSX1 DFFPOSX1_2095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_33__14_), .Q(data_129__14_) );
DFFPOSX1 DFFPOSX1_2096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_33__15_), .Q(data_129__15_) );
DFFPOSX1 DFFPOSX1_2097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_35__0_), .Q(data_130__0_) );
DFFPOSX1 DFFPOSX1_2098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_35__1_), .Q(data_130__1_) );
DFFPOSX1 DFFPOSX1_2099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_35__2_), .Q(data_130__2_) );
DFFPOSX1 DFFPOSX1_2100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_35__3_), .Q(data_130__3_) );
DFFPOSX1 DFFPOSX1_2101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_35__4_), .Q(data_130__4_) );
DFFPOSX1 DFFPOSX1_2102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_35__5_), .Q(data_130__5_) );
DFFPOSX1 DFFPOSX1_2103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_35__6_), .Q(data_130__6_) );
DFFPOSX1 DFFPOSX1_2104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_35__7_), .Q(data_130__7_) );
DFFPOSX1 DFFPOSX1_2105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_35__8_), .Q(data_130__8_) );
DFFPOSX1 DFFPOSX1_2106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_35__9_), .Q(data_130__9_) );
DFFPOSX1 DFFPOSX1_2107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_35__10_), .Q(data_130__10_) );
DFFPOSX1 DFFPOSX1_2108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_35__11_), .Q(data_130__11_) );
DFFPOSX1 DFFPOSX1_2109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_35__12_), .Q(data_130__12_) );
DFFPOSX1 DFFPOSX1_2110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_35__13_), .Q(data_130__13_) );
DFFPOSX1 DFFPOSX1_2111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_35__14_), .Q(data_130__14_) );
DFFPOSX1 DFFPOSX1_2112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_35__15_), .Q(data_130__15_) );
DFFPOSX1 DFFPOSX1_2113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_36__0_), .Q(data_131__0_) );
DFFPOSX1 DFFPOSX1_2114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_36__1_), .Q(data_131__1_) );
DFFPOSX1 DFFPOSX1_2115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_36__2_), .Q(data_131__2_) );
DFFPOSX1 DFFPOSX1_2116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_36__3_), .Q(data_131__3_) );
DFFPOSX1 DFFPOSX1_2117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_36__4_), .Q(data_131__4_) );
DFFPOSX1 DFFPOSX1_2118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_36__5_), .Q(data_131__5_) );
DFFPOSX1 DFFPOSX1_2119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_36__6_), .Q(data_131__6_) );
DFFPOSX1 DFFPOSX1_2120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_36__7_), .Q(data_131__7_) );
DFFPOSX1 DFFPOSX1_2121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_36__8_), .Q(data_131__8_) );
DFFPOSX1 DFFPOSX1_2122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_36__9_), .Q(data_131__9_) );
DFFPOSX1 DFFPOSX1_2123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_36__10_), .Q(data_131__10_) );
DFFPOSX1 DFFPOSX1_2124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_36__11_), .Q(data_131__11_) );
DFFPOSX1 DFFPOSX1_2125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_36__12_), .Q(data_131__12_) );
DFFPOSX1 DFFPOSX1_2126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_36__13_), .Q(data_131__13_) );
DFFPOSX1 DFFPOSX1_2127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_36__14_), .Q(data_131__14_) );
DFFPOSX1 DFFPOSX1_2128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_36__15_), .Q(data_131__15_) );
DFFPOSX1 DFFPOSX1_2129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_37__0_), .Q(data_132__0_) );
DFFPOSX1 DFFPOSX1_2130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_37__1_), .Q(data_132__1_) );
DFFPOSX1 DFFPOSX1_2131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_37__2_), .Q(data_132__2_) );
DFFPOSX1 DFFPOSX1_2132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_37__3_), .Q(data_132__3_) );
DFFPOSX1 DFFPOSX1_2133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_37__4_), .Q(data_132__4_) );
DFFPOSX1 DFFPOSX1_2134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_37__5_), .Q(data_132__5_) );
DFFPOSX1 DFFPOSX1_2135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_37__6_), .Q(data_132__6_) );
DFFPOSX1 DFFPOSX1_2136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_37__7_), .Q(data_132__7_) );
DFFPOSX1 DFFPOSX1_2137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_37__8_), .Q(data_132__8_) );
DFFPOSX1 DFFPOSX1_2138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_37__9_), .Q(data_132__9_) );
DFFPOSX1 DFFPOSX1_2139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_37__10_), .Q(data_132__10_) );
DFFPOSX1 DFFPOSX1_2140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_37__11_), .Q(data_132__11_) );
DFFPOSX1 DFFPOSX1_2141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_37__12_), .Q(data_132__12_) );
DFFPOSX1 DFFPOSX1_2142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_37__13_), .Q(data_132__13_) );
DFFPOSX1 DFFPOSX1_2143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_37__14_), .Q(data_132__14_) );
DFFPOSX1 DFFPOSX1_2144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_37__15_), .Q(data_132__15_) );
DFFPOSX1 DFFPOSX1_2145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_38__0_), .Q(data_133__0_) );
DFFPOSX1 DFFPOSX1_2146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_38__1_), .Q(data_133__1_) );
DFFPOSX1 DFFPOSX1_2147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_38__2_), .Q(data_133__2_) );
DFFPOSX1 DFFPOSX1_2148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_38__3_), .Q(data_133__3_) );
DFFPOSX1 DFFPOSX1_2149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_38__4_), .Q(data_133__4_) );
DFFPOSX1 DFFPOSX1_2150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_38__5_), .Q(data_133__5_) );
DFFPOSX1 DFFPOSX1_2151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_38__6_), .Q(data_133__6_) );
DFFPOSX1 DFFPOSX1_2152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_38__7_), .Q(data_133__7_) );
DFFPOSX1 DFFPOSX1_2153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_38__8_), .Q(data_133__8_) );
DFFPOSX1 DFFPOSX1_2154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_38__9_), .Q(data_133__9_) );
DFFPOSX1 DFFPOSX1_2155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_38__10_), .Q(data_133__10_) );
DFFPOSX1 DFFPOSX1_2156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_38__11_), .Q(data_133__11_) );
DFFPOSX1 DFFPOSX1_2157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_38__12_), .Q(data_133__12_) );
DFFPOSX1 DFFPOSX1_2158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_38__13_), .Q(data_133__13_) );
DFFPOSX1 DFFPOSX1_2159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_38__14_), .Q(data_133__14_) );
DFFPOSX1 DFFPOSX1_2160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_38__15_), .Q(data_133__15_) );
DFFPOSX1 DFFPOSX1_2161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_39__0_), .Q(data_134__0_) );
DFFPOSX1 DFFPOSX1_2162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_39__1_), .Q(data_134__1_) );
DFFPOSX1 DFFPOSX1_2163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_39__2_), .Q(data_134__2_) );
DFFPOSX1 DFFPOSX1_2164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_39__3_), .Q(data_134__3_) );
DFFPOSX1 DFFPOSX1_2165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_39__4_), .Q(data_134__4_) );
DFFPOSX1 DFFPOSX1_2166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_39__5_), .Q(data_134__5_) );
DFFPOSX1 DFFPOSX1_2167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_39__6_), .Q(data_134__6_) );
DFFPOSX1 DFFPOSX1_2168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_39__7_), .Q(data_134__7_) );
DFFPOSX1 DFFPOSX1_2169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_39__8_), .Q(data_134__8_) );
DFFPOSX1 DFFPOSX1_2170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_39__9_), .Q(data_134__9_) );
DFFPOSX1 DFFPOSX1_2171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_39__10_), .Q(data_134__10_) );
DFFPOSX1 DFFPOSX1_2172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_39__11_), .Q(data_134__11_) );
DFFPOSX1 DFFPOSX1_2173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_39__12_), .Q(data_134__12_) );
DFFPOSX1 DFFPOSX1_2174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_39__13_), .Q(data_134__13_) );
DFFPOSX1 DFFPOSX1_2175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_39__14_), .Q(data_134__14_) );
DFFPOSX1 DFFPOSX1_2176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_39__15_), .Q(data_134__15_) );
DFFPOSX1 DFFPOSX1_2177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_40__0_), .Q(data_135__0_) );
DFFPOSX1 DFFPOSX1_2178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_40__1_), .Q(data_135__1_) );
DFFPOSX1 DFFPOSX1_2179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_40__2_), .Q(data_135__2_) );
DFFPOSX1 DFFPOSX1_2180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_40__3_), .Q(data_135__3_) );
DFFPOSX1 DFFPOSX1_2181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_40__4_), .Q(data_135__4_) );
DFFPOSX1 DFFPOSX1_2182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_40__5_), .Q(data_135__5_) );
DFFPOSX1 DFFPOSX1_2183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_40__6_), .Q(data_135__6_) );
DFFPOSX1 DFFPOSX1_2184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_40__7_), .Q(data_135__7_) );
DFFPOSX1 DFFPOSX1_2185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_40__8_), .Q(data_135__8_) );
DFFPOSX1 DFFPOSX1_2186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_40__9_), .Q(data_135__9_) );
DFFPOSX1 DFFPOSX1_2187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_40__10_), .Q(data_135__10_) );
DFFPOSX1 DFFPOSX1_2188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_40__11_), .Q(data_135__11_) );
DFFPOSX1 DFFPOSX1_2189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_40__12_), .Q(data_135__12_) );
DFFPOSX1 DFFPOSX1_2190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_40__13_), .Q(data_135__13_) );
DFFPOSX1 DFFPOSX1_2191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_40__14_), .Q(data_135__14_) );
DFFPOSX1 DFFPOSX1_2192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_40__15_), .Q(data_135__15_) );
DFFPOSX1 DFFPOSX1_2193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_41__0_), .Q(data_136__0_) );
DFFPOSX1 DFFPOSX1_2194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_41__1_), .Q(data_136__1_) );
DFFPOSX1 DFFPOSX1_2195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_41__2_), .Q(data_136__2_) );
DFFPOSX1 DFFPOSX1_2196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_41__3_), .Q(data_136__3_) );
DFFPOSX1 DFFPOSX1_2197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_41__4_), .Q(data_136__4_) );
DFFPOSX1 DFFPOSX1_2198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_41__5_), .Q(data_136__5_) );
DFFPOSX1 DFFPOSX1_2199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_41__6_), .Q(data_136__6_) );
DFFPOSX1 DFFPOSX1_2200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_41__7_), .Q(data_136__7_) );
DFFPOSX1 DFFPOSX1_2201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_41__8_), .Q(data_136__8_) );
DFFPOSX1 DFFPOSX1_2202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_41__9_), .Q(data_136__9_) );
DFFPOSX1 DFFPOSX1_2203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_41__10_), .Q(data_136__10_) );
DFFPOSX1 DFFPOSX1_2204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_41__11_), .Q(data_136__11_) );
DFFPOSX1 DFFPOSX1_2205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_41__12_), .Q(data_136__12_) );
DFFPOSX1 DFFPOSX1_2206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_41__13_), .Q(data_136__13_) );
DFFPOSX1 DFFPOSX1_2207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_41__14_), .Q(data_136__14_) );
DFFPOSX1 DFFPOSX1_2208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_41__15_), .Q(data_136__15_) );
DFFPOSX1 DFFPOSX1_2209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_42__0_), .Q(data_137__0_) );
DFFPOSX1 DFFPOSX1_2210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_42__1_), .Q(data_137__1_) );
DFFPOSX1 DFFPOSX1_2211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_42__2_), .Q(data_137__2_) );
DFFPOSX1 DFFPOSX1_2212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_42__3_), .Q(data_137__3_) );
DFFPOSX1 DFFPOSX1_2213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_42__4_), .Q(data_137__4_) );
DFFPOSX1 DFFPOSX1_2214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_42__5_), .Q(data_137__5_) );
DFFPOSX1 DFFPOSX1_2215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_42__6_), .Q(data_137__6_) );
DFFPOSX1 DFFPOSX1_2216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_42__7_), .Q(data_137__7_) );
DFFPOSX1 DFFPOSX1_2217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_42__8_), .Q(data_137__8_) );
DFFPOSX1 DFFPOSX1_2218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_42__9_), .Q(data_137__9_) );
DFFPOSX1 DFFPOSX1_2219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_42__10_), .Q(data_137__10_) );
DFFPOSX1 DFFPOSX1_2220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_42__11_), .Q(data_137__11_) );
DFFPOSX1 DFFPOSX1_2221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_42__12_), .Q(data_137__12_) );
DFFPOSX1 DFFPOSX1_2222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_42__13_), .Q(data_137__13_) );
DFFPOSX1 DFFPOSX1_2223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_42__14_), .Q(data_137__14_) );
DFFPOSX1 DFFPOSX1_2224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_42__15_), .Q(data_137__15_) );
DFFPOSX1 DFFPOSX1_2225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_43__0_), .Q(data_138__0_) );
DFFPOSX1 DFFPOSX1_2226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_43__1_), .Q(data_138__1_) );
DFFPOSX1 DFFPOSX1_2227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_43__2_), .Q(data_138__2_) );
DFFPOSX1 DFFPOSX1_2228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_43__3_), .Q(data_138__3_) );
DFFPOSX1 DFFPOSX1_2229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_43__4_), .Q(data_138__4_) );
DFFPOSX1 DFFPOSX1_2230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_43__5_), .Q(data_138__5_) );
DFFPOSX1 DFFPOSX1_2231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_43__6_), .Q(data_138__6_) );
DFFPOSX1 DFFPOSX1_2232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_43__7_), .Q(data_138__7_) );
DFFPOSX1 DFFPOSX1_2233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_43__8_), .Q(data_138__8_) );
DFFPOSX1 DFFPOSX1_2234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_43__9_), .Q(data_138__9_) );
DFFPOSX1 DFFPOSX1_2235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_43__10_), .Q(data_138__10_) );
DFFPOSX1 DFFPOSX1_2236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_43__11_), .Q(data_138__11_) );
DFFPOSX1 DFFPOSX1_2237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_43__12_), .Q(data_138__12_) );
DFFPOSX1 DFFPOSX1_2238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_43__13_), .Q(data_138__13_) );
DFFPOSX1 DFFPOSX1_2239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_43__14_), .Q(data_138__14_) );
DFFPOSX1 DFFPOSX1_2240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_43__15_), .Q(data_138__15_) );
DFFPOSX1 DFFPOSX1_2241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_44__0_), .Q(data_139__0_) );
DFFPOSX1 DFFPOSX1_2242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_44__1_), .Q(data_139__1_) );
DFFPOSX1 DFFPOSX1_2243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_44__2_), .Q(data_139__2_) );
DFFPOSX1 DFFPOSX1_2244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_44__3_), .Q(data_139__3_) );
DFFPOSX1 DFFPOSX1_2245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_44__4_), .Q(data_139__4_) );
DFFPOSX1 DFFPOSX1_2246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_44__5_), .Q(data_139__5_) );
DFFPOSX1 DFFPOSX1_2247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_44__6_), .Q(data_139__6_) );
DFFPOSX1 DFFPOSX1_2248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_44__7_), .Q(data_139__7_) );
DFFPOSX1 DFFPOSX1_2249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_44__8_), .Q(data_139__8_) );
DFFPOSX1 DFFPOSX1_2250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_44__9_), .Q(data_139__9_) );
DFFPOSX1 DFFPOSX1_2251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_44__10_), .Q(data_139__10_) );
DFFPOSX1 DFFPOSX1_2252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_44__11_), .Q(data_139__11_) );
DFFPOSX1 DFFPOSX1_2253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_44__12_), .Q(data_139__12_) );
DFFPOSX1 DFFPOSX1_2254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_44__13_), .Q(data_139__13_) );
DFFPOSX1 DFFPOSX1_2255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_44__14_), .Q(data_139__14_) );
DFFPOSX1 DFFPOSX1_2256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_44__15_), .Q(data_139__15_) );
DFFPOSX1 DFFPOSX1_2257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_46__0_), .Q(data_140__0_) );
DFFPOSX1 DFFPOSX1_2258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_46__1_), .Q(data_140__1_) );
DFFPOSX1 DFFPOSX1_2259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_46__2_), .Q(data_140__2_) );
DFFPOSX1 DFFPOSX1_2260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_46__3_), .Q(data_140__3_) );
DFFPOSX1 DFFPOSX1_2261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_46__4_), .Q(data_140__4_) );
DFFPOSX1 DFFPOSX1_2262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_46__5_), .Q(data_140__5_) );
DFFPOSX1 DFFPOSX1_2263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_46__6_), .Q(data_140__6_) );
DFFPOSX1 DFFPOSX1_2264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_46__7_), .Q(data_140__7_) );
DFFPOSX1 DFFPOSX1_2265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_46__8_), .Q(data_140__8_) );
DFFPOSX1 DFFPOSX1_2266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_46__9_), .Q(data_140__9_) );
DFFPOSX1 DFFPOSX1_2267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_46__10_), .Q(data_140__10_) );
DFFPOSX1 DFFPOSX1_2268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_46__11_), .Q(data_140__11_) );
DFFPOSX1 DFFPOSX1_2269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_46__12_), .Q(data_140__12_) );
DFFPOSX1 DFFPOSX1_2270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_46__13_), .Q(data_140__13_) );
DFFPOSX1 DFFPOSX1_2271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_46__14_), .Q(data_140__14_) );
DFFPOSX1 DFFPOSX1_2272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_46__15_), .Q(data_140__15_) );
DFFPOSX1 DFFPOSX1_2273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_47__0_), .Q(data_141__0_) );
DFFPOSX1 DFFPOSX1_2274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_47__1_), .Q(data_141__1_) );
DFFPOSX1 DFFPOSX1_2275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_47__2_), .Q(data_141__2_) );
DFFPOSX1 DFFPOSX1_2276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_47__3_), .Q(data_141__3_) );
DFFPOSX1 DFFPOSX1_2277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_47__4_), .Q(data_141__4_) );
DFFPOSX1 DFFPOSX1_2278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_47__5_), .Q(data_141__5_) );
DFFPOSX1 DFFPOSX1_2279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_47__6_), .Q(data_141__6_) );
DFFPOSX1 DFFPOSX1_2280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_47__7_), .Q(data_141__7_) );
DFFPOSX1 DFFPOSX1_2281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_47__8_), .Q(data_141__8_) );
DFFPOSX1 DFFPOSX1_2282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_47__9_), .Q(data_141__9_) );
DFFPOSX1 DFFPOSX1_2283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_47__10_), .Q(data_141__10_) );
DFFPOSX1 DFFPOSX1_2284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_47__11_), .Q(data_141__11_) );
DFFPOSX1 DFFPOSX1_2285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_47__12_), .Q(data_141__12_) );
DFFPOSX1 DFFPOSX1_2286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_47__13_), .Q(data_141__13_) );
DFFPOSX1 DFFPOSX1_2287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_47__14_), .Q(data_141__14_) );
DFFPOSX1 DFFPOSX1_2288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_47__15_), .Q(data_141__15_) );
DFFPOSX1 DFFPOSX1_2289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_48__0_), .Q(data_142__0_) );
DFFPOSX1 DFFPOSX1_2290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_48__1_), .Q(data_142__1_) );
DFFPOSX1 DFFPOSX1_2291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_48__2_), .Q(data_142__2_) );
DFFPOSX1 DFFPOSX1_2292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_48__3_), .Q(data_142__3_) );
DFFPOSX1 DFFPOSX1_2293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_48__4_), .Q(data_142__4_) );
DFFPOSX1 DFFPOSX1_2294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_48__5_), .Q(data_142__5_) );
DFFPOSX1 DFFPOSX1_2295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_48__6_), .Q(data_142__6_) );
DFFPOSX1 DFFPOSX1_2296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_48__7_), .Q(data_142__7_) );
DFFPOSX1 DFFPOSX1_2297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_48__8_), .Q(data_142__8_) );
DFFPOSX1 DFFPOSX1_2298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_48__9_), .Q(data_142__9_) );
DFFPOSX1 DFFPOSX1_2299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_48__10_), .Q(data_142__10_) );
DFFPOSX1 DFFPOSX1_2300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_48__11_), .Q(data_142__11_) );
DFFPOSX1 DFFPOSX1_2301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_48__12_), .Q(data_142__12_) );
DFFPOSX1 DFFPOSX1_2302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_48__13_), .Q(data_142__13_) );
DFFPOSX1 DFFPOSX1_2303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_48__14_), .Q(data_142__14_) );
DFFPOSX1 DFFPOSX1_2304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_48__15_), .Q(data_142__15_) );
DFFPOSX1 DFFPOSX1_2305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf2), .D(_49__0_), .Q(data_143__0_) );
DFFPOSX1 DFFPOSX1_2306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf2), .D(_49__1_), .Q(data_143__1_) );
DFFPOSX1 DFFPOSX1_2307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf2), .D(_49__2_), .Q(data_143__2_) );
DFFPOSX1 DFFPOSX1_2308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf2), .D(_49__3_), .Q(data_143__3_) );
DFFPOSX1 DFFPOSX1_2309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf2), .D(_49__4_), .Q(data_143__4_) );
DFFPOSX1 DFFPOSX1_2310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf2), .D(_49__5_), .Q(data_143__5_) );
DFFPOSX1 DFFPOSX1_2311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf2), .D(_49__6_), .Q(data_143__6_) );
DFFPOSX1 DFFPOSX1_2312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf2), .D(_49__7_), .Q(data_143__7_) );
DFFPOSX1 DFFPOSX1_2313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf2), .D(_49__8_), .Q(data_143__8_) );
DFFPOSX1 DFFPOSX1_2314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf2), .D(_49__9_), .Q(data_143__9_) );
DFFPOSX1 DFFPOSX1_2315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf2), .D(_49__10_), .Q(data_143__10_) );
DFFPOSX1 DFFPOSX1_2316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf2), .D(_49__11_), .Q(data_143__11_) );
DFFPOSX1 DFFPOSX1_2317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf2), .D(_49__12_), .Q(data_143__12_) );
DFFPOSX1 DFFPOSX1_2318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf2), .D(_49__13_), .Q(data_143__13_) );
DFFPOSX1 DFFPOSX1_2319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf2), .D(_49__14_), .Q(data_143__14_) );
DFFPOSX1 DFFPOSX1_2320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf2), .D(_49__15_), .Q(data_143__15_) );
DFFPOSX1 DFFPOSX1_2321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_50__0_), .Q(data_144__0_) );
DFFPOSX1 DFFPOSX1_2322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_50__1_), .Q(data_144__1_) );
DFFPOSX1 DFFPOSX1_2323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_50__2_), .Q(data_144__2_) );
DFFPOSX1 DFFPOSX1_2324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_50__3_), .Q(data_144__3_) );
DFFPOSX1 DFFPOSX1_2325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_50__4_), .Q(data_144__4_) );
DFFPOSX1 DFFPOSX1_2326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_50__5_), .Q(data_144__5_) );
DFFPOSX1 DFFPOSX1_2327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_50__6_), .Q(data_144__6_) );
DFFPOSX1 DFFPOSX1_2328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_50__7_), .Q(data_144__7_) );
DFFPOSX1 DFFPOSX1_2329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_50__8_), .Q(data_144__8_) );
DFFPOSX1 DFFPOSX1_2330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_50__9_), .Q(data_144__9_) );
DFFPOSX1 DFFPOSX1_2331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_50__10_), .Q(data_144__10_) );
DFFPOSX1 DFFPOSX1_2332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_50__11_), .Q(data_144__11_) );
DFFPOSX1 DFFPOSX1_2333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_50__12_), .Q(data_144__12_) );
DFFPOSX1 DFFPOSX1_2334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_50__13_), .Q(data_144__13_) );
DFFPOSX1 DFFPOSX1_2335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_50__14_), .Q(data_144__14_) );
DFFPOSX1 DFFPOSX1_2336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_50__15_), .Q(data_144__15_) );
DFFPOSX1 DFFPOSX1_2337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_51__0_), .Q(data_145__0_) );
DFFPOSX1 DFFPOSX1_2338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_51__1_), .Q(data_145__1_) );
DFFPOSX1 DFFPOSX1_2339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_51__2_), .Q(data_145__2_) );
DFFPOSX1 DFFPOSX1_2340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_51__3_), .Q(data_145__3_) );
DFFPOSX1 DFFPOSX1_2341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_51__4_), .Q(data_145__4_) );
DFFPOSX1 DFFPOSX1_2342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_51__5_), .Q(data_145__5_) );
DFFPOSX1 DFFPOSX1_2343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_51__6_), .Q(data_145__6_) );
DFFPOSX1 DFFPOSX1_2344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_51__7_), .Q(data_145__7_) );
DFFPOSX1 DFFPOSX1_2345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_51__8_), .Q(data_145__8_) );
DFFPOSX1 DFFPOSX1_2346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_51__9_), .Q(data_145__9_) );
DFFPOSX1 DFFPOSX1_2347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_51__10_), .Q(data_145__10_) );
DFFPOSX1 DFFPOSX1_2348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_51__11_), .Q(data_145__11_) );
DFFPOSX1 DFFPOSX1_2349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_51__12_), .Q(data_145__12_) );
DFFPOSX1 DFFPOSX1_2350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_51__13_), .Q(data_145__13_) );
DFFPOSX1 DFFPOSX1_2351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_51__14_), .Q(data_145__14_) );
DFFPOSX1 DFFPOSX1_2352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_51__15_), .Q(data_145__15_) );
DFFPOSX1 DFFPOSX1_2353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_52__0_), .Q(data_146__0_) );
DFFPOSX1 DFFPOSX1_2354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_52__1_), .Q(data_146__1_) );
DFFPOSX1 DFFPOSX1_2355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_52__2_), .Q(data_146__2_) );
DFFPOSX1 DFFPOSX1_2356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_52__3_), .Q(data_146__3_) );
DFFPOSX1 DFFPOSX1_2357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_52__4_), .Q(data_146__4_) );
DFFPOSX1 DFFPOSX1_2358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_52__5_), .Q(data_146__5_) );
DFFPOSX1 DFFPOSX1_2359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_52__6_), .Q(data_146__6_) );
DFFPOSX1 DFFPOSX1_2360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_52__7_), .Q(data_146__7_) );
DFFPOSX1 DFFPOSX1_2361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_52__8_), .Q(data_146__8_) );
DFFPOSX1 DFFPOSX1_2362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_52__9_), .Q(data_146__9_) );
DFFPOSX1 DFFPOSX1_2363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_52__10_), .Q(data_146__10_) );
DFFPOSX1 DFFPOSX1_2364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_52__11_), .Q(data_146__11_) );
DFFPOSX1 DFFPOSX1_2365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_52__12_), .Q(data_146__12_) );
DFFPOSX1 DFFPOSX1_2366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_52__13_), .Q(data_146__13_) );
DFFPOSX1 DFFPOSX1_2367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_52__14_), .Q(data_146__14_) );
DFFPOSX1 DFFPOSX1_2368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_52__15_), .Q(data_146__15_) );
DFFPOSX1 DFFPOSX1_2369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_53__0_), .Q(data_147__0_) );
DFFPOSX1 DFFPOSX1_2370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_53__1_), .Q(data_147__1_) );
DFFPOSX1 DFFPOSX1_2371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_53__2_), .Q(data_147__2_) );
DFFPOSX1 DFFPOSX1_2372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_53__3_), .Q(data_147__3_) );
DFFPOSX1 DFFPOSX1_2373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_53__4_), .Q(data_147__4_) );
DFFPOSX1 DFFPOSX1_2374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_53__5_), .Q(data_147__5_) );
DFFPOSX1 DFFPOSX1_2375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_53__6_), .Q(data_147__6_) );
DFFPOSX1 DFFPOSX1_2376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_53__7_), .Q(data_147__7_) );
DFFPOSX1 DFFPOSX1_2377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_53__8_), .Q(data_147__8_) );
DFFPOSX1 DFFPOSX1_2378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_53__9_), .Q(data_147__9_) );
DFFPOSX1 DFFPOSX1_2379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_53__10_), .Q(data_147__10_) );
DFFPOSX1 DFFPOSX1_2380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_53__11_), .Q(data_147__11_) );
DFFPOSX1 DFFPOSX1_2381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_53__12_), .Q(data_147__12_) );
DFFPOSX1 DFFPOSX1_2382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_53__13_), .Q(data_147__13_) );
DFFPOSX1 DFFPOSX1_2383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_53__14_), .Q(data_147__14_) );
DFFPOSX1 DFFPOSX1_2384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_53__15_), .Q(data_147__15_) );
DFFPOSX1 DFFPOSX1_2385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_54__0_), .Q(data_148__0_) );
DFFPOSX1 DFFPOSX1_2386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_54__1_), .Q(data_148__1_) );
DFFPOSX1 DFFPOSX1_2387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_54__2_), .Q(data_148__2_) );
DFFPOSX1 DFFPOSX1_2388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_54__3_), .Q(data_148__3_) );
DFFPOSX1 DFFPOSX1_2389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_54__4_), .Q(data_148__4_) );
DFFPOSX1 DFFPOSX1_2390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_54__5_), .Q(data_148__5_) );
DFFPOSX1 DFFPOSX1_2391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_54__6_), .Q(data_148__6_) );
DFFPOSX1 DFFPOSX1_2392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_54__7_), .Q(data_148__7_) );
DFFPOSX1 DFFPOSX1_2393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_54__8_), .Q(data_148__8_) );
DFFPOSX1 DFFPOSX1_2394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_54__9_), .Q(data_148__9_) );
DFFPOSX1 DFFPOSX1_2395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_54__10_), .Q(data_148__10_) );
DFFPOSX1 DFFPOSX1_2396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_54__11_), .Q(data_148__11_) );
DFFPOSX1 DFFPOSX1_2397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_54__12_), .Q(data_148__12_) );
DFFPOSX1 DFFPOSX1_2398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_54__13_), .Q(data_148__13_) );
DFFPOSX1 DFFPOSX1_2399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_54__14_), .Q(data_148__14_) );
DFFPOSX1 DFFPOSX1_2400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_54__15_), .Q(data_148__15_) );
DFFPOSX1 DFFPOSX1_2401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_55__0_), .Q(data_149__0_) );
DFFPOSX1 DFFPOSX1_2402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_55__1_), .Q(data_149__1_) );
DFFPOSX1 DFFPOSX1_2403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_55__2_), .Q(data_149__2_) );
DFFPOSX1 DFFPOSX1_2404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_55__3_), .Q(data_149__3_) );
DFFPOSX1 DFFPOSX1_2405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_55__4_), .Q(data_149__4_) );
DFFPOSX1 DFFPOSX1_2406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_55__5_), .Q(data_149__5_) );
DFFPOSX1 DFFPOSX1_2407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_55__6_), .Q(data_149__6_) );
DFFPOSX1 DFFPOSX1_2408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_55__7_), .Q(data_149__7_) );
DFFPOSX1 DFFPOSX1_2409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_55__8_), .Q(data_149__8_) );
DFFPOSX1 DFFPOSX1_2410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_55__9_), .Q(data_149__9_) );
DFFPOSX1 DFFPOSX1_2411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_55__10_), .Q(data_149__10_) );
DFFPOSX1 DFFPOSX1_2412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_55__11_), .Q(data_149__11_) );
DFFPOSX1 DFFPOSX1_2413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_55__12_), .Q(data_149__12_) );
DFFPOSX1 DFFPOSX1_2414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_55__13_), .Q(data_149__13_) );
DFFPOSX1 DFFPOSX1_2415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_55__14_), .Q(data_149__14_) );
DFFPOSX1 DFFPOSX1_2416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_55__15_), .Q(data_149__15_) );
DFFPOSX1 DFFPOSX1_2417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_57__0_), .Q(data_150__0_) );
DFFPOSX1 DFFPOSX1_2418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_57__1_), .Q(data_150__1_) );
DFFPOSX1 DFFPOSX1_2419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_57__2_), .Q(data_150__2_) );
DFFPOSX1 DFFPOSX1_2420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_57__3_), .Q(data_150__3_) );
DFFPOSX1 DFFPOSX1_2421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_57__4_), .Q(data_150__4_) );
DFFPOSX1 DFFPOSX1_2422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_57__5_), .Q(data_150__5_) );
DFFPOSX1 DFFPOSX1_2423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_57__6_), .Q(data_150__6_) );
DFFPOSX1 DFFPOSX1_2424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_57__7_), .Q(data_150__7_) );
DFFPOSX1 DFFPOSX1_2425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_57__8_), .Q(data_150__8_) );
DFFPOSX1 DFFPOSX1_2426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_57__9_), .Q(data_150__9_) );
DFFPOSX1 DFFPOSX1_2427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_57__10_), .Q(data_150__10_) );
DFFPOSX1 DFFPOSX1_2428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_57__11_), .Q(data_150__11_) );
DFFPOSX1 DFFPOSX1_2429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_57__12_), .Q(data_150__12_) );
DFFPOSX1 DFFPOSX1_2430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_57__13_), .Q(data_150__13_) );
DFFPOSX1 DFFPOSX1_2431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_57__14_), .Q(data_150__14_) );
DFFPOSX1 DFFPOSX1_2432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_57__15_), .Q(data_150__15_) );
DFFPOSX1 DFFPOSX1_2433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_58__0_), .Q(data_151__0_) );
DFFPOSX1 DFFPOSX1_2434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_58__1_), .Q(data_151__1_) );
DFFPOSX1 DFFPOSX1_2435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_58__2_), .Q(data_151__2_) );
DFFPOSX1 DFFPOSX1_2436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_58__3_), .Q(data_151__3_) );
DFFPOSX1 DFFPOSX1_2437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_58__4_), .Q(data_151__4_) );
DFFPOSX1 DFFPOSX1_2438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_58__5_), .Q(data_151__5_) );
DFFPOSX1 DFFPOSX1_2439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_58__6_), .Q(data_151__6_) );
DFFPOSX1 DFFPOSX1_2440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_58__7_), .Q(data_151__7_) );
DFFPOSX1 DFFPOSX1_2441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_58__8_), .Q(data_151__8_) );
DFFPOSX1 DFFPOSX1_2442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_58__9_), .Q(data_151__9_) );
DFFPOSX1 DFFPOSX1_2443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_58__10_), .Q(data_151__10_) );
DFFPOSX1 DFFPOSX1_2444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_58__11_), .Q(data_151__11_) );
DFFPOSX1 DFFPOSX1_2445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_58__12_), .Q(data_151__12_) );
DFFPOSX1 DFFPOSX1_2446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_58__13_), .Q(data_151__13_) );
DFFPOSX1 DFFPOSX1_2447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_58__14_), .Q(data_151__14_) );
DFFPOSX1 DFFPOSX1_2448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_58__15_), .Q(data_151__15_) );
DFFPOSX1 DFFPOSX1_2449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_59__0_), .Q(data_152__0_) );
DFFPOSX1 DFFPOSX1_2450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_59__1_), .Q(data_152__1_) );
DFFPOSX1 DFFPOSX1_2451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_59__2_), .Q(data_152__2_) );
DFFPOSX1 DFFPOSX1_2452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_59__3_), .Q(data_152__3_) );
DFFPOSX1 DFFPOSX1_2453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_59__4_), .Q(data_152__4_) );
DFFPOSX1 DFFPOSX1_2454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_59__5_), .Q(data_152__5_) );
DFFPOSX1 DFFPOSX1_2455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_59__6_), .Q(data_152__6_) );
DFFPOSX1 DFFPOSX1_2456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_59__7_), .Q(data_152__7_) );
DFFPOSX1 DFFPOSX1_2457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_59__8_), .Q(data_152__8_) );
DFFPOSX1 DFFPOSX1_2458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_59__9_), .Q(data_152__9_) );
DFFPOSX1 DFFPOSX1_2459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_59__10_), .Q(data_152__10_) );
DFFPOSX1 DFFPOSX1_2460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_59__11_), .Q(data_152__11_) );
DFFPOSX1 DFFPOSX1_2461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_59__12_), .Q(data_152__12_) );
DFFPOSX1 DFFPOSX1_2462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_59__13_), .Q(data_152__13_) );
DFFPOSX1 DFFPOSX1_2463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_59__14_), .Q(data_152__14_) );
DFFPOSX1 DFFPOSX1_2464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_59__15_), .Q(data_152__15_) );
DFFPOSX1 DFFPOSX1_2465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_60__0_), .Q(data_153__0_) );
DFFPOSX1 DFFPOSX1_2466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_60__1_), .Q(data_153__1_) );
DFFPOSX1 DFFPOSX1_2467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_60__2_), .Q(data_153__2_) );
DFFPOSX1 DFFPOSX1_2468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_60__3_), .Q(data_153__3_) );
DFFPOSX1 DFFPOSX1_2469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_60__4_), .Q(data_153__4_) );
DFFPOSX1 DFFPOSX1_2470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_60__5_), .Q(data_153__5_) );
DFFPOSX1 DFFPOSX1_2471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_60__6_), .Q(data_153__6_) );
DFFPOSX1 DFFPOSX1_2472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_60__7_), .Q(data_153__7_) );
DFFPOSX1 DFFPOSX1_2473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_60__8_), .Q(data_153__8_) );
DFFPOSX1 DFFPOSX1_2474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_60__9_), .Q(data_153__9_) );
DFFPOSX1 DFFPOSX1_2475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_60__10_), .Q(data_153__10_) );
DFFPOSX1 DFFPOSX1_2476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_60__11_), .Q(data_153__11_) );
DFFPOSX1 DFFPOSX1_2477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_60__12_), .Q(data_153__12_) );
DFFPOSX1 DFFPOSX1_2478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_60__13_), .Q(data_153__13_) );
DFFPOSX1 DFFPOSX1_2479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_60__14_), .Q(data_153__14_) );
DFFPOSX1 DFFPOSX1_2480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_60__15_), .Q(data_153__15_) );
DFFPOSX1 DFFPOSX1_2481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_61__0_), .Q(data_154__0_) );
DFFPOSX1 DFFPOSX1_2482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_61__1_), .Q(data_154__1_) );
DFFPOSX1 DFFPOSX1_2483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_61__2_), .Q(data_154__2_) );
DFFPOSX1 DFFPOSX1_2484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_61__3_), .Q(data_154__3_) );
DFFPOSX1 DFFPOSX1_2485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_61__4_), .Q(data_154__4_) );
DFFPOSX1 DFFPOSX1_2486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_61__5_), .Q(data_154__5_) );
DFFPOSX1 DFFPOSX1_2487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_61__6_), .Q(data_154__6_) );
DFFPOSX1 DFFPOSX1_2488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_61__7_), .Q(data_154__7_) );
DFFPOSX1 DFFPOSX1_2489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_61__8_), .Q(data_154__8_) );
DFFPOSX1 DFFPOSX1_2490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_61__9_), .Q(data_154__9_) );
DFFPOSX1 DFFPOSX1_2491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_61__10_), .Q(data_154__10_) );
DFFPOSX1 DFFPOSX1_2492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_61__11_), .Q(data_154__11_) );
DFFPOSX1 DFFPOSX1_2493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_61__12_), .Q(data_154__12_) );
DFFPOSX1 DFFPOSX1_2494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_61__13_), .Q(data_154__13_) );
DFFPOSX1 DFFPOSX1_2495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_61__14_), .Q(data_154__14_) );
DFFPOSX1 DFFPOSX1_2496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_61__15_), .Q(data_154__15_) );
DFFPOSX1 DFFPOSX1_2497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_62__0_), .Q(data_155__0_) );
DFFPOSX1 DFFPOSX1_2498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_62__1_), .Q(data_155__1_) );
DFFPOSX1 DFFPOSX1_2499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_62__2_), .Q(data_155__2_) );
DFFPOSX1 DFFPOSX1_2500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_62__3_), .Q(data_155__3_) );
DFFPOSX1 DFFPOSX1_2501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_62__4_), .Q(data_155__4_) );
DFFPOSX1 DFFPOSX1_2502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_62__5_), .Q(data_155__5_) );
DFFPOSX1 DFFPOSX1_2503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_62__6_), .Q(data_155__6_) );
DFFPOSX1 DFFPOSX1_2504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_62__7_), .Q(data_155__7_) );
DFFPOSX1 DFFPOSX1_2505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_62__8_), .Q(data_155__8_) );
DFFPOSX1 DFFPOSX1_2506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_62__9_), .Q(data_155__9_) );
DFFPOSX1 DFFPOSX1_2507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_62__10_), .Q(data_155__10_) );
DFFPOSX1 DFFPOSX1_2508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_62__11_), .Q(data_155__11_) );
DFFPOSX1 DFFPOSX1_2509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_62__12_), .Q(data_155__12_) );
DFFPOSX1 DFFPOSX1_2510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_62__13_), .Q(data_155__13_) );
DFFPOSX1 DFFPOSX1_2511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_62__14_), .Q(data_155__14_) );
DFFPOSX1 DFFPOSX1_2512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_62__15_), .Q(data_155__15_) );
DFFPOSX1 DFFPOSX1_2513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_63__0_), .Q(data_156__0_) );
DFFPOSX1 DFFPOSX1_2514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_63__1_), .Q(data_156__1_) );
DFFPOSX1 DFFPOSX1_2515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_63__2_), .Q(data_156__2_) );
DFFPOSX1 DFFPOSX1_2516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_63__3_), .Q(data_156__3_) );
DFFPOSX1 DFFPOSX1_2517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_63__4_), .Q(data_156__4_) );
DFFPOSX1 DFFPOSX1_2518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_63__5_), .Q(data_156__5_) );
DFFPOSX1 DFFPOSX1_2519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_63__6_), .Q(data_156__6_) );
DFFPOSX1 DFFPOSX1_2520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_63__7_), .Q(data_156__7_) );
DFFPOSX1 DFFPOSX1_2521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_63__8_), .Q(data_156__8_) );
DFFPOSX1 DFFPOSX1_2522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_63__9_), .Q(data_156__9_) );
DFFPOSX1 DFFPOSX1_2523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_63__10_), .Q(data_156__10_) );
DFFPOSX1 DFFPOSX1_2524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_63__11_), .Q(data_156__11_) );
DFFPOSX1 DFFPOSX1_2525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_63__12_), .Q(data_156__12_) );
DFFPOSX1 DFFPOSX1_2526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_63__13_), .Q(data_156__13_) );
DFFPOSX1 DFFPOSX1_2527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_63__14_), .Q(data_156__14_) );
DFFPOSX1 DFFPOSX1_2528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_63__15_), .Q(data_156__15_) );
DFFPOSX1 DFFPOSX1_2529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_64__0_), .Q(data_157__0_) );
DFFPOSX1 DFFPOSX1_2530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_64__1_), .Q(data_157__1_) );
DFFPOSX1 DFFPOSX1_2531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_64__2_), .Q(data_157__2_) );
DFFPOSX1 DFFPOSX1_2532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_64__3_), .Q(data_157__3_) );
DFFPOSX1 DFFPOSX1_2533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_64__4_), .Q(data_157__4_) );
DFFPOSX1 DFFPOSX1_2534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_64__5_), .Q(data_157__5_) );
DFFPOSX1 DFFPOSX1_2535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_64__6_), .Q(data_157__6_) );
DFFPOSX1 DFFPOSX1_2536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_64__7_), .Q(data_157__7_) );
DFFPOSX1 DFFPOSX1_2537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_64__8_), .Q(data_157__8_) );
DFFPOSX1 DFFPOSX1_2538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_64__9_), .Q(data_157__9_) );
DFFPOSX1 DFFPOSX1_2539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_64__10_), .Q(data_157__10_) );
DFFPOSX1 DFFPOSX1_2540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_64__11_), .Q(data_157__11_) );
DFFPOSX1 DFFPOSX1_2541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_64__12_), .Q(data_157__12_) );
DFFPOSX1 DFFPOSX1_2542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_64__13_), .Q(data_157__13_) );
DFFPOSX1 DFFPOSX1_2543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_64__14_), .Q(data_157__14_) );
DFFPOSX1 DFFPOSX1_2544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_64__15_), .Q(data_157__15_) );
DFFPOSX1 DFFPOSX1_2545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_65__0_), .Q(data_158__0_) );
DFFPOSX1 DFFPOSX1_2546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_65__1_), .Q(data_158__1_) );
DFFPOSX1 DFFPOSX1_2547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_65__2_), .Q(data_158__2_) );
DFFPOSX1 DFFPOSX1_2548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_65__3_), .Q(data_158__3_) );
DFFPOSX1 DFFPOSX1_2549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_65__4_), .Q(data_158__4_) );
DFFPOSX1 DFFPOSX1_2550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_65__5_), .Q(data_158__5_) );
DFFPOSX1 DFFPOSX1_2551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_65__6_), .Q(data_158__6_) );
DFFPOSX1 DFFPOSX1_2552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_65__7_), .Q(data_158__7_) );
DFFPOSX1 DFFPOSX1_2553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_65__8_), .Q(data_158__8_) );
DFFPOSX1 DFFPOSX1_2554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_65__9_), .Q(data_158__9_) );
DFFPOSX1 DFFPOSX1_2555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_65__10_), .Q(data_158__10_) );
DFFPOSX1 DFFPOSX1_2556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_65__11_), .Q(data_158__11_) );
DFFPOSX1 DFFPOSX1_2557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_65__12_), .Q(data_158__12_) );
DFFPOSX1 DFFPOSX1_2558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_65__13_), .Q(data_158__13_) );
DFFPOSX1 DFFPOSX1_2559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_65__14_), .Q(data_158__14_) );
DFFPOSX1 DFFPOSX1_2560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_65__15_), .Q(data_158__15_) );
DFFPOSX1 DFFPOSX1_2561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf1), .D(_66__0_), .Q(data_159__0_) );
DFFPOSX1 DFFPOSX1_2562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf1), .D(_66__1_), .Q(data_159__1_) );
DFFPOSX1 DFFPOSX1_2563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf1), .D(_66__2_), .Q(data_159__2_) );
DFFPOSX1 DFFPOSX1_2564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf1), .D(_66__3_), .Q(data_159__3_) );
DFFPOSX1 DFFPOSX1_2565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf1), .D(_66__4_), .Q(data_159__4_) );
DFFPOSX1 DFFPOSX1_2566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf1), .D(_66__5_), .Q(data_159__5_) );
DFFPOSX1 DFFPOSX1_2567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf1), .D(_66__6_), .Q(data_159__6_) );
DFFPOSX1 DFFPOSX1_2568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf1), .D(_66__7_), .Q(data_159__7_) );
DFFPOSX1 DFFPOSX1_2569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf1), .D(_66__8_), .Q(data_159__8_) );
DFFPOSX1 DFFPOSX1_2570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf1), .D(_66__9_), .Q(data_159__9_) );
DFFPOSX1 DFFPOSX1_2571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf1), .D(_66__10_), .Q(data_159__10_) );
DFFPOSX1 DFFPOSX1_2572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf1), .D(_66__11_), .Q(data_159__11_) );
DFFPOSX1 DFFPOSX1_2573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf1), .D(_66__12_), .Q(data_159__12_) );
DFFPOSX1 DFFPOSX1_2574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf1), .D(_66__13_), .Q(data_159__13_) );
DFFPOSX1 DFFPOSX1_2575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf1), .D(_66__14_), .Q(data_159__14_) );
DFFPOSX1 DFFPOSX1_2576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf1), .D(_66__15_), .Q(data_159__15_) );
DFFPOSX1 DFFPOSX1_2577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_68__0_), .Q(data_160__0_) );
DFFPOSX1 DFFPOSX1_2578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_68__1_), .Q(data_160__1_) );
DFFPOSX1 DFFPOSX1_2579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_68__2_), .Q(data_160__2_) );
DFFPOSX1 DFFPOSX1_2580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_68__3_), .Q(data_160__3_) );
DFFPOSX1 DFFPOSX1_2581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_68__4_), .Q(data_160__4_) );
DFFPOSX1 DFFPOSX1_2582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_68__5_), .Q(data_160__5_) );
DFFPOSX1 DFFPOSX1_2583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_68__6_), .Q(data_160__6_) );
DFFPOSX1 DFFPOSX1_2584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_68__7_), .Q(data_160__7_) );
DFFPOSX1 DFFPOSX1_2585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_68__8_), .Q(data_160__8_) );
DFFPOSX1 DFFPOSX1_2586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_68__9_), .Q(data_160__9_) );
DFFPOSX1 DFFPOSX1_2587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_68__10_), .Q(data_160__10_) );
DFFPOSX1 DFFPOSX1_2588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_68__11_), .Q(data_160__11_) );
DFFPOSX1 DFFPOSX1_2589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_68__12_), .Q(data_160__12_) );
DFFPOSX1 DFFPOSX1_2590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_68__13_), .Q(data_160__13_) );
DFFPOSX1 DFFPOSX1_2591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_68__14_), .Q(data_160__14_) );
DFFPOSX1 DFFPOSX1_2592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_68__15_), .Q(data_160__15_) );
DFFPOSX1 DFFPOSX1_2593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_69__0_), .Q(data_161__0_) );
DFFPOSX1 DFFPOSX1_2594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_69__1_), .Q(data_161__1_) );
DFFPOSX1 DFFPOSX1_2595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_69__2_), .Q(data_161__2_) );
DFFPOSX1 DFFPOSX1_2596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_69__3_), .Q(data_161__3_) );
DFFPOSX1 DFFPOSX1_2597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_69__4_), .Q(data_161__4_) );
DFFPOSX1 DFFPOSX1_2598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_69__5_), .Q(data_161__5_) );
DFFPOSX1 DFFPOSX1_2599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_69__6_), .Q(data_161__6_) );
DFFPOSX1 DFFPOSX1_2600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_69__7_), .Q(data_161__7_) );
DFFPOSX1 DFFPOSX1_2601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_69__8_), .Q(data_161__8_) );
DFFPOSX1 DFFPOSX1_2602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_69__9_), .Q(data_161__9_) );
DFFPOSX1 DFFPOSX1_2603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_69__10_), .Q(data_161__10_) );
DFFPOSX1 DFFPOSX1_2604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_69__11_), .Q(data_161__11_) );
DFFPOSX1 DFFPOSX1_2605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_69__12_), .Q(data_161__12_) );
DFFPOSX1 DFFPOSX1_2606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_69__13_), .Q(data_161__13_) );
DFFPOSX1 DFFPOSX1_2607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_69__14_), .Q(data_161__14_) );
DFFPOSX1 DFFPOSX1_2608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_69__15_), .Q(data_161__15_) );
DFFPOSX1 DFFPOSX1_2609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_70__0_), .Q(data_162__0_) );
DFFPOSX1 DFFPOSX1_2610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_70__1_), .Q(data_162__1_) );
DFFPOSX1 DFFPOSX1_2611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_70__2_), .Q(data_162__2_) );
DFFPOSX1 DFFPOSX1_2612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_70__3_), .Q(data_162__3_) );
DFFPOSX1 DFFPOSX1_2613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_70__4_), .Q(data_162__4_) );
DFFPOSX1 DFFPOSX1_2614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_70__5_), .Q(data_162__5_) );
DFFPOSX1 DFFPOSX1_2615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_70__6_), .Q(data_162__6_) );
DFFPOSX1 DFFPOSX1_2616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_70__7_), .Q(data_162__7_) );
DFFPOSX1 DFFPOSX1_2617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_70__8_), .Q(data_162__8_) );
DFFPOSX1 DFFPOSX1_2618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_70__9_), .Q(data_162__9_) );
DFFPOSX1 DFFPOSX1_2619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_70__10_), .Q(data_162__10_) );
DFFPOSX1 DFFPOSX1_2620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_70__11_), .Q(data_162__11_) );
DFFPOSX1 DFFPOSX1_2621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_70__12_), .Q(data_162__12_) );
DFFPOSX1 DFFPOSX1_2622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_70__13_), .Q(data_162__13_) );
DFFPOSX1 DFFPOSX1_2623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_70__14_), .Q(data_162__14_) );
DFFPOSX1 DFFPOSX1_2624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_70__15_), .Q(data_162__15_) );
DFFPOSX1 DFFPOSX1_2625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_71__0_), .Q(data_163__0_) );
DFFPOSX1 DFFPOSX1_2626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_71__1_), .Q(data_163__1_) );
DFFPOSX1 DFFPOSX1_2627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_71__2_), .Q(data_163__2_) );
DFFPOSX1 DFFPOSX1_2628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_71__3_), .Q(data_163__3_) );
DFFPOSX1 DFFPOSX1_2629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_71__4_), .Q(data_163__4_) );
DFFPOSX1 DFFPOSX1_2630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_71__5_), .Q(data_163__5_) );
DFFPOSX1 DFFPOSX1_2631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_71__6_), .Q(data_163__6_) );
DFFPOSX1 DFFPOSX1_2632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_71__7_), .Q(data_163__7_) );
DFFPOSX1 DFFPOSX1_2633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_71__8_), .Q(data_163__8_) );
DFFPOSX1 DFFPOSX1_2634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_71__9_), .Q(data_163__9_) );
DFFPOSX1 DFFPOSX1_2635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_71__10_), .Q(data_163__10_) );
DFFPOSX1 DFFPOSX1_2636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_71__11_), .Q(data_163__11_) );
DFFPOSX1 DFFPOSX1_2637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_71__12_), .Q(data_163__12_) );
DFFPOSX1 DFFPOSX1_2638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_71__13_), .Q(data_163__13_) );
DFFPOSX1 DFFPOSX1_2639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_71__14_), .Q(data_163__14_) );
DFFPOSX1 DFFPOSX1_2640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_71__15_), .Q(data_163__15_) );
DFFPOSX1 DFFPOSX1_2641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_72__0_), .Q(data_164__0_) );
DFFPOSX1 DFFPOSX1_2642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_72__1_), .Q(data_164__1_) );
DFFPOSX1 DFFPOSX1_2643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_72__2_), .Q(data_164__2_) );
DFFPOSX1 DFFPOSX1_2644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_72__3_), .Q(data_164__3_) );
DFFPOSX1 DFFPOSX1_2645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_72__4_), .Q(data_164__4_) );
DFFPOSX1 DFFPOSX1_2646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_72__5_), .Q(data_164__5_) );
DFFPOSX1 DFFPOSX1_2647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_72__6_), .Q(data_164__6_) );
DFFPOSX1 DFFPOSX1_2648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_72__7_), .Q(data_164__7_) );
DFFPOSX1 DFFPOSX1_2649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_72__8_), .Q(data_164__8_) );
DFFPOSX1 DFFPOSX1_2650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_72__9_), .Q(data_164__9_) );
DFFPOSX1 DFFPOSX1_2651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_72__10_), .Q(data_164__10_) );
DFFPOSX1 DFFPOSX1_2652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_72__11_), .Q(data_164__11_) );
DFFPOSX1 DFFPOSX1_2653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_72__12_), .Q(data_164__12_) );
DFFPOSX1 DFFPOSX1_2654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_72__13_), .Q(data_164__13_) );
DFFPOSX1 DFFPOSX1_2655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_72__14_), .Q(data_164__14_) );
DFFPOSX1 DFFPOSX1_2656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_72__15_), .Q(data_164__15_) );
DFFPOSX1 DFFPOSX1_2657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_73__0_), .Q(data_165__0_) );
DFFPOSX1 DFFPOSX1_2658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_73__1_), .Q(data_165__1_) );
DFFPOSX1 DFFPOSX1_2659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_73__2_), .Q(data_165__2_) );
DFFPOSX1 DFFPOSX1_2660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_73__3_), .Q(data_165__3_) );
DFFPOSX1 DFFPOSX1_2661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_73__4_), .Q(data_165__4_) );
DFFPOSX1 DFFPOSX1_2662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_73__5_), .Q(data_165__5_) );
DFFPOSX1 DFFPOSX1_2663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_73__6_), .Q(data_165__6_) );
DFFPOSX1 DFFPOSX1_2664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_73__7_), .Q(data_165__7_) );
DFFPOSX1 DFFPOSX1_2665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_73__8_), .Q(data_165__8_) );
DFFPOSX1 DFFPOSX1_2666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_73__9_), .Q(data_165__9_) );
DFFPOSX1 DFFPOSX1_2667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_73__10_), .Q(data_165__10_) );
DFFPOSX1 DFFPOSX1_2668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_73__11_), .Q(data_165__11_) );
DFFPOSX1 DFFPOSX1_2669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_73__12_), .Q(data_165__12_) );
DFFPOSX1 DFFPOSX1_2670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_73__13_), .Q(data_165__13_) );
DFFPOSX1 DFFPOSX1_2671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_73__14_), .Q(data_165__14_) );
DFFPOSX1 DFFPOSX1_2672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_73__15_), .Q(data_165__15_) );
DFFPOSX1 DFFPOSX1_2673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_74__0_), .Q(data_166__0_) );
DFFPOSX1 DFFPOSX1_2674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_74__1_), .Q(data_166__1_) );
DFFPOSX1 DFFPOSX1_2675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_74__2_), .Q(data_166__2_) );
DFFPOSX1 DFFPOSX1_2676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_74__3_), .Q(data_166__3_) );
DFFPOSX1 DFFPOSX1_2677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_74__4_), .Q(data_166__4_) );
DFFPOSX1 DFFPOSX1_2678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_74__5_), .Q(data_166__5_) );
DFFPOSX1 DFFPOSX1_2679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_74__6_), .Q(data_166__6_) );
DFFPOSX1 DFFPOSX1_2680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_74__7_), .Q(data_166__7_) );
DFFPOSX1 DFFPOSX1_2681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_74__8_), .Q(data_166__8_) );
DFFPOSX1 DFFPOSX1_2682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_74__9_), .Q(data_166__9_) );
DFFPOSX1 DFFPOSX1_2683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_74__10_), .Q(data_166__10_) );
DFFPOSX1 DFFPOSX1_2684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_74__11_), .Q(data_166__11_) );
DFFPOSX1 DFFPOSX1_2685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_74__12_), .Q(data_166__12_) );
DFFPOSX1 DFFPOSX1_2686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_74__13_), .Q(data_166__13_) );
DFFPOSX1 DFFPOSX1_2687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_74__14_), .Q(data_166__14_) );
DFFPOSX1 DFFPOSX1_2688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_74__15_), .Q(data_166__15_) );
DFFPOSX1 DFFPOSX1_2689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_75__0_), .Q(data_167__0_) );
DFFPOSX1 DFFPOSX1_2690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_75__1_), .Q(data_167__1_) );
DFFPOSX1 DFFPOSX1_2691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_75__2_), .Q(data_167__2_) );
DFFPOSX1 DFFPOSX1_2692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_75__3_), .Q(data_167__3_) );
DFFPOSX1 DFFPOSX1_2693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_75__4_), .Q(data_167__4_) );
DFFPOSX1 DFFPOSX1_2694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_75__5_), .Q(data_167__5_) );
DFFPOSX1 DFFPOSX1_2695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_75__6_), .Q(data_167__6_) );
DFFPOSX1 DFFPOSX1_2696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_75__7_), .Q(data_167__7_) );
DFFPOSX1 DFFPOSX1_2697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_75__8_), .Q(data_167__8_) );
DFFPOSX1 DFFPOSX1_2698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_75__9_), .Q(data_167__9_) );
DFFPOSX1 DFFPOSX1_2699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_75__10_), .Q(data_167__10_) );
DFFPOSX1 DFFPOSX1_2700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_75__11_), .Q(data_167__11_) );
DFFPOSX1 DFFPOSX1_2701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_75__12_), .Q(data_167__12_) );
DFFPOSX1 DFFPOSX1_2702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_75__13_), .Q(data_167__13_) );
DFFPOSX1 DFFPOSX1_2703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_75__14_), .Q(data_167__14_) );
DFFPOSX1 DFFPOSX1_2704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_75__15_), .Q(data_167__15_) );
DFFPOSX1 DFFPOSX1_2705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_76__0_), .Q(data_168__0_) );
DFFPOSX1 DFFPOSX1_2706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_76__1_), .Q(data_168__1_) );
DFFPOSX1 DFFPOSX1_2707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_76__2_), .Q(data_168__2_) );
DFFPOSX1 DFFPOSX1_2708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_76__3_), .Q(data_168__3_) );
DFFPOSX1 DFFPOSX1_2709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_76__4_), .Q(data_168__4_) );
DFFPOSX1 DFFPOSX1_2710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_76__5_), .Q(data_168__5_) );
DFFPOSX1 DFFPOSX1_2711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_76__6_), .Q(data_168__6_) );
DFFPOSX1 DFFPOSX1_2712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_76__7_), .Q(data_168__7_) );
DFFPOSX1 DFFPOSX1_2713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_76__8_), .Q(data_168__8_) );
DFFPOSX1 DFFPOSX1_2714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_76__9_), .Q(data_168__9_) );
DFFPOSX1 DFFPOSX1_2715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_76__10_), .Q(data_168__10_) );
DFFPOSX1 DFFPOSX1_2716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_76__11_), .Q(data_168__11_) );
DFFPOSX1 DFFPOSX1_2717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_76__12_), .Q(data_168__12_) );
DFFPOSX1 DFFPOSX1_2718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_76__13_), .Q(data_168__13_) );
DFFPOSX1 DFFPOSX1_2719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_76__14_), .Q(data_168__14_) );
DFFPOSX1 DFFPOSX1_2720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_76__15_), .Q(data_168__15_) );
DFFPOSX1 DFFPOSX1_2721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_77__0_), .Q(data_169__0_) );
DFFPOSX1 DFFPOSX1_2722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_77__1_), .Q(data_169__1_) );
DFFPOSX1 DFFPOSX1_2723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_77__2_), .Q(data_169__2_) );
DFFPOSX1 DFFPOSX1_2724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_77__3_), .Q(data_169__3_) );
DFFPOSX1 DFFPOSX1_2725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_77__4_), .Q(data_169__4_) );
DFFPOSX1 DFFPOSX1_2726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_77__5_), .Q(data_169__5_) );
DFFPOSX1 DFFPOSX1_2727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_77__6_), .Q(data_169__6_) );
DFFPOSX1 DFFPOSX1_2728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_77__7_), .Q(data_169__7_) );
DFFPOSX1 DFFPOSX1_2729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_77__8_), .Q(data_169__8_) );
DFFPOSX1 DFFPOSX1_2730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_77__9_), .Q(data_169__9_) );
DFFPOSX1 DFFPOSX1_2731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_77__10_), .Q(data_169__10_) );
DFFPOSX1 DFFPOSX1_2732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_77__11_), .Q(data_169__11_) );
DFFPOSX1 DFFPOSX1_2733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_77__12_), .Q(data_169__12_) );
DFFPOSX1 DFFPOSX1_2734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_77__13_), .Q(data_169__13_) );
DFFPOSX1 DFFPOSX1_2735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_77__14_), .Q(data_169__14_) );
DFFPOSX1 DFFPOSX1_2736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_77__15_), .Q(data_169__15_) );
DFFPOSX1 DFFPOSX1_2737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_79__0_), .Q(data_170__0_) );
DFFPOSX1 DFFPOSX1_2738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_79__1_), .Q(data_170__1_) );
DFFPOSX1 DFFPOSX1_2739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_79__2_), .Q(data_170__2_) );
DFFPOSX1 DFFPOSX1_2740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_79__3_), .Q(data_170__3_) );
DFFPOSX1 DFFPOSX1_2741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_79__4_), .Q(data_170__4_) );
DFFPOSX1 DFFPOSX1_2742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_79__5_), .Q(data_170__5_) );
DFFPOSX1 DFFPOSX1_2743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_79__6_), .Q(data_170__6_) );
DFFPOSX1 DFFPOSX1_2744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_79__7_), .Q(data_170__7_) );
DFFPOSX1 DFFPOSX1_2745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_79__8_), .Q(data_170__8_) );
DFFPOSX1 DFFPOSX1_2746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_79__9_), .Q(data_170__9_) );
DFFPOSX1 DFFPOSX1_2747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_79__10_), .Q(data_170__10_) );
DFFPOSX1 DFFPOSX1_2748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_79__11_), .Q(data_170__11_) );
DFFPOSX1 DFFPOSX1_2749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_79__12_), .Q(data_170__12_) );
DFFPOSX1 DFFPOSX1_2750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_79__13_), .Q(data_170__13_) );
DFFPOSX1 DFFPOSX1_2751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_79__14_), .Q(data_170__14_) );
DFFPOSX1 DFFPOSX1_2752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_79__15_), .Q(data_170__15_) );
DFFPOSX1 DFFPOSX1_2753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_80__0_), .Q(data_171__0_) );
DFFPOSX1 DFFPOSX1_2754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_80__1_), .Q(data_171__1_) );
DFFPOSX1 DFFPOSX1_2755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_80__2_), .Q(data_171__2_) );
DFFPOSX1 DFFPOSX1_2756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_80__3_), .Q(data_171__3_) );
DFFPOSX1 DFFPOSX1_2757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_80__4_), .Q(data_171__4_) );
DFFPOSX1 DFFPOSX1_2758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_80__5_), .Q(data_171__5_) );
DFFPOSX1 DFFPOSX1_2759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_80__6_), .Q(data_171__6_) );
DFFPOSX1 DFFPOSX1_2760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_80__7_), .Q(data_171__7_) );
DFFPOSX1 DFFPOSX1_2761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_80__8_), .Q(data_171__8_) );
DFFPOSX1 DFFPOSX1_2762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_80__9_), .Q(data_171__9_) );
DFFPOSX1 DFFPOSX1_2763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_80__10_), .Q(data_171__10_) );
DFFPOSX1 DFFPOSX1_2764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_80__11_), .Q(data_171__11_) );
DFFPOSX1 DFFPOSX1_2765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_80__12_), .Q(data_171__12_) );
DFFPOSX1 DFFPOSX1_2766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_80__13_), .Q(data_171__13_) );
DFFPOSX1 DFFPOSX1_2767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_80__14_), .Q(data_171__14_) );
DFFPOSX1 DFFPOSX1_2768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_80__15_), .Q(data_171__15_) );
DFFPOSX1 DFFPOSX1_2769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_81__0_), .Q(data_172__0_) );
DFFPOSX1 DFFPOSX1_2770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_81__1_), .Q(data_172__1_) );
DFFPOSX1 DFFPOSX1_2771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_81__2_), .Q(data_172__2_) );
DFFPOSX1 DFFPOSX1_2772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_81__3_), .Q(data_172__3_) );
DFFPOSX1 DFFPOSX1_2773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_81__4_), .Q(data_172__4_) );
DFFPOSX1 DFFPOSX1_2774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_81__5_), .Q(data_172__5_) );
DFFPOSX1 DFFPOSX1_2775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_81__6_), .Q(data_172__6_) );
DFFPOSX1 DFFPOSX1_2776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_81__7_), .Q(data_172__7_) );
DFFPOSX1 DFFPOSX1_2777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_81__8_), .Q(data_172__8_) );
DFFPOSX1 DFFPOSX1_2778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_81__9_), .Q(data_172__9_) );
DFFPOSX1 DFFPOSX1_2779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_81__10_), .Q(data_172__10_) );
DFFPOSX1 DFFPOSX1_2780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_81__11_), .Q(data_172__11_) );
DFFPOSX1 DFFPOSX1_2781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_81__12_), .Q(data_172__12_) );
DFFPOSX1 DFFPOSX1_2782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_81__13_), .Q(data_172__13_) );
DFFPOSX1 DFFPOSX1_2783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_81__14_), .Q(data_172__14_) );
DFFPOSX1 DFFPOSX1_2784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_81__15_), .Q(data_172__15_) );
DFFPOSX1 DFFPOSX1_2785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_82__0_), .Q(data_173__0_) );
DFFPOSX1 DFFPOSX1_2786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_82__1_), .Q(data_173__1_) );
DFFPOSX1 DFFPOSX1_2787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_82__2_), .Q(data_173__2_) );
DFFPOSX1 DFFPOSX1_2788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_82__3_), .Q(data_173__3_) );
DFFPOSX1 DFFPOSX1_2789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_82__4_), .Q(data_173__4_) );
DFFPOSX1 DFFPOSX1_2790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_82__5_), .Q(data_173__5_) );
DFFPOSX1 DFFPOSX1_2791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_82__6_), .Q(data_173__6_) );
DFFPOSX1 DFFPOSX1_2792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_82__7_), .Q(data_173__7_) );
DFFPOSX1 DFFPOSX1_2793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_82__8_), .Q(data_173__8_) );
DFFPOSX1 DFFPOSX1_2794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_82__9_), .Q(data_173__9_) );
DFFPOSX1 DFFPOSX1_2795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_82__10_), .Q(data_173__10_) );
DFFPOSX1 DFFPOSX1_2796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_82__11_), .Q(data_173__11_) );
DFFPOSX1 DFFPOSX1_2797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_82__12_), .Q(data_173__12_) );
DFFPOSX1 DFFPOSX1_2798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_82__13_), .Q(data_173__13_) );
DFFPOSX1 DFFPOSX1_2799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_82__14_), .Q(data_173__14_) );
DFFPOSX1 DFFPOSX1_2800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_82__15_), .Q(data_173__15_) );
DFFPOSX1 DFFPOSX1_2801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_83__0_), .Q(data_174__0_) );
DFFPOSX1 DFFPOSX1_2802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_83__1_), .Q(data_174__1_) );
DFFPOSX1 DFFPOSX1_2803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_83__2_), .Q(data_174__2_) );
DFFPOSX1 DFFPOSX1_2804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_83__3_), .Q(data_174__3_) );
DFFPOSX1 DFFPOSX1_2805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_83__4_), .Q(data_174__4_) );
DFFPOSX1 DFFPOSX1_2806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_83__5_), .Q(data_174__5_) );
DFFPOSX1 DFFPOSX1_2807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_83__6_), .Q(data_174__6_) );
DFFPOSX1 DFFPOSX1_2808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_83__7_), .Q(data_174__7_) );
DFFPOSX1 DFFPOSX1_2809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_83__8_), .Q(data_174__8_) );
DFFPOSX1 DFFPOSX1_2810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_83__9_), .Q(data_174__9_) );
DFFPOSX1 DFFPOSX1_2811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_83__10_), .Q(data_174__10_) );
DFFPOSX1 DFFPOSX1_2812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_83__11_), .Q(data_174__11_) );
DFFPOSX1 DFFPOSX1_2813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_83__12_), .Q(data_174__12_) );
DFFPOSX1 DFFPOSX1_2814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_83__13_), .Q(data_174__13_) );
DFFPOSX1 DFFPOSX1_2815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_83__14_), .Q(data_174__14_) );
DFFPOSX1 DFFPOSX1_2816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_83__15_), .Q(data_174__15_) );
DFFPOSX1 DFFPOSX1_2817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf0), .D(_84__0_), .Q(data_175__0_) );
DFFPOSX1 DFFPOSX1_2818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf0), .D(_84__1_), .Q(data_175__1_) );
DFFPOSX1 DFFPOSX1_2819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf0), .D(_84__2_), .Q(data_175__2_) );
DFFPOSX1 DFFPOSX1_2820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf0), .D(_84__3_), .Q(data_175__3_) );
DFFPOSX1 DFFPOSX1_2821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf0), .D(_84__4_), .Q(data_175__4_) );
DFFPOSX1 DFFPOSX1_2822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf0), .D(_84__5_), .Q(data_175__5_) );
DFFPOSX1 DFFPOSX1_2823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf0), .D(_84__6_), .Q(data_175__6_) );
DFFPOSX1 DFFPOSX1_2824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf0), .D(_84__7_), .Q(data_175__7_) );
DFFPOSX1 DFFPOSX1_2825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf0), .D(_84__8_), .Q(data_175__8_) );
DFFPOSX1 DFFPOSX1_2826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf0), .D(_84__9_), .Q(data_175__9_) );
DFFPOSX1 DFFPOSX1_2827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf0), .D(_84__10_), .Q(data_175__10_) );
DFFPOSX1 DFFPOSX1_2828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf0), .D(_84__11_), .Q(data_175__11_) );
DFFPOSX1 DFFPOSX1_2829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf0), .D(_84__12_), .Q(data_175__12_) );
DFFPOSX1 DFFPOSX1_2830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf0), .D(_84__13_), .Q(data_175__13_) );
DFFPOSX1 DFFPOSX1_2831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf0), .D(_84__14_), .Q(data_175__14_) );
DFFPOSX1 DFFPOSX1_2832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf0), .D(_84__15_), .Q(data_175__15_) );
DFFPOSX1 DFFPOSX1_2833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_85__0_), .Q(data_176__0_) );
DFFPOSX1 DFFPOSX1_2834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_85__1_), .Q(data_176__1_) );
DFFPOSX1 DFFPOSX1_2835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_85__2_), .Q(data_176__2_) );
DFFPOSX1 DFFPOSX1_2836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_85__3_), .Q(data_176__3_) );
DFFPOSX1 DFFPOSX1_2837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_85__4_), .Q(data_176__4_) );
DFFPOSX1 DFFPOSX1_2838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_85__5_), .Q(data_176__5_) );
DFFPOSX1 DFFPOSX1_2839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_85__6_), .Q(data_176__6_) );
DFFPOSX1 DFFPOSX1_2840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_85__7_), .Q(data_176__7_) );
DFFPOSX1 DFFPOSX1_2841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_85__8_), .Q(data_176__8_) );
DFFPOSX1 DFFPOSX1_2842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_85__9_), .Q(data_176__9_) );
DFFPOSX1 DFFPOSX1_2843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_85__10_), .Q(data_176__10_) );
DFFPOSX1 DFFPOSX1_2844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_85__11_), .Q(data_176__11_) );
DFFPOSX1 DFFPOSX1_2845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_85__12_), .Q(data_176__12_) );
DFFPOSX1 DFFPOSX1_2846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_85__13_), .Q(data_176__13_) );
DFFPOSX1 DFFPOSX1_2847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_85__14_), .Q(data_176__14_) );
DFFPOSX1 DFFPOSX1_2848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_85__15_), .Q(data_176__15_) );
DFFPOSX1 DFFPOSX1_2849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_86__0_), .Q(data_177__0_) );
DFFPOSX1 DFFPOSX1_2850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_86__1_), .Q(data_177__1_) );
DFFPOSX1 DFFPOSX1_2851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_86__2_), .Q(data_177__2_) );
DFFPOSX1 DFFPOSX1_2852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_86__3_), .Q(data_177__3_) );
DFFPOSX1 DFFPOSX1_2853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_86__4_), .Q(data_177__4_) );
DFFPOSX1 DFFPOSX1_2854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_86__5_), .Q(data_177__5_) );
DFFPOSX1 DFFPOSX1_2855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_86__6_), .Q(data_177__6_) );
DFFPOSX1 DFFPOSX1_2856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_86__7_), .Q(data_177__7_) );
DFFPOSX1 DFFPOSX1_2857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_86__8_), .Q(data_177__8_) );
DFFPOSX1 DFFPOSX1_2858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_86__9_), .Q(data_177__9_) );
DFFPOSX1 DFFPOSX1_2859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_86__10_), .Q(data_177__10_) );
DFFPOSX1 DFFPOSX1_2860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_86__11_), .Q(data_177__11_) );
DFFPOSX1 DFFPOSX1_2861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_86__12_), .Q(data_177__12_) );
DFFPOSX1 DFFPOSX1_2862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_86__13_), .Q(data_177__13_) );
DFFPOSX1 DFFPOSX1_2863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_86__14_), .Q(data_177__14_) );
DFFPOSX1 DFFPOSX1_2864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_86__15_), .Q(data_177__15_) );
DFFPOSX1 DFFPOSX1_2865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_87__0_), .Q(data_178__0_) );
DFFPOSX1 DFFPOSX1_2866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_87__1_), .Q(data_178__1_) );
DFFPOSX1 DFFPOSX1_2867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_87__2_), .Q(data_178__2_) );
DFFPOSX1 DFFPOSX1_2868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_87__3_), .Q(data_178__3_) );
DFFPOSX1 DFFPOSX1_2869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_87__4_), .Q(data_178__4_) );
DFFPOSX1 DFFPOSX1_2870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_87__5_), .Q(data_178__5_) );
DFFPOSX1 DFFPOSX1_2871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_87__6_), .Q(data_178__6_) );
DFFPOSX1 DFFPOSX1_2872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_87__7_), .Q(data_178__7_) );
DFFPOSX1 DFFPOSX1_2873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_87__8_), .Q(data_178__8_) );
DFFPOSX1 DFFPOSX1_2874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_87__9_), .Q(data_178__9_) );
DFFPOSX1 DFFPOSX1_2875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_87__10_), .Q(data_178__10_) );
DFFPOSX1 DFFPOSX1_2876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_87__11_), .Q(data_178__11_) );
DFFPOSX1 DFFPOSX1_2877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_87__12_), .Q(data_178__12_) );
DFFPOSX1 DFFPOSX1_2878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_87__13_), .Q(data_178__13_) );
DFFPOSX1 DFFPOSX1_2879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_87__14_), .Q(data_178__14_) );
DFFPOSX1 DFFPOSX1_2880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_87__15_), .Q(data_178__15_) );
DFFPOSX1 DFFPOSX1_2881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_88__0_), .Q(data_179__0_) );
DFFPOSX1 DFFPOSX1_2882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_88__1_), .Q(data_179__1_) );
DFFPOSX1 DFFPOSX1_2883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_88__2_), .Q(data_179__2_) );
DFFPOSX1 DFFPOSX1_2884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_88__3_), .Q(data_179__3_) );
DFFPOSX1 DFFPOSX1_2885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_88__4_), .Q(data_179__4_) );
DFFPOSX1 DFFPOSX1_2886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_88__5_), .Q(data_179__5_) );
DFFPOSX1 DFFPOSX1_2887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_88__6_), .Q(data_179__6_) );
DFFPOSX1 DFFPOSX1_2888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_88__7_), .Q(data_179__7_) );
DFFPOSX1 DFFPOSX1_2889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_88__8_), .Q(data_179__8_) );
DFFPOSX1 DFFPOSX1_2890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_88__9_), .Q(data_179__9_) );
DFFPOSX1 DFFPOSX1_2891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_88__10_), .Q(data_179__10_) );
DFFPOSX1 DFFPOSX1_2892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_88__11_), .Q(data_179__11_) );
DFFPOSX1 DFFPOSX1_2893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_88__12_), .Q(data_179__12_) );
DFFPOSX1 DFFPOSX1_2894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_88__13_), .Q(data_179__13_) );
DFFPOSX1 DFFPOSX1_2895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_88__14_), .Q(data_179__14_) );
DFFPOSX1 DFFPOSX1_2896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_88__15_), .Q(data_179__15_) );
DFFPOSX1 DFFPOSX1_2897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_90__0_), .Q(data_180__0_) );
DFFPOSX1 DFFPOSX1_2898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_90__1_), .Q(data_180__1_) );
DFFPOSX1 DFFPOSX1_2899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_90__2_), .Q(data_180__2_) );
DFFPOSX1 DFFPOSX1_2900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_90__3_), .Q(data_180__3_) );
DFFPOSX1 DFFPOSX1_2901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_90__4_), .Q(data_180__4_) );
DFFPOSX1 DFFPOSX1_2902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_90__5_), .Q(data_180__5_) );
DFFPOSX1 DFFPOSX1_2903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_90__6_), .Q(data_180__6_) );
DFFPOSX1 DFFPOSX1_2904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_90__7_), .Q(data_180__7_) );
DFFPOSX1 DFFPOSX1_2905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_90__8_), .Q(data_180__8_) );
DFFPOSX1 DFFPOSX1_2906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_90__9_), .Q(data_180__9_) );
DFFPOSX1 DFFPOSX1_2907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_90__10_), .Q(data_180__10_) );
DFFPOSX1 DFFPOSX1_2908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_90__11_), .Q(data_180__11_) );
DFFPOSX1 DFFPOSX1_2909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_90__12_), .Q(data_180__12_) );
DFFPOSX1 DFFPOSX1_2910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_90__13_), .Q(data_180__13_) );
DFFPOSX1 DFFPOSX1_2911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_90__14_), .Q(data_180__14_) );
DFFPOSX1 DFFPOSX1_2912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_90__15_), .Q(data_180__15_) );
DFFPOSX1 DFFPOSX1_2913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_91__0_), .Q(data_181__0_) );
DFFPOSX1 DFFPOSX1_2914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_91__1_), .Q(data_181__1_) );
DFFPOSX1 DFFPOSX1_2915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_91__2_), .Q(data_181__2_) );
DFFPOSX1 DFFPOSX1_2916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_91__3_), .Q(data_181__3_) );
DFFPOSX1 DFFPOSX1_2917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_91__4_), .Q(data_181__4_) );
DFFPOSX1 DFFPOSX1_2918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_91__5_), .Q(data_181__5_) );
DFFPOSX1 DFFPOSX1_2919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_91__6_), .Q(data_181__6_) );
DFFPOSX1 DFFPOSX1_2920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_91__7_), .Q(data_181__7_) );
DFFPOSX1 DFFPOSX1_2921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_91__8_), .Q(data_181__8_) );
DFFPOSX1 DFFPOSX1_2922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_91__9_), .Q(data_181__9_) );
DFFPOSX1 DFFPOSX1_2923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_91__10_), .Q(data_181__10_) );
DFFPOSX1 DFFPOSX1_2924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_91__11_), .Q(data_181__11_) );
DFFPOSX1 DFFPOSX1_2925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_91__12_), .Q(data_181__12_) );
DFFPOSX1 DFFPOSX1_2926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_91__13_), .Q(data_181__13_) );
DFFPOSX1 DFFPOSX1_2927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_91__14_), .Q(data_181__14_) );
DFFPOSX1 DFFPOSX1_2928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_91__15_), .Q(data_181__15_) );
DFFPOSX1 DFFPOSX1_2929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_92__0_), .Q(data_182__0_) );
DFFPOSX1 DFFPOSX1_2930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_92__1_), .Q(data_182__1_) );
DFFPOSX1 DFFPOSX1_2931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_92__2_), .Q(data_182__2_) );
DFFPOSX1 DFFPOSX1_2932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_92__3_), .Q(data_182__3_) );
DFFPOSX1 DFFPOSX1_2933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_92__4_), .Q(data_182__4_) );
DFFPOSX1 DFFPOSX1_2934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_92__5_), .Q(data_182__5_) );
DFFPOSX1 DFFPOSX1_2935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_92__6_), .Q(data_182__6_) );
DFFPOSX1 DFFPOSX1_2936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_92__7_), .Q(data_182__7_) );
DFFPOSX1 DFFPOSX1_2937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_92__8_), .Q(data_182__8_) );
DFFPOSX1 DFFPOSX1_2938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_92__9_), .Q(data_182__9_) );
DFFPOSX1 DFFPOSX1_2939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_92__10_), .Q(data_182__10_) );
DFFPOSX1 DFFPOSX1_2940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_92__11_), .Q(data_182__11_) );
DFFPOSX1 DFFPOSX1_2941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_92__12_), .Q(data_182__12_) );
DFFPOSX1 DFFPOSX1_2942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_92__13_), .Q(data_182__13_) );
DFFPOSX1 DFFPOSX1_2943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_92__14_), .Q(data_182__14_) );
DFFPOSX1 DFFPOSX1_2944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_92__15_), .Q(data_182__15_) );
DFFPOSX1 DFFPOSX1_2945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_93__0_), .Q(data_183__0_) );
DFFPOSX1 DFFPOSX1_2946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_93__1_), .Q(data_183__1_) );
DFFPOSX1 DFFPOSX1_2947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_93__2_), .Q(data_183__2_) );
DFFPOSX1 DFFPOSX1_2948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_93__3_), .Q(data_183__3_) );
DFFPOSX1 DFFPOSX1_2949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_93__4_), .Q(data_183__4_) );
DFFPOSX1 DFFPOSX1_2950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_93__5_), .Q(data_183__5_) );
DFFPOSX1 DFFPOSX1_2951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_93__6_), .Q(data_183__6_) );
DFFPOSX1 DFFPOSX1_2952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_93__7_), .Q(data_183__7_) );
DFFPOSX1 DFFPOSX1_2953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_93__8_), .Q(data_183__8_) );
DFFPOSX1 DFFPOSX1_2954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_93__9_), .Q(data_183__9_) );
DFFPOSX1 DFFPOSX1_2955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_93__10_), .Q(data_183__10_) );
DFFPOSX1 DFFPOSX1_2956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_93__11_), .Q(data_183__11_) );
DFFPOSX1 DFFPOSX1_2957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_93__12_), .Q(data_183__12_) );
DFFPOSX1 DFFPOSX1_2958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_93__13_), .Q(data_183__13_) );
DFFPOSX1 DFFPOSX1_2959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_93__14_), .Q(data_183__14_) );
DFFPOSX1 DFFPOSX1_2960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_93__15_), .Q(data_183__15_) );
DFFPOSX1 DFFPOSX1_2961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_94__0_), .Q(data_184__0_) );
DFFPOSX1 DFFPOSX1_2962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_94__1_), .Q(data_184__1_) );
DFFPOSX1 DFFPOSX1_2963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_94__2_), .Q(data_184__2_) );
DFFPOSX1 DFFPOSX1_2964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_94__3_), .Q(data_184__3_) );
DFFPOSX1 DFFPOSX1_2965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_94__4_), .Q(data_184__4_) );
DFFPOSX1 DFFPOSX1_2966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_94__5_), .Q(data_184__5_) );
DFFPOSX1 DFFPOSX1_2967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_94__6_), .Q(data_184__6_) );
DFFPOSX1 DFFPOSX1_2968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_94__7_), .Q(data_184__7_) );
DFFPOSX1 DFFPOSX1_2969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_94__8_), .Q(data_184__8_) );
DFFPOSX1 DFFPOSX1_2970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_94__9_), .Q(data_184__9_) );
DFFPOSX1 DFFPOSX1_2971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_94__10_), .Q(data_184__10_) );
DFFPOSX1 DFFPOSX1_2972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_94__11_), .Q(data_184__11_) );
DFFPOSX1 DFFPOSX1_2973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_94__12_), .Q(data_184__12_) );
DFFPOSX1 DFFPOSX1_2974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_94__13_), .Q(data_184__13_) );
DFFPOSX1 DFFPOSX1_2975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_94__14_), .Q(data_184__14_) );
DFFPOSX1 DFFPOSX1_2976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_94__15_), .Q(data_184__15_) );
DFFPOSX1 DFFPOSX1_2977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_95__0_), .Q(data_185__0_) );
DFFPOSX1 DFFPOSX1_2978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_95__1_), .Q(data_185__1_) );
DFFPOSX1 DFFPOSX1_2979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_95__2_), .Q(data_185__2_) );
DFFPOSX1 DFFPOSX1_2980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_95__3_), .Q(data_185__3_) );
DFFPOSX1 DFFPOSX1_2981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_95__4_), .Q(data_185__4_) );
DFFPOSX1 DFFPOSX1_2982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_95__5_), .Q(data_185__5_) );
DFFPOSX1 DFFPOSX1_2983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_95__6_), .Q(data_185__6_) );
DFFPOSX1 DFFPOSX1_2984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_95__7_), .Q(data_185__7_) );
DFFPOSX1 DFFPOSX1_2985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_95__8_), .Q(data_185__8_) );
DFFPOSX1 DFFPOSX1_2986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_95__9_), .Q(data_185__9_) );
DFFPOSX1 DFFPOSX1_2987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_95__10_), .Q(data_185__10_) );
DFFPOSX1 DFFPOSX1_2988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_95__11_), .Q(data_185__11_) );
DFFPOSX1 DFFPOSX1_2989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_95__12_), .Q(data_185__12_) );
DFFPOSX1 DFFPOSX1_2990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_95__13_), .Q(data_185__13_) );
DFFPOSX1 DFFPOSX1_2991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_95__14_), .Q(data_185__14_) );
DFFPOSX1 DFFPOSX1_2992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_95__15_), .Q(data_185__15_) );
DFFPOSX1 DFFPOSX1_2993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_96__0_), .Q(data_186__0_) );
DFFPOSX1 DFFPOSX1_2994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_96__1_), .Q(data_186__1_) );
DFFPOSX1 DFFPOSX1_2995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_96__2_), .Q(data_186__2_) );
DFFPOSX1 DFFPOSX1_2996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_96__3_), .Q(data_186__3_) );
DFFPOSX1 DFFPOSX1_2997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_96__4_), .Q(data_186__4_) );
DFFPOSX1 DFFPOSX1_2998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_96__5_), .Q(data_186__5_) );
DFFPOSX1 DFFPOSX1_2999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_96__6_), .Q(data_186__6_) );
DFFPOSX1 DFFPOSX1_3000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_96__7_), .Q(data_186__7_) );
DFFPOSX1 DFFPOSX1_3001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_96__8_), .Q(data_186__8_) );
DFFPOSX1 DFFPOSX1_3002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_96__9_), .Q(data_186__9_) );
DFFPOSX1 DFFPOSX1_3003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_96__10_), .Q(data_186__10_) );
DFFPOSX1 DFFPOSX1_3004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_96__11_), .Q(data_186__11_) );
DFFPOSX1 DFFPOSX1_3005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_96__12_), .Q(data_186__12_) );
DFFPOSX1 DFFPOSX1_3006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_96__13_), .Q(data_186__13_) );
DFFPOSX1 DFFPOSX1_3007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_96__14_), .Q(data_186__14_) );
DFFPOSX1 DFFPOSX1_3008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_96__15_), .Q(data_186__15_) );
DFFPOSX1 DFFPOSX1_3009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_97__0_), .Q(data_187__0_) );
DFFPOSX1 DFFPOSX1_3010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_97__1_), .Q(data_187__1_) );
DFFPOSX1 DFFPOSX1_3011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_97__2_), .Q(data_187__2_) );
DFFPOSX1 DFFPOSX1_3012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_97__3_), .Q(data_187__3_) );
DFFPOSX1 DFFPOSX1_3013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_97__4_), .Q(data_187__4_) );
DFFPOSX1 DFFPOSX1_3014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_97__5_), .Q(data_187__5_) );
DFFPOSX1 DFFPOSX1_3015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_97__6_), .Q(data_187__6_) );
DFFPOSX1 DFFPOSX1_3016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_97__7_), .Q(data_187__7_) );
DFFPOSX1 DFFPOSX1_3017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_97__8_), .Q(data_187__8_) );
DFFPOSX1 DFFPOSX1_3018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_97__9_), .Q(data_187__9_) );
DFFPOSX1 DFFPOSX1_3019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_97__10_), .Q(data_187__10_) );
DFFPOSX1 DFFPOSX1_3020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_97__11_), .Q(data_187__11_) );
DFFPOSX1 DFFPOSX1_3021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_97__12_), .Q(data_187__12_) );
DFFPOSX1 DFFPOSX1_3022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_97__13_), .Q(data_187__13_) );
DFFPOSX1 DFFPOSX1_3023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_97__14_), .Q(data_187__14_) );
DFFPOSX1 DFFPOSX1_3024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_97__15_), .Q(data_187__15_) );
DFFPOSX1 DFFPOSX1_3025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_98__0_), .Q(data_188__0_) );
DFFPOSX1 DFFPOSX1_3026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_98__1_), .Q(data_188__1_) );
DFFPOSX1 DFFPOSX1_3027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_98__2_), .Q(data_188__2_) );
DFFPOSX1 DFFPOSX1_3028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_98__3_), .Q(data_188__3_) );
DFFPOSX1 DFFPOSX1_3029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_98__4_), .Q(data_188__4_) );
DFFPOSX1 DFFPOSX1_3030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_98__5_), .Q(data_188__5_) );
DFFPOSX1 DFFPOSX1_3031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_98__6_), .Q(data_188__6_) );
DFFPOSX1 DFFPOSX1_3032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_98__7_), .Q(data_188__7_) );
DFFPOSX1 DFFPOSX1_3033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_98__8_), .Q(data_188__8_) );
DFFPOSX1 DFFPOSX1_3034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_98__9_), .Q(data_188__9_) );
DFFPOSX1 DFFPOSX1_3035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_98__10_), .Q(data_188__10_) );
DFFPOSX1 DFFPOSX1_3036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_98__11_), .Q(data_188__11_) );
DFFPOSX1 DFFPOSX1_3037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_98__12_), .Q(data_188__12_) );
DFFPOSX1 DFFPOSX1_3038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_98__13_), .Q(data_188__13_) );
DFFPOSX1 DFFPOSX1_3039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_98__14_), .Q(data_188__14_) );
DFFPOSX1 DFFPOSX1_3040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_98__15_), .Q(data_188__15_) );
DFFPOSX1 DFFPOSX1_3041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_99__0_), .Q(data_189__0_) );
DFFPOSX1 DFFPOSX1_3042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_99__1_), .Q(data_189__1_) );
DFFPOSX1 DFFPOSX1_3043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_99__2_), .Q(data_189__2_) );
DFFPOSX1 DFFPOSX1_3044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_99__3_), .Q(data_189__3_) );
DFFPOSX1 DFFPOSX1_3045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_99__4_), .Q(data_189__4_) );
DFFPOSX1 DFFPOSX1_3046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_99__5_), .Q(data_189__5_) );
DFFPOSX1 DFFPOSX1_3047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_99__6_), .Q(data_189__6_) );
DFFPOSX1 DFFPOSX1_3048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_99__7_), .Q(data_189__7_) );
DFFPOSX1 DFFPOSX1_3049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_99__8_), .Q(data_189__8_) );
DFFPOSX1 DFFPOSX1_3050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_99__9_), .Q(data_189__9_) );
DFFPOSX1 DFFPOSX1_3051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_99__10_), .Q(data_189__10_) );
DFFPOSX1 DFFPOSX1_3052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_99__11_), .Q(data_189__11_) );
DFFPOSX1 DFFPOSX1_3053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_99__12_), .Q(data_189__12_) );
DFFPOSX1 DFFPOSX1_3054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_99__13_), .Q(data_189__13_) );
DFFPOSX1 DFFPOSX1_3055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_99__14_), .Q(data_189__14_) );
DFFPOSX1 DFFPOSX1_3056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_99__15_), .Q(data_189__15_) );
DFFPOSX1 DFFPOSX1_3057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_101__0_), .Q(data_190__0_) );
DFFPOSX1 DFFPOSX1_3058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_101__1_), .Q(data_190__1_) );
DFFPOSX1 DFFPOSX1_3059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_101__2_), .Q(data_190__2_) );
DFFPOSX1 DFFPOSX1_3060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_101__3_), .Q(data_190__3_) );
DFFPOSX1 DFFPOSX1_3061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_101__4_), .Q(data_190__4_) );
DFFPOSX1 DFFPOSX1_3062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_101__5_), .Q(data_190__5_) );
DFFPOSX1 DFFPOSX1_3063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_101__6_), .Q(data_190__6_) );
DFFPOSX1 DFFPOSX1_3064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_101__7_), .Q(data_190__7_) );
DFFPOSX1 DFFPOSX1_3065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_101__8_), .Q(data_190__8_) );
DFFPOSX1 DFFPOSX1_3066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_101__9_), .Q(data_190__9_) );
DFFPOSX1 DFFPOSX1_3067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_101__10_), .Q(data_190__10_) );
DFFPOSX1 DFFPOSX1_3068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_101__11_), .Q(data_190__11_) );
DFFPOSX1 DFFPOSX1_3069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_101__12_), .Q(data_190__12_) );
DFFPOSX1 DFFPOSX1_3070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_101__13_), .Q(data_190__13_) );
DFFPOSX1 DFFPOSX1_3071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_101__14_), .Q(data_190__14_) );
DFFPOSX1 DFFPOSX1_3072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_101__15_), .Q(data_190__15_) );
DFFPOSX1 DFFPOSX1_3073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf3), .D(_102__0_), .Q(data_191__0_) );
DFFPOSX1 DFFPOSX1_3074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf3), .D(_102__1_), .Q(data_191__1_) );
DFFPOSX1 DFFPOSX1_3075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf3), .D(_102__2_), .Q(data_191__2_) );
DFFPOSX1 DFFPOSX1_3076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf3), .D(_102__3_), .Q(data_191__3_) );
DFFPOSX1 DFFPOSX1_3077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf3), .D(_102__4_), .Q(data_191__4_) );
DFFPOSX1 DFFPOSX1_3078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf3), .D(_102__5_), .Q(data_191__5_) );
DFFPOSX1 DFFPOSX1_3079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf3), .D(_102__6_), .Q(data_191__6_) );
DFFPOSX1 DFFPOSX1_3080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf3), .D(_102__7_), .Q(data_191__7_) );
DFFPOSX1 DFFPOSX1_3081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf3), .D(_102__8_), .Q(data_191__8_) );
DFFPOSX1 DFFPOSX1_3082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf3), .D(_102__9_), .Q(data_191__9_) );
DFFPOSX1 DFFPOSX1_3083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf3), .D(_102__10_), .Q(data_191__10_) );
DFFPOSX1 DFFPOSX1_3084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf3), .D(_102__11_), .Q(data_191__11_) );
DFFPOSX1 DFFPOSX1_3085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf3), .D(_102__12_), .Q(data_191__12_) );
DFFPOSX1 DFFPOSX1_3086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf3), .D(_102__13_), .Q(data_191__13_) );
DFFPOSX1 DFFPOSX1_3087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf3), .D(_102__14_), .Q(data_191__14_) );
DFFPOSX1 DFFPOSX1_3088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf3), .D(_102__15_), .Q(data_191__15_) );
DFFPOSX1 DFFPOSX1_3089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_103__0_), .Q(data_192__0_) );
DFFPOSX1 DFFPOSX1_3090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_103__1_), .Q(data_192__1_) );
DFFPOSX1 DFFPOSX1_3091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_103__2_), .Q(data_192__2_) );
DFFPOSX1 DFFPOSX1_3092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_103__3_), .Q(data_192__3_) );
DFFPOSX1 DFFPOSX1_3093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_103__4_), .Q(data_192__4_) );
DFFPOSX1 DFFPOSX1_3094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_103__5_), .Q(data_192__5_) );
DFFPOSX1 DFFPOSX1_3095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_103__6_), .Q(data_192__6_) );
DFFPOSX1 DFFPOSX1_3096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_103__7_), .Q(data_192__7_) );
DFFPOSX1 DFFPOSX1_3097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_103__8_), .Q(data_192__8_) );
DFFPOSX1 DFFPOSX1_3098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_103__9_), .Q(data_192__9_) );
DFFPOSX1 DFFPOSX1_3099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_103__10_), .Q(data_192__10_) );
DFFPOSX1 DFFPOSX1_3100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_103__11_), .Q(data_192__11_) );
DFFPOSX1 DFFPOSX1_3101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_103__12_), .Q(data_192__12_) );
DFFPOSX1 DFFPOSX1_3102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_103__13_), .Q(data_192__13_) );
DFFPOSX1 DFFPOSX1_3103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_103__14_), .Q(data_192__14_) );
DFFPOSX1 DFFPOSX1_3104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_103__15_), .Q(data_192__15_) );
DFFPOSX1 DFFPOSX1_3105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_104__0_), .Q(data_193__0_) );
DFFPOSX1 DFFPOSX1_3106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_104__1_), .Q(data_193__1_) );
DFFPOSX1 DFFPOSX1_3107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_104__2_), .Q(data_193__2_) );
DFFPOSX1 DFFPOSX1_3108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_104__3_), .Q(data_193__3_) );
DFFPOSX1 DFFPOSX1_3109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_104__4_), .Q(data_193__4_) );
DFFPOSX1 DFFPOSX1_3110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_104__5_), .Q(data_193__5_) );
DFFPOSX1 DFFPOSX1_3111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_104__6_), .Q(data_193__6_) );
DFFPOSX1 DFFPOSX1_3112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_104__7_), .Q(data_193__7_) );
DFFPOSX1 DFFPOSX1_3113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_104__8_), .Q(data_193__8_) );
DFFPOSX1 DFFPOSX1_3114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_104__9_), .Q(data_193__9_) );
DFFPOSX1 DFFPOSX1_3115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_104__10_), .Q(data_193__10_) );
DFFPOSX1 DFFPOSX1_3116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_104__11_), .Q(data_193__11_) );
DFFPOSX1 DFFPOSX1_3117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_104__12_), .Q(data_193__12_) );
DFFPOSX1 DFFPOSX1_3118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_104__13_), .Q(data_193__13_) );
DFFPOSX1 DFFPOSX1_3119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_104__14_), .Q(data_193__14_) );
DFFPOSX1 DFFPOSX1_3120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_104__15_), .Q(data_193__15_) );
DFFPOSX1 DFFPOSX1_3121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_105__0_), .Q(data_194__0_) );
DFFPOSX1 DFFPOSX1_3122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_105__1_), .Q(data_194__1_) );
DFFPOSX1 DFFPOSX1_3123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_105__2_), .Q(data_194__2_) );
DFFPOSX1 DFFPOSX1_3124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_105__3_), .Q(data_194__3_) );
DFFPOSX1 DFFPOSX1_3125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_105__4_), .Q(data_194__4_) );
DFFPOSX1 DFFPOSX1_3126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_105__5_), .Q(data_194__5_) );
DFFPOSX1 DFFPOSX1_3127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_105__6_), .Q(data_194__6_) );
DFFPOSX1 DFFPOSX1_3128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_105__7_), .Q(data_194__7_) );
DFFPOSX1 DFFPOSX1_3129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_105__8_), .Q(data_194__8_) );
DFFPOSX1 DFFPOSX1_3130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_105__9_), .Q(data_194__9_) );
DFFPOSX1 DFFPOSX1_3131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_105__10_), .Q(data_194__10_) );
DFFPOSX1 DFFPOSX1_3132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_105__11_), .Q(data_194__11_) );
DFFPOSX1 DFFPOSX1_3133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_105__12_), .Q(data_194__12_) );
DFFPOSX1 DFFPOSX1_3134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_105__13_), .Q(data_194__13_) );
DFFPOSX1 DFFPOSX1_3135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_105__14_), .Q(data_194__14_) );
DFFPOSX1 DFFPOSX1_3136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_105__15_), .Q(data_194__15_) );
DFFPOSX1 DFFPOSX1_3137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_106__0_), .Q(data_195__0_) );
DFFPOSX1 DFFPOSX1_3138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_106__1_), .Q(data_195__1_) );
DFFPOSX1 DFFPOSX1_3139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_106__2_), .Q(data_195__2_) );
DFFPOSX1 DFFPOSX1_3140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_106__3_), .Q(data_195__3_) );
DFFPOSX1 DFFPOSX1_3141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_106__4_), .Q(data_195__4_) );
DFFPOSX1 DFFPOSX1_3142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_106__5_), .Q(data_195__5_) );
DFFPOSX1 DFFPOSX1_3143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_106__6_), .Q(data_195__6_) );
DFFPOSX1 DFFPOSX1_3144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_106__7_), .Q(data_195__7_) );
DFFPOSX1 DFFPOSX1_3145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_106__8_), .Q(data_195__8_) );
DFFPOSX1 DFFPOSX1_3146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_106__9_), .Q(data_195__9_) );
DFFPOSX1 DFFPOSX1_3147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_106__10_), .Q(data_195__10_) );
DFFPOSX1 DFFPOSX1_3148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_106__11_), .Q(data_195__11_) );
DFFPOSX1 DFFPOSX1_3149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_106__12_), .Q(data_195__12_) );
DFFPOSX1 DFFPOSX1_3150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_106__13_), .Q(data_195__13_) );
DFFPOSX1 DFFPOSX1_3151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_106__14_), .Q(data_195__14_) );
DFFPOSX1 DFFPOSX1_3152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_106__15_), .Q(data_195__15_) );
DFFPOSX1 DFFPOSX1_3153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_107__0_), .Q(data_196__0_) );
DFFPOSX1 DFFPOSX1_3154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_107__1_), .Q(data_196__1_) );
DFFPOSX1 DFFPOSX1_3155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_107__2_), .Q(data_196__2_) );
DFFPOSX1 DFFPOSX1_3156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_107__3_), .Q(data_196__3_) );
DFFPOSX1 DFFPOSX1_3157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_107__4_), .Q(data_196__4_) );
DFFPOSX1 DFFPOSX1_3158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_107__5_), .Q(data_196__5_) );
DFFPOSX1 DFFPOSX1_3159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_107__6_), .Q(data_196__6_) );
DFFPOSX1 DFFPOSX1_3160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_107__7_), .Q(data_196__7_) );
DFFPOSX1 DFFPOSX1_3161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_107__8_), .Q(data_196__8_) );
DFFPOSX1 DFFPOSX1_3162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_107__9_), .Q(data_196__9_) );
DFFPOSX1 DFFPOSX1_3163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_107__10_), .Q(data_196__10_) );
DFFPOSX1 DFFPOSX1_3164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_107__11_), .Q(data_196__11_) );
DFFPOSX1 DFFPOSX1_3165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_107__12_), .Q(data_196__12_) );
DFFPOSX1 DFFPOSX1_3166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_107__13_), .Q(data_196__13_) );
DFFPOSX1 DFFPOSX1_3167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_107__14_), .Q(data_196__14_) );
DFFPOSX1 DFFPOSX1_3168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_107__15_), .Q(data_196__15_) );
DFFPOSX1 DFFPOSX1_3169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_108__0_), .Q(data_197__0_) );
DFFPOSX1 DFFPOSX1_3170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_108__1_), .Q(data_197__1_) );
DFFPOSX1 DFFPOSX1_3171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_108__2_), .Q(data_197__2_) );
DFFPOSX1 DFFPOSX1_3172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_108__3_), .Q(data_197__3_) );
DFFPOSX1 DFFPOSX1_3173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_108__4_), .Q(data_197__4_) );
DFFPOSX1 DFFPOSX1_3174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_108__5_), .Q(data_197__5_) );
DFFPOSX1 DFFPOSX1_3175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_108__6_), .Q(data_197__6_) );
DFFPOSX1 DFFPOSX1_3176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_108__7_), .Q(data_197__7_) );
DFFPOSX1 DFFPOSX1_3177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_108__8_), .Q(data_197__8_) );
DFFPOSX1 DFFPOSX1_3178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_108__9_), .Q(data_197__9_) );
DFFPOSX1 DFFPOSX1_3179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_108__10_), .Q(data_197__10_) );
DFFPOSX1 DFFPOSX1_3180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_108__11_), .Q(data_197__11_) );
DFFPOSX1 DFFPOSX1_3181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_108__12_), .Q(data_197__12_) );
DFFPOSX1 DFFPOSX1_3182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_108__13_), .Q(data_197__13_) );
DFFPOSX1 DFFPOSX1_3183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_108__14_), .Q(data_197__14_) );
DFFPOSX1 DFFPOSX1_3184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_108__15_), .Q(data_197__15_) );
DFFPOSX1 DFFPOSX1_3185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_109__0_), .Q(data_198__0_) );
DFFPOSX1 DFFPOSX1_3186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_109__1_), .Q(data_198__1_) );
DFFPOSX1 DFFPOSX1_3187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_109__2_), .Q(data_198__2_) );
DFFPOSX1 DFFPOSX1_3188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_109__3_), .Q(data_198__3_) );
DFFPOSX1 DFFPOSX1_3189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_109__4_), .Q(data_198__4_) );
DFFPOSX1 DFFPOSX1_3190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_109__5_), .Q(data_198__5_) );
DFFPOSX1 DFFPOSX1_3191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_109__6_), .Q(data_198__6_) );
DFFPOSX1 DFFPOSX1_3192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_109__7_), .Q(data_198__7_) );
DFFPOSX1 DFFPOSX1_3193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_109__8_), .Q(data_198__8_) );
DFFPOSX1 DFFPOSX1_3194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_109__9_), .Q(data_198__9_) );
DFFPOSX1 DFFPOSX1_3195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_109__10_), .Q(data_198__10_) );
DFFPOSX1 DFFPOSX1_3196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_109__11_), .Q(data_198__11_) );
DFFPOSX1 DFFPOSX1_3197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_109__12_), .Q(data_198__12_) );
DFFPOSX1 DFFPOSX1_3198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_109__13_), .Q(data_198__13_) );
DFFPOSX1 DFFPOSX1_3199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_109__14_), .Q(data_198__14_) );
DFFPOSX1 DFFPOSX1_3200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_109__15_), .Q(data_198__15_) );
DFFPOSX1 DFFPOSX1_3201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_110__0_), .Q(data_199__0_) );
DFFPOSX1 DFFPOSX1_3202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_110__1_), .Q(data_199__1_) );
DFFPOSX1 DFFPOSX1_3203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_110__2_), .Q(data_199__2_) );
DFFPOSX1 DFFPOSX1_3204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_110__3_), .Q(data_199__3_) );
DFFPOSX1 DFFPOSX1_3205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_110__4_), .Q(data_199__4_) );
DFFPOSX1 DFFPOSX1_3206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_110__5_), .Q(data_199__5_) );
DFFPOSX1 DFFPOSX1_3207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_110__6_), .Q(data_199__6_) );
DFFPOSX1 DFFPOSX1_3208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_110__7_), .Q(data_199__7_) );
DFFPOSX1 DFFPOSX1_3209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_110__8_), .Q(data_199__8_) );
DFFPOSX1 DFFPOSX1_3210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_110__9_), .Q(data_199__9_) );
DFFPOSX1 DFFPOSX1_3211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_110__10_), .Q(data_199__10_) );
DFFPOSX1 DFFPOSX1_3212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_110__11_), .Q(data_199__11_) );
DFFPOSX1 DFFPOSX1_3213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_110__12_), .Q(data_199__12_) );
DFFPOSX1 DFFPOSX1_3214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_110__13_), .Q(data_199__13_) );
DFFPOSX1 DFFPOSX1_3215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_110__14_), .Q(data_199__14_) );
DFFPOSX1 DFFPOSX1_3216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_110__15_), .Q(data_199__15_) );
DFFPOSX1 DFFPOSX1_3217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_113__0_), .Q(data_200__0_) );
DFFPOSX1 DFFPOSX1_3218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_113__1_), .Q(data_200__1_) );
DFFPOSX1 DFFPOSX1_3219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_113__2_), .Q(data_200__2_) );
DFFPOSX1 DFFPOSX1_3220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_113__3_), .Q(data_200__3_) );
DFFPOSX1 DFFPOSX1_3221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_113__4_), .Q(data_200__4_) );
DFFPOSX1 DFFPOSX1_3222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_113__5_), .Q(data_200__5_) );
DFFPOSX1 DFFPOSX1_3223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_113__6_), .Q(data_200__6_) );
DFFPOSX1 DFFPOSX1_3224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_113__7_), .Q(data_200__7_) );
DFFPOSX1 DFFPOSX1_3225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_113__8_), .Q(data_200__8_) );
DFFPOSX1 DFFPOSX1_3226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_113__9_), .Q(data_200__9_) );
DFFPOSX1 DFFPOSX1_3227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_113__10_), .Q(data_200__10_) );
DFFPOSX1 DFFPOSX1_3228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_113__11_), .Q(data_200__11_) );
DFFPOSX1 DFFPOSX1_3229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_113__12_), .Q(data_200__12_) );
DFFPOSX1 DFFPOSX1_3230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_113__13_), .Q(data_200__13_) );
DFFPOSX1 DFFPOSX1_3231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_113__14_), .Q(data_200__14_) );
DFFPOSX1 DFFPOSX1_3232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_113__15_), .Q(data_200__15_) );
DFFPOSX1 DFFPOSX1_3233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_114__0_), .Q(data_201__0_) );
DFFPOSX1 DFFPOSX1_3234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_114__1_), .Q(data_201__1_) );
DFFPOSX1 DFFPOSX1_3235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_114__2_), .Q(data_201__2_) );
DFFPOSX1 DFFPOSX1_3236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_114__3_), .Q(data_201__3_) );
DFFPOSX1 DFFPOSX1_3237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_114__4_), .Q(data_201__4_) );
DFFPOSX1 DFFPOSX1_3238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_114__5_), .Q(data_201__5_) );
DFFPOSX1 DFFPOSX1_3239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_114__6_), .Q(data_201__6_) );
DFFPOSX1 DFFPOSX1_3240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_114__7_), .Q(data_201__7_) );
DFFPOSX1 DFFPOSX1_3241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_114__8_), .Q(data_201__8_) );
DFFPOSX1 DFFPOSX1_3242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_114__9_), .Q(data_201__9_) );
DFFPOSX1 DFFPOSX1_3243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_114__10_), .Q(data_201__10_) );
DFFPOSX1 DFFPOSX1_3244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_114__11_), .Q(data_201__11_) );
DFFPOSX1 DFFPOSX1_3245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_114__12_), .Q(data_201__12_) );
DFFPOSX1 DFFPOSX1_3246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_114__13_), .Q(data_201__13_) );
DFFPOSX1 DFFPOSX1_3247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_114__14_), .Q(data_201__14_) );
DFFPOSX1 DFFPOSX1_3248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_114__15_), .Q(data_201__15_) );
DFFPOSX1 DFFPOSX1_3249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_115__0_), .Q(data_202__0_) );
DFFPOSX1 DFFPOSX1_3250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_115__1_), .Q(data_202__1_) );
DFFPOSX1 DFFPOSX1_3251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_115__2_), .Q(data_202__2_) );
DFFPOSX1 DFFPOSX1_3252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_115__3_), .Q(data_202__3_) );
DFFPOSX1 DFFPOSX1_3253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_115__4_), .Q(data_202__4_) );
DFFPOSX1 DFFPOSX1_3254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_115__5_), .Q(data_202__5_) );
DFFPOSX1 DFFPOSX1_3255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_115__6_), .Q(data_202__6_) );
DFFPOSX1 DFFPOSX1_3256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_115__7_), .Q(data_202__7_) );
DFFPOSX1 DFFPOSX1_3257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_115__8_), .Q(data_202__8_) );
DFFPOSX1 DFFPOSX1_3258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_115__9_), .Q(data_202__9_) );
DFFPOSX1 DFFPOSX1_3259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_115__10_), .Q(data_202__10_) );
DFFPOSX1 DFFPOSX1_3260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_115__11_), .Q(data_202__11_) );
DFFPOSX1 DFFPOSX1_3261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_115__12_), .Q(data_202__12_) );
DFFPOSX1 DFFPOSX1_3262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_115__13_), .Q(data_202__13_) );
DFFPOSX1 DFFPOSX1_3263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_115__14_), .Q(data_202__14_) );
DFFPOSX1 DFFPOSX1_3264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_115__15_), .Q(data_202__15_) );
DFFPOSX1 DFFPOSX1_3265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_116__0_), .Q(data_203__0_) );
DFFPOSX1 DFFPOSX1_3266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_116__1_), .Q(data_203__1_) );
DFFPOSX1 DFFPOSX1_3267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_116__2_), .Q(data_203__2_) );
DFFPOSX1 DFFPOSX1_3268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_116__3_), .Q(data_203__3_) );
DFFPOSX1 DFFPOSX1_3269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_116__4_), .Q(data_203__4_) );
DFFPOSX1 DFFPOSX1_3270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_116__5_), .Q(data_203__5_) );
DFFPOSX1 DFFPOSX1_3271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_116__6_), .Q(data_203__6_) );
DFFPOSX1 DFFPOSX1_3272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_116__7_), .Q(data_203__7_) );
DFFPOSX1 DFFPOSX1_3273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_116__8_), .Q(data_203__8_) );
DFFPOSX1 DFFPOSX1_3274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_116__9_), .Q(data_203__9_) );
DFFPOSX1 DFFPOSX1_3275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_116__10_), .Q(data_203__10_) );
DFFPOSX1 DFFPOSX1_3276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_116__11_), .Q(data_203__11_) );
DFFPOSX1 DFFPOSX1_3277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_116__12_), .Q(data_203__12_) );
DFFPOSX1 DFFPOSX1_3278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_116__13_), .Q(data_203__13_) );
DFFPOSX1 DFFPOSX1_3279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_116__14_), .Q(data_203__14_) );
DFFPOSX1 DFFPOSX1_3280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_116__15_), .Q(data_203__15_) );
DFFPOSX1 DFFPOSX1_3281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_117__0_), .Q(data_204__0_) );
DFFPOSX1 DFFPOSX1_3282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_117__1_), .Q(data_204__1_) );
DFFPOSX1 DFFPOSX1_3283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_117__2_), .Q(data_204__2_) );
DFFPOSX1 DFFPOSX1_3284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_117__3_), .Q(data_204__3_) );
DFFPOSX1 DFFPOSX1_3285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_117__4_), .Q(data_204__4_) );
DFFPOSX1 DFFPOSX1_3286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_117__5_), .Q(data_204__5_) );
DFFPOSX1 DFFPOSX1_3287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_117__6_), .Q(data_204__6_) );
DFFPOSX1 DFFPOSX1_3288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_117__7_), .Q(data_204__7_) );
DFFPOSX1 DFFPOSX1_3289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_117__8_), .Q(data_204__8_) );
DFFPOSX1 DFFPOSX1_3290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_117__9_), .Q(data_204__9_) );
DFFPOSX1 DFFPOSX1_3291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_117__10_), .Q(data_204__10_) );
DFFPOSX1 DFFPOSX1_3292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_117__11_), .Q(data_204__11_) );
DFFPOSX1 DFFPOSX1_3293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_117__12_), .Q(data_204__12_) );
DFFPOSX1 DFFPOSX1_3294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_117__13_), .Q(data_204__13_) );
DFFPOSX1 DFFPOSX1_3295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_117__14_), .Q(data_204__14_) );
DFFPOSX1 DFFPOSX1_3296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_117__15_), .Q(data_204__15_) );
DFFPOSX1 DFFPOSX1_3297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_118__0_), .Q(data_205__0_) );
DFFPOSX1 DFFPOSX1_3298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_118__1_), .Q(data_205__1_) );
DFFPOSX1 DFFPOSX1_3299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_118__2_), .Q(data_205__2_) );
DFFPOSX1 DFFPOSX1_3300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_118__3_), .Q(data_205__3_) );
DFFPOSX1 DFFPOSX1_3301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_118__4_), .Q(data_205__4_) );
DFFPOSX1 DFFPOSX1_3302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_118__5_), .Q(data_205__5_) );
DFFPOSX1 DFFPOSX1_3303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_118__6_), .Q(data_205__6_) );
DFFPOSX1 DFFPOSX1_3304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_118__7_), .Q(data_205__7_) );
DFFPOSX1 DFFPOSX1_3305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_118__8_), .Q(data_205__8_) );
DFFPOSX1 DFFPOSX1_3306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_118__9_), .Q(data_205__9_) );
DFFPOSX1 DFFPOSX1_3307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_118__10_), .Q(data_205__10_) );
DFFPOSX1 DFFPOSX1_3308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_118__11_), .Q(data_205__11_) );
DFFPOSX1 DFFPOSX1_3309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_118__12_), .Q(data_205__12_) );
DFFPOSX1 DFFPOSX1_3310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_118__13_), .Q(data_205__13_) );
DFFPOSX1 DFFPOSX1_3311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_118__14_), .Q(data_205__14_) );
DFFPOSX1 DFFPOSX1_3312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_118__15_), .Q(data_205__15_) );
DFFPOSX1 DFFPOSX1_3313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_119__0_), .Q(data_206__0_) );
DFFPOSX1 DFFPOSX1_3314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_119__1_), .Q(data_206__1_) );
DFFPOSX1 DFFPOSX1_3315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_119__2_), .Q(data_206__2_) );
DFFPOSX1 DFFPOSX1_3316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_119__3_), .Q(data_206__3_) );
DFFPOSX1 DFFPOSX1_3317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_119__4_), .Q(data_206__4_) );
DFFPOSX1 DFFPOSX1_3318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_119__5_), .Q(data_206__5_) );
DFFPOSX1 DFFPOSX1_3319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_119__6_), .Q(data_206__6_) );
DFFPOSX1 DFFPOSX1_3320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_119__7_), .Q(data_206__7_) );
DFFPOSX1 DFFPOSX1_3321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_119__8_), .Q(data_206__8_) );
DFFPOSX1 DFFPOSX1_3322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_119__9_), .Q(data_206__9_) );
DFFPOSX1 DFFPOSX1_3323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_119__10_), .Q(data_206__10_) );
DFFPOSX1 DFFPOSX1_3324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_119__11_), .Q(data_206__11_) );
DFFPOSX1 DFFPOSX1_3325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_119__12_), .Q(data_206__12_) );
DFFPOSX1 DFFPOSX1_3326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_119__13_), .Q(data_206__13_) );
DFFPOSX1 DFFPOSX1_3327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_119__14_), .Q(data_206__14_) );
DFFPOSX1 DFFPOSX1_3328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_119__15_), .Q(data_206__15_) );
DFFPOSX1 DFFPOSX1_3329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf2), .D(_120__0_), .Q(data_207__0_) );
DFFPOSX1 DFFPOSX1_3330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf2), .D(_120__1_), .Q(data_207__1_) );
DFFPOSX1 DFFPOSX1_3331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf2), .D(_120__2_), .Q(data_207__2_) );
DFFPOSX1 DFFPOSX1_3332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf2), .D(_120__3_), .Q(data_207__3_) );
DFFPOSX1 DFFPOSX1_3333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf2), .D(_120__4_), .Q(data_207__4_) );
DFFPOSX1 DFFPOSX1_3334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf2), .D(_120__5_), .Q(data_207__5_) );
DFFPOSX1 DFFPOSX1_3335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf2), .D(_120__6_), .Q(data_207__6_) );
DFFPOSX1 DFFPOSX1_3336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf2), .D(_120__7_), .Q(data_207__7_) );
DFFPOSX1 DFFPOSX1_3337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf2), .D(_120__8_), .Q(data_207__8_) );
DFFPOSX1 DFFPOSX1_3338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf2), .D(_120__9_), .Q(data_207__9_) );
DFFPOSX1 DFFPOSX1_3339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf2), .D(_120__10_), .Q(data_207__10_) );
DFFPOSX1 DFFPOSX1_3340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf2), .D(_120__11_), .Q(data_207__11_) );
DFFPOSX1 DFFPOSX1_3341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf2), .D(_120__12_), .Q(data_207__12_) );
DFFPOSX1 DFFPOSX1_3342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf2), .D(_120__13_), .Q(data_207__13_) );
DFFPOSX1 DFFPOSX1_3343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf2), .D(_120__14_), .Q(data_207__14_) );
DFFPOSX1 DFFPOSX1_3344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf2), .D(_120__15_), .Q(data_207__15_) );
DFFPOSX1 DFFPOSX1_3345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_121__0_), .Q(data_208__0_) );
DFFPOSX1 DFFPOSX1_3346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_121__1_), .Q(data_208__1_) );
DFFPOSX1 DFFPOSX1_3347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_121__2_), .Q(data_208__2_) );
DFFPOSX1 DFFPOSX1_3348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_121__3_), .Q(data_208__3_) );
DFFPOSX1 DFFPOSX1_3349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_121__4_), .Q(data_208__4_) );
DFFPOSX1 DFFPOSX1_3350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_121__5_), .Q(data_208__5_) );
DFFPOSX1 DFFPOSX1_3351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_121__6_), .Q(data_208__6_) );
DFFPOSX1 DFFPOSX1_3352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_121__7_), .Q(data_208__7_) );
DFFPOSX1 DFFPOSX1_3353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_121__8_), .Q(data_208__8_) );
DFFPOSX1 DFFPOSX1_3354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_121__9_), .Q(data_208__9_) );
DFFPOSX1 DFFPOSX1_3355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_121__10_), .Q(data_208__10_) );
DFFPOSX1 DFFPOSX1_3356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_121__11_), .Q(data_208__11_) );
DFFPOSX1 DFFPOSX1_3357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_121__12_), .Q(data_208__12_) );
DFFPOSX1 DFFPOSX1_3358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_121__13_), .Q(data_208__13_) );
DFFPOSX1 DFFPOSX1_3359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_121__14_), .Q(data_208__14_) );
DFFPOSX1 DFFPOSX1_3360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_121__15_), .Q(data_208__15_) );
DFFPOSX1 DFFPOSX1_3361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_122__0_), .Q(data_209__0_) );
DFFPOSX1 DFFPOSX1_3362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_122__1_), .Q(data_209__1_) );
DFFPOSX1 DFFPOSX1_3363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_122__2_), .Q(data_209__2_) );
DFFPOSX1 DFFPOSX1_3364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_122__3_), .Q(data_209__3_) );
DFFPOSX1 DFFPOSX1_3365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_122__4_), .Q(data_209__4_) );
DFFPOSX1 DFFPOSX1_3366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_122__5_), .Q(data_209__5_) );
DFFPOSX1 DFFPOSX1_3367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_122__6_), .Q(data_209__6_) );
DFFPOSX1 DFFPOSX1_3368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_122__7_), .Q(data_209__7_) );
DFFPOSX1 DFFPOSX1_3369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_122__8_), .Q(data_209__8_) );
DFFPOSX1 DFFPOSX1_3370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_122__9_), .Q(data_209__9_) );
DFFPOSX1 DFFPOSX1_3371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_122__10_), .Q(data_209__10_) );
DFFPOSX1 DFFPOSX1_3372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_122__11_), .Q(data_209__11_) );
DFFPOSX1 DFFPOSX1_3373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_122__12_), .Q(data_209__12_) );
DFFPOSX1 DFFPOSX1_3374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_122__13_), .Q(data_209__13_) );
DFFPOSX1 DFFPOSX1_3375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_122__14_), .Q(data_209__14_) );
DFFPOSX1 DFFPOSX1_3376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_122__15_), .Q(data_209__15_) );
DFFPOSX1 DFFPOSX1_3377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_124__0_), .Q(data_210__0_) );
DFFPOSX1 DFFPOSX1_3378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_124__1_), .Q(data_210__1_) );
DFFPOSX1 DFFPOSX1_3379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_124__2_), .Q(data_210__2_) );
DFFPOSX1 DFFPOSX1_3380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_124__3_), .Q(data_210__3_) );
DFFPOSX1 DFFPOSX1_3381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_124__4_), .Q(data_210__4_) );
DFFPOSX1 DFFPOSX1_3382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_124__5_), .Q(data_210__5_) );
DFFPOSX1 DFFPOSX1_3383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_124__6_), .Q(data_210__6_) );
DFFPOSX1 DFFPOSX1_3384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_124__7_), .Q(data_210__7_) );
DFFPOSX1 DFFPOSX1_3385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_124__8_), .Q(data_210__8_) );
DFFPOSX1 DFFPOSX1_3386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_124__9_), .Q(data_210__9_) );
DFFPOSX1 DFFPOSX1_3387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_124__10_), .Q(data_210__10_) );
DFFPOSX1 DFFPOSX1_3388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_124__11_), .Q(data_210__11_) );
DFFPOSX1 DFFPOSX1_3389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_124__12_), .Q(data_210__12_) );
DFFPOSX1 DFFPOSX1_3390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_124__13_), .Q(data_210__13_) );
DFFPOSX1 DFFPOSX1_3391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_124__14_), .Q(data_210__14_) );
DFFPOSX1 DFFPOSX1_3392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_124__15_), .Q(data_210__15_) );
DFFPOSX1 DFFPOSX1_3393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_125__0_), .Q(data_211__0_) );
DFFPOSX1 DFFPOSX1_3394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_125__1_), .Q(data_211__1_) );
DFFPOSX1 DFFPOSX1_3395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_125__2_), .Q(data_211__2_) );
DFFPOSX1 DFFPOSX1_3396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_125__3_), .Q(data_211__3_) );
DFFPOSX1 DFFPOSX1_3397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_125__4_), .Q(data_211__4_) );
DFFPOSX1 DFFPOSX1_3398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_125__5_), .Q(data_211__5_) );
DFFPOSX1 DFFPOSX1_3399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_125__6_), .Q(data_211__6_) );
DFFPOSX1 DFFPOSX1_3400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_125__7_), .Q(data_211__7_) );
DFFPOSX1 DFFPOSX1_3401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_125__8_), .Q(data_211__8_) );
DFFPOSX1 DFFPOSX1_3402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_125__9_), .Q(data_211__9_) );
DFFPOSX1 DFFPOSX1_3403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_125__10_), .Q(data_211__10_) );
DFFPOSX1 DFFPOSX1_3404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_125__11_), .Q(data_211__11_) );
DFFPOSX1 DFFPOSX1_3405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_125__12_), .Q(data_211__12_) );
DFFPOSX1 DFFPOSX1_3406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_125__13_), .Q(data_211__13_) );
DFFPOSX1 DFFPOSX1_3407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_125__14_), .Q(data_211__14_) );
DFFPOSX1 DFFPOSX1_3408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_125__15_), .Q(data_211__15_) );
DFFPOSX1 DFFPOSX1_3409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_126__0_), .Q(data_212__0_) );
DFFPOSX1 DFFPOSX1_3410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_126__1_), .Q(data_212__1_) );
DFFPOSX1 DFFPOSX1_3411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_126__2_), .Q(data_212__2_) );
DFFPOSX1 DFFPOSX1_3412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_126__3_), .Q(data_212__3_) );
DFFPOSX1 DFFPOSX1_3413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_126__4_), .Q(data_212__4_) );
DFFPOSX1 DFFPOSX1_3414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_126__5_), .Q(data_212__5_) );
DFFPOSX1 DFFPOSX1_3415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_126__6_), .Q(data_212__6_) );
DFFPOSX1 DFFPOSX1_3416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_126__7_), .Q(data_212__7_) );
DFFPOSX1 DFFPOSX1_3417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_126__8_), .Q(data_212__8_) );
DFFPOSX1 DFFPOSX1_3418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_126__9_), .Q(data_212__9_) );
DFFPOSX1 DFFPOSX1_3419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_126__10_), .Q(data_212__10_) );
DFFPOSX1 DFFPOSX1_3420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_126__11_), .Q(data_212__11_) );
DFFPOSX1 DFFPOSX1_3421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_126__12_), .Q(data_212__12_) );
DFFPOSX1 DFFPOSX1_3422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_126__13_), .Q(data_212__13_) );
DFFPOSX1 DFFPOSX1_3423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_126__14_), .Q(data_212__14_) );
DFFPOSX1 DFFPOSX1_3424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_126__15_), .Q(data_212__15_) );
DFFPOSX1 DFFPOSX1_3425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_127__0_), .Q(data_213__0_) );
DFFPOSX1 DFFPOSX1_3426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_127__1_), .Q(data_213__1_) );
DFFPOSX1 DFFPOSX1_3427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_127__2_), .Q(data_213__2_) );
DFFPOSX1 DFFPOSX1_3428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_127__3_), .Q(data_213__3_) );
DFFPOSX1 DFFPOSX1_3429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_127__4_), .Q(data_213__4_) );
DFFPOSX1 DFFPOSX1_3430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_127__5_), .Q(data_213__5_) );
DFFPOSX1 DFFPOSX1_3431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_127__6_), .Q(data_213__6_) );
DFFPOSX1 DFFPOSX1_3432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_127__7_), .Q(data_213__7_) );
DFFPOSX1 DFFPOSX1_3433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_127__8_), .Q(data_213__8_) );
DFFPOSX1 DFFPOSX1_3434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_127__9_), .Q(data_213__9_) );
DFFPOSX1 DFFPOSX1_3435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_127__10_), .Q(data_213__10_) );
DFFPOSX1 DFFPOSX1_3436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_127__11_), .Q(data_213__11_) );
DFFPOSX1 DFFPOSX1_3437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_127__12_), .Q(data_213__12_) );
DFFPOSX1 DFFPOSX1_3438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_127__13_), .Q(data_213__13_) );
DFFPOSX1 DFFPOSX1_3439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_127__14_), .Q(data_213__14_) );
DFFPOSX1 DFFPOSX1_3440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_127__15_), .Q(data_213__15_) );
DFFPOSX1 DFFPOSX1_3441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_128__0_), .Q(data_214__0_) );
DFFPOSX1 DFFPOSX1_3442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_128__1_), .Q(data_214__1_) );
DFFPOSX1 DFFPOSX1_3443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_128__2_), .Q(data_214__2_) );
DFFPOSX1 DFFPOSX1_3444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_128__3_), .Q(data_214__3_) );
DFFPOSX1 DFFPOSX1_3445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_128__4_), .Q(data_214__4_) );
DFFPOSX1 DFFPOSX1_3446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_128__5_), .Q(data_214__5_) );
DFFPOSX1 DFFPOSX1_3447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_128__6_), .Q(data_214__6_) );
DFFPOSX1 DFFPOSX1_3448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_128__7_), .Q(data_214__7_) );
DFFPOSX1 DFFPOSX1_3449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_128__8_), .Q(data_214__8_) );
DFFPOSX1 DFFPOSX1_3450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_128__9_), .Q(data_214__9_) );
DFFPOSX1 DFFPOSX1_3451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_128__10_), .Q(data_214__10_) );
DFFPOSX1 DFFPOSX1_3452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_128__11_), .Q(data_214__11_) );
DFFPOSX1 DFFPOSX1_3453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_128__12_), .Q(data_214__12_) );
DFFPOSX1 DFFPOSX1_3454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_128__13_), .Q(data_214__13_) );
DFFPOSX1 DFFPOSX1_3455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_128__14_), .Q(data_214__14_) );
DFFPOSX1 DFFPOSX1_3456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_128__15_), .Q(data_214__15_) );
DFFPOSX1 DFFPOSX1_3457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_129__0_), .Q(data_215__0_) );
DFFPOSX1 DFFPOSX1_3458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_129__1_), .Q(data_215__1_) );
DFFPOSX1 DFFPOSX1_3459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_129__2_), .Q(data_215__2_) );
DFFPOSX1 DFFPOSX1_3460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_129__3_), .Q(data_215__3_) );
DFFPOSX1 DFFPOSX1_3461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_129__4_), .Q(data_215__4_) );
DFFPOSX1 DFFPOSX1_3462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_129__5_), .Q(data_215__5_) );
DFFPOSX1 DFFPOSX1_3463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_129__6_), .Q(data_215__6_) );
DFFPOSX1 DFFPOSX1_3464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_129__7_), .Q(data_215__7_) );
DFFPOSX1 DFFPOSX1_3465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_129__8_), .Q(data_215__8_) );
DFFPOSX1 DFFPOSX1_3466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_129__9_), .Q(data_215__9_) );
DFFPOSX1 DFFPOSX1_3467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_129__10_), .Q(data_215__10_) );
DFFPOSX1 DFFPOSX1_3468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_129__11_), .Q(data_215__11_) );
DFFPOSX1 DFFPOSX1_3469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_129__12_), .Q(data_215__12_) );
DFFPOSX1 DFFPOSX1_3470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_129__13_), .Q(data_215__13_) );
DFFPOSX1 DFFPOSX1_3471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_129__14_), .Q(data_215__14_) );
DFFPOSX1 DFFPOSX1_3472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_129__15_), .Q(data_215__15_) );
DFFPOSX1 DFFPOSX1_3473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_130__0_), .Q(data_216__0_) );
DFFPOSX1 DFFPOSX1_3474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_130__1_), .Q(data_216__1_) );
DFFPOSX1 DFFPOSX1_3475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_130__2_), .Q(data_216__2_) );
DFFPOSX1 DFFPOSX1_3476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_130__3_), .Q(data_216__3_) );
DFFPOSX1 DFFPOSX1_3477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_130__4_), .Q(data_216__4_) );
DFFPOSX1 DFFPOSX1_3478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_130__5_), .Q(data_216__5_) );
DFFPOSX1 DFFPOSX1_3479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_130__6_), .Q(data_216__6_) );
DFFPOSX1 DFFPOSX1_3480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_130__7_), .Q(data_216__7_) );
DFFPOSX1 DFFPOSX1_3481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_130__8_), .Q(data_216__8_) );
DFFPOSX1 DFFPOSX1_3482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_130__9_), .Q(data_216__9_) );
DFFPOSX1 DFFPOSX1_3483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_130__10_), .Q(data_216__10_) );
DFFPOSX1 DFFPOSX1_3484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_130__11_), .Q(data_216__11_) );
DFFPOSX1 DFFPOSX1_3485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_130__12_), .Q(data_216__12_) );
DFFPOSX1 DFFPOSX1_3486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_130__13_), .Q(data_216__13_) );
DFFPOSX1 DFFPOSX1_3487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_130__14_), .Q(data_216__14_) );
DFFPOSX1 DFFPOSX1_3488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_130__15_), .Q(data_216__15_) );
DFFPOSX1 DFFPOSX1_3489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_131__0_), .Q(data_217__0_) );
DFFPOSX1 DFFPOSX1_3490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_131__1_), .Q(data_217__1_) );
DFFPOSX1 DFFPOSX1_3491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_131__2_), .Q(data_217__2_) );
DFFPOSX1 DFFPOSX1_3492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_131__3_), .Q(data_217__3_) );
DFFPOSX1 DFFPOSX1_3493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_131__4_), .Q(data_217__4_) );
DFFPOSX1 DFFPOSX1_3494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_131__5_), .Q(data_217__5_) );
DFFPOSX1 DFFPOSX1_3495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_131__6_), .Q(data_217__6_) );
DFFPOSX1 DFFPOSX1_3496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_131__7_), .Q(data_217__7_) );
DFFPOSX1 DFFPOSX1_3497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_131__8_), .Q(data_217__8_) );
DFFPOSX1 DFFPOSX1_3498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_131__9_), .Q(data_217__9_) );
DFFPOSX1 DFFPOSX1_3499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_131__10_), .Q(data_217__10_) );
DFFPOSX1 DFFPOSX1_3500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_131__11_), .Q(data_217__11_) );
DFFPOSX1 DFFPOSX1_3501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_131__12_), .Q(data_217__12_) );
DFFPOSX1 DFFPOSX1_3502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_131__13_), .Q(data_217__13_) );
DFFPOSX1 DFFPOSX1_3503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_131__14_), .Q(data_217__14_) );
DFFPOSX1 DFFPOSX1_3504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_131__15_), .Q(data_217__15_) );
DFFPOSX1 DFFPOSX1_3505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_132__0_), .Q(data_218__0_) );
DFFPOSX1 DFFPOSX1_3506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_132__1_), .Q(data_218__1_) );
DFFPOSX1 DFFPOSX1_3507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_132__2_), .Q(data_218__2_) );
DFFPOSX1 DFFPOSX1_3508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_132__3_), .Q(data_218__3_) );
DFFPOSX1 DFFPOSX1_3509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_132__4_), .Q(data_218__4_) );
DFFPOSX1 DFFPOSX1_3510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_132__5_), .Q(data_218__5_) );
DFFPOSX1 DFFPOSX1_3511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_132__6_), .Q(data_218__6_) );
DFFPOSX1 DFFPOSX1_3512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_132__7_), .Q(data_218__7_) );
DFFPOSX1 DFFPOSX1_3513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_132__8_), .Q(data_218__8_) );
DFFPOSX1 DFFPOSX1_3514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_132__9_), .Q(data_218__9_) );
DFFPOSX1 DFFPOSX1_3515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_132__10_), .Q(data_218__10_) );
DFFPOSX1 DFFPOSX1_3516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_132__11_), .Q(data_218__11_) );
DFFPOSX1 DFFPOSX1_3517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_132__12_), .Q(data_218__12_) );
DFFPOSX1 DFFPOSX1_3518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_132__13_), .Q(data_218__13_) );
DFFPOSX1 DFFPOSX1_3519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_132__14_), .Q(data_218__14_) );
DFFPOSX1 DFFPOSX1_3520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_132__15_), .Q(data_218__15_) );
DFFPOSX1 DFFPOSX1_3521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_133__0_), .Q(data_219__0_) );
DFFPOSX1 DFFPOSX1_3522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_133__1_), .Q(data_219__1_) );
DFFPOSX1 DFFPOSX1_3523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_133__2_), .Q(data_219__2_) );
DFFPOSX1 DFFPOSX1_3524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_133__3_), .Q(data_219__3_) );
DFFPOSX1 DFFPOSX1_3525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_133__4_), .Q(data_219__4_) );
DFFPOSX1 DFFPOSX1_3526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_133__5_), .Q(data_219__5_) );
DFFPOSX1 DFFPOSX1_3527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_133__6_), .Q(data_219__6_) );
DFFPOSX1 DFFPOSX1_3528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_133__7_), .Q(data_219__7_) );
DFFPOSX1 DFFPOSX1_3529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_133__8_), .Q(data_219__8_) );
DFFPOSX1 DFFPOSX1_3530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_133__9_), .Q(data_219__9_) );
DFFPOSX1 DFFPOSX1_3531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_133__10_), .Q(data_219__10_) );
DFFPOSX1 DFFPOSX1_3532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_133__11_), .Q(data_219__11_) );
DFFPOSX1 DFFPOSX1_3533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_133__12_), .Q(data_219__12_) );
DFFPOSX1 DFFPOSX1_3534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_133__13_), .Q(data_219__13_) );
DFFPOSX1 DFFPOSX1_3535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_133__14_), .Q(data_219__14_) );
DFFPOSX1 DFFPOSX1_3536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_133__15_), .Q(data_219__15_) );
DFFPOSX1 DFFPOSX1_3537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_135__0_), .Q(data_220__0_) );
DFFPOSX1 DFFPOSX1_3538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_135__1_), .Q(data_220__1_) );
DFFPOSX1 DFFPOSX1_3539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_135__2_), .Q(data_220__2_) );
DFFPOSX1 DFFPOSX1_3540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_135__3_), .Q(data_220__3_) );
DFFPOSX1 DFFPOSX1_3541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_135__4_), .Q(data_220__4_) );
DFFPOSX1 DFFPOSX1_3542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_135__5_), .Q(data_220__5_) );
DFFPOSX1 DFFPOSX1_3543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_135__6_), .Q(data_220__6_) );
DFFPOSX1 DFFPOSX1_3544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_135__7_), .Q(data_220__7_) );
DFFPOSX1 DFFPOSX1_3545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_135__8_), .Q(data_220__8_) );
DFFPOSX1 DFFPOSX1_3546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_135__9_), .Q(data_220__9_) );
DFFPOSX1 DFFPOSX1_3547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_135__10_), .Q(data_220__10_) );
DFFPOSX1 DFFPOSX1_3548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_135__11_), .Q(data_220__11_) );
DFFPOSX1 DFFPOSX1_3549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_135__12_), .Q(data_220__12_) );
DFFPOSX1 DFFPOSX1_3550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_135__13_), .Q(data_220__13_) );
DFFPOSX1 DFFPOSX1_3551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_135__14_), .Q(data_220__14_) );
DFFPOSX1 DFFPOSX1_3552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_135__15_), .Q(data_220__15_) );
DFFPOSX1 DFFPOSX1_3553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_136__0_), .Q(data_221__0_) );
DFFPOSX1 DFFPOSX1_3554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_136__1_), .Q(data_221__1_) );
DFFPOSX1 DFFPOSX1_3555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_136__2_), .Q(data_221__2_) );
DFFPOSX1 DFFPOSX1_3556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_136__3_), .Q(data_221__3_) );
DFFPOSX1 DFFPOSX1_3557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_136__4_), .Q(data_221__4_) );
DFFPOSX1 DFFPOSX1_3558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_136__5_), .Q(data_221__5_) );
DFFPOSX1 DFFPOSX1_3559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_136__6_), .Q(data_221__6_) );
DFFPOSX1 DFFPOSX1_3560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_136__7_), .Q(data_221__7_) );
DFFPOSX1 DFFPOSX1_3561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_136__8_), .Q(data_221__8_) );
DFFPOSX1 DFFPOSX1_3562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_136__9_), .Q(data_221__9_) );
DFFPOSX1 DFFPOSX1_3563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_136__10_), .Q(data_221__10_) );
DFFPOSX1 DFFPOSX1_3564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_136__11_), .Q(data_221__11_) );
DFFPOSX1 DFFPOSX1_3565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_136__12_), .Q(data_221__12_) );
DFFPOSX1 DFFPOSX1_3566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_136__13_), .Q(data_221__13_) );
DFFPOSX1 DFFPOSX1_3567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_136__14_), .Q(data_221__14_) );
DFFPOSX1 DFFPOSX1_3568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_136__15_), .Q(data_221__15_) );
DFFPOSX1 DFFPOSX1_3569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_137__0_), .Q(data_222__0_) );
DFFPOSX1 DFFPOSX1_3570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_137__1_), .Q(data_222__1_) );
DFFPOSX1 DFFPOSX1_3571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_137__2_), .Q(data_222__2_) );
DFFPOSX1 DFFPOSX1_3572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_137__3_), .Q(data_222__3_) );
DFFPOSX1 DFFPOSX1_3573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_137__4_), .Q(data_222__4_) );
DFFPOSX1 DFFPOSX1_3574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_137__5_), .Q(data_222__5_) );
DFFPOSX1 DFFPOSX1_3575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_137__6_), .Q(data_222__6_) );
DFFPOSX1 DFFPOSX1_3576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_137__7_), .Q(data_222__7_) );
DFFPOSX1 DFFPOSX1_3577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_137__8_), .Q(data_222__8_) );
DFFPOSX1 DFFPOSX1_3578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_137__9_), .Q(data_222__9_) );
DFFPOSX1 DFFPOSX1_3579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_137__10_), .Q(data_222__10_) );
DFFPOSX1 DFFPOSX1_3580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_137__11_), .Q(data_222__11_) );
DFFPOSX1 DFFPOSX1_3581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_137__12_), .Q(data_222__12_) );
DFFPOSX1 DFFPOSX1_3582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_137__13_), .Q(data_222__13_) );
DFFPOSX1 DFFPOSX1_3583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_137__14_), .Q(data_222__14_) );
DFFPOSX1 DFFPOSX1_3584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_137__15_), .Q(data_222__15_) );
DFFPOSX1 DFFPOSX1_3585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf1), .D(_138__0_), .Q(data_223__0_) );
DFFPOSX1 DFFPOSX1_3586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf1), .D(_138__1_), .Q(data_223__1_) );
DFFPOSX1 DFFPOSX1_3587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf1), .D(_138__2_), .Q(data_223__2_) );
DFFPOSX1 DFFPOSX1_3588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf1), .D(_138__3_), .Q(data_223__3_) );
DFFPOSX1 DFFPOSX1_3589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf1), .D(_138__4_), .Q(data_223__4_) );
DFFPOSX1 DFFPOSX1_3590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf1), .D(_138__5_), .Q(data_223__5_) );
DFFPOSX1 DFFPOSX1_3591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf1), .D(_138__6_), .Q(data_223__6_) );
DFFPOSX1 DFFPOSX1_3592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf1), .D(_138__7_), .Q(data_223__7_) );
DFFPOSX1 DFFPOSX1_3593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf1), .D(_138__8_), .Q(data_223__8_) );
DFFPOSX1 DFFPOSX1_3594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf1), .D(_138__9_), .Q(data_223__9_) );
DFFPOSX1 DFFPOSX1_3595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf1), .D(_138__10_), .Q(data_223__10_) );
DFFPOSX1 DFFPOSX1_3596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf1), .D(_138__11_), .Q(data_223__11_) );
DFFPOSX1 DFFPOSX1_3597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf1), .D(_138__12_), .Q(data_223__12_) );
DFFPOSX1 DFFPOSX1_3598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf1), .D(_138__13_), .Q(data_223__13_) );
DFFPOSX1 DFFPOSX1_3599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf1), .D(_138__14_), .Q(data_223__14_) );
DFFPOSX1 DFFPOSX1_3600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf1), .D(_138__15_), .Q(data_223__15_) );
DFFPOSX1 DFFPOSX1_3601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_139__0_), .Q(data_224__0_) );
DFFPOSX1 DFFPOSX1_3602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_139__1_), .Q(data_224__1_) );
DFFPOSX1 DFFPOSX1_3603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_139__2_), .Q(data_224__2_) );
DFFPOSX1 DFFPOSX1_3604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_139__3_), .Q(data_224__3_) );
DFFPOSX1 DFFPOSX1_3605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_139__4_), .Q(data_224__4_) );
DFFPOSX1 DFFPOSX1_3606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_139__5_), .Q(data_224__5_) );
DFFPOSX1 DFFPOSX1_3607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_139__6_), .Q(data_224__6_) );
DFFPOSX1 DFFPOSX1_3608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_139__7_), .Q(data_224__7_) );
DFFPOSX1 DFFPOSX1_3609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_139__8_), .Q(data_224__8_) );
DFFPOSX1 DFFPOSX1_3610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_139__9_), .Q(data_224__9_) );
DFFPOSX1 DFFPOSX1_3611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_139__10_), .Q(data_224__10_) );
DFFPOSX1 DFFPOSX1_3612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_139__11_), .Q(data_224__11_) );
DFFPOSX1 DFFPOSX1_3613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_139__12_), .Q(data_224__12_) );
DFFPOSX1 DFFPOSX1_3614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_139__13_), .Q(data_224__13_) );
DFFPOSX1 DFFPOSX1_3615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_139__14_), .Q(data_224__14_) );
DFFPOSX1 DFFPOSX1_3616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_139__15_), .Q(data_224__15_) );
DFFPOSX1 DFFPOSX1_3617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_140__0_), .Q(data_225__0_) );
DFFPOSX1 DFFPOSX1_3618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_140__1_), .Q(data_225__1_) );
DFFPOSX1 DFFPOSX1_3619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_140__2_), .Q(data_225__2_) );
DFFPOSX1 DFFPOSX1_3620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_140__3_), .Q(data_225__3_) );
DFFPOSX1 DFFPOSX1_3621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_140__4_), .Q(data_225__4_) );
DFFPOSX1 DFFPOSX1_3622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_140__5_), .Q(data_225__5_) );
DFFPOSX1 DFFPOSX1_3623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_140__6_), .Q(data_225__6_) );
DFFPOSX1 DFFPOSX1_3624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_140__7_), .Q(data_225__7_) );
DFFPOSX1 DFFPOSX1_3625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_140__8_), .Q(data_225__8_) );
DFFPOSX1 DFFPOSX1_3626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_140__9_), .Q(data_225__9_) );
DFFPOSX1 DFFPOSX1_3627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_140__10_), .Q(data_225__10_) );
DFFPOSX1 DFFPOSX1_3628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_140__11_), .Q(data_225__11_) );
DFFPOSX1 DFFPOSX1_3629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_140__12_), .Q(data_225__12_) );
DFFPOSX1 DFFPOSX1_3630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_140__13_), .Q(data_225__13_) );
DFFPOSX1 DFFPOSX1_3631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_140__14_), .Q(data_225__14_) );
DFFPOSX1 DFFPOSX1_3632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_140__15_), .Q(data_225__15_) );
DFFPOSX1 DFFPOSX1_3633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_141__0_), .Q(data_226__0_) );
DFFPOSX1 DFFPOSX1_3634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_141__1_), .Q(data_226__1_) );
DFFPOSX1 DFFPOSX1_3635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_141__2_), .Q(data_226__2_) );
DFFPOSX1 DFFPOSX1_3636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_141__3_), .Q(data_226__3_) );
DFFPOSX1 DFFPOSX1_3637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_141__4_), .Q(data_226__4_) );
DFFPOSX1 DFFPOSX1_3638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_141__5_), .Q(data_226__5_) );
DFFPOSX1 DFFPOSX1_3639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_141__6_), .Q(data_226__6_) );
DFFPOSX1 DFFPOSX1_3640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_141__7_), .Q(data_226__7_) );
DFFPOSX1 DFFPOSX1_3641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_141__8_), .Q(data_226__8_) );
DFFPOSX1 DFFPOSX1_3642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_141__9_), .Q(data_226__9_) );
DFFPOSX1 DFFPOSX1_3643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_141__10_), .Q(data_226__10_) );
DFFPOSX1 DFFPOSX1_3644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_141__11_), .Q(data_226__11_) );
DFFPOSX1 DFFPOSX1_3645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_141__12_), .Q(data_226__12_) );
DFFPOSX1 DFFPOSX1_3646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_141__13_), .Q(data_226__13_) );
DFFPOSX1 DFFPOSX1_3647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_141__14_), .Q(data_226__14_) );
DFFPOSX1 DFFPOSX1_3648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_141__15_), .Q(data_226__15_) );
DFFPOSX1 DFFPOSX1_3649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_142__0_), .Q(data_227__0_) );
DFFPOSX1 DFFPOSX1_3650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_142__1_), .Q(data_227__1_) );
DFFPOSX1 DFFPOSX1_3651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_142__2_), .Q(data_227__2_) );
DFFPOSX1 DFFPOSX1_3652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_142__3_), .Q(data_227__3_) );
DFFPOSX1 DFFPOSX1_3653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_142__4_), .Q(data_227__4_) );
DFFPOSX1 DFFPOSX1_3654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_142__5_), .Q(data_227__5_) );
DFFPOSX1 DFFPOSX1_3655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_142__6_), .Q(data_227__6_) );
DFFPOSX1 DFFPOSX1_3656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_142__7_), .Q(data_227__7_) );
DFFPOSX1 DFFPOSX1_3657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_142__8_), .Q(data_227__8_) );
DFFPOSX1 DFFPOSX1_3658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_142__9_), .Q(data_227__9_) );
DFFPOSX1 DFFPOSX1_3659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_142__10_), .Q(data_227__10_) );
DFFPOSX1 DFFPOSX1_3660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_142__11_), .Q(data_227__11_) );
DFFPOSX1 DFFPOSX1_3661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_142__12_), .Q(data_227__12_) );
DFFPOSX1 DFFPOSX1_3662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_142__13_), .Q(data_227__13_) );
DFFPOSX1 DFFPOSX1_3663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_142__14_), .Q(data_227__14_) );
DFFPOSX1 DFFPOSX1_3664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_142__15_), .Q(data_227__15_) );
DFFPOSX1 DFFPOSX1_3665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_143__0_), .Q(data_228__0_) );
DFFPOSX1 DFFPOSX1_3666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_143__1_), .Q(data_228__1_) );
DFFPOSX1 DFFPOSX1_3667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_143__2_), .Q(data_228__2_) );
DFFPOSX1 DFFPOSX1_3668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_143__3_), .Q(data_228__3_) );
DFFPOSX1 DFFPOSX1_3669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_143__4_), .Q(data_228__4_) );
DFFPOSX1 DFFPOSX1_3670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_143__5_), .Q(data_228__5_) );
DFFPOSX1 DFFPOSX1_3671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_143__6_), .Q(data_228__6_) );
DFFPOSX1 DFFPOSX1_3672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_143__7_), .Q(data_228__7_) );
DFFPOSX1 DFFPOSX1_3673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_143__8_), .Q(data_228__8_) );
DFFPOSX1 DFFPOSX1_3674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_143__9_), .Q(data_228__9_) );
DFFPOSX1 DFFPOSX1_3675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_143__10_), .Q(data_228__10_) );
DFFPOSX1 DFFPOSX1_3676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_143__11_), .Q(data_228__11_) );
DFFPOSX1 DFFPOSX1_3677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_143__12_), .Q(data_228__12_) );
DFFPOSX1 DFFPOSX1_3678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_143__13_), .Q(data_228__13_) );
DFFPOSX1 DFFPOSX1_3679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_143__14_), .Q(data_228__14_) );
DFFPOSX1 DFFPOSX1_3680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_143__15_), .Q(data_228__15_) );
DFFPOSX1 DFFPOSX1_3681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_144__0_), .Q(data_229__0_) );
DFFPOSX1 DFFPOSX1_3682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_144__1_), .Q(data_229__1_) );
DFFPOSX1 DFFPOSX1_3683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_144__2_), .Q(data_229__2_) );
DFFPOSX1 DFFPOSX1_3684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_144__3_), .Q(data_229__3_) );
DFFPOSX1 DFFPOSX1_3685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_144__4_), .Q(data_229__4_) );
DFFPOSX1 DFFPOSX1_3686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_144__5_), .Q(data_229__5_) );
DFFPOSX1 DFFPOSX1_3687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_144__6_), .Q(data_229__6_) );
DFFPOSX1 DFFPOSX1_3688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_144__7_), .Q(data_229__7_) );
DFFPOSX1 DFFPOSX1_3689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_144__8_), .Q(data_229__8_) );
DFFPOSX1 DFFPOSX1_3690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_144__9_), .Q(data_229__9_) );
DFFPOSX1 DFFPOSX1_3691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_144__10_), .Q(data_229__10_) );
DFFPOSX1 DFFPOSX1_3692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_144__11_), .Q(data_229__11_) );
DFFPOSX1 DFFPOSX1_3693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_144__12_), .Q(data_229__12_) );
DFFPOSX1 DFFPOSX1_3694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_144__13_), .Q(data_229__13_) );
DFFPOSX1 DFFPOSX1_3695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_144__14_), .Q(data_229__14_) );
DFFPOSX1 DFFPOSX1_3696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_144__15_), .Q(data_229__15_) );
DFFPOSX1 DFFPOSX1_3697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_146__0_), .Q(data_230__0_) );
DFFPOSX1 DFFPOSX1_3698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_146__1_), .Q(data_230__1_) );
DFFPOSX1 DFFPOSX1_3699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_146__2_), .Q(data_230__2_) );
DFFPOSX1 DFFPOSX1_3700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_146__3_), .Q(data_230__3_) );
DFFPOSX1 DFFPOSX1_3701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_146__4_), .Q(data_230__4_) );
DFFPOSX1 DFFPOSX1_3702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_146__5_), .Q(data_230__5_) );
DFFPOSX1 DFFPOSX1_3703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_146__6_), .Q(data_230__6_) );
DFFPOSX1 DFFPOSX1_3704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_146__7_), .Q(data_230__7_) );
DFFPOSX1 DFFPOSX1_3705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_146__8_), .Q(data_230__8_) );
DFFPOSX1 DFFPOSX1_3706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_146__9_), .Q(data_230__9_) );
DFFPOSX1 DFFPOSX1_3707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_146__10_), .Q(data_230__10_) );
DFFPOSX1 DFFPOSX1_3708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_146__11_), .Q(data_230__11_) );
DFFPOSX1 DFFPOSX1_3709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_146__12_), .Q(data_230__12_) );
DFFPOSX1 DFFPOSX1_3710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_146__13_), .Q(data_230__13_) );
DFFPOSX1 DFFPOSX1_3711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_146__14_), .Q(data_230__14_) );
DFFPOSX1 DFFPOSX1_3712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_146__15_), .Q(data_230__15_) );
DFFPOSX1 DFFPOSX1_3713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_147__0_), .Q(data_231__0_) );
DFFPOSX1 DFFPOSX1_3714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_147__1_), .Q(data_231__1_) );
DFFPOSX1 DFFPOSX1_3715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_147__2_), .Q(data_231__2_) );
DFFPOSX1 DFFPOSX1_3716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_147__3_), .Q(data_231__3_) );
DFFPOSX1 DFFPOSX1_3717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_147__4_), .Q(data_231__4_) );
DFFPOSX1 DFFPOSX1_3718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_147__5_), .Q(data_231__5_) );
DFFPOSX1 DFFPOSX1_3719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_147__6_), .Q(data_231__6_) );
DFFPOSX1 DFFPOSX1_3720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_147__7_), .Q(data_231__7_) );
DFFPOSX1 DFFPOSX1_3721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_147__8_), .Q(data_231__8_) );
DFFPOSX1 DFFPOSX1_3722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_147__9_), .Q(data_231__9_) );
DFFPOSX1 DFFPOSX1_3723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_147__10_), .Q(data_231__10_) );
DFFPOSX1 DFFPOSX1_3724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_147__11_), .Q(data_231__11_) );
DFFPOSX1 DFFPOSX1_3725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_147__12_), .Q(data_231__12_) );
DFFPOSX1 DFFPOSX1_3726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_147__13_), .Q(data_231__13_) );
DFFPOSX1 DFFPOSX1_3727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_147__14_), .Q(data_231__14_) );
DFFPOSX1 DFFPOSX1_3728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_147__15_), .Q(data_231__15_) );
DFFPOSX1 DFFPOSX1_3729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_148__0_), .Q(data_232__0_) );
DFFPOSX1 DFFPOSX1_3730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_148__1_), .Q(data_232__1_) );
DFFPOSX1 DFFPOSX1_3731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_148__2_), .Q(data_232__2_) );
DFFPOSX1 DFFPOSX1_3732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_148__3_), .Q(data_232__3_) );
DFFPOSX1 DFFPOSX1_3733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_148__4_), .Q(data_232__4_) );
DFFPOSX1 DFFPOSX1_3734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_148__5_), .Q(data_232__5_) );
DFFPOSX1 DFFPOSX1_3735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_148__6_), .Q(data_232__6_) );
DFFPOSX1 DFFPOSX1_3736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_148__7_), .Q(data_232__7_) );
DFFPOSX1 DFFPOSX1_3737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_148__8_), .Q(data_232__8_) );
DFFPOSX1 DFFPOSX1_3738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_148__9_), .Q(data_232__9_) );
DFFPOSX1 DFFPOSX1_3739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_148__10_), .Q(data_232__10_) );
DFFPOSX1 DFFPOSX1_3740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_148__11_), .Q(data_232__11_) );
DFFPOSX1 DFFPOSX1_3741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_148__12_), .Q(data_232__12_) );
DFFPOSX1 DFFPOSX1_3742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_148__13_), .Q(data_232__13_) );
DFFPOSX1 DFFPOSX1_3743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_148__14_), .Q(data_232__14_) );
DFFPOSX1 DFFPOSX1_3744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_148__15_), .Q(data_232__15_) );
DFFPOSX1 DFFPOSX1_3745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_149__0_), .Q(data_233__0_) );
DFFPOSX1 DFFPOSX1_3746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_149__1_), .Q(data_233__1_) );
DFFPOSX1 DFFPOSX1_3747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_149__2_), .Q(data_233__2_) );
DFFPOSX1 DFFPOSX1_3748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_149__3_), .Q(data_233__3_) );
DFFPOSX1 DFFPOSX1_3749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_149__4_), .Q(data_233__4_) );
DFFPOSX1 DFFPOSX1_3750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_149__5_), .Q(data_233__5_) );
DFFPOSX1 DFFPOSX1_3751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_149__6_), .Q(data_233__6_) );
DFFPOSX1 DFFPOSX1_3752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_149__7_), .Q(data_233__7_) );
DFFPOSX1 DFFPOSX1_3753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_149__8_), .Q(data_233__8_) );
DFFPOSX1 DFFPOSX1_3754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_149__9_), .Q(data_233__9_) );
DFFPOSX1 DFFPOSX1_3755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_149__10_), .Q(data_233__10_) );
DFFPOSX1 DFFPOSX1_3756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_149__11_), .Q(data_233__11_) );
DFFPOSX1 DFFPOSX1_3757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_149__12_), .Q(data_233__12_) );
DFFPOSX1 DFFPOSX1_3758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_149__13_), .Q(data_233__13_) );
DFFPOSX1 DFFPOSX1_3759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_149__14_), .Q(data_233__14_) );
DFFPOSX1 DFFPOSX1_3760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_149__15_), .Q(data_233__15_) );
DFFPOSX1 DFFPOSX1_3761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_150__0_), .Q(data_234__0_) );
DFFPOSX1 DFFPOSX1_3762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_150__1_), .Q(data_234__1_) );
DFFPOSX1 DFFPOSX1_3763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_150__2_), .Q(data_234__2_) );
DFFPOSX1 DFFPOSX1_3764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_150__3_), .Q(data_234__3_) );
DFFPOSX1 DFFPOSX1_3765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_150__4_), .Q(data_234__4_) );
DFFPOSX1 DFFPOSX1_3766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_150__5_), .Q(data_234__5_) );
DFFPOSX1 DFFPOSX1_3767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_150__6_), .Q(data_234__6_) );
DFFPOSX1 DFFPOSX1_3768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_150__7_), .Q(data_234__7_) );
DFFPOSX1 DFFPOSX1_3769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_150__8_), .Q(data_234__8_) );
DFFPOSX1 DFFPOSX1_3770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_150__9_), .Q(data_234__9_) );
DFFPOSX1 DFFPOSX1_3771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_150__10_), .Q(data_234__10_) );
DFFPOSX1 DFFPOSX1_3772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_150__11_), .Q(data_234__11_) );
DFFPOSX1 DFFPOSX1_3773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_150__12_), .Q(data_234__12_) );
DFFPOSX1 DFFPOSX1_3774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_150__13_), .Q(data_234__13_) );
DFFPOSX1 DFFPOSX1_3775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_150__14_), .Q(data_234__14_) );
DFFPOSX1 DFFPOSX1_3776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_150__15_), .Q(data_234__15_) );
DFFPOSX1 DFFPOSX1_3777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_151__0_), .Q(data_235__0_) );
DFFPOSX1 DFFPOSX1_3778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_151__1_), .Q(data_235__1_) );
DFFPOSX1 DFFPOSX1_3779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_151__2_), .Q(data_235__2_) );
DFFPOSX1 DFFPOSX1_3780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_151__3_), .Q(data_235__3_) );
DFFPOSX1 DFFPOSX1_3781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_151__4_), .Q(data_235__4_) );
DFFPOSX1 DFFPOSX1_3782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_151__5_), .Q(data_235__5_) );
DFFPOSX1 DFFPOSX1_3783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_151__6_), .Q(data_235__6_) );
DFFPOSX1 DFFPOSX1_3784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_151__7_), .Q(data_235__7_) );
DFFPOSX1 DFFPOSX1_3785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_151__8_), .Q(data_235__8_) );
DFFPOSX1 DFFPOSX1_3786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_151__9_), .Q(data_235__9_) );
DFFPOSX1 DFFPOSX1_3787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_151__10_), .Q(data_235__10_) );
DFFPOSX1 DFFPOSX1_3788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_151__11_), .Q(data_235__11_) );
DFFPOSX1 DFFPOSX1_3789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_151__12_), .Q(data_235__12_) );
DFFPOSX1 DFFPOSX1_3790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_151__13_), .Q(data_235__13_) );
DFFPOSX1 DFFPOSX1_3791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_151__14_), .Q(data_235__14_) );
DFFPOSX1 DFFPOSX1_3792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_151__15_), .Q(data_235__15_) );
DFFPOSX1 DFFPOSX1_3793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_152__0_), .Q(data_236__0_) );
DFFPOSX1 DFFPOSX1_3794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_152__1_), .Q(data_236__1_) );
DFFPOSX1 DFFPOSX1_3795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_152__2_), .Q(data_236__2_) );
DFFPOSX1 DFFPOSX1_3796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_152__3_), .Q(data_236__3_) );
DFFPOSX1 DFFPOSX1_3797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_152__4_), .Q(data_236__4_) );
DFFPOSX1 DFFPOSX1_3798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_152__5_), .Q(data_236__5_) );
DFFPOSX1 DFFPOSX1_3799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_152__6_), .Q(data_236__6_) );
DFFPOSX1 DFFPOSX1_3800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_152__7_), .Q(data_236__7_) );
DFFPOSX1 DFFPOSX1_3801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_152__8_), .Q(data_236__8_) );
DFFPOSX1 DFFPOSX1_3802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_152__9_), .Q(data_236__9_) );
DFFPOSX1 DFFPOSX1_3803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_152__10_), .Q(data_236__10_) );
DFFPOSX1 DFFPOSX1_3804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_152__11_), .Q(data_236__11_) );
DFFPOSX1 DFFPOSX1_3805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_152__12_), .Q(data_236__12_) );
DFFPOSX1 DFFPOSX1_3806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_152__13_), .Q(data_236__13_) );
DFFPOSX1 DFFPOSX1_3807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_152__14_), .Q(data_236__14_) );
DFFPOSX1 DFFPOSX1_3808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_152__15_), .Q(data_236__15_) );
DFFPOSX1 DFFPOSX1_3809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_153__0_), .Q(data_237__0_) );
DFFPOSX1 DFFPOSX1_3810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_153__1_), .Q(data_237__1_) );
DFFPOSX1 DFFPOSX1_3811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_153__2_), .Q(data_237__2_) );
DFFPOSX1 DFFPOSX1_3812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_153__3_), .Q(data_237__3_) );
DFFPOSX1 DFFPOSX1_3813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_153__4_), .Q(data_237__4_) );
DFFPOSX1 DFFPOSX1_3814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_153__5_), .Q(data_237__5_) );
DFFPOSX1 DFFPOSX1_3815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_153__6_), .Q(data_237__6_) );
DFFPOSX1 DFFPOSX1_3816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_153__7_), .Q(data_237__7_) );
DFFPOSX1 DFFPOSX1_3817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_153__8_), .Q(data_237__8_) );
DFFPOSX1 DFFPOSX1_3818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_153__9_), .Q(data_237__9_) );
DFFPOSX1 DFFPOSX1_3819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_153__10_), .Q(data_237__10_) );
DFFPOSX1 DFFPOSX1_3820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_153__11_), .Q(data_237__11_) );
DFFPOSX1 DFFPOSX1_3821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_153__12_), .Q(data_237__12_) );
DFFPOSX1 DFFPOSX1_3822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_153__13_), .Q(data_237__13_) );
DFFPOSX1 DFFPOSX1_3823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_153__14_), .Q(data_237__14_) );
DFFPOSX1 DFFPOSX1_3824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_153__15_), .Q(data_237__15_) );
DFFPOSX1 DFFPOSX1_3825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_154__0_), .Q(data_238__0_) );
DFFPOSX1 DFFPOSX1_3826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_154__1_), .Q(data_238__1_) );
DFFPOSX1 DFFPOSX1_3827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_154__2_), .Q(data_238__2_) );
DFFPOSX1 DFFPOSX1_3828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_154__3_), .Q(data_238__3_) );
DFFPOSX1 DFFPOSX1_3829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_154__4_), .Q(data_238__4_) );
DFFPOSX1 DFFPOSX1_3830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_154__5_), .Q(data_238__5_) );
DFFPOSX1 DFFPOSX1_3831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_154__6_), .Q(data_238__6_) );
DFFPOSX1 DFFPOSX1_3832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_154__7_), .Q(data_238__7_) );
DFFPOSX1 DFFPOSX1_3833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_154__8_), .Q(data_238__8_) );
DFFPOSX1 DFFPOSX1_3834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_154__9_), .Q(data_238__9_) );
DFFPOSX1 DFFPOSX1_3835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_154__10_), .Q(data_238__10_) );
DFFPOSX1 DFFPOSX1_3836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_154__11_), .Q(data_238__11_) );
DFFPOSX1 DFFPOSX1_3837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_154__12_), .Q(data_238__12_) );
DFFPOSX1 DFFPOSX1_3838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_154__13_), .Q(data_238__13_) );
DFFPOSX1 DFFPOSX1_3839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_154__14_), .Q(data_238__14_) );
DFFPOSX1 DFFPOSX1_3840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_154__15_), .Q(data_238__15_) );
DFFPOSX1 DFFPOSX1_3841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf0), .D(_155__0_), .Q(data_239__0_) );
DFFPOSX1 DFFPOSX1_3842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf0), .D(_155__1_), .Q(data_239__1_) );
DFFPOSX1 DFFPOSX1_3843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf0), .D(_155__2_), .Q(data_239__2_) );
DFFPOSX1 DFFPOSX1_3844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf0), .D(_155__3_), .Q(data_239__3_) );
DFFPOSX1 DFFPOSX1_3845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf0), .D(_155__4_), .Q(data_239__4_) );
DFFPOSX1 DFFPOSX1_3846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf0), .D(_155__5_), .Q(data_239__5_) );
DFFPOSX1 DFFPOSX1_3847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf0), .D(_155__6_), .Q(data_239__6_) );
DFFPOSX1 DFFPOSX1_3848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf0), .D(_155__7_), .Q(data_239__7_) );
DFFPOSX1 DFFPOSX1_3849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf0), .D(_155__8_), .Q(data_239__8_) );
DFFPOSX1 DFFPOSX1_3850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf0), .D(_155__9_), .Q(data_239__9_) );
DFFPOSX1 DFFPOSX1_3851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf0), .D(_155__10_), .Q(data_239__10_) );
DFFPOSX1 DFFPOSX1_3852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf0), .D(_155__11_), .Q(data_239__11_) );
DFFPOSX1 DFFPOSX1_3853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf0), .D(_155__12_), .Q(data_239__12_) );
DFFPOSX1 DFFPOSX1_3854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf0), .D(_155__13_), .Q(data_239__13_) );
DFFPOSX1 DFFPOSX1_3855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf0), .D(_155__14_), .Q(data_239__14_) );
DFFPOSX1 DFFPOSX1_3856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf0), .D(_155__15_), .Q(data_239__15_) );
DFFPOSX1 DFFPOSX1_3857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf239), .D(_157__0_), .Q(data_240__0_) );
DFFPOSX1 DFFPOSX1_3858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf238), .D(_157__1_), .Q(data_240__1_) );
DFFPOSX1 DFFPOSX1_3859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf237), .D(_157__2_), .Q(data_240__2_) );
DFFPOSX1 DFFPOSX1_3860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf236), .D(_157__3_), .Q(data_240__3_) );
DFFPOSX1 DFFPOSX1_3861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf235), .D(_157__4_), .Q(data_240__4_) );
DFFPOSX1 DFFPOSX1_3862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf234), .D(_157__5_), .Q(data_240__5_) );
DFFPOSX1 DFFPOSX1_3863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf233), .D(_157__6_), .Q(data_240__6_) );
DFFPOSX1 DFFPOSX1_3864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf232), .D(_157__7_), .Q(data_240__7_) );
DFFPOSX1 DFFPOSX1_3865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf231), .D(_157__8_), .Q(data_240__8_) );
DFFPOSX1 DFFPOSX1_3866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf230), .D(_157__9_), .Q(data_240__9_) );
DFFPOSX1 DFFPOSX1_3867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf229), .D(_157__10_), .Q(data_240__10_) );
DFFPOSX1 DFFPOSX1_3868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf228), .D(_157__11_), .Q(data_240__11_) );
DFFPOSX1 DFFPOSX1_3869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf227), .D(_157__12_), .Q(data_240__12_) );
DFFPOSX1 DFFPOSX1_3870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf226), .D(_157__13_), .Q(data_240__13_) );
DFFPOSX1 DFFPOSX1_3871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf225), .D(_157__14_), .Q(data_240__14_) );
DFFPOSX1 DFFPOSX1_3872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf224), .D(_157__15_), .Q(data_240__15_) );
DFFPOSX1 DFFPOSX1_3873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf223), .D(_158__0_), .Q(data_241__0_) );
DFFPOSX1 DFFPOSX1_3874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf222), .D(_158__1_), .Q(data_241__1_) );
DFFPOSX1 DFFPOSX1_3875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf221), .D(_158__2_), .Q(data_241__2_) );
DFFPOSX1 DFFPOSX1_3876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf220), .D(_158__3_), .Q(data_241__3_) );
DFFPOSX1 DFFPOSX1_3877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf219), .D(_158__4_), .Q(data_241__4_) );
DFFPOSX1 DFFPOSX1_3878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf218), .D(_158__5_), .Q(data_241__5_) );
DFFPOSX1 DFFPOSX1_3879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf217), .D(_158__6_), .Q(data_241__6_) );
DFFPOSX1 DFFPOSX1_3880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf216), .D(_158__7_), .Q(data_241__7_) );
DFFPOSX1 DFFPOSX1_3881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf215), .D(_158__8_), .Q(data_241__8_) );
DFFPOSX1 DFFPOSX1_3882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf214), .D(_158__9_), .Q(data_241__9_) );
DFFPOSX1 DFFPOSX1_3883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf213), .D(_158__10_), .Q(data_241__10_) );
DFFPOSX1 DFFPOSX1_3884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf212), .D(_158__11_), .Q(data_241__11_) );
DFFPOSX1 DFFPOSX1_3885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf211), .D(_158__12_), .Q(data_241__12_) );
DFFPOSX1 DFFPOSX1_3886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf210), .D(_158__13_), .Q(data_241__13_) );
DFFPOSX1 DFFPOSX1_3887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf209), .D(_158__14_), .Q(data_241__14_) );
DFFPOSX1 DFFPOSX1_3888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf208), .D(_158__15_), .Q(data_241__15_) );
DFFPOSX1 DFFPOSX1_3889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf207), .D(_159__0_), .Q(data_242__0_) );
DFFPOSX1 DFFPOSX1_3890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf206), .D(_159__1_), .Q(data_242__1_) );
DFFPOSX1 DFFPOSX1_3891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf205), .D(_159__2_), .Q(data_242__2_) );
DFFPOSX1 DFFPOSX1_3892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf204), .D(_159__3_), .Q(data_242__3_) );
DFFPOSX1 DFFPOSX1_3893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf203), .D(_159__4_), .Q(data_242__4_) );
DFFPOSX1 DFFPOSX1_3894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf202), .D(_159__5_), .Q(data_242__5_) );
DFFPOSX1 DFFPOSX1_3895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf201), .D(_159__6_), .Q(data_242__6_) );
DFFPOSX1 DFFPOSX1_3896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf200), .D(_159__7_), .Q(data_242__7_) );
DFFPOSX1 DFFPOSX1_3897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf199), .D(_159__8_), .Q(data_242__8_) );
DFFPOSX1 DFFPOSX1_3898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf198), .D(_159__9_), .Q(data_242__9_) );
DFFPOSX1 DFFPOSX1_3899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf197), .D(_159__10_), .Q(data_242__10_) );
DFFPOSX1 DFFPOSX1_3900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf196), .D(_159__11_), .Q(data_242__11_) );
DFFPOSX1 DFFPOSX1_3901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf195), .D(_159__12_), .Q(data_242__12_) );
DFFPOSX1 DFFPOSX1_3902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf194), .D(_159__13_), .Q(data_242__13_) );
DFFPOSX1 DFFPOSX1_3903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf193), .D(_159__14_), .Q(data_242__14_) );
DFFPOSX1 DFFPOSX1_3904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf192), .D(_159__15_), .Q(data_242__15_) );
DFFPOSX1 DFFPOSX1_3905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf191), .D(_160__0_), .Q(data_243__0_) );
DFFPOSX1 DFFPOSX1_3906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf190), .D(_160__1_), .Q(data_243__1_) );
DFFPOSX1 DFFPOSX1_3907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf189), .D(_160__2_), .Q(data_243__2_) );
DFFPOSX1 DFFPOSX1_3908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf188), .D(_160__3_), .Q(data_243__3_) );
DFFPOSX1 DFFPOSX1_3909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf187), .D(_160__4_), .Q(data_243__4_) );
DFFPOSX1 DFFPOSX1_3910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf186), .D(_160__5_), .Q(data_243__5_) );
DFFPOSX1 DFFPOSX1_3911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf185), .D(_160__6_), .Q(data_243__6_) );
DFFPOSX1 DFFPOSX1_3912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf184), .D(_160__7_), .Q(data_243__7_) );
DFFPOSX1 DFFPOSX1_3913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf183), .D(_160__8_), .Q(data_243__8_) );
DFFPOSX1 DFFPOSX1_3914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf182), .D(_160__9_), .Q(data_243__9_) );
DFFPOSX1 DFFPOSX1_3915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf181), .D(_160__10_), .Q(data_243__10_) );
DFFPOSX1 DFFPOSX1_3916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf180), .D(_160__11_), .Q(data_243__11_) );
DFFPOSX1 DFFPOSX1_3917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf179), .D(_160__12_), .Q(data_243__12_) );
DFFPOSX1 DFFPOSX1_3918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf178), .D(_160__13_), .Q(data_243__13_) );
DFFPOSX1 DFFPOSX1_3919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf177), .D(_160__14_), .Q(data_243__14_) );
DFFPOSX1 DFFPOSX1_3920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf176), .D(_160__15_), .Q(data_243__15_) );
DFFPOSX1 DFFPOSX1_3921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf175), .D(_161__0_), .Q(data_244__0_) );
DFFPOSX1 DFFPOSX1_3922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf174), .D(_161__1_), .Q(data_244__1_) );
DFFPOSX1 DFFPOSX1_3923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf173), .D(_161__2_), .Q(data_244__2_) );
DFFPOSX1 DFFPOSX1_3924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf172), .D(_161__3_), .Q(data_244__3_) );
DFFPOSX1 DFFPOSX1_3925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf171), .D(_161__4_), .Q(data_244__4_) );
DFFPOSX1 DFFPOSX1_3926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf170), .D(_161__5_), .Q(data_244__5_) );
DFFPOSX1 DFFPOSX1_3927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf169), .D(_161__6_), .Q(data_244__6_) );
DFFPOSX1 DFFPOSX1_3928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf168), .D(_161__7_), .Q(data_244__7_) );
DFFPOSX1 DFFPOSX1_3929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf167), .D(_161__8_), .Q(data_244__8_) );
DFFPOSX1 DFFPOSX1_3930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf166), .D(_161__9_), .Q(data_244__9_) );
DFFPOSX1 DFFPOSX1_3931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf165), .D(_161__10_), .Q(data_244__10_) );
DFFPOSX1 DFFPOSX1_3932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf164), .D(_161__11_), .Q(data_244__11_) );
DFFPOSX1 DFFPOSX1_3933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf163), .D(_161__12_), .Q(data_244__12_) );
DFFPOSX1 DFFPOSX1_3934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf162), .D(_161__13_), .Q(data_244__13_) );
DFFPOSX1 DFFPOSX1_3935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf161), .D(_161__14_), .Q(data_244__14_) );
DFFPOSX1 DFFPOSX1_3936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf160), .D(_161__15_), .Q(data_244__15_) );
DFFPOSX1 DFFPOSX1_3937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf159), .D(_162__0_), .Q(data_245__0_) );
DFFPOSX1 DFFPOSX1_3938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf158), .D(_162__1_), .Q(data_245__1_) );
DFFPOSX1 DFFPOSX1_3939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf157), .D(_162__2_), .Q(data_245__2_) );
DFFPOSX1 DFFPOSX1_3940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf156), .D(_162__3_), .Q(data_245__3_) );
DFFPOSX1 DFFPOSX1_3941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf155), .D(_162__4_), .Q(data_245__4_) );
DFFPOSX1 DFFPOSX1_3942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf154), .D(_162__5_), .Q(data_245__5_) );
DFFPOSX1 DFFPOSX1_3943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf153), .D(_162__6_), .Q(data_245__6_) );
DFFPOSX1 DFFPOSX1_3944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf152), .D(_162__7_), .Q(data_245__7_) );
DFFPOSX1 DFFPOSX1_3945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf151), .D(_162__8_), .Q(data_245__8_) );
DFFPOSX1 DFFPOSX1_3946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf150), .D(_162__9_), .Q(data_245__9_) );
DFFPOSX1 DFFPOSX1_3947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf149), .D(_162__10_), .Q(data_245__10_) );
DFFPOSX1 DFFPOSX1_3948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf148), .D(_162__11_), .Q(data_245__11_) );
DFFPOSX1 DFFPOSX1_3949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf147), .D(_162__12_), .Q(data_245__12_) );
DFFPOSX1 DFFPOSX1_3950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf146), .D(_162__13_), .Q(data_245__13_) );
DFFPOSX1 DFFPOSX1_3951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf145), .D(_162__14_), .Q(data_245__14_) );
DFFPOSX1 DFFPOSX1_3952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf144), .D(_162__15_), .Q(data_245__15_) );
DFFPOSX1 DFFPOSX1_3953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf143), .D(_163__0_), .Q(data_246__0_) );
DFFPOSX1 DFFPOSX1_3954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf142), .D(_163__1_), .Q(data_246__1_) );
DFFPOSX1 DFFPOSX1_3955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf141), .D(_163__2_), .Q(data_246__2_) );
DFFPOSX1 DFFPOSX1_3956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf140), .D(_163__3_), .Q(data_246__3_) );
DFFPOSX1 DFFPOSX1_3957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf139), .D(_163__4_), .Q(data_246__4_) );
DFFPOSX1 DFFPOSX1_3958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf138), .D(_163__5_), .Q(data_246__5_) );
DFFPOSX1 DFFPOSX1_3959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf137), .D(_163__6_), .Q(data_246__6_) );
DFFPOSX1 DFFPOSX1_3960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf136), .D(_163__7_), .Q(data_246__7_) );
DFFPOSX1 DFFPOSX1_3961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf135), .D(_163__8_), .Q(data_246__8_) );
DFFPOSX1 DFFPOSX1_3962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf134), .D(_163__9_), .Q(data_246__9_) );
DFFPOSX1 DFFPOSX1_3963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf133), .D(_163__10_), .Q(data_246__10_) );
DFFPOSX1 DFFPOSX1_3964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf132), .D(_163__11_), .Q(data_246__11_) );
DFFPOSX1 DFFPOSX1_3965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf131), .D(_163__12_), .Q(data_246__12_) );
DFFPOSX1 DFFPOSX1_3966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf130), .D(_163__13_), .Q(data_246__13_) );
DFFPOSX1 DFFPOSX1_3967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf129), .D(_163__14_), .Q(data_246__14_) );
DFFPOSX1 DFFPOSX1_3968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf128), .D(_163__15_), .Q(data_246__15_) );
DFFPOSX1 DFFPOSX1_3969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf127), .D(_164__0_), .Q(data_247__0_) );
DFFPOSX1 DFFPOSX1_3970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf126), .D(_164__1_), .Q(data_247__1_) );
DFFPOSX1 DFFPOSX1_3971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf125), .D(_164__2_), .Q(data_247__2_) );
DFFPOSX1 DFFPOSX1_3972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf124), .D(_164__3_), .Q(data_247__3_) );
DFFPOSX1 DFFPOSX1_3973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf123), .D(_164__4_), .Q(data_247__4_) );
DFFPOSX1 DFFPOSX1_3974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf122), .D(_164__5_), .Q(data_247__5_) );
DFFPOSX1 DFFPOSX1_3975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf121), .D(_164__6_), .Q(data_247__6_) );
DFFPOSX1 DFFPOSX1_3976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf120), .D(_164__7_), .Q(data_247__7_) );
DFFPOSX1 DFFPOSX1_3977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf119), .D(_164__8_), .Q(data_247__8_) );
DFFPOSX1 DFFPOSX1_3978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf118), .D(_164__9_), .Q(data_247__9_) );
DFFPOSX1 DFFPOSX1_3979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf117), .D(_164__10_), .Q(data_247__10_) );
DFFPOSX1 DFFPOSX1_3980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf116), .D(_164__11_), .Q(data_247__11_) );
DFFPOSX1 DFFPOSX1_3981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf115), .D(_164__12_), .Q(data_247__12_) );
DFFPOSX1 DFFPOSX1_3982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf114), .D(_164__13_), .Q(data_247__13_) );
DFFPOSX1 DFFPOSX1_3983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf113), .D(_164__14_), .Q(data_247__14_) );
DFFPOSX1 DFFPOSX1_3984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf112), .D(_164__15_), .Q(data_247__15_) );
DFFPOSX1 DFFPOSX1_3985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf111), .D(_165__0_), .Q(data_248__0_) );
DFFPOSX1 DFFPOSX1_3986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf110), .D(_165__1_), .Q(data_248__1_) );
DFFPOSX1 DFFPOSX1_3987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf109), .D(_165__2_), .Q(data_248__2_) );
DFFPOSX1 DFFPOSX1_3988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf108), .D(_165__3_), .Q(data_248__3_) );
DFFPOSX1 DFFPOSX1_3989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf107), .D(_165__4_), .Q(data_248__4_) );
DFFPOSX1 DFFPOSX1_3990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf106), .D(_165__5_), .Q(data_248__5_) );
DFFPOSX1 DFFPOSX1_3991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf105), .D(_165__6_), .Q(data_248__6_) );
DFFPOSX1 DFFPOSX1_3992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf104), .D(_165__7_), .Q(data_248__7_) );
DFFPOSX1 DFFPOSX1_3993 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf103), .D(_165__8_), .Q(data_248__8_) );
DFFPOSX1 DFFPOSX1_3994 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf102), .D(_165__9_), .Q(data_248__9_) );
DFFPOSX1 DFFPOSX1_3995 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf101), .D(_165__10_), .Q(data_248__10_) );
DFFPOSX1 DFFPOSX1_3996 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf100), .D(_165__11_), .Q(data_248__11_) );
DFFPOSX1 DFFPOSX1_3997 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf99), .D(_165__12_), .Q(data_248__12_) );
DFFPOSX1 DFFPOSX1_3998 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_165__13_), .Q(data_248__13_) );
DFFPOSX1 DFFPOSX1_3999 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_165__14_), .Q(data_248__14_) );
DFFPOSX1 DFFPOSX1_4000 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_165__15_), .Q(data_248__15_) );
DFFPOSX1 DFFPOSX1_4001 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_166__0_), .Q(data_249__0_) );
DFFPOSX1 DFFPOSX1_4002 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_166__1_), .Q(data_249__1_) );
DFFPOSX1 DFFPOSX1_4003 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_166__2_), .Q(data_249__2_) );
DFFPOSX1 DFFPOSX1_4004 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_166__3_), .Q(data_249__3_) );
DFFPOSX1 DFFPOSX1_4005 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_166__4_), .Q(data_249__4_) );
DFFPOSX1 DFFPOSX1_4006 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_166__5_), .Q(data_249__5_) );
DFFPOSX1 DFFPOSX1_4007 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_166__6_), .Q(data_249__6_) );
DFFPOSX1 DFFPOSX1_4008 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_166__7_), .Q(data_249__7_) );
DFFPOSX1 DFFPOSX1_4009 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_166__8_), .Q(data_249__8_) );
DFFPOSX1 DFFPOSX1_4010 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_166__9_), .Q(data_249__9_) );
DFFPOSX1 DFFPOSX1_4011 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_166__10_), .Q(data_249__10_) );
DFFPOSX1 DFFPOSX1_4012 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_166__11_), .Q(data_249__11_) );
DFFPOSX1 DFFPOSX1_4013 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_166__12_), .Q(data_249__12_) );
DFFPOSX1 DFFPOSX1_4014 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_166__13_), .Q(data_249__13_) );
DFFPOSX1 DFFPOSX1_4015 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_166__14_), .Q(data_249__14_) );
DFFPOSX1 DFFPOSX1_4016 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_166__15_), .Q(data_249__15_) );
DFFPOSX1 DFFPOSX1_4017 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_168__0_), .Q(data_250__0_) );
DFFPOSX1 DFFPOSX1_4018 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_168__1_), .Q(data_250__1_) );
DFFPOSX1 DFFPOSX1_4019 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_168__2_), .Q(data_250__2_) );
DFFPOSX1 DFFPOSX1_4020 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_168__3_), .Q(data_250__3_) );
DFFPOSX1 DFFPOSX1_4021 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_168__4_), .Q(data_250__4_) );
DFFPOSX1 DFFPOSX1_4022 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_168__5_), .Q(data_250__5_) );
DFFPOSX1 DFFPOSX1_4023 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_168__6_), .Q(data_250__6_) );
DFFPOSX1 DFFPOSX1_4024 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_168__7_), .Q(data_250__7_) );
DFFPOSX1 DFFPOSX1_4025 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_168__8_), .Q(data_250__8_) );
DFFPOSX1 DFFPOSX1_4026 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_168__9_), .Q(data_250__9_) );
DFFPOSX1 DFFPOSX1_4027 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_168__10_), .Q(data_250__10_) );
DFFPOSX1 DFFPOSX1_4028 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_168__11_), .Q(data_250__11_) );
DFFPOSX1 DFFPOSX1_4029 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_168__12_), .Q(data_250__12_) );
DFFPOSX1 DFFPOSX1_4030 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_168__13_), .Q(data_250__13_) );
DFFPOSX1 DFFPOSX1_4031 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_168__14_), .Q(data_250__14_) );
DFFPOSX1 DFFPOSX1_4032 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_168__15_), .Q(data_250__15_) );
DFFPOSX1 DFFPOSX1_4033 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_169__0_), .Q(data_251__0_) );
DFFPOSX1 DFFPOSX1_4034 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_169__1_), .Q(data_251__1_) );
DFFPOSX1 DFFPOSX1_4035 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_169__2_), .Q(data_251__2_) );
DFFPOSX1 DFFPOSX1_4036 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_169__3_), .Q(data_251__3_) );
DFFPOSX1 DFFPOSX1_4037 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_169__4_), .Q(data_251__4_) );
DFFPOSX1 DFFPOSX1_4038 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_169__5_), .Q(data_251__5_) );
DFFPOSX1 DFFPOSX1_4039 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_169__6_), .Q(data_251__6_) );
DFFPOSX1 DFFPOSX1_4040 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_169__7_), .Q(data_251__7_) );
DFFPOSX1 DFFPOSX1_4041 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_169__8_), .Q(data_251__8_) );
DFFPOSX1 DFFPOSX1_4042 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_169__9_), .Q(data_251__9_) );
DFFPOSX1 DFFPOSX1_4043 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_169__10_), .Q(data_251__10_) );
DFFPOSX1 DFFPOSX1_4044 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_169__11_), .Q(data_251__11_) );
DFFPOSX1 DFFPOSX1_4045 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_169__12_), .Q(data_251__12_) );
DFFPOSX1 DFFPOSX1_4046 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_169__13_), .Q(data_251__13_) );
DFFPOSX1 DFFPOSX1_4047 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_169__14_), .Q(data_251__14_) );
DFFPOSX1 DFFPOSX1_4048 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_169__15_), .Q(data_251__15_) );
DFFPOSX1 DFFPOSX1_4049 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_170__0_), .Q(data_252__0_) );
DFFPOSX1 DFFPOSX1_4050 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_170__1_), .Q(data_252__1_) );
DFFPOSX1 DFFPOSX1_4051 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_170__2_), .Q(data_252__2_) );
DFFPOSX1 DFFPOSX1_4052 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_170__3_), .Q(data_252__3_) );
DFFPOSX1 DFFPOSX1_4053 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_170__4_), .Q(data_252__4_) );
DFFPOSX1 DFFPOSX1_4054 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_170__5_), .Q(data_252__5_) );
DFFPOSX1 DFFPOSX1_4055 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_170__6_), .Q(data_252__6_) );
DFFPOSX1 DFFPOSX1_4056 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_170__7_), .Q(data_252__7_) );
DFFPOSX1 DFFPOSX1_4057 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_170__8_), .Q(data_252__8_) );
DFFPOSX1 DFFPOSX1_4058 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_170__9_), .Q(data_252__9_) );
DFFPOSX1 DFFPOSX1_4059 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_170__10_), .Q(data_252__10_) );
DFFPOSX1 DFFPOSX1_4060 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_170__11_), .Q(data_252__11_) );
DFFPOSX1 DFFPOSX1_4061 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_170__12_), .Q(data_252__12_) );
DFFPOSX1 DFFPOSX1_4062 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_170__13_), .Q(data_252__13_) );
DFFPOSX1 DFFPOSX1_4063 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_170__14_), .Q(data_252__14_) );
DFFPOSX1 DFFPOSX1_4064 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_170__15_), .Q(data_252__15_) );
DFFPOSX1 DFFPOSX1_4065 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_171__0_), .Q(data_253__0_) );
DFFPOSX1 DFFPOSX1_4066 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_171__1_), .Q(data_253__1_) );
DFFPOSX1 DFFPOSX1_4067 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_171__2_), .Q(data_253__2_) );
DFFPOSX1 DFFPOSX1_4068 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_171__3_), .Q(data_253__3_) );
DFFPOSX1 DFFPOSX1_4069 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_171__4_), .Q(data_253__4_) );
DFFPOSX1 DFFPOSX1_4070 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_171__5_), .Q(data_253__5_) );
DFFPOSX1 DFFPOSX1_4071 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_171__6_), .Q(data_253__6_) );
DFFPOSX1 DFFPOSX1_4072 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_171__7_), .Q(data_253__7_) );
DFFPOSX1 DFFPOSX1_4073 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_171__8_), .Q(data_253__8_) );
DFFPOSX1 DFFPOSX1_4074 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_171__9_), .Q(data_253__9_) );
DFFPOSX1 DFFPOSX1_4075 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_171__10_), .Q(data_253__10_) );
DFFPOSX1 DFFPOSX1_4076 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_171__11_), .Q(data_253__11_) );
DFFPOSX1 DFFPOSX1_4077 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_171__12_), .Q(data_253__12_) );
DFFPOSX1 DFFPOSX1_4078 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_171__13_), .Q(data_253__13_) );
DFFPOSX1 DFFPOSX1_4079 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_171__14_), .Q(data_253__14_) );
DFFPOSX1 DFFPOSX1_4080 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_171__15_), .Q(data_253__15_) );
DFFPOSX1 DFFPOSX1_4081 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_172__0_), .Q(data_254__0_) );
DFFPOSX1 DFFPOSX1_4082 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_172__1_), .Q(data_254__1_) );
DFFPOSX1 DFFPOSX1_4083 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_172__2_), .Q(data_254__2_) );
DFFPOSX1 DFFPOSX1_4084 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_172__3_), .Q(data_254__3_) );
DFFPOSX1 DFFPOSX1_4085 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_172__4_), .Q(data_254__4_) );
DFFPOSX1 DFFPOSX1_4086 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_172__5_), .Q(data_254__5_) );
DFFPOSX1 DFFPOSX1_4087 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_172__6_), .Q(data_254__6_) );
DFFPOSX1 DFFPOSX1_4088 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_172__7_), .Q(data_254__7_) );
DFFPOSX1 DFFPOSX1_4089 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_172__8_), .Q(data_254__8_) );
DFFPOSX1 DFFPOSX1_4090 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_172__9_), .Q(data_254__9_) );
DFFPOSX1 DFFPOSX1_4091 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_172__10_), .Q(data_254__10_) );
DFFPOSX1 DFFPOSX1_4092 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_172__11_), .Q(data_254__11_) );
DFFPOSX1 DFFPOSX1_4093 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_172__12_), .Q(data_254__12_) );
DFFPOSX1 DFFPOSX1_4094 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_172__13_), .Q(data_254__13_) );
DFFPOSX1 DFFPOSX1_4095 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_172__14_), .Q(data_254__14_) );
DFFPOSX1 DFFPOSX1_4096 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_172__15_), .Q(data_254__15_) );
DFFPOSX1 DFFPOSX1_4097 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf255_bF_buf3), .D(_173__0_), .Q(data_255__0_) );
DFFPOSX1 DFFPOSX1_4098 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf254_bF_buf3), .D(_173__1_), .Q(data_255__1_) );
DFFPOSX1 DFFPOSX1_4099 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf253_bF_buf3), .D(_173__2_), .Q(data_255__2_) );
DFFPOSX1 DFFPOSX1_4100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf252_bF_buf3), .D(_173__3_), .Q(data_255__3_) );
DFFPOSX1 DFFPOSX1_4101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf251_bF_buf3), .D(_173__4_), .Q(data_255__4_) );
DFFPOSX1 DFFPOSX1_4102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf250_bF_buf3), .D(_173__5_), .Q(data_255__5_) );
DFFPOSX1 DFFPOSX1_4103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf249_bF_buf3), .D(_173__6_), .Q(data_255__6_) );
DFFPOSX1 DFFPOSX1_4104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf248_bF_buf3), .D(_173__7_), .Q(data_255__7_) );
DFFPOSX1 DFFPOSX1_4105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf247_bF_buf3), .D(_173__8_), .Q(data_255__8_) );
DFFPOSX1 DFFPOSX1_4106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf246_bF_buf3), .D(_173__9_), .Q(data_255__9_) );
DFFPOSX1 DFFPOSX1_4107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf245_bF_buf3), .D(_173__10_), .Q(data_255__10_) );
DFFPOSX1 DFFPOSX1_4108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf244_bF_buf3), .D(_173__11_), .Q(data_255__11_) );
DFFPOSX1 DFFPOSX1_4109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf243_bF_buf3), .D(_173__12_), .Q(data_255__12_) );
DFFPOSX1 DFFPOSX1_4110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf242_bF_buf3), .D(_173__13_), .Q(data_255__13_) );
DFFPOSX1 DFFPOSX1_4111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf241_bF_buf3), .D(_173__14_), .Q(data_255__14_) );
DFFPOSX1 DFFPOSX1_4112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf240_bF_buf3), .D(_173__15_), .Q(data_255__15_) );
endmodule
