module NRISC_UP (IDATA_CORE_out, DDATA_CORE_out, CORE_ctrl, INTERRUPT_ch, INTERRUPT_flag, clk, rst, IDATA_CORE_addr, IDATA_CORE_clk, DDATA_CORE_addr, DDATA_CORE_in, DDATA_CORE_load, DDATA_CORE_write, DDATA_CORE_ctrl);

input INTERRUPT_flag;
input clk;
input rst;
output IDATA_CORE_clk;
output DDATA_CORE_load;
output DDATA_CORE_write;
input [31:0] IDATA_CORE_out;
input [31:0] DDATA_CORE_out;
input [2:0] CORE_ctrl;
input [7:0] INTERRUPT_ch;
output [7:0] IDATA_CORE_addr;
output [7:0] DDATA_CORE_addr;
output [31:0] DDATA_CORE_in;
output [2:0] DDATA_CORE_ctrl;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX2 BUFX2_2 ( .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX2 BUFX2_3 ( .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX2 BUFX2_4 ( .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX2 BUFX2_5 ( .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX2 BUFX2_6 ( .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX2 BUFX2_7 ( .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX2 BUFX2_8 ( .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX2 BUFX2_9 ( .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX2 BUFX2_10 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf10_bF_buf3) );
BUFX2 BUFX2_11 ( .A(INTERRUPT_flag_bF_buf6), .Y(INTERRUPT_flag_bF_buf10_bF_buf2) );
BUFX2 BUFX2_12 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf10_bF_buf1) );
BUFX2 BUFX2_13 ( .A(INTERRUPT_flag_bF_buf3), .Y(INTERRUPT_flag_bF_buf10_bF_buf0) );
BUFX2 BUFX2_14 ( .A(INTERRUPT_flag_bF_buf2), .Y(INTERRUPT_flag_bF_buf11_bF_buf3) );
BUFX2 BUFX2_15 ( .A(INTERRUPT_flag_bF_buf5), .Y(INTERRUPT_flag_bF_buf11_bF_buf2) );
BUFX2 BUFX2_16 ( .A(INTERRUPT_flag_bF_buf1), .Y(INTERRUPT_flag_bF_buf11_bF_buf1) );
BUFX2 BUFX2_17 ( .A(INTERRUPT_flag_bF_buf14), .Y(INTERRUPT_flag_bF_buf11_bF_buf0) );
BUFX2 BUFX2_18 ( .A(INTERRUPT_flag_bF_buf3), .Y(INTERRUPT_flag_bF_buf12_bF_buf3) );
BUFX2 BUFX2_19 ( .A(INTERRUPT_flag_bF_buf1), .Y(INTERRUPT_flag_bF_buf12_bF_buf2) );
BUFX2 BUFX2_20 ( .A(INTERRUPT_flag_bF_buf9), .Y(INTERRUPT_flag_bF_buf12_bF_buf1) );
BUFX2 BUFX2_21 ( .A(INTERRUPT_flag_bF_buf2), .Y(INTERRUPT_flag_bF_buf12_bF_buf0) );
BUFX2 BUFX2_22 ( .A(INTERRUPT_flag_bF_buf2), .Y(INTERRUPT_flag_bF_buf13_bF_buf3) );
BUFX2 BUFX2_23 ( .A(INTERRUPT_flag_bF_buf3), .Y(INTERRUPT_flag_bF_buf13_bF_buf2) );
BUFX2 BUFX2_24 ( .A(INTERRUPT_flag_bF_buf5), .Y(INTERRUPT_flag_bF_buf13_bF_buf1) );
BUFX2 BUFX2_25 ( .A(INTERRUPT_flag_bF_buf1), .Y(INTERRUPT_flag_bF_buf13_bF_buf0) );
BUFX2 BUFX2_26 ( .A(INTERRUPT_flag_bF_buf1), .Y(INTERRUPT_flag_bF_buf14_bF_buf3) );
BUFX2 BUFX2_27 ( .A(INTERRUPT_flag_bF_buf12), .Y(INTERRUPT_flag_bF_buf14_bF_buf2) );
BUFX2 BUFX2_28 ( .A(INTERRUPT_flag_bF_buf5), .Y(INTERRUPT_flag_bF_buf14_bF_buf1) );
BUFX2 BUFX2_29 ( .A(INTERRUPT_flag_bF_buf5), .Y(INTERRUPT_flag_bF_buf14_bF_buf0) );
BUFX2 BUFX2_30 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf15_bF_buf3) );
BUFX2 BUFX2_31 ( .A(INTERRUPT_flag_bF_buf10), .Y(INTERRUPT_flag_bF_buf15_bF_buf2) );
BUFX2 BUFX2_32 ( .A(INTERRUPT_flag_bF_buf6), .Y(INTERRUPT_flag_bF_buf15_bF_buf1) );
BUFX2 BUFX2_33 ( .A(INTERRUPT_flag_bF_buf3), .Y(INTERRUPT_flag_bF_buf15_bF_buf0) );
BUFX2 BUFX2_34 ( .A(_1568__bF_buf2), .Y(_1568__bF_buf15_bF_buf3) );
BUFX2 BUFX2_35 ( .A(_1568__bF_buf6), .Y(_1568__bF_buf15_bF_buf2) );
BUFX2 BUFX2_36 ( .A(_1568__bF_buf6), .Y(_1568__bF_buf15_bF_buf1) );
BUFX2 BUFX2_37 ( .A(_1568__bF_buf3), .Y(_1568__bF_buf15_bF_buf0) );
BUFX2 BUFX2_38 ( .A(_1573_), .Y(_1573__hier0_bF_buf7) );
BUFX2 BUFX2_39 ( .A(_1573_), .Y(_1573__hier0_bF_buf6) );
BUFX2 BUFX2_40 ( .A(_1573_), .Y(_1573__hier0_bF_buf5) );
BUFX2 BUFX2_41 ( .A(_1573_), .Y(_1573__hier0_bF_buf4) );
BUFX2 BUFX2_42 ( .A(_1573_), .Y(_1573__hier0_bF_buf3) );
BUFX2 BUFX2_43 ( .A(_1573_), .Y(_1573__hier0_bF_buf2) );
BUFX2 BUFX2_44 ( .A(_1573_), .Y(_1573__hier0_bF_buf1) );
BUFX2 BUFX2_45 ( .A(_1573_), .Y(_1573__hier0_bF_buf0) );
BUFX2 BUFX2_46 ( .A(INTERRUPT_flag_bF_buf6), .Y(INTERRUPT_flag_bF_buf7_bF_buf3) );
BUFX2 BUFX2_47 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf7_bF_buf2) );
BUFX2 BUFX2_48 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf7_bF_buf1) );
BUFX2 BUFX2_49 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf7_bF_buf0) );
BUFX2 BUFX2_50 ( .A(INTERRUPT_flag_bF_buf6), .Y(INTERRUPT_flag_bF_buf8_bF_buf3) );
BUFX2 BUFX2_51 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf8_bF_buf2) );
BUFX2 BUFX2_52 ( .A(INTERRUPT_flag_bF_buf3), .Y(INTERRUPT_flag_bF_buf8_bF_buf1) );
BUFX2 BUFX2_53 ( .A(INTERRUPT_flag_bF_buf4), .Y(INTERRUPT_flag_bF_buf8_bF_buf0) );
BUFX2 BUFX2_54 ( .A(INTERRUPT_flag_bF_buf3), .Y(INTERRUPT_flag_bF_buf9_bF_buf3) );
BUFX2 BUFX2_55 ( .A(INTERRUPT_flag_bF_buf12), .Y(INTERRUPT_flag_bF_buf9_bF_buf2) );
BUFX2 BUFX2_56 ( .A(INTERRUPT_flag_bF_buf6), .Y(INTERRUPT_flag_bF_buf9_bF_buf1) );
BUFX2 BUFX2_57 ( .A(INTERRUPT_flag_bF_buf1), .Y(INTERRUPT_flag_bF_buf9_bF_buf0) );
BUFX2 BUFX2_58 ( .A(_3403_), .Y(_3403__bF_buf4) );
BUFX2 BUFX2_59 ( .A(_3403_), .Y(_3403__bF_buf3) );
BUFX2 BUFX2_60 ( .A(_3403_), .Y(_3403__bF_buf2) );
BUFX2 BUFX2_61 ( .A(_3403_), .Y(_3403__bF_buf1) );
BUFX2 BUFX2_62 ( .A(_3403_), .Y(_3403__bF_buf0) );
BUFX2 BUFX2_63 ( .A(_4361_), .Y(_4361__bF_buf4) );
BUFX2 BUFX2_64 ( .A(_4361_), .Y(_4361__bF_buf3) );
BUFX2 BUFX2_65 ( .A(_4361_), .Y(_4361__bF_buf2) );
BUFX2 BUFX2_66 ( .A(_4361_), .Y(_4361__bF_buf1) );
BUFX2 BUFX2_67 ( .A(_4361_), .Y(_4361__bF_buf0) );
BUFX2 BUFX2_68 ( .A(_1601_), .Y(_1601__bF_buf3) );
BUFX2 BUFX2_69 ( .A(_1601_), .Y(_1601__bF_buf2) );
BUFX2 BUFX2_70 ( .A(_1601_), .Y(_1601__bF_buf1) );
BUFX2 BUFX2_71 ( .A(_1601_), .Y(_1601__bF_buf0) );
BUFX2 BUFX2_72 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf7) );
BUFX2 BUFX2_73 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf6) );
BUFX2 BUFX2_74 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf5) );
BUFX2 BUFX2_75 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf4) );
BUFX2 BUFX2_76 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf3) );
BUFX2 BUFX2_77 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf2) );
BUFX2 BUFX2_78 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf1) );
BUFX2 BUFX2_79 ( .A(ULA_B_1_), .Y(ULA_B_1_bF_buf0) );
BUFX2 BUFX2_80 ( .A(_5945_), .Y(_5945__bF_buf3) );
BUFX2 BUFX2_81 ( .A(_5945_), .Y(_5945__bF_buf2) );
BUFX2 BUFX2_82 ( .A(_5945_), .Y(_5945__bF_buf1) );
BUFX2 BUFX2_83 ( .A(_5945_), .Y(_5945__bF_buf0) );
BUFX2 BUFX2_84 ( .A(_776_), .Y(_776__bF_buf3) );
BUFX2 BUFX2_85 ( .A(_776_), .Y(_776__bF_buf2) );
BUFX2 BUFX2_86 ( .A(_776_), .Y(_776__bF_buf1) );
BUFX2 BUFX2_87 ( .A(_776_), .Y(_776__bF_buf0) );
BUFX2 BUFX2_88 ( .A(_1577_), .Y(_1577__bF_buf3) );
BUFX2 BUFX2_89 ( .A(_1577_), .Y(_1577__bF_buf2) );
BUFX2 BUFX2_90 ( .A(_1577_), .Y(_1577__bF_buf1) );
BUFX2 BUFX2_91 ( .A(_1577_), .Y(_1577__bF_buf0) );
BUFX2 BUFX2_92 ( .A(_1730_), .Y(_1730__bF_buf4) );
BUFX2 BUFX2_93 ( .A(_1730_), .Y(_1730__bF_buf3) );
BUFX2 BUFX2_94 ( .A(_1730_), .Y(_1730__bF_buf2) );
BUFX2 BUFX2_95 ( .A(_1730_), .Y(_1730__bF_buf1) );
BUFX2 BUFX2_96 ( .A(_1730_), .Y(_1730__bF_buf0) );
BUFX2 BUFX2_97 ( .A(_1633_), .Y(_1633__bF_buf3) );
BUFX2 BUFX2_98 ( .A(_1633_), .Y(_1633__bF_buf2) );
BUFX2 BUFX2_99 ( .A(_1633_), .Y(_1633__bF_buf1) );
BUFX2 BUFX2_100 ( .A(_1633_), .Y(_1633__bF_buf0) );
BUFX2 BUFX2_101 ( .A(_409_), .Y(_409__bF_buf5) );
BUFX2 BUFX2_102 ( .A(_409_), .Y(_409__bF_buf4) );
BUFX2 BUFX2_103 ( .A(_409_), .Y(_409__bF_buf3) );
BUFX2 BUFX2_104 ( .A(_409_), .Y(_409__bF_buf2) );
BUFX2 BUFX2_105 ( .A(_409_), .Y(_409__bF_buf1) );
BUFX2 BUFX2_106 ( .A(_409_), .Y(_409__bF_buf0) );
BUFX2 BUFX2_107 ( .A(_3373_), .Y(_3373__bF_buf4) );
BUFX2 BUFX2_108 ( .A(_3373_), .Y(_3373__bF_buf3) );
BUFX2 BUFX2_109 ( .A(_3373_), .Y(_3373__bF_buf2) );
BUFX2 BUFX2_110 ( .A(_3373_), .Y(_3373__bF_buf1) );
BUFX2 BUFX2_111 ( .A(_3373_), .Y(_3373__bF_buf0) );
BUFX2 BUFX2_112 ( .A(_1627_), .Y(_1627__bF_buf3) );
BUFX2 BUFX2_113 ( .A(_1627_), .Y(_1627__bF_buf2) );
BUFX2 BUFX2_114 ( .A(_1627_), .Y(_1627__bF_buf1) );
BUFX2 BUFX2_115 ( .A(_1627_), .Y(_1627__bF_buf0) );
BUFX2 BUFX2_116 ( .A(_1568_), .Y(_1568__bF_buf15) );
BUFX2 BUFX2_117 ( .A(_1568_), .Y(_1568__bF_buf14) );
BUFX2 BUFX2_118 ( .A(_1568_), .Y(_1568__bF_buf13) );
BUFX2 BUFX2_119 ( .A(_1568_), .Y(_1568__bF_buf12) );
BUFX2 BUFX2_120 ( .A(_1568_), .Y(_1568__bF_buf11) );
BUFX2 BUFX2_121 ( .A(_1568_), .Y(_1568__bF_buf10) );
BUFX2 BUFX2_122 ( .A(_1568_), .Y(_1568__bF_buf9) );
BUFX2 BUFX2_123 ( .A(_1568_), .Y(_1568__bF_buf8) );
BUFX2 BUFX2_124 ( .A(_1568_), .Y(_1568__bF_buf7) );
BUFX2 BUFX2_125 ( .A(_1568_), .Y(_1568__bF_buf6) );
BUFX2 BUFX2_126 ( .A(_1568_), .Y(_1568__bF_buf5) );
BUFX2 BUFX2_127 ( .A(_1568_), .Y(_1568__bF_buf4) );
BUFX2 BUFX2_128 ( .A(_1568_), .Y(_1568__bF_buf3) );
BUFX2 BUFX2_129 ( .A(_1568_), .Y(_1568__bF_buf2) );
BUFX2 BUFX2_130 ( .A(_1568_), .Y(_1568__bF_buf1) );
BUFX2 BUFX2_131 ( .A(_1568_), .Y(_1568__bF_buf0) );
BUFX2 BUFX2_132 ( .A(_4728_), .Y(_4728__bF_buf4) );
BUFX2 BUFX2_133 ( .A(_4728_), .Y(_4728__bF_buf3) );
BUFX2 BUFX2_134 ( .A(_4728_), .Y(_4728__bF_buf2) );
BUFX2 BUFX2_135 ( .A(_4728_), .Y(_4728__bF_buf1) );
BUFX2 BUFX2_136 ( .A(_4728_), .Y(_4728__bF_buf0) );
BUFX2 BUFX2_137 ( .A(_1721_), .Y(_1721__bF_buf4) );
BUFX2 BUFX2_138 ( .A(_1721_), .Y(_1721__bF_buf3) );
BUFX2 BUFX2_139 ( .A(_1721_), .Y(_1721__bF_buf2) );
BUFX2 BUFX2_140 ( .A(_1721_), .Y(_1721__bF_buf1) );
BUFX2 BUFX2_141 ( .A(_1721_), .Y(_1721__bF_buf0) );
BUFX2 BUFX2_142 ( .A(_4860_), .Y(_4860__bF_buf4) );
BUFX2 BUFX2_143 ( .A(_4860_), .Y(_4860__bF_buf3) );
BUFX2 BUFX2_144 ( .A(_4860_), .Y(_4860__bF_buf2) );
BUFX2 BUFX2_145 ( .A(_4860_), .Y(_4860__bF_buf1) );
BUFX2 BUFX2_146 ( .A(_4860_), .Y(_4860__bF_buf0) );
BUFX2 BUFX2_147 ( .A(_5739_), .Y(_5739__bF_buf7) );
BUFX2 BUFX2_148 ( .A(_5739_), .Y(_5739__bF_buf6) );
BUFX2 BUFX2_149 ( .A(_5739_), .Y(_5739__bF_buf5) );
BUFX2 BUFX2_150 ( .A(_5739_), .Y(_5739__bF_buf4) );
BUFX2 BUFX2_151 ( .A(_5739_), .Y(_5739__bF_buf3) );
BUFX2 BUFX2_152 ( .A(_5739_), .Y(_5739__bF_buf2) );
BUFX2 BUFX2_153 ( .A(_5739_), .Y(_5739__bF_buf1) );
BUFX2 BUFX2_154 ( .A(_5739_), .Y(_5739__bF_buf0) );
BUFX2 BUFX2_155 ( .A(_1697_), .Y(_1697__bF_buf4) );
BUFX2 BUFX2_156 ( .A(_1697_), .Y(_1697__bF_buf3) );
BUFX2 BUFX2_157 ( .A(_1697_), .Y(_1697__bF_buf2) );
BUFX2 BUFX2_158 ( .A(_1697_), .Y(_1697__bF_buf1) );
BUFX2 BUFX2_159 ( .A(_1697_), .Y(_1697__bF_buf0) );
BUFX2 BUFX2_160 ( .A(_1621_), .Y(_1621__bF_buf3) );
BUFX2 BUFX2_161 ( .A(_1621_), .Y(_1621__bF_buf2) );
BUFX2 BUFX2_162 ( .A(_1621_), .Y(_1621__bF_buf1) );
BUFX2 BUFX2_163 ( .A(_1621_), .Y(_1621__bF_buf0) );
BUFX2 BUFX2_164 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf88) );
BUFX2 BUFX2_165 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf87) );
BUFX2 BUFX2_166 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf86) );
BUFX2 BUFX2_167 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf85) );
BUFX2 BUFX2_168 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf84) );
BUFX2 BUFX2_169 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf83) );
BUFX2 BUFX2_170 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf82) );
BUFX2 BUFX2_171 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf81) );
BUFX2 BUFX2_172 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf80) );
BUFX2 BUFX2_173 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf79) );
BUFX2 BUFX2_174 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf78) );
BUFX2 BUFX2_175 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf77) );
BUFX2 BUFX2_176 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf76) );
BUFX2 BUFX2_177 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf75) );
BUFX2 BUFX2_178 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf74) );
BUFX2 BUFX2_179 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf73) );
BUFX2 BUFX2_180 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf72) );
BUFX2 BUFX2_181 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf71) );
BUFX2 BUFX2_182 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf70) );
BUFX2 BUFX2_183 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf69) );
BUFX2 BUFX2_184 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf68) );
BUFX2 BUFX2_185 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf67) );
BUFX2 BUFX2_186 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf66) );
BUFX2 BUFX2_187 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf65) );
BUFX2 BUFX2_188 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf64) );
BUFX2 BUFX2_189 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf63) );
BUFX2 BUFX2_190 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf62) );
BUFX2 BUFX2_191 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf61) );
BUFX2 BUFX2_192 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf60) );
BUFX2 BUFX2_193 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf59) );
BUFX2 BUFX2_194 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf58) );
BUFX2 BUFX2_195 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf57) );
BUFX2 BUFX2_196 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf56) );
BUFX2 BUFX2_197 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf55) );
BUFX2 BUFX2_198 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf54) );
BUFX2 BUFX2_199 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf53) );
BUFX2 BUFX2_200 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf52) );
BUFX2 BUFX2_201 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf51) );
BUFX2 BUFX2_202 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf50) );
BUFX2 BUFX2_203 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf49) );
BUFX2 BUFX2_204 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf48) );
BUFX2 BUFX2_205 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf47) );
BUFX2 BUFX2_206 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf46) );
BUFX2 BUFX2_207 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf45) );
BUFX2 BUFX2_208 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf44) );
BUFX2 BUFX2_209 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf43) );
BUFX2 BUFX2_210 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf42) );
BUFX2 BUFX2_211 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf41) );
BUFX2 BUFX2_212 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf40) );
BUFX2 BUFX2_213 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf39) );
BUFX2 BUFX2_214 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf38) );
BUFX2 BUFX2_215 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf37) );
BUFX2 BUFX2_216 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf36) );
BUFX2 BUFX2_217 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf35) );
BUFX2 BUFX2_218 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf34) );
BUFX2 BUFX2_219 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf33) );
BUFX2 BUFX2_220 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf32) );
BUFX2 BUFX2_221 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf31) );
BUFX2 BUFX2_222 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf30) );
BUFX2 BUFX2_223 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf29) );
BUFX2 BUFX2_224 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28) );
BUFX2 BUFX2_225 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf27) );
BUFX2 BUFX2_226 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf26) );
BUFX2 BUFX2_227 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf25) );
BUFX2 BUFX2_228 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf24) );
BUFX2 BUFX2_229 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf23) );
BUFX2 BUFX2_230 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf22) );
BUFX2 BUFX2_231 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf21) );
BUFX2 BUFX2_232 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf20) );
BUFX2 BUFX2_233 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf19) );
BUFX2 BUFX2_234 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf18) );
BUFX2 BUFX2_235 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf17) );
BUFX2 BUFX2_236 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf16) );
BUFX2 BUFX2_237 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf15) );
BUFX2 BUFX2_238 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf14) );
BUFX2 BUFX2_239 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf13) );
BUFX2 BUFX2_240 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf12) );
BUFX2 BUFX2_241 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf11) );
BUFX2 BUFX2_242 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf10) );
BUFX2 BUFX2_243 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf9) );
BUFX2 BUFX2_244 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf8) );
BUFX2 BUFX2_245 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf7) );
BUFX2 BUFX2_246 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf6) );
BUFX2 BUFX2_247 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf5) );
BUFX2 BUFX2_248 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf4) );
BUFX2 BUFX2_249 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf3) );
BUFX2 BUFX2_250 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf2) );
BUFX2 BUFX2_251 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf1) );
BUFX2 BUFX2_252 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf0) );
BUFX2 BUFX2_253 ( .A(_626_), .Y(_626__bF_buf3) );
BUFX2 BUFX2_254 ( .A(_626_), .Y(_626__bF_buf2) );
BUFX2 BUFX2_255 ( .A(_626_), .Y(_626__bF_buf1) );
BUFX2 BUFX2_256 ( .A(_626_), .Y(_626__bF_buf0) );
BUFX2 BUFX2_257 ( .A(_473_), .Y(_473__bF_buf3) );
BUFX2 BUFX2_258 ( .A(_473_), .Y(_473__bF_buf2) );
BUFX2 BUFX2_259 ( .A(_473_), .Y(_473__bF_buf1) );
BUFX2 BUFX2_260 ( .A(_473_), .Y(_473__bF_buf0) );
BUFX2 BUFX2_261 ( .A(_1597_), .Y(_1597__bF_buf3) );
BUFX2 BUFX2_262 ( .A(_1597_), .Y(_1597__bF_buf2) );
BUFX2 BUFX2_263 ( .A(_1597_), .Y(_1597__bF_buf1) );
BUFX2 BUFX2_264 ( .A(_1597_), .Y(_1597__bF_buf0) );
BUFX2 BUFX2_265 ( .A(_470_), .Y(_470__bF_buf3) );
BUFX2 BUFX2_266 ( .A(_470_), .Y(_470__bF_buf2) );
BUFX2 BUFX2_267 ( .A(_470_), .Y(_470__bF_buf1) );
BUFX2 BUFX2_268 ( .A(_470_), .Y(_470__bF_buf0) );
BUFX2 BUFX2_269 ( .A(_1615_), .Y(_1615__bF_buf3) );
BUFX2 BUFX2_270 ( .A(_1615_), .Y(_1615__bF_buf2) );
BUFX2 BUFX2_271 ( .A(_1615_), .Y(_1615__bF_buf1) );
BUFX2 BUFX2_272 ( .A(_1615_), .Y(_1615__bF_buf0) );
BUFX2 BUFX2_273 ( .A(_3396_), .Y(_3396__bF_buf4) );
BUFX2 BUFX2_274 ( .A(_3396_), .Y(_3396__bF_buf3) );
BUFX2 BUFX2_275 ( .A(_3396_), .Y(_3396__bF_buf2) );
BUFX2 BUFX2_276 ( .A(_3396_), .Y(_3396__bF_buf1) );
BUFX2 BUFX2_277 ( .A(_3396_), .Y(_3396__bF_buf0) );
BUFX2 BUFX2_278 ( .A(_4563_), .Y(_4563__bF_buf4) );
BUFX2 BUFX2_279 ( .A(_4563_), .Y(_4563__bF_buf3) );
BUFX2 BUFX2_280 ( .A(_4563_), .Y(_4563__bF_buf2) );
BUFX2 BUFX2_281 ( .A(_4563_), .Y(_4563__bF_buf1) );
BUFX2 BUFX2_282 ( .A(_4563_), .Y(_4563__bF_buf0) );
BUFX2 BUFX2_283 ( .A(_3414_), .Y(_3414__bF_buf4) );
BUFX2 BUFX2_284 ( .A(_3414_), .Y(_3414__bF_buf3) );
BUFX2 BUFX2_285 ( .A(_3414_), .Y(_3414__bF_buf2) );
BUFX2 BUFX2_286 ( .A(_3414_), .Y(_3414__bF_buf1) );
BUFX2 BUFX2_287 ( .A(_3414_), .Y(_3414__bF_buf0) );
BUFX2 BUFX2_288 ( .A(_4695_), .Y(_4695__bF_buf4) );
BUFX2 BUFX2_289 ( .A(_4695_), .Y(_4695__bF_buf3) );
BUFX2 BUFX2_290 ( .A(_4695_), .Y(_4695__bF_buf2) );
BUFX2 BUFX2_291 ( .A(_4695_), .Y(_4695__bF_buf1) );
BUFX2 BUFX2_292 ( .A(_4695_), .Y(_4695__bF_buf0) );
BUFX2 BUFX2_293 ( .A(_5289_), .Y(_5289__bF_buf6) );
BUFX2 BUFX2_294 ( .A(_5289_), .Y(_5289__bF_buf5) );
BUFX2 BUFX2_295 ( .A(_5289_), .Y(_5289__bF_buf4) );
BUFX2 BUFX2_296 ( .A(_5289_), .Y(_5289__bF_buf3) );
BUFX2 BUFX2_297 ( .A(_5289_), .Y(_5289__bF_buf2) );
BUFX2 BUFX2_298 ( .A(_5289_), .Y(_5289__bF_buf1) );
BUFX2 BUFX2_299 ( .A(_5289_), .Y(_5289__bF_buf0) );
BUFX2 BUFX2_300 ( .A(_5730_), .Y(_5730__bF_buf3) );
BUFX2 BUFX2_301 ( .A(_5730_), .Y(_5730__bF_buf2) );
BUFX2 BUFX2_302 ( .A(_5730_), .Y(_5730__bF_buf1) );
BUFX2 BUFX2_303 ( .A(_5730_), .Y(_5730__bF_buf0) );
BUFX2 BUFX2_304 ( .A(_617_), .Y(_617__bF_buf3) );
BUFX2 BUFX2_305 ( .A(_617_), .Y(_617__bF_buf2) );
BUFX2 BUFX2_306 ( .A(_617_), .Y(_617__bF_buf1) );
BUFX2 BUFX2_307 ( .A(_617_), .Y(_617__bF_buf0) );
BUFX2 BUFX2_308 ( .A(_1609_), .Y(_1609__bF_buf3) );
BUFX2 BUFX2_309 ( .A(_1609_), .Y(_1609__bF_buf2) );
BUFX2 BUFX2_310 ( .A(_1609_), .Y(_1609__bF_buf1) );
BUFX2 BUFX2_311 ( .A(_1609_), .Y(_1609__bF_buf0) );
BUFX2 BUFX2_312 ( .A(_1591_), .Y(_1591__bF_buf3) );
BUFX2 BUFX2_313 ( .A(_1591_), .Y(_1591__bF_buf2) );
BUFX2 BUFX2_314 ( .A(_1591_), .Y(_1591__bF_buf1) );
BUFX2 BUFX2_315 ( .A(_1591_), .Y(_1591__bF_buf0) );
BUFX2 BUFX2_316 ( .A(CORE_ULA_REGB_Stall), .Y(CORE_ULA_REGB_Stall_bF_buf4) );
BUFX2 BUFX2_317 ( .A(CORE_ULA_REGB_Stall), .Y(CORE_ULA_REGB_Stall_bF_buf3) );
BUFX2 BUFX2_318 ( .A(CORE_ULA_REGB_Stall), .Y(CORE_ULA_REGB_Stall_bF_buf2) );
BUFX2 BUFX2_319 ( .A(CORE_ULA_REGB_Stall), .Y(CORE_ULA_REGB_Stall_bF_buf1) );
BUFX2 BUFX2_320 ( .A(CORE_ULA_REGB_Stall), .Y(CORE_ULA_REGB_Stall_bF_buf0) );
BUFX2 BUFX2_321 ( .A(_3411_), .Y(_3411__bF_buf4) );
BUFX2 BUFX2_322 ( .A(_3411_), .Y(_3411__bF_buf3) );
BUFX2 BUFX2_323 ( .A(_3411_), .Y(_3411__bF_buf2) );
BUFX2 BUFX2_324 ( .A(_3411_), .Y(_3411__bF_buf1) );
BUFX2 BUFX2_325 ( .A(_3411_), .Y(_3411__bF_buf0) );
BUFX2 BUFX2_326 ( .A(_3390_), .Y(_3390__bF_buf4) );
BUFX2 BUFX2_327 ( .A(_3390_), .Y(_3390__bF_buf3) );
BUFX2 BUFX2_328 ( .A(_3390_), .Y(_3390__bF_buf2) );
BUFX2 BUFX2_329 ( .A(_3390_), .Y(_3390__bF_buf1) );
BUFX2 BUFX2_330 ( .A(_3390_), .Y(_3390__bF_buf0) );
BUFX2 BUFX2_331 ( .A(_1741_), .Y(_1741__bF_buf4) );
BUFX2 BUFX2_332 ( .A(_1741_), .Y(_1741__bF_buf3) );
BUFX2 BUFX2_333 ( .A(_1741_), .Y(_1741__bF_buf2) );
BUFX2 BUFX2_334 ( .A(_1741_), .Y(_1741__bF_buf1) );
BUFX2 BUFX2_335 ( .A(_1741_), .Y(_1741__bF_buf0) );
BUFX2 BUFX2_336 ( .A(_1682_), .Y(_1682__bF_buf4) );
BUFX2 BUFX2_337 ( .A(_1682_), .Y(_1682__bF_buf3) );
BUFX2 BUFX2_338 ( .A(_1682_), .Y(_1682__bF_buf2) );
BUFX2 BUFX2_339 ( .A(_1682_), .Y(_1682__bF_buf1) );
BUFX2 BUFX2_340 ( .A(_1682_), .Y(_1682__bF_buf0) );
BUFX2 BUFX2_341 ( .A(_1585_), .Y(_1585__bF_buf3) );
BUFX2 BUFX2_342 ( .A(_1585_), .Y(_1585__bF_buf2) );
BUFX2 BUFX2_343 ( .A(_1585_), .Y(_1585__bF_buf1) );
BUFX2 BUFX2_344 ( .A(_1585_), .Y(_1585__bF_buf0) );
BUFX2 BUFX2_345 ( .A(_4325_), .Y(_4325__bF_buf4) );
BUFX2 BUFX2_346 ( .A(_4325_), .Y(_4325__bF_buf3) );
BUFX2 BUFX2_347 ( .A(_4325_), .Y(_4325__bF_buf2) );
BUFX2 BUFX2_348 ( .A(_4325_), .Y(_4325__bF_buf1) );
BUFX2 BUFX2_349 ( .A(_4325_), .Y(_4325__bF_buf0) );
BUFX2 BUFX2_350 ( .A(_1603_), .Y(_1603__bF_buf3) );
BUFX2 BUFX2_351 ( .A(_1603_), .Y(_1603__bF_buf2) );
BUFX2 BUFX2_352 ( .A(_1603_), .Y(_1603__bF_buf1) );
BUFX2 BUFX2_353 ( .A(_1603_), .Y(_1603__bF_buf0) );
BUFX2 BUFX2_354 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf7) );
BUFX2 BUFX2_355 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf6) );
BUFX2 BUFX2_356 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf5) );
BUFX2 BUFX2_357 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf4) );
BUFX2 BUFX2_358 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf3) );
BUFX2 BUFX2_359 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf2) );
BUFX2 BUFX2_360 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf1) );
BUFX2 BUFX2_361 ( .A(ULA_B_3_), .Y(ULA_B_3_bF_buf0) );
BUFX2 BUFX2_362 ( .A(_1735_), .Y(_1735__bF_buf4) );
BUFX2 BUFX2_363 ( .A(_1735_), .Y(_1735__bF_buf3) );
BUFX2 BUFX2_364 ( .A(_1735_), .Y(_1735__bF_buf2) );
BUFX2 BUFX2_365 ( .A(_1735_), .Y(_1735__bF_buf1) );
BUFX2 BUFX2_366 ( .A(_1735_), .Y(_1735__bF_buf0) );
BUFX2 BUFX2_367 ( .A(_1579_), .Y(_1579__bF_buf3) );
BUFX2 BUFX2_368 ( .A(_1579_), .Y(_1579__bF_buf2) );
BUFX2 BUFX2_369 ( .A(_1579_), .Y(_1579__bF_buf1) );
BUFX2 BUFX2_370 ( .A(_1579_), .Y(_1579__bF_buf0) );
BUFX2 BUFX2_371 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf7) );
BUFX2 BUFX2_372 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf6) );
BUFX2 BUFX2_373 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf5) );
BUFX2 BUFX2_374 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf4) );
BUFX2 BUFX2_375 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf3) );
BUFX2 BUFX2_376 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf2) );
BUFX2 BUFX2_377 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf1) );
BUFX2 BUFX2_378 ( .A(ULA_B_0_), .Y(ULA_B_0_bF_buf0) );
BUFX2 BUFX2_379 ( .A(_3381_), .Y(_3381__bF_buf4) );
BUFX2 BUFX2_380 ( .A(_3381_), .Y(_3381__bF_buf3) );
BUFX2 BUFX2_381 ( .A(_3381_), .Y(_3381__bF_buf2) );
BUFX2 BUFX2_382 ( .A(_3381_), .Y(_3381__bF_buf1) );
BUFX2 BUFX2_383 ( .A(_3381_), .Y(_3381__bF_buf0) );
BUFX2 BUFX2_384 ( .A(_4395_), .Y(_4395__bF_buf4) );
BUFX2 BUFX2_385 ( .A(_4395_), .Y(_4395__bF_buf3) );
BUFX2 BUFX2_386 ( .A(_4395_), .Y(_4395__bF_buf2) );
BUFX2 BUFX2_387 ( .A(_4395_), .Y(_4395__bF_buf1) );
BUFX2 BUFX2_388 ( .A(_4395_), .Y(_4395__bF_buf0) );
BUFX2 BUFX2_389 ( .A(_1635_), .Y(_1635__bF_buf3) );
BUFX2 BUFX2_390 ( .A(_1635_), .Y(_1635__bF_buf2) );
BUFX2 BUFX2_391 ( .A(_1635_), .Y(_1635__bF_buf1) );
BUFX2 BUFX2_392 ( .A(_1635_), .Y(_1635__bF_buf0) );
BUFX2 BUFX2_393 ( .A(_3378_), .Y(_3378__bF_buf4) );
BUFX2 BUFX2_394 ( .A(_3378_), .Y(_3378__bF_buf3) );
BUFX2 BUFX2_395 ( .A(_3378_), .Y(_3378__bF_buf2) );
BUFX2 BUFX2_396 ( .A(_3378_), .Y(_3378__bF_buf1) );
BUFX2 BUFX2_397 ( .A(_3378_), .Y(_3378__bF_buf0) );
BUFX2 BUFX2_398 ( .A(_5524_), .Y(_5524__bF_buf3) );
BUFX2 BUFX2_399 ( .A(_5524_), .Y(_5524__bF_buf2) );
BUFX2 BUFX2_400 ( .A(_5524_), .Y(_5524__bF_buf1) );
BUFX2 BUFX2_401 ( .A(_5524_), .Y(_5524__bF_buf0) );
BUFX2 BUFX2_402 ( .A(_487_), .Y(_487__bF_buf3) );
BUFX2 BUFX2_403 ( .A(_487_), .Y(_487__bF_buf2) );
BUFX2 BUFX2_404 ( .A(_487_), .Y(_487__bF_buf1) );
BUFX2 BUFX2_405 ( .A(_487_), .Y(_487__bF_buf0) );
BUFX2 BUFX2_406 ( .A(_505_), .Y(_505__bF_buf3) );
BUFX2 BUFX2_407 ( .A(_505_), .Y(_505__bF_buf2) );
BUFX2 BUFX2_408 ( .A(_505_), .Y(_505__bF_buf1) );
BUFX2 BUFX2_409 ( .A(_505_), .Y(_505__bF_buf0) );
BUFX2 BUFX2_410 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf78) );
BUFX2 BUFX2_411 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf77) );
BUFX2 BUFX2_412 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf76) );
BUFX2 BUFX2_413 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf75) );
BUFX2 BUFX2_414 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf74) );
BUFX2 BUFX2_415 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf73) );
BUFX2 BUFX2_416 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf72) );
BUFX2 BUFX2_417 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf71) );
BUFX2 BUFX2_418 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf70) );
BUFX2 BUFX2_419 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf69) );
BUFX2 BUFX2_420 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf68) );
BUFX2 BUFX2_421 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf67) );
BUFX2 BUFX2_422 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf66) );
BUFX2 BUFX2_423 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf65) );
BUFX2 BUFX2_424 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf64) );
BUFX2 BUFX2_425 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf63) );
BUFX2 BUFX2_426 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf62) );
BUFX2 BUFX2_427 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf61) );
BUFX2 BUFX2_428 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf60) );
BUFX2 BUFX2_429 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf59) );
BUFX2 BUFX2_430 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf58) );
BUFX2 BUFX2_431 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf57) );
BUFX2 BUFX2_432 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf56) );
BUFX2 BUFX2_433 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf55) );
BUFX2 BUFX2_434 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf54) );
BUFX2 BUFX2_435 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf53) );
BUFX2 BUFX2_436 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf52) );
BUFX2 BUFX2_437 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf51) );
BUFX2 BUFX2_438 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf50) );
BUFX2 BUFX2_439 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf49) );
BUFX2 BUFX2_440 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf48) );
BUFX2 BUFX2_441 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf47) );
BUFX2 BUFX2_442 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf46) );
BUFX2 BUFX2_443 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf45) );
BUFX2 BUFX2_444 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf44) );
BUFX2 BUFX2_445 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf43) );
BUFX2 BUFX2_446 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf42) );
BUFX2 BUFX2_447 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf41) );
BUFX2 BUFX2_448 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf40) );
BUFX2 BUFX2_449 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf39) );
BUFX2 BUFX2_450 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf38) );
BUFX2 BUFX2_451 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf37) );
BUFX2 BUFX2_452 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf36) );
BUFX2 BUFX2_453 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf35) );
BUFX2 BUFX2_454 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf34) );
BUFX2 BUFX2_455 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf33) );
BUFX2 BUFX2_456 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf32) );
BUFX2 BUFX2_457 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf31) );
BUFX2 BUFX2_458 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf30) );
BUFX2 BUFX2_459 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf29) );
BUFX2 BUFX2_460 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf28) );
BUFX2 BUFX2_461 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf27) );
BUFX2 BUFX2_462 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf26) );
BUFX2 BUFX2_463 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf25) );
BUFX2 BUFX2_464 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf24) );
BUFX2 BUFX2_465 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf23) );
BUFX2 BUFX2_466 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf22) );
BUFX2 BUFX2_467 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf21) );
BUFX2 BUFX2_468 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf20) );
BUFX2 BUFX2_469 ( .A(_1573__hier0_bF_buf5), .Y(_1573__bF_buf19) );
BUFX2 BUFX2_470 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf18) );
BUFX2 BUFX2_471 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf17) );
BUFX2 BUFX2_472 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf16) );
BUFX2 BUFX2_473 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf15) );
BUFX2 BUFX2_474 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf14) );
BUFX2 BUFX2_475 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf13) );
BUFX2 BUFX2_476 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf12) );
BUFX2 BUFX2_477 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf11) );
BUFX2 BUFX2_478 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf10) );
BUFX2 BUFX2_479 ( .A(_1573__hier0_bF_buf7), .Y(_1573__bF_buf9) );
BUFX2 BUFX2_480 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf8) );
BUFX2 BUFX2_481 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf7) );
BUFX2 BUFX2_482 ( .A(_1573__hier0_bF_buf6), .Y(_1573__bF_buf6) );
BUFX2 BUFX2_483 ( .A(_1573__hier0_bF_buf4), .Y(_1573__bF_buf5) );
BUFX2 BUFX2_484 ( .A(_1573__hier0_bF_buf0), .Y(_1573__bF_buf4) );
BUFX2 BUFX2_485 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf3) );
BUFX2 BUFX2_486 ( .A(_1573__hier0_bF_buf1), .Y(_1573__bF_buf2) );
BUFX2 BUFX2_487 ( .A(_1573__hier0_bF_buf2), .Y(_1573__bF_buf1) );
BUFX2 BUFX2_488 ( .A(_1573__hier0_bF_buf3), .Y(_1573__bF_buf0) );
BUFX2 BUFX2_489 ( .A(_484_), .Y(_484__bF_buf3) );
BUFX2 BUFX2_490 ( .A(_484_), .Y(_484__bF_buf2) );
BUFX2 BUFX2_491 ( .A(_484_), .Y(_484__bF_buf1) );
BUFX2 BUFX2_492 ( .A(_484_), .Y(_484__bF_buf0) );
BUFX2 BUFX2_493 ( .A(_1629_), .Y(_1629__bF_buf3) );
BUFX2 BUFX2_494 ( .A(_1629_), .Y(_1629__bF_buf2) );
BUFX2 BUFX2_495 ( .A(_1629_), .Y(_1629__bF_buf1) );
BUFX2 BUFX2_496 ( .A(_1629_), .Y(_1629__bF_buf0) );
BUFX2 BUFX2_497 ( .A(_4827_), .Y(_4827__bF_buf4) );
BUFX2 BUFX2_498 ( .A(_4827_), .Y(_4827__bF_buf3) );
BUFX2 BUFX2_499 ( .A(_4827_), .Y(_4827__bF_buf2) );
BUFX2 BUFX2_500 ( .A(_4827_), .Y(_4827__bF_buf1) );
BUFX2 BUFX2_501 ( .A(_4827_), .Y(_4827__bF_buf0) );
BUFX2 BUFX2_502 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf15) );
BUFX2 BUFX2_503 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf14) );
BUFX2 BUFX2_504 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf13) );
BUFX2 BUFX2_505 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf12) );
BUFX2 BUFX2_506 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf11) );
BUFX2 BUFX2_507 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf10) );
BUFX2 BUFX2_508 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf9) );
BUFX2 BUFX2_509 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf8) );
BUFX2 BUFX2_510 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf7) );
BUFX2 BUFX2_511 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf6) );
BUFX2 BUFX2_512 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf5) );
BUFX2 BUFX2_513 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf4) );
BUFX2 BUFX2_514 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf3) );
BUFX2 BUFX2_515 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf2) );
BUFX2 BUFX2_516 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf1) );
BUFX2 BUFX2_517 ( .A(INTERRUPT_flag), .Y(INTERRUPT_flag_bF_buf0) );
BUFX2 BUFX2_518 ( .A(rst), .Y(rst_bF_buf4) );
BUFX2 BUFX2_519 ( .A(rst), .Y(rst_bF_buf3) );
BUFX2 BUFX2_520 ( .A(rst), .Y(rst_bF_buf2) );
BUFX2 BUFX2_521 ( .A(rst), .Y(rst_bF_buf1) );
BUFX2 BUFX2_522 ( .A(rst), .Y(rst_bF_buf0) );
BUFX2 BUFX2_523 ( .A(_3369_), .Y(_3369__bF_buf4) );
BUFX2 BUFX2_524 ( .A(_3369_), .Y(_3369__bF_buf3) );
BUFX2 BUFX2_525 ( .A(_3369_), .Y(_3369__bF_buf2) );
BUFX2 BUFX2_526 ( .A(_3369_), .Y(_3369__bF_buf1) );
BUFX2 BUFX2_527 ( .A(_3369_), .Y(_3369__bF_buf0) );
BUFX2 BUFX2_528 ( .A(_1567_), .Y(_1567__bF_buf3) );
BUFX2 BUFX2_529 ( .A(_1567_), .Y(_1567__bF_buf2) );
BUFX2 BUFX2_530 ( .A(_1567_), .Y(_1567__bF_buf1) );
BUFX2 BUFX2_531 ( .A(_1567_), .Y(_1567__bF_buf0) );
BUFX2 BUFX2_532 ( .A(_1699_), .Y(_1699__bF_buf4) );
BUFX2 BUFX2_533 ( .A(_1699_), .Y(_1699__bF_buf3) );
BUFX2 BUFX2_534 ( .A(_1699_), .Y(_1699__bF_buf2) );
BUFX2 BUFX2_535 ( .A(_1699_), .Y(_1699__bF_buf1) );
BUFX2 BUFX2_536 ( .A(_1699_), .Y(_1699__bF_buf0) );
BUFX2 BUFX2_537 ( .A(_1623_), .Y(_1623__bF_buf3) );
BUFX2 BUFX2_538 ( .A(_1623_), .Y(_1623__bF_buf2) );
BUFX2 BUFX2_539 ( .A(_1623_), .Y(_1623__bF_buf1) );
BUFX2 BUFX2_540 ( .A(_1623_), .Y(_1623__bF_buf0) );
BUFX2 BUFX2_541 ( .A(_5682_), .Y(_5682__bF_buf6) );
BUFX2 BUFX2_542 ( .A(_5682_), .Y(_5682__bF_buf5) );
BUFX2 BUFX2_543 ( .A(_5682_), .Y(_5682__bF_buf4) );
BUFX2 BUFX2_544 ( .A(_5682_), .Y(_5682__bF_buf3) );
BUFX2 BUFX2_545 ( .A(_5682_), .Y(_5682__bF_buf2) );
BUFX2 BUFX2_546 ( .A(_5682_), .Y(_5682__bF_buf1) );
BUFX2 BUFX2_547 ( .A(_5682_), .Y(_5682__bF_buf0) );
BUFX2 BUFX2_548 ( .A(_1599_), .Y(_1599__bF_buf3) );
BUFX2 BUFX2_549 ( .A(_1599_), .Y(_1599__bF_buf2) );
BUFX2 BUFX2_550 ( .A(_1599_), .Y(_1599__bF_buf1) );
BUFX2 BUFX2_551 ( .A(_1599_), .Y(_1599__bF_buf0) );
BUFX2 BUFX2_552 ( .A(_1617_), .Y(_1617__bF_buf3) );
BUFX2 BUFX2_553 ( .A(_1617_), .Y(_1617__bF_buf2) );
BUFX2 BUFX2_554 ( .A(_1617_), .Y(_1617__bF_buf1) );
BUFX2 BUFX2_555 ( .A(_1617_), .Y(_1617__bF_buf0) );
BUFX2 BUFX2_556 ( .A(_4530_), .Y(_4530__bF_buf4) );
BUFX2 BUFX2_557 ( .A(_4530_), .Y(_4530__bF_buf3) );
BUFX2 BUFX2_558 ( .A(_4530_), .Y(_4530__bF_buf2) );
BUFX2 BUFX2_559 ( .A(_4530_), .Y(_4530__bF_buf1) );
BUFX2 BUFX2_560 ( .A(_4530_), .Y(_4530__bF_buf0) );
BUFX2 BUFX2_561 ( .A(_5735_), .Y(_5735__bF_buf4) );
BUFX2 BUFX2_562 ( .A(_5735_), .Y(_5735__bF_buf3) );
BUFX2 BUFX2_563 ( .A(_5735_), .Y(_5735__bF_buf2) );
BUFX2 BUFX2_564 ( .A(_5735_), .Y(_5735__bF_buf1) );
BUFX2 BUFX2_565 ( .A(_5735_), .Y(_5735__bF_buf0) );
BUFX2 BUFX2_566 ( .A(_3398_), .Y(_3398__bF_buf4) );
BUFX2 BUFX2_567 ( .A(_3398_), .Y(_3398__bF_buf3) );
BUFX2 BUFX2_568 ( .A(_3398_), .Y(_3398__bF_buf2) );
BUFX2 BUFX2_569 ( .A(_3398_), .Y(_3398__bF_buf1) );
BUFX2 BUFX2_570 ( .A(_3398_), .Y(_3398__bF_buf0) );
BUFX2 BUFX2_571 ( .A(_5353_), .Y(_5353__bF_buf4) );
BUFX2 BUFX2_572 ( .A(_5353_), .Y(_5353__bF_buf3) );
BUFX2 BUFX2_573 ( .A(_5353_), .Y(_5353__bF_buf2) );
BUFX2 BUFX2_574 ( .A(_5353_), .Y(_5353__bF_buf1) );
BUFX2 BUFX2_575 ( .A(_5353_), .Y(_5353__bF_buf0) );
BUFX2 BUFX2_576 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf7) );
BUFX2 BUFX2_577 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf6) );
BUFX2 BUFX2_578 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf5) );
BUFX2 BUFX2_579 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf4) );
BUFX2 BUFX2_580 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf3) );
BUFX2 BUFX2_581 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf2) );
BUFX2 BUFX2_582 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf1) );
BUFX2 BUFX2_583 ( .A(CORE_DATA_REGMux_exec_pipe), .Y(CORE_DATA_REGMux_exec_pipe_bF_buf0) );
BUFX2 BUFX2_584 ( .A(_4662_), .Y(_4662__bF_buf4) );
BUFX2 BUFX2_585 ( .A(_4662_), .Y(_4662__bF_buf3) );
BUFX2 BUFX2_586 ( .A(_4662_), .Y(_4662__bF_buf2) );
BUFX2 BUFX2_587 ( .A(_4662_), .Y(_4662__bF_buf1) );
BUFX2 BUFX2_588 ( .A(_4662_), .Y(_4662__bF_buf0) );
BUFX2 BUFX2_589 ( .A(_3416_), .Y(_3416__bF_buf4) );
BUFX2 BUFX2_590 ( .A(_3416_), .Y(_3416__bF_buf3) );
BUFX2 BUFX2_591 ( .A(_3416_), .Y(_3416__bF_buf2) );
BUFX2 BUFX2_592 ( .A(_3416_), .Y(_3416__bF_buf1) );
BUFX2 BUFX2_593 ( .A(_3416_), .Y(_3416__bF_buf0) );
BUFX2 BUFX2_594 ( .A(_4794_), .Y(_4794__bF_buf4) );
BUFX2 BUFX2_595 ( .A(_4794_), .Y(_4794__bF_buf3) );
BUFX2 BUFX2_596 ( .A(_4794_), .Y(_4794__bF_buf2) );
BUFX2 BUFX2_597 ( .A(_4794_), .Y(_4794__bF_buf1) );
BUFX2 BUFX2_598 ( .A(_4794_), .Y(_4794__bF_buf0) );
BUFX2 BUFX2_599 ( .A(_1690_), .Y(_1690__bF_buf4) );
BUFX2 BUFX2_600 ( .A(_1690_), .Y(_1690__bF_buf3) );
BUFX2 BUFX2_601 ( .A(_1690_), .Y(_1690__bF_buf2) );
BUFX2 BUFX2_602 ( .A(_1690_), .Y(_1690__bF_buf1) );
BUFX2 BUFX2_603 ( .A(_1690_), .Y(_1690__bF_buf0) );
BUFX2 BUFX2_604 ( .A(_1746_), .Y(_1746__bF_buf4) );
BUFX2 BUFX2_605 ( .A(_1746_), .Y(_1746__bF_buf3) );
BUFX2 BUFX2_606 ( .A(_1746_), .Y(_1746__bF_buf2) );
BUFX2 BUFX2_607 ( .A(_1746_), .Y(_1746__bF_buf1) );
BUFX2 BUFX2_608 ( .A(_1746_), .Y(_1746__bF_buf0) );
BUFX2 BUFX2_609 ( .A(_466_), .Y(_466__bF_buf3) );
BUFX2 BUFX2_610 ( .A(_466_), .Y(_466__bF_buf2) );
BUFX2 BUFX2_611 ( .A(_466_), .Y(_466__bF_buf1) );
BUFX2 BUFX2_612 ( .A(_466_), .Y(_466__bF_buf0) );
BUFX2 BUFX2_613 ( .A(_1593_), .Y(_1593__bF_buf3) );
BUFX2 BUFX2_614 ( .A(_1593_), .Y(_1593__bF_buf2) );
BUFX2 BUFX2_615 ( .A(_1593_), .Y(_1593__bF_buf1) );
BUFX2 BUFX2_616 ( .A(_1593_), .Y(_1593__bF_buf0) );
BUFX2 BUFX2_617 ( .A(_1687_), .Y(_1687__bF_buf4) );
BUFX2 BUFX2_618 ( .A(_1687_), .Y(_1687__bF_buf3) );
BUFX2 BUFX2_619 ( .A(_1687_), .Y(_1687__bF_buf2) );
BUFX2 BUFX2_620 ( .A(_1687_), .Y(_1687__bF_buf1) );
BUFX2 BUFX2_621 ( .A(_1687_), .Y(_1687__bF_buf0) );
BUFX2 BUFX2_622 ( .A(ULA_cin), .Y(ULA_cin_bF_buf7) );
BUFX2 BUFX2_623 ( .A(ULA_cin), .Y(ULA_cin_bF_buf6) );
BUFX2 BUFX2_624 ( .A(ULA_cin), .Y(ULA_cin_bF_buf5) );
BUFX2 BUFX2_625 ( .A(ULA_cin), .Y(ULA_cin_bF_buf4) );
BUFX2 BUFX2_626 ( .A(ULA_cin), .Y(ULA_cin_bF_buf3) );
BUFX2 BUFX2_627 ( .A(ULA_cin), .Y(ULA_cin_bF_buf2) );
BUFX2 BUFX2_628 ( .A(ULA_cin), .Y(ULA_cin_bF_buf1) );
BUFX2 BUFX2_629 ( .A(ULA_cin), .Y(ULA_cin_bF_buf0) );
BUFX2 BUFX2_630 ( .A(_1611_), .Y(_1611__bF_buf3) );
BUFX2 BUFX2_631 ( .A(_1611_), .Y(_1611__bF_buf2) );
BUFX2 BUFX2_632 ( .A(_1611_), .Y(_1611__bF_buf1) );
BUFX2 BUFX2_633 ( .A(_1611_), .Y(_1611__bF_buf0) );
BUFX2 BUFX2_634 ( .A(_1705_), .Y(_1705__bF_buf4) );
BUFX2 BUFX2_635 ( .A(_1705_), .Y(_1705__bF_buf3) );
BUFX2 BUFX2_636 ( .A(_1705_), .Y(_1705__bF_buf2) );
BUFX2 BUFX2_637 ( .A(_1705_), .Y(_1705__bF_buf1) );
BUFX2 BUFX2_638 ( .A(_1705_), .Y(_1705__bF_buf0) );
BUFX2 BUFX2_639 ( .A(_5438_), .Y(_5438__bF_buf3) );
BUFX2 BUFX2_640 ( .A(_5438_), .Y(_5438__bF_buf2) );
BUFX2 BUFX2_641 ( .A(_5438_), .Y(_5438__bF_buf1) );
BUFX2 BUFX2_642 ( .A(_5438_), .Y(_5438__bF_buf0) );
BUFX2 BUFX2_643 ( .A(_4462_), .Y(_4462__bF_buf4) );
BUFX2 BUFX2_644 ( .A(_4462_), .Y(_4462__bF_buf3) );
BUFX2 BUFX2_645 ( .A(_4462_), .Y(_4462__bF_buf2) );
BUFX2 BUFX2_646 ( .A(_4462_), .Y(_4462__bF_buf1) );
BUFX2 BUFX2_647 ( .A(_4462_), .Y(_4462__bF_buf0) );
BUFX2 BUFX2_648 ( .A(_1587_), .Y(_1587__bF_buf3) );
BUFX2 BUFX2_649 ( .A(_1587_), .Y(_1587__bF_buf2) );
BUFX2 BUFX2_650 ( .A(_1587_), .Y(_1587__bF_buf1) );
BUFX2 BUFX2_651 ( .A(_1587_), .Y(_1587__bF_buf0) );
BUFX2 BUFX2_652 ( .A(_1605_), .Y(_1605__bF_buf3) );
BUFX2 BUFX2_653 ( .A(_1605_), .Y(_1605__bF_buf2) );
BUFX2 BUFX2_654 ( .A(_1605_), .Y(_1605__bF_buf1) );
BUFX2 BUFX2_655 ( .A(_1605_), .Y(_1605__bF_buf0) );
BUFX2 BUFX2_656 ( .A(_3386_), .Y(_3386__bF_buf4) );
BUFX2 BUFX2_657 ( .A(_3386_), .Y(_3386__bF_buf3) );
BUFX2 BUFX2_658 ( .A(_3386_), .Y(_3386__bF_buf2) );
BUFX2 BUFX2_659 ( .A(_3386_), .Y(_3386__bF_buf1) );
BUFX2 BUFX2_660 ( .A(_3386_), .Y(_3386__bF_buf0) );
BUFX2 BUFX2_661 ( .A(_1678_), .Y(_1678__bF_buf4) );
BUFX2 BUFX2_662 ( .A(_1678_), .Y(_1678__bF_buf3) );
BUFX2 BUFX2_663 ( .A(_1678_), .Y(_1678__bF_buf2) );
BUFX2 BUFX2_664 ( .A(_1678_), .Y(_1678__bF_buf1) );
BUFX2 BUFX2_665 ( .A(_1678_), .Y(_1678__bF_buf0) );
BUFX2 BUFX2_666 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf7) );
BUFX2 BUFX2_667 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf6) );
BUFX2 BUFX2_668 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf5) );
BUFX2 BUFX2_669 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf4) );
BUFX2 BUFX2_670 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf3) );
BUFX2 BUFX2_671 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf2) );
BUFX2 BUFX2_672 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf1) );
BUFX2 BUFX2_673 ( .A(ULA_B_2_), .Y(ULA_B_2_bF_buf0) );
BUFX2 BUFX2_674 ( .A(_1581_), .Y(_1581__bF_buf3) );
BUFX2 BUFX2_675 ( .A(_1581_), .Y(_1581__bF_buf2) );
BUFX2 BUFX2_676 ( .A(_1581_), .Y(_1581__bF_buf1) );
BUFX2 BUFX2_677 ( .A(_1581_), .Y(_1581__bF_buf0) );
BUFX2 BUFX2_678 ( .A(_5470_), .Y(_5470__bF_buf3) );
BUFX2 BUFX2_679 ( .A(_5470_), .Y(_5470__bF_buf2) );
BUFX2 BUFX2_680 ( .A(_5470_), .Y(_5470__bF_buf1) );
BUFX2 BUFX2_681 ( .A(_5470_), .Y(_5470__bF_buf0) );
BUFX2 BUFX2_682 ( .A(_3401_), .Y(_3401__bF_buf4) );
BUFX2 BUFX2_683 ( .A(_3401_), .Y(_3401__bF_buf3) );
BUFX2 BUFX2_684 ( .A(_3401_), .Y(_3401__bF_buf2) );
BUFX2 BUFX2_685 ( .A(_3401_), .Y(_3401__bF_buf1) );
BUFX2 BUFX2_686 ( .A(_3401_), .Y(_3401__bF_buf0) );
BUFX2 BUFX2_687 ( .A(_5620_), .Y(_5620__bF_buf3) );
BUFX2 BUFX2_688 ( .A(_5620_), .Y(_5620__bF_buf2) );
BUFX2 BUFX2_689 ( .A(_5620_), .Y(_5620__bF_buf1) );
BUFX2 BUFX2_690 ( .A(_5620_), .Y(_5620__bF_buf0) );
BUFX2 BUFX2_691 ( .A(_451_), .Y(_451__bF_buf3) );
BUFX2 BUFX2_692 ( .A(_451_), .Y(_451__bF_buf2) );
BUFX2 BUFX2_693 ( .A(_451_), .Y(_451__bF_buf1) );
BUFX2 BUFX2_694 ( .A(_451_), .Y(_451__bF_buf0) );
BUFX2 BUFX2_695 ( .A(_5332_), .Y(_5332__bF_buf3) );
BUFX2 BUFX2_696 ( .A(_5332_), .Y(_5332__bF_buf2) );
BUFX2 BUFX2_697 ( .A(_5332_), .Y(_5332__bF_buf1) );
BUFX2 BUFX2_698 ( .A(_5332_), .Y(_5332__bF_buf0) );
BUFX2 BUFX2_699 ( .A(_1575_), .Y(_1575__bF_buf3) );
BUFX2 BUFX2_700 ( .A(_1575_), .Y(_1575__bF_buf2) );
BUFX2 BUFX2_701 ( .A(_1575_), .Y(_1575__bF_buf1) );
BUFX2 BUFX2_702 ( .A(_1575_), .Y(_1575__bF_buf0) );
BUFX2 BUFX2_703 ( .A(_4926_), .Y(_4926__bF_buf4) );
BUFX2 BUFX2_704 ( .A(_4926_), .Y(_4926__bF_buf3) );
BUFX2 BUFX2_705 ( .A(_4926_), .Y(_4926__bF_buf2) );
BUFX2 BUFX2_706 ( .A(_4926_), .Y(_4926__bF_buf1) );
BUFX2 BUFX2_707 ( .A(_4926_), .Y(_4926__bF_buf0) );
BUFX2 BUFX2_708 ( .A(_601_), .Y(_601__bF_buf3) );
BUFX2 BUFX2_709 ( .A(_601_), .Y(_601__bF_buf2) );
BUFX2 BUFX2_710 ( .A(_601_), .Y(_601__bF_buf1) );
BUFX2 BUFX2_711 ( .A(_601_), .Y(_601__bF_buf0) );
BUFX2 BUFX2_712 ( .A(_1631_), .Y(_1631__bF_buf3) );
BUFX2 BUFX2_713 ( .A(_1631_), .Y(_1631__bF_buf2) );
BUFX2 BUFX2_714 ( .A(_1631_), .Y(_1631__bF_buf1) );
BUFX2 BUFX2_715 ( .A(_1631_), .Y(_1631__bF_buf0) );
BUFX2 BUFX2_716 ( .A(_1572_), .Y(_1572__bF_buf4) );
BUFX2 BUFX2_717 ( .A(_1572_), .Y(_1572__bF_buf3) );
BUFX2 BUFX2_718 ( .A(_1572_), .Y(_1572__bF_buf2) );
BUFX2 BUFX2_719 ( .A(_1572_), .Y(_1572__bF_buf1) );
BUFX2 BUFX2_720 ( .A(_1572_), .Y(_1572__bF_buf0) );
BUFX2 BUFX2_721 ( .A(_4291_), .Y(_4291__bF_buf4) );
BUFX2 BUFX2_722 ( .A(_4291_), .Y(_4291__bF_buf3) );
BUFX2 BUFX2_723 ( .A(_4291_), .Y(_4291__bF_buf2) );
BUFX2 BUFX2_724 ( .A(_4291_), .Y(_4291__bF_buf1) );
BUFX2 BUFX2_725 ( .A(_4291_), .Y(_4291__bF_buf0) );
BUFX2 BUFX2_726 ( .A(_1625_), .Y(_1625__bF_buf3) );
BUFX2 BUFX2_727 ( .A(_1625_), .Y(_1625__bF_buf2) );
BUFX2 BUFX2_728 ( .A(_1625_), .Y(_1625__bF_buf1) );
BUFX2 BUFX2_729 ( .A(_1625_), .Y(_1625__bF_buf0) );
BUFX2 BUFX2_730 ( .A(_5417_), .Y(_5417__bF_buf5) );
BUFX2 BUFX2_731 ( .A(_5417_), .Y(_5417__bF_buf4) );
BUFX2 BUFX2_732 ( .A(_5417_), .Y(_5417__bF_buf3) );
BUFX2 BUFX2_733 ( .A(_5417_), .Y(_5417__bF_buf2) );
BUFX2 BUFX2_734 ( .A(_5417_), .Y(_5417__bF_buf1) );
BUFX2 BUFX2_735 ( .A(_5417_), .Y(_5417__bF_buf0) );
BUFX2 BUFX2_736 ( .A(_4629_), .Y(_4629__bF_buf4) );
BUFX2 BUFX2_737 ( .A(_4629_), .Y(_4629__bF_buf3) );
BUFX2 BUFX2_738 ( .A(_4629_), .Y(_4629__bF_buf2) );
BUFX2 BUFX2_739 ( .A(_4629_), .Y(_4629__bF_buf1) );
BUFX2 BUFX2_740 ( .A(_4629_), .Y(_4629__bF_buf0) );
BUFX2 BUFX2_741 ( .A(_5740_), .Y(_5740__bF_buf3) );
BUFX2 BUFX2_742 ( .A(_5740_), .Y(_5740__bF_buf2) );
BUFX2 BUFX2_743 ( .A(_5740_), .Y(_5740__bF_buf1) );
BUFX2 BUFX2_744 ( .A(_5740_), .Y(_5740__bF_buf0) );
BUFX2 BUFX2_745 ( .A(_1716_), .Y(_1716__bF_buf4) );
BUFX2 BUFX2_746 ( .A(_1716_), .Y(_1716__bF_buf3) );
BUFX2 BUFX2_747 ( .A(_1716_), .Y(_1716__bF_buf2) );
BUFX2 BUFX2_748 ( .A(_1716_), .Y(_1716__bF_buf1) );
BUFX2 BUFX2_749 ( .A(_1716_), .Y(_1716__bF_buf0) );
BUFX2 BUFX2_750 ( .A(_1619_), .Y(_1619__bF_buf3) );
BUFX2 BUFX2_751 ( .A(_1619_), .Y(_1619__bF_buf2) );
BUFX2 BUFX2_752 ( .A(_1619_), .Y(_1619__bF_buf1) );
BUFX2 BUFX2_753 ( .A(_1619_), .Y(_1619__bF_buf0) );
BUFX2 BUFX2_754 ( .A(_5681_), .Y(_5681__bF_buf6) );
BUFX2 BUFX2_755 ( .A(_5681_), .Y(_5681__bF_buf5) );
BUFX2 BUFX2_756 ( .A(_5681_), .Y(_5681__bF_buf4) );
BUFX2 BUFX2_757 ( .A(_5681_), .Y(_5681__bF_buf3) );
BUFX2 BUFX2_758 ( .A(_5681_), .Y(_5681__bF_buf2) );
BUFX2 BUFX2_759 ( .A(_5681_), .Y(_5681__bF_buf1) );
BUFX2 BUFX2_760 ( .A(_5681_), .Y(_5681__bF_buf0) );
BUFX2 BUFX2_761 ( .A(_4761_), .Y(_4761__bF_buf4) );
BUFX2 BUFX2_762 ( .A(_4761_), .Y(_4761__bF_buf3) );
BUFX2 BUFX2_763 ( .A(_4761_), .Y(_4761__bF_buf2) );
BUFX2 BUFX2_764 ( .A(_4761_), .Y(_4761__bF_buf1) );
BUFX2 BUFX2_765 ( .A(_4761_), .Y(_4761__bF_buf0) );
BUFX2 BUFX2_766 ( .A(_1695_), .Y(_1695__bF_buf4) );
BUFX2 BUFX2_767 ( .A(_1695_), .Y(_1695__bF_buf3) );
BUFX2 BUFX2_768 ( .A(_1695_), .Y(_1695__bF_buf2) );
BUFX2 BUFX2_769 ( .A(_1695_), .Y(_1695__bF_buf1) );
BUFX2 BUFX2_770 ( .A(_1695_), .Y(_1695__bF_buf0) );
BUFX2 BUFX2_771 ( .A(_4893_), .Y(_4893__bF_buf4) );
BUFX2 BUFX2_772 ( .A(_4893_), .Y(_4893__bF_buf3) );
BUFX2 BUFX2_773 ( .A(_4893_), .Y(_4893__bF_buf2) );
BUFX2 BUFX2_774 ( .A(_4893_), .Y(_4893__bF_buf1) );
BUFX2 BUFX2_775 ( .A(_4893_), .Y(_4893__bF_buf0) );
BUFX2 BUFX2_776 ( .A(_110_), .Y(_110__bF_buf4) );
BUFX2 BUFX2_777 ( .A(_110_), .Y(_110__bF_buf3) );
BUFX2 BUFX2_778 ( .A(_110_), .Y(_110__bF_buf2) );
BUFX2 BUFX2_779 ( .A(_110_), .Y(_110__bF_buf1) );
BUFX2 BUFX2_780 ( .A(_110_), .Y(_110__bF_buf0) );
BUFX2 BUFX2_781 ( .A(_107_), .Y(_107__bF_buf3) );
BUFX2 BUFX2_782 ( .A(_107_), .Y(_107__bF_buf2) );
BUFX2 BUFX2_783 ( .A(_107_), .Y(_107__bF_buf1) );
BUFX2 BUFX2_784 ( .A(_107_), .Y(_107__bF_buf0) );
BUFX2 BUFX2_785 ( .A(_5734_), .Y(_5734__bF_buf4) );
BUFX2 BUFX2_786 ( .A(_5734_), .Y(_5734__bF_buf3) );
BUFX2 BUFX2_787 ( .A(_5734_), .Y(_5734__bF_buf2) );
BUFX2 BUFX2_788 ( .A(_5734_), .Y(_5734__bF_buf1) );
BUFX2 BUFX2_789 ( .A(_5734_), .Y(_5734__bF_buf0) );
BUFX2 BUFX2_790 ( .A(_1595_), .Y(_1595__bF_buf3) );
BUFX2 BUFX2_791 ( .A(_1595_), .Y(_1595__bF_buf2) );
BUFX2 BUFX2_792 ( .A(_1595_), .Y(_1595__bF_buf1) );
BUFX2 BUFX2_793 ( .A(_1595_), .Y(_1595__bF_buf0) );
BUFX2 BUFX2_794 ( .A(_4429_), .Y(_4429__bF_buf4) );
BUFX2 BUFX2_795 ( .A(_4429_), .Y(_4429__bF_buf3) );
BUFX2 BUFX2_796 ( .A(_4429_), .Y(_4429__bF_buf2) );
BUFX2 BUFX2_797 ( .A(_4429_), .Y(_4429__bF_buf1) );
BUFX2 BUFX2_798 ( .A(_4429_), .Y(_4429__bF_buf0) );
BUFX2 BUFX2_799 ( .A(_1710_), .Y(_1710__bF_buf4) );
BUFX2 BUFX2_800 ( .A(_1710_), .Y(_1710__bF_buf3) );
BUFX2 BUFX2_801 ( .A(_1710_), .Y(_1710__bF_buf2) );
BUFX2 BUFX2_802 ( .A(_1710_), .Y(_1710__bF_buf1) );
BUFX2 BUFX2_803 ( .A(_1710_), .Y(_1710__bF_buf0) );
BUFX2 BUFX2_804 ( .A(_1613_), .Y(_1613__bF_buf3) );
BUFX2 BUFX2_805 ( .A(_1613_), .Y(_1613__bF_buf2) );
BUFX2 BUFX2_806 ( .A(_1613_), .Y(_1613__bF_buf1) );
BUFX2 BUFX2_807 ( .A(_1613_), .Y(_1613__bF_buf0) );
BUFX2 BUFX2_808 ( .A(_5669_), .Y(_5669__bF_buf3) );
BUFX2 BUFX2_809 ( .A(_5669_), .Y(_5669__bF_buf2) );
BUFX2 BUFX2_810 ( .A(_5669_), .Y(_5669__bF_buf1) );
BUFX2 BUFX2_811 ( .A(_5669_), .Y(_5669__bF_buf0) );
BUFX2 BUFX2_812 ( .A(_1589_), .Y(_1589__bF_buf3) );
BUFX2 BUFX2_813 ( .A(_1589_), .Y(_1589__bF_buf2) );
BUFX2 BUFX2_814 ( .A(_1589_), .Y(_1589__bF_buf1) );
BUFX2 BUFX2_815 ( .A(_1589_), .Y(_1589__bF_buf0) );
BUFX2 BUFX2_816 ( .A(_3409_), .Y(_3409__bF_buf4) );
BUFX2 BUFX2_817 ( .A(_3409_), .Y(_3409__bF_buf3) );
BUFX2 BUFX2_818 ( .A(_3409_), .Y(_3409__bF_buf2) );
BUFX2 BUFX2_819 ( .A(_3409_), .Y(_3409__bF_buf1) );
BUFX2 BUFX2_820 ( .A(_3409_), .Y(_3409__bF_buf0) );
BUFX2 BUFX2_821 ( .A(_4596_), .Y(_4596__bF_buf4) );
BUFX2 BUFX2_822 ( .A(_4596_), .Y(_4596__bF_buf3) );
BUFX2 BUFX2_823 ( .A(_4596_), .Y(_4596__bF_buf2) );
BUFX2 BUFX2_824 ( .A(_4596_), .Y(_4596__bF_buf1) );
BUFX2 BUFX2_825 ( .A(_4596_), .Y(_4596__bF_buf0) );
BUFX2 BUFX2_826 ( .A(_1607_), .Y(_1607__bF_buf3) );
BUFX2 BUFX2_827 ( .A(_1607_), .Y(_1607__bF_buf2) );
BUFX2 BUFX2_828 ( .A(_1607_), .Y(_1607__bF_buf1) );
BUFX2 BUFX2_829 ( .A(_1607_), .Y(_1607__bF_buf0) );
BUFX2 BUFX2_830 ( .A(_3388_), .Y(_3388__bF_buf4) );
BUFX2 BUFX2_831 ( .A(_3388_), .Y(_3388__bF_buf3) );
BUFX2 BUFX2_832 ( .A(_3388_), .Y(_3388__bF_buf2) );
BUFX2 BUFX2_833 ( .A(_3388_), .Y(_3388__bF_buf1) );
BUFX2 BUFX2_834 ( .A(_3388_), .Y(_3388__bF_buf0) );
BUFX2 BUFX2_835 ( .A(_4496_), .Y(_4496__bF_buf4) );
BUFX2 BUFX2_836 ( .A(_4496_), .Y(_4496__bF_buf3) );
BUFX2 BUFX2_837 ( .A(_4496_), .Y(_4496__bF_buf2) );
BUFX2 BUFX2_838 ( .A(_4496_), .Y(_4496__bF_buf1) );
BUFX2 BUFX2_839 ( .A(_4496_), .Y(_4496__bF_buf0) );
BUFX2 BUFX2_840 ( .A(ULA_B_4_), .Y(ULA_B_4_bF_buf3) );
BUFX2 BUFX2_841 ( .A(ULA_B_4_), .Y(ULA_B_4_bF_buf2) );
BUFX2 BUFX2_842 ( .A(ULA_B_4_), .Y(ULA_B_4_bF_buf1) );
BUFX2 BUFX2_843 ( .A(ULA_B_4_), .Y(ULA_B_4_bF_buf0) );
BUFX2 BUFX2_844 ( .A(_1642_), .Y(_1642__bF_buf4) );
BUFX2 BUFX2_845 ( .A(_1642_), .Y(_1642__bF_buf3) );
BUFX2 BUFX2_846 ( .A(_1642_), .Y(_1642__bF_buf2) );
BUFX2 BUFX2_847 ( .A(_1642_), .Y(_1642__bF_buf1) );
BUFX2 BUFX2_848 ( .A(_1642_), .Y(_1642__bF_buf0) );
BUFX2 BUFX2_849 ( .A(_98_), .Y(_98__bF_buf4) );
BUFX2 BUFX2_850 ( .A(_98_), .Y(_98__bF_buf3) );
BUFX2 BUFX2_851 ( .A(_98_), .Y(_98__bF_buf2) );
BUFX2 BUFX2_852 ( .A(_98_), .Y(_98__bF_buf1) );
BUFX2 BUFX2_853 ( .A(_98_), .Y(_98__bF_buf0) );
BUFX2 BUFX2_854 ( .A(_456_), .Y(_456__bF_buf3) );
BUFX2 BUFX2_855 ( .A(_456_), .Y(_456__bF_buf2) );
BUFX2 BUFX2_856 ( .A(_456_), .Y(_456__bF_buf1) );
BUFX2 BUFX2_857 ( .A(_456_), .Y(_456__bF_buf0) );
BUFX2 BUFX2_858 ( .A(_1583_), .Y(_1583__bF_buf3) );
BUFX2 BUFX2_859 ( .A(_1583_), .Y(_1583__bF_buf2) );
BUFX2 BUFX2_860 ( .A(_1583_), .Y(_1583__bF_buf1) );
BUFX2 BUFX2_861 ( .A(_1583_), .Y(_1583__bF_buf0) );
AND2X2 AND2X2_1 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__3_), .Y(_3486_) );
OR2X2 OR2X2_1 ( .A(_3485_), .B(_3486_), .Y(_3487_) );
OR2X2 OR2X2_2 ( .A(_3484_), .B(_3487_), .Y(_3488_) );
OR2X2 OR2X2_3 ( .A(_3488_), .B(_3483_), .Y(_3489_) );
AND2X2 AND2X2_2 ( .A(_1873_), .B(_3396__bF_buf1), .Y(_3490_) );
AND2X2 AND2X2_3 ( .A(_1877_), .B(_3398__bF_buf3), .Y(_3491_) );
OR2X2 OR2X2_4 ( .A(_3491_), .B(_3490_), .Y(_3492_) );
AND2X2 AND2X2_4 ( .A(_1882_), .B(_3401__bF_buf3), .Y(_3493_) );
AND2X2 AND2X2_5 ( .A(_1886_), .B(_3403__bF_buf2), .Y(_3494_) );
OR2X2 OR2X2_5 ( .A(_3494_), .B(_3493_), .Y(_3495_) );
OR2X2 OR2X2_6 ( .A(_3492_), .B(_3495_), .Y(_3496_) );
AND2X2 AND2X2_6 ( .A(_3409__bF_buf1), .B(_1892_), .Y(_3497_) );
AND2X2 AND2X2_7 ( .A(_3411__bF_buf0), .B(_1896_), .Y(_3498_) );
OR2X2 OR2X2_7 ( .A(_3497_), .B(_3498_), .Y(_3499_) );
AND2X2 AND2X2_8 ( .A(_1901_), .B(_3414__bF_buf3), .Y(_3500_) );
AND2X2 AND2X2_9 ( .A(_3416__bF_buf0), .B(_1905_), .Y(_3501_) );
OR2X2 OR2X2_8 ( .A(_3500_), .B(_3501_), .Y(_3502_) );
OR2X2 OR2X2_9 ( .A(_3502_), .B(_3499_), .Y(_3503_) );
OR2X2 OR2X2_10 ( .A(_3496_), .B(_3503_), .Y(_3504_) );
OR2X2 OR2X2_11 ( .A(_3489_), .B(_3504_), .Y(REG_A_3_) );
AND2X2 AND2X2_10 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__4_), .Y(_3505_) );
AND2X2 AND2X2_11 ( .A(_3373__bF_buf1), .B(REGs_REGS_5__4_), .Y(_3506_) );
OR2X2 OR2X2_12 ( .A(_3505_), .B(_3506_), .Y(_3507_) );
AND2X2 AND2X2_12 ( .A(_3378__bF_buf0), .B(REGs_REGS_6__4_), .Y(_3508_) );
AND2X2 AND2X2_13 ( .A(_3381__bF_buf1), .B(REGs_REGS_7__4_), .Y(_3509_) );
OR2X2 OR2X2_13 ( .A(_3509_), .B(_3508_), .Y(_3510_) );
OR2X2 OR2X2_14 ( .A(_3507_), .B(_3510_), .Y(_3511_) );
AND2X2 AND2X2_14 ( .A(_3386__bF_buf4), .B(PC_ADDR_stack_1__4_), .Y(_3512_) );
AND2X2 AND2X2_15 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__4_), .Y(_3513_) );
AND2X2 AND2X2_16 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__4_), .Y(_3514_) );
OR2X2 OR2X2_15 ( .A(_3513_), .B(_3514_), .Y(_3515_) );
OR2X2 OR2X2_16 ( .A(_3512_), .B(_3515_), .Y(_3516_) );
OR2X2 OR2X2_17 ( .A(_3516_), .B(_3511_), .Y(_3517_) );
AND2X2 AND2X2_17 ( .A(_1925_), .B(_3396__bF_buf1), .Y(_3518_) );
AND2X2 AND2X2_18 ( .A(_1929_), .B(_3398__bF_buf3), .Y(_3519_) );
OR2X2 OR2X2_18 ( .A(_3519_), .B(_3518_), .Y(_3520_) );
AND2X2 AND2X2_19 ( .A(_1934_), .B(_3401__bF_buf3), .Y(_3521_) );
AND2X2 AND2X2_20 ( .A(_1938_), .B(_3403__bF_buf2), .Y(_3522_) );
OR2X2 OR2X2_19 ( .A(_3522_), .B(_3521_), .Y(_3523_) );
OR2X2 OR2X2_20 ( .A(_3520_), .B(_3523_), .Y(_3524_) );
AND2X2 AND2X2_21 ( .A(_3409__bF_buf1), .B(_1944_), .Y(_3525_) );
AND2X2 AND2X2_22 ( .A(_3411__bF_buf0), .B(_1948_), .Y(_3526_) );
OR2X2 OR2X2_21 ( .A(_3525_), .B(_3526_), .Y(_3527_) );
AND2X2 AND2X2_23 ( .A(_1953_), .B(_3414__bF_buf3), .Y(_3528_) );
AND2X2 AND2X2_24 ( .A(_3416__bF_buf0), .B(_1957_), .Y(_3529_) );
OR2X2 OR2X2_22 ( .A(_3528_), .B(_3529_), .Y(_3530_) );
OR2X2 OR2X2_23 ( .A(_3530_), .B(_3527_), .Y(_3531_) );
OR2X2 OR2X2_24 ( .A(_3524_), .B(_3531_), .Y(_3532_) );
OR2X2 OR2X2_25 ( .A(_3517_), .B(_3532_), .Y(REG_A_4_) );
AND2X2 AND2X2_25 ( .A(_3369__bF_buf2), .B(REGs_REGS_4__5_), .Y(_3533_) );
AND2X2 AND2X2_26 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__5_), .Y(_3534_) );
OR2X2 OR2X2_26 ( .A(_3533_), .B(_3534_), .Y(_3535_) );
AND2X2 AND2X2_27 ( .A(_3378__bF_buf1), .B(REGs_REGS_6__5_), .Y(_3536_) );
AND2X2 AND2X2_28 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__5_), .Y(_3537_) );
OR2X2 OR2X2_27 ( .A(_3537_), .B(_3536_), .Y(_3538_) );
OR2X2 OR2X2_28 ( .A(_3535_), .B(_3538_), .Y(_3539_) );
AND2X2 AND2X2_29 ( .A(_3386__bF_buf0), .B(PC_ADDR_stack_1__5_), .Y(_3540_) );
AND2X2 AND2X2_30 ( .A(_3388__bF_buf2), .B(REGs_REGS_3__5_), .Y(_3541_) );
AND2X2 AND2X2_31 ( .A(_3390__bF_buf0), .B(REGs_REGS_2__5_), .Y(_3542_) );
OR2X2 OR2X2_29 ( .A(_3541_), .B(_3542_), .Y(_3543_) );
OR2X2 OR2X2_30 ( .A(_3540_), .B(_3543_), .Y(_3544_) );
OR2X2 OR2X2_31 ( .A(_3544_), .B(_3539_), .Y(_3545_) );
AND2X2 AND2X2_32 ( .A(_1977_), .B(_3396__bF_buf3), .Y(_3546_) );
AND2X2 AND2X2_33 ( .A(_1981_), .B(_3398__bF_buf0), .Y(_3547_) );
OR2X2 OR2X2_32 ( .A(_3547_), .B(_3546_), .Y(_3548_) );
AND2X2 AND2X2_34 ( .A(_1986_), .B(_3401__bF_buf1), .Y(_3549_) );
AND2X2 AND2X2_35 ( .A(_1990_), .B(_3403__bF_buf4), .Y(_3550_) );
OR2X2 OR2X2_33 ( .A(_3550_), .B(_3549_), .Y(_3551_) );
OR2X2 OR2X2_34 ( .A(_3548_), .B(_3551_), .Y(_3552_) );
AND2X2 AND2X2_36 ( .A(_3409__bF_buf2), .B(_1996_), .Y(_3553_) );
AND2X2 AND2X2_37 ( .A(_3411__bF_buf1), .B(_2000_), .Y(_3554_) );
OR2X2 OR2X2_35 ( .A(_3553_), .B(_3554_), .Y(_3555_) );
AND2X2 AND2X2_38 ( .A(_2005_), .B(_3414__bF_buf2), .Y(_3556_) );
AND2X2 AND2X2_39 ( .A(_3416__bF_buf2), .B(_2009_), .Y(_3557_) );
OR2X2 OR2X2_36 ( .A(_3556_), .B(_3557_), .Y(_3558_) );
OR2X2 OR2X2_37 ( .A(_3558_), .B(_3555_), .Y(_3559_) );
OR2X2 OR2X2_38 ( .A(_3552_), .B(_3559_), .Y(_3560_) );
OR2X2 OR2X2_39 ( .A(_3545_), .B(_3560_), .Y(REG_A_5_) );
AND2X2 AND2X2_40 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__6_), .Y(_3561_) );
AND2X2 AND2X2_41 ( .A(_3373__bF_buf1), .B(REGs_REGS_5__6_), .Y(_3562_) );
OR2X2 OR2X2_40 ( .A(_3561_), .B(_3562_), .Y(_3563_) );
AND2X2 AND2X2_42 ( .A(_3378__bF_buf0), .B(REGs_REGS_6__6_), .Y(_3564_) );
AND2X2 AND2X2_43 ( .A(_3381__bF_buf1), .B(REGs_REGS_7__6_), .Y(_3565_) );
OR2X2 OR2X2_41 ( .A(_3565_), .B(_3564_), .Y(_3566_) );
OR2X2 OR2X2_42 ( .A(_3563_), .B(_3566_), .Y(_3567_) );
AND2X2 AND2X2_44 ( .A(_3386__bF_buf4), .B(PC_ADDR_stack_1__6_), .Y(_3568_) );
AND2X2 AND2X2_45 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__6_), .Y(_3569_) );
AND2X2 AND2X2_46 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__6_), .Y(_3570_) );
OR2X2 OR2X2_43 ( .A(_3569_), .B(_3570_), .Y(_3571_) );
OR2X2 OR2X2_44 ( .A(_3568_), .B(_3571_), .Y(_3572_) );
OR2X2 OR2X2_45 ( .A(_3572_), .B(_3567_), .Y(_3573_) );
AND2X2 AND2X2_47 ( .A(_2029_), .B(_3396__bF_buf1), .Y(_3574_) );
AND2X2 AND2X2_48 ( .A(_2033_), .B(_3398__bF_buf3), .Y(_3575_) );
OR2X2 OR2X2_46 ( .A(_3575_), .B(_3574_), .Y(_3576_) );
AND2X2 AND2X2_49 ( .A(_2038_), .B(_3401__bF_buf3), .Y(_3577_) );
AND2X2 AND2X2_50 ( .A(_2042_), .B(_3403__bF_buf2), .Y(_3578_) );
OR2X2 OR2X2_47 ( .A(_3578_), .B(_3577_), .Y(_3579_) );
OR2X2 OR2X2_48 ( .A(_3576_), .B(_3579_), .Y(_3580_) );
AND2X2 AND2X2_51 ( .A(_3409__bF_buf1), .B(_2048_), .Y(_3581_) );
AND2X2 AND2X2_52 ( .A(_3411__bF_buf0), .B(_2052_), .Y(_3582_) );
OR2X2 OR2X2_49 ( .A(_3581_), .B(_3582_), .Y(_3583_) );
AND2X2 AND2X2_53 ( .A(_2057_), .B(_3414__bF_buf3), .Y(_3584_) );
AND2X2 AND2X2_54 ( .A(_3416__bF_buf0), .B(_2061_), .Y(_3585_) );
OR2X2 OR2X2_50 ( .A(_3584_), .B(_3585_), .Y(_3586_) );
OR2X2 OR2X2_51 ( .A(_3586_), .B(_3583_), .Y(_3587_) );
OR2X2 OR2X2_52 ( .A(_3580_), .B(_3587_), .Y(_3588_) );
OR2X2 OR2X2_53 ( .A(_3573_), .B(_3588_), .Y(REG_A_6_) );
AND2X2 AND2X2_55 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__7_), .Y(_3589_) );
AND2X2 AND2X2_56 ( .A(_3373__bF_buf1), .B(REGs_REGS_5__7_), .Y(_3590_) );
OR2X2 OR2X2_54 ( .A(_3589_), .B(_3590_), .Y(_3591_) );
AND2X2 AND2X2_57 ( .A(_3378__bF_buf0), .B(REGs_REGS_6__7_), .Y(_3592_) );
AND2X2 AND2X2_58 ( .A(_3381__bF_buf1), .B(REGs_REGS_7__7_), .Y(_3593_) );
OR2X2 OR2X2_55 ( .A(_3593_), .B(_3592_), .Y(_3594_) );
OR2X2 OR2X2_56 ( .A(_3591_), .B(_3594_), .Y(_3595_) );
AND2X2 AND2X2_59 ( .A(_3386__bF_buf4), .B(PC_ADDR_stack_1__7_), .Y(_3596_) );
AND2X2 AND2X2_60 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__7_), .Y(_3597_) );
AND2X2 AND2X2_61 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__7_), .Y(_3598_) );
OR2X2 OR2X2_57 ( .A(_3597_), .B(_3598_), .Y(_3599_) );
OR2X2 OR2X2_58 ( .A(_3596_), .B(_3599_), .Y(_3600_) );
OR2X2 OR2X2_59 ( .A(_3600_), .B(_3595_), .Y(_3601_) );
AND2X2 AND2X2_62 ( .A(_2081_), .B(_3396__bF_buf2), .Y(_3602_) );
AND2X2 AND2X2_63 ( .A(_2085_), .B(_3398__bF_buf1), .Y(_3603_) );
OR2X2 OR2X2_60 ( .A(_3603_), .B(_3602_), .Y(_3604_) );
AND2X2 AND2X2_64 ( .A(_2090_), .B(_3401__bF_buf0), .Y(_3605_) );
AND2X2 AND2X2_65 ( .A(_2094_), .B(_3403__bF_buf3), .Y(_3606_) );
OR2X2 OR2X2_61 ( .A(_3606_), .B(_3605_), .Y(_3607_) );
OR2X2 OR2X2_62 ( .A(_3604_), .B(_3607_), .Y(_3608_) );
AND2X2 AND2X2_66 ( .A(_3409__bF_buf4), .B(_2100_), .Y(_3609_) );
AND2X2 AND2X2_67 ( .A(_3411__bF_buf2), .B(_2104_), .Y(_3610_) );
OR2X2 OR2X2_63 ( .A(_3609_), .B(_3610_), .Y(_3611_) );
AND2X2 AND2X2_68 ( .A(_2109_), .B(_3414__bF_buf4), .Y(_3612_) );
AND2X2 AND2X2_69 ( .A(_3416__bF_buf4), .B(_2113_), .Y(_3613_) );
OR2X2 OR2X2_64 ( .A(_3612_), .B(_3613_), .Y(_3614_) );
OR2X2 OR2X2_65 ( .A(_3614_), .B(_3611_), .Y(_3615_) );
OR2X2 OR2X2_66 ( .A(_3608_), .B(_3615_), .Y(_3616_) );
OR2X2 OR2X2_67 ( .A(_3601_), .B(_3616_), .Y(REG_A_7_) );
AND2X2 AND2X2_70 ( .A(_3369__bF_buf2), .B(REGs_REGS_4__8_), .Y(_3617_) );
AND2X2 AND2X2_71 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__8_), .Y(_3618_) );
OR2X2 OR2X2_68 ( .A(_3617_), .B(_3618_), .Y(_3619_) );
AND2X2 AND2X2_72 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__8_), .Y(_3620_) );
AND2X2 AND2X2_73 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__8_), .Y(_3621_) );
OR2X2 OR2X2_69 ( .A(_3621_), .B(_3620_), .Y(_3622_) );
OR2X2 OR2X2_70 ( .A(_3619_), .B(_3622_), .Y(_3623_) );
AND2X2 AND2X2_74 ( .A(_3386__bF_buf3), .B(gnd), .Y(_3624_) );
AND2X2 AND2X2_75 ( .A(_3388__bF_buf2), .B(REGs_REGS_3__8_), .Y(_3625_) );
AND2X2 AND2X2_76 ( .A(_3390__bF_buf0), .B(REGs_REGS_2__8_), .Y(_3626_) );
OR2X2 OR2X2_71 ( .A(_3625_), .B(_3626_), .Y(_3627_) );
OR2X2 OR2X2_72 ( .A(_3624_), .B(_3627_), .Y(_3628_) );
OR2X2 OR2X2_73 ( .A(_3628_), .B(_3623_), .Y(_3629_) );
AND2X2 AND2X2_77 ( .A(_2133_), .B(_3396__bF_buf0), .Y(_3630_) );
AND2X2 AND2X2_78 ( .A(_2137_), .B(_3398__bF_buf4), .Y(_3631_) );
OR2X2 OR2X2_74 ( .A(_3631_), .B(_3630_), .Y(_3632_) );
AND2X2 AND2X2_79 ( .A(_2142_), .B(_3401__bF_buf2), .Y(_3633_) );
AND2X2 AND2X2_80 ( .A(_2146_), .B(_3403__bF_buf0), .Y(_3634_) );
OR2X2 OR2X2_75 ( .A(_3634_), .B(_3633_), .Y(_3635_) );
OR2X2 OR2X2_76 ( .A(_3632_), .B(_3635_), .Y(_3636_) );
AND2X2 AND2X2_81 ( .A(_3409__bF_buf2), .B(_2152_), .Y(_3637_) );
AND2X2 AND2X2_82 ( .A(_3411__bF_buf1), .B(_2156_), .Y(_3638_) );
OR2X2 OR2X2_77 ( .A(_3637_), .B(_3638_), .Y(_3639_) );
AND2X2 AND2X2_83 ( .A(_2161_), .B(_3414__bF_buf0), .Y(_3640_) );
AND2X2 AND2X2_84 ( .A(_3416__bF_buf2), .B(_2165_), .Y(_3641_) );
OR2X2 OR2X2_78 ( .A(_3640_), .B(_3641_), .Y(_3642_) );
OR2X2 OR2X2_79 ( .A(_3642_), .B(_3639_), .Y(_3643_) );
OR2X2 OR2X2_80 ( .A(_3636_), .B(_3643_), .Y(_3644_) );
OR2X2 OR2X2_81 ( .A(_3629_), .B(_3644_), .Y(REG_A_8_) );
AND2X2 AND2X2_85 ( .A(_3369__bF_buf1), .B(REGs_REGS_4__9_), .Y(_3645_) );
AND2X2 AND2X2_86 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__9_), .Y(_3646_) );
OR2X2 OR2X2_82 ( .A(_3645_), .B(_3646_), .Y(_3647_) );
AND2X2 AND2X2_87 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__9_), .Y(_3648_) );
AND2X2 AND2X2_88 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__9_), .Y(_3649_) );
OR2X2 OR2X2_83 ( .A(_3649_), .B(_3648_), .Y(_3650_) );
OR2X2 OR2X2_84 ( .A(_3647_), .B(_3650_), .Y(_3651_) );
AND2X2 AND2X2_89 ( .A(_3386__bF_buf3), .B(gnd), .Y(_3652_) );
AND2X2 AND2X2_90 ( .A(_3388__bF_buf1), .B(REGs_REGS_3__9_), .Y(_3653_) );
AND2X2 AND2X2_91 ( .A(_3390__bF_buf1), .B(REGs_REGS_2__9_), .Y(_3654_) );
OR2X2 OR2X2_85 ( .A(_3653_), .B(_3654_), .Y(_3655_) );
OR2X2 OR2X2_86 ( .A(_3652_), .B(_3655_), .Y(_3656_) );
OR2X2 OR2X2_87 ( .A(_3656_), .B(_3651_), .Y(_3657_) );
AND2X2 AND2X2_92 ( .A(_2185_), .B(_3396__bF_buf3), .Y(_3658_) );
AND2X2 AND2X2_93 ( .A(_2189_), .B(_3398__bF_buf0), .Y(_3659_) );
OR2X2 OR2X2_88 ( .A(_3659_), .B(_3658_), .Y(_3660_) );
AND2X2 AND2X2_94 ( .A(_2194_), .B(_3401__bF_buf1), .Y(_3661_) );
AND2X2 AND2X2_95 ( .A(_2198_), .B(_3403__bF_buf4), .Y(_3662_) );
OR2X2 OR2X2_89 ( .A(_3662_), .B(_3661_), .Y(_3663_) );
OR2X2 OR2X2_90 ( .A(_3660_), .B(_3663_), .Y(_3664_) );
AND2X2 AND2X2_96 ( .A(_3409__bF_buf3), .B(_2204_), .Y(_3665_) );
AND2X2 AND2X2_97 ( .A(_3411__bF_buf3), .B(_2208_), .Y(_3666_) );
OR2X2 OR2X2_91 ( .A(_3665_), .B(_3666_), .Y(_3667_) );
AND2X2 AND2X2_98 ( .A(_2213_), .B(_3414__bF_buf2), .Y(_3668_) );
AND2X2 AND2X2_99 ( .A(_3416__bF_buf3), .B(_2217_), .Y(_3669_) );
OR2X2 OR2X2_92 ( .A(_3668_), .B(_3669_), .Y(_3670_) );
OR2X2 OR2X2_93 ( .A(_3670_), .B(_3667_), .Y(_3671_) );
OR2X2 OR2X2_94 ( .A(_3664_), .B(_3671_), .Y(_3672_) );
OR2X2 OR2X2_95 ( .A(_3657_), .B(_3672_), .Y(REG_A_9_) );
AND2X2 AND2X2_100 ( .A(_3369__bF_buf1), .B(REGs_REGS_4__10_), .Y(_3673_) );
AND2X2 AND2X2_101 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__10_), .Y(_3674_) );
OR2X2 OR2X2_96 ( .A(_3673_), .B(_3674_), .Y(_3675_) );
AND2X2 AND2X2_102 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__10_), .Y(_3676_) );
AND2X2 AND2X2_103 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__10_), .Y(_3677_) );
OR2X2 OR2X2_97 ( .A(_3677_), .B(_3676_), .Y(_3678_) );
OR2X2 OR2X2_98 ( .A(_3675_), .B(_3678_), .Y(_3679_) );
AND2X2 AND2X2_104 ( .A(_3386__bF_buf3), .B(gnd), .Y(_3680_) );
AND2X2 AND2X2_105 ( .A(_3388__bF_buf1), .B(REGs_REGS_3__10_), .Y(_3681_) );
AND2X2 AND2X2_106 ( .A(_3390__bF_buf1), .B(REGs_REGS_2__10_), .Y(_3682_) );
OR2X2 OR2X2_99 ( .A(_3681_), .B(_3682_), .Y(_3683_) );
OR2X2 OR2X2_100 ( .A(_3680_), .B(_3683_), .Y(_3684_) );
OR2X2 OR2X2_101 ( .A(_3684_), .B(_3679_), .Y(_3685_) );
AND2X2 AND2X2_107 ( .A(_2237_), .B(_3396__bF_buf3), .Y(_3686_) );
AND2X2 AND2X2_108 ( .A(_2241_), .B(_3398__bF_buf0), .Y(_3687_) );
OR2X2 OR2X2_102 ( .A(_3687_), .B(_3686_), .Y(_3688_) );
AND2X2 AND2X2_109 ( .A(_2246_), .B(_3401__bF_buf1), .Y(_3689_) );
AND2X2 AND2X2_110 ( .A(_2250_), .B(_3403__bF_buf4), .Y(_3690_) );
OR2X2 OR2X2_103 ( .A(_3690_), .B(_3689_), .Y(_3691_) );
OR2X2 OR2X2_104 ( .A(_3688_), .B(_3691_), .Y(_3692_) );
AND2X2 AND2X2_111 ( .A(_3409__bF_buf3), .B(_2256_), .Y(_3693_) );
AND2X2 AND2X2_112 ( .A(_3411__bF_buf3), .B(_2260_), .Y(_3694_) );
OR2X2 OR2X2_105 ( .A(_3693_), .B(_3694_), .Y(_3695_) );
AND2X2 AND2X2_113 ( .A(_2265_), .B(_3414__bF_buf1), .Y(_3696_) );
AND2X2 AND2X2_114 ( .A(_3416__bF_buf3), .B(_2269_), .Y(_3697_) );
OR2X2 OR2X2_106 ( .A(_3696_), .B(_3697_), .Y(_3698_) );
OR2X2 OR2X2_107 ( .A(_3698_), .B(_3695_), .Y(_3699_) );
OR2X2 OR2X2_108 ( .A(_3692_), .B(_3699_), .Y(_3700_) );
OR2X2 OR2X2_109 ( .A(_3685_), .B(_3700_), .Y(REG_A_10_) );
AND2X2 AND2X2_115 ( .A(_3369__bF_buf2), .B(REGs_REGS_4__11_), .Y(_3701_) );
AND2X2 AND2X2_116 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__11_), .Y(_3702_) );
OR2X2 OR2X2_110 ( .A(_3701_), .B(_3702_), .Y(_3703_) );
AND2X2 AND2X2_117 ( .A(_3378__bF_buf1), .B(REGs_REGS_6__11_), .Y(_3704_) );
AND2X2 AND2X2_118 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__11_), .Y(_3705_) );
OR2X2 OR2X2_111 ( .A(_3705_), .B(_3704_), .Y(_3706_) );
OR2X2 OR2X2_112 ( .A(_3703_), .B(_3706_), .Y(_3707_) );
AND2X2 AND2X2_119 ( .A(_3386__bF_buf0), .B(gnd), .Y(_3708_) );
AND2X2 AND2X2_120 ( .A(_3388__bF_buf2), .B(REGs_REGS_3__11_), .Y(_3709_) );
AND2X2 AND2X2_121 ( .A(_3390__bF_buf0), .B(REGs_REGS_2__11_), .Y(_3710_) );
OR2X2 OR2X2_113 ( .A(_3709_), .B(_3710_), .Y(_3711_) );
OR2X2 OR2X2_114 ( .A(_3708_), .B(_3711_), .Y(_3712_) );
OR2X2 OR2X2_115 ( .A(_3712_), .B(_3707_), .Y(_3713_) );
AND2X2 AND2X2_122 ( .A(_2289_), .B(_3396__bF_buf0), .Y(_3714_) );
AND2X2 AND2X2_123 ( .A(_2293_), .B(_3398__bF_buf4), .Y(_3715_) );
OR2X2 OR2X2_116 ( .A(_3715_), .B(_3714_), .Y(_3716_) );
AND2X2 AND2X2_124 ( .A(_2298_), .B(_3401__bF_buf4), .Y(_3717_) );
AND2X2 AND2X2_125 ( .A(_2302_), .B(_3403__bF_buf1), .Y(_3718_) );
OR2X2 OR2X2_117 ( .A(_3718_), .B(_3717_), .Y(_3719_) );
OR2X2 OR2X2_118 ( .A(_3716_), .B(_3719_), .Y(_3720_) );
AND2X2 AND2X2_126 ( .A(_3409__bF_buf2), .B(_2308_), .Y(_3721_) );
AND2X2 AND2X2_127 ( .A(_3411__bF_buf1), .B(_2312_), .Y(_3722_) );
OR2X2 OR2X2_119 ( .A(_3721_), .B(_3722_), .Y(_3723_) );
AND2X2 AND2X2_128 ( .A(_2317_), .B(_3414__bF_buf2), .Y(_3724_) );
AND2X2 AND2X2_129 ( .A(_3416__bF_buf1), .B(_2321_), .Y(_3725_) );
OR2X2 OR2X2_120 ( .A(_3724_), .B(_3725_), .Y(_3726_) );
OR2X2 OR2X2_121 ( .A(_3726_), .B(_3723_), .Y(_3727_) );
OR2X2 OR2X2_122 ( .A(_3720_), .B(_3727_), .Y(_3728_) );
OR2X2 OR2X2_123 ( .A(_3713_), .B(_3728_), .Y(REG_A_11_) );
AND2X2 AND2X2_130 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__12_), .Y(_3729_) );
AND2X2 AND2X2_131 ( .A(_3373__bF_buf1), .B(REGs_REGS_5__12_), .Y(_3730_) );
OR2X2 OR2X2_124 ( .A(_3729_), .B(_3730_), .Y(_3731_) );
AND2X2 AND2X2_132 ( .A(_3378__bF_buf0), .B(REGs_REGS_6__12_), .Y(_3732_) );
AND2X2 AND2X2_133 ( .A(_3381__bF_buf1), .B(REGs_REGS_7__12_), .Y(_3733_) );
OR2X2 OR2X2_125 ( .A(_3733_), .B(_3732_), .Y(_3734_) );
OR2X2 OR2X2_126 ( .A(_3731_), .B(_3734_), .Y(_3735_) );
AND2X2 AND2X2_134 ( .A(_3386__bF_buf4), .B(gnd), .Y(_3736_) );
AND2X2 AND2X2_135 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__12_), .Y(_3737_) );
AND2X2 AND2X2_136 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__12_), .Y(_3738_) );
OR2X2 OR2X2_127 ( .A(_3737_), .B(_3738_), .Y(_3739_) );
OR2X2 OR2X2_128 ( .A(_3736_), .B(_3739_), .Y(_3740_) );
OR2X2 OR2X2_129 ( .A(_3740_), .B(_3735_), .Y(_3741_) );
AND2X2 AND2X2_137 ( .A(_2341_), .B(_3396__bF_buf1), .Y(_3742_) );
AND2X2 AND2X2_138 ( .A(_2345_), .B(_3398__bF_buf3), .Y(_3743_) );
OR2X2 OR2X2_130 ( .A(_3743_), .B(_3742_), .Y(_3744_) );
AND2X2 AND2X2_139 ( .A(_2350_), .B(_3401__bF_buf3), .Y(_3745_) );
AND2X2 AND2X2_140 ( .A(_2354_), .B(_3403__bF_buf2), .Y(_3746_) );
OR2X2 OR2X2_131 ( .A(_3746_), .B(_3745_), .Y(_3747_) );
OR2X2 OR2X2_132 ( .A(_3744_), .B(_3747_), .Y(_3748_) );
AND2X2 AND2X2_141 ( .A(_3409__bF_buf1), .B(_2360_), .Y(_3749_) );
AND2X2 AND2X2_142 ( .A(_3411__bF_buf0), .B(_2364_), .Y(_3750_) );
OR2X2 OR2X2_133 ( .A(_3749_), .B(_3750_), .Y(_3751_) );
AND2X2 AND2X2_143 ( .A(_2369_), .B(_3414__bF_buf3), .Y(_3752_) );
AND2X2 AND2X2_144 ( .A(_3416__bF_buf0), .B(_2373_), .Y(_3753_) );
OR2X2 OR2X2_134 ( .A(_3752_), .B(_3753_), .Y(_3754_) );
OR2X2 OR2X2_135 ( .A(_3754_), .B(_3751_), .Y(_3755_) );
OR2X2 OR2X2_136 ( .A(_3748_), .B(_3755_), .Y(_3756_) );
OR2X2 OR2X2_137 ( .A(_3741_), .B(_3756_), .Y(REG_A_12_) );
AND2X2 AND2X2_145 ( .A(_3369__bF_buf0), .B(REGs_REGS_4__13_), .Y(_3757_) );
AND2X2 AND2X2_146 ( .A(_3373__bF_buf2), .B(REGs_REGS_5__13_), .Y(_3758_) );
OR2X2 OR2X2_138 ( .A(_3757_), .B(_3758_), .Y(_3759_) );
AND2X2 AND2X2_147 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__13_), .Y(_3760_) );
AND2X2 AND2X2_148 ( .A(_3381__bF_buf0), .B(REGs_REGS_7__13_), .Y(_3761_) );
OR2X2 OR2X2_139 ( .A(_3761_), .B(_3760_), .Y(_3762_) );
OR2X2 OR2X2_140 ( .A(_3759_), .B(_3762_), .Y(_3763_) );
AND2X2 AND2X2_149 ( .A(_3386__bF_buf1), .B(gnd), .Y(_3764_) );
AND2X2 AND2X2_150 ( .A(_3388__bF_buf0), .B(REGs_REGS_3__13_), .Y(_3765_) );
AND2X2 AND2X2_151 ( .A(_3390__bF_buf2), .B(REGs_REGS_2__13_), .Y(_3766_) );
OR2X2 OR2X2_141 ( .A(_3765_), .B(_3766_), .Y(_3767_) );
OR2X2 OR2X2_142 ( .A(_3764_), .B(_3767_), .Y(_3768_) );
OR2X2 OR2X2_143 ( .A(_3768_), .B(_3763_), .Y(_3769_) );
AND2X2 AND2X2_152 ( .A(_2393_), .B(_3396__bF_buf4), .Y(_3770_) );
AND2X2 AND2X2_153 ( .A(_2397_), .B(_3398__bF_buf2), .Y(_3771_) );
OR2X2 OR2X2_144 ( .A(_3771_), .B(_3770_), .Y(_3772_) );
AND2X2 AND2X2_154 ( .A(_2402_), .B(_3401__bF_buf2), .Y(_3773_) );
AND2X2 AND2X2_155 ( .A(_2406_), .B(_3403__bF_buf0), .Y(_3774_) );
OR2X2 OR2X2_145 ( .A(_3774_), .B(_3773_), .Y(_3775_) );
OR2X2 OR2X2_146 ( .A(_3772_), .B(_3775_), .Y(_3776_) );
AND2X2 AND2X2_156 ( .A(_3409__bF_buf0), .B(_2412_), .Y(_3777_) );
AND2X2 AND2X2_157 ( .A(_3411__bF_buf4), .B(_2416_), .Y(_3778_) );
OR2X2 OR2X2_147 ( .A(_3777_), .B(_3778_), .Y(_3779_) );
AND2X2 AND2X2_158 ( .A(_2421_), .B(_3414__bF_buf4), .Y(_3780_) );
AND2X2 AND2X2_159 ( .A(_3416__bF_buf4), .B(_2425_), .Y(_3781_) );
OR2X2 OR2X2_148 ( .A(_3780_), .B(_3781_), .Y(_3782_) );
OR2X2 OR2X2_149 ( .A(_3782_), .B(_3779_), .Y(_3783_) );
OR2X2 OR2X2_150 ( .A(_3776_), .B(_3783_), .Y(_3784_) );
OR2X2 OR2X2_151 ( .A(_3769_), .B(_3784_), .Y(REG_A_13_) );
AND2X2 AND2X2_160 ( .A(_3369__bF_buf1), .B(REGs_REGS_4__14_), .Y(_3785_) );
AND2X2 AND2X2_161 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__14_), .Y(_3786_) );
OR2X2 OR2X2_152 ( .A(_3785_), .B(_3786_), .Y(_3787_) );
AND2X2 AND2X2_162 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__14_), .Y(_3788_) );
AND2X2 AND2X2_163 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__14_), .Y(_3789_) );
OR2X2 OR2X2_153 ( .A(_3789_), .B(_3788_), .Y(_3790_) );
OR2X2 OR2X2_154 ( .A(_3787_), .B(_3790_), .Y(_3791_) );
AND2X2 AND2X2_164 ( .A(_3386__bF_buf3), .B(gnd), .Y(_3792_) );
AND2X2 AND2X2_165 ( .A(_3388__bF_buf1), .B(REGs_REGS_3__14_), .Y(_3793_) );
AND2X2 AND2X2_166 ( .A(_3390__bF_buf1), .B(REGs_REGS_2__14_), .Y(_3794_) );
OR2X2 OR2X2_155 ( .A(_3793_), .B(_3794_), .Y(_3795_) );
OR2X2 OR2X2_156 ( .A(_3792_), .B(_3795_), .Y(_3796_) );
OR2X2 OR2X2_157 ( .A(_3796_), .B(_3791_), .Y(_3797_) );
AND2X2 AND2X2_167 ( .A(_2445_), .B(_3396__bF_buf3), .Y(_3798_) );
AND2X2 AND2X2_168 ( .A(_2449_), .B(_3398__bF_buf0), .Y(_3799_) );
OR2X2 OR2X2_158 ( .A(_3799_), .B(_3798_), .Y(_3800_) );
AND2X2 AND2X2_169 ( .A(_2454_), .B(_3401__bF_buf1), .Y(_3801_) );
AND2X2 AND2X2_170 ( .A(_2458_), .B(_3403__bF_buf4), .Y(_3802_) );
OR2X2 OR2X2_159 ( .A(_3802_), .B(_3801_), .Y(_3803_) );
OR2X2 OR2X2_160 ( .A(_3800_), .B(_3803_), .Y(_3804_) );
AND2X2 AND2X2_171 ( .A(_3409__bF_buf3), .B(_2464_), .Y(_3805_) );
AND2X2 AND2X2_172 ( .A(_3411__bF_buf3), .B(_2468_), .Y(_3806_) );
OR2X2 OR2X2_161 ( .A(_3805_), .B(_3806_), .Y(_3807_) );
AND2X2 AND2X2_173 ( .A(_2473_), .B(_3414__bF_buf1), .Y(_3808_) );
AND2X2 AND2X2_174 ( .A(_3416__bF_buf3), .B(_2477_), .Y(_3809_) );
OR2X2 OR2X2_162 ( .A(_3808_), .B(_3809_), .Y(_3810_) );
OR2X2 OR2X2_163 ( .A(_3810_), .B(_3807_), .Y(_3811_) );
OR2X2 OR2X2_164 ( .A(_3804_), .B(_3811_), .Y(_3812_) );
OR2X2 OR2X2_165 ( .A(_3797_), .B(_3812_), .Y(REG_A_14_) );
AND2X2 AND2X2_175 ( .A(_3369__bF_buf1), .B(REGs_REGS_4__15_), .Y(_3813_) );
AND2X2 AND2X2_176 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__15_), .Y(_3814_) );
OR2X2 OR2X2_166 ( .A(_3813_), .B(_3814_), .Y(_3815_) );
AND2X2 AND2X2_177 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__15_), .Y(_3816_) );
AND2X2 AND2X2_178 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__15_), .Y(_3817_) );
OR2X2 OR2X2_167 ( .A(_3817_), .B(_3816_), .Y(_3818_) );
OR2X2 OR2X2_168 ( .A(_3815_), .B(_3818_), .Y(_3819_) );
AND2X2 AND2X2_179 ( .A(_3386__bF_buf3), .B(gnd), .Y(_3820_) );
AND2X2 AND2X2_180 ( .A(_3388__bF_buf1), .B(REGs_REGS_3__15_), .Y(_3821_) );
AND2X2 AND2X2_181 ( .A(_3390__bF_buf1), .B(REGs_REGS_2__15_), .Y(_3822_) );
OR2X2 OR2X2_169 ( .A(_3821_), .B(_3822_), .Y(_3823_) );
OR2X2 OR2X2_170 ( .A(_3820_), .B(_3823_), .Y(_3824_) );
OR2X2 OR2X2_171 ( .A(_3824_), .B(_3819_), .Y(_3825_) );
AND2X2 AND2X2_182 ( .A(_2497_), .B(_3396__bF_buf3), .Y(_3826_) );
AND2X2 AND2X2_183 ( .A(_2501_), .B(_3398__bF_buf0), .Y(_3827_) );
OR2X2 OR2X2_172 ( .A(_3827_), .B(_3826_), .Y(_3828_) );
AND2X2 AND2X2_184 ( .A(_2506_), .B(_3401__bF_buf1), .Y(_3829_) );
AND2X2 AND2X2_185 ( .A(_2510_), .B(_3403__bF_buf4), .Y(_3830_) );
OR2X2 OR2X2_173 ( .A(_3830_), .B(_3829_), .Y(_3831_) );
OR2X2 OR2X2_174 ( .A(_3828_), .B(_3831_), .Y(_3832_) );
AND2X2 AND2X2_186 ( .A(_3409__bF_buf3), .B(_2516_), .Y(_3833_) );
AND2X2 AND2X2_187 ( .A(_3411__bF_buf3), .B(_2520_), .Y(_3834_) );
OR2X2 OR2X2_175 ( .A(_3833_), .B(_3834_), .Y(_3835_) );
AND2X2 AND2X2_188 ( .A(_2525_), .B(_3414__bF_buf1), .Y(_3836_) );
AND2X2 AND2X2_189 ( .A(_3416__bF_buf3), .B(_2529_), .Y(_3837_) );
OR2X2 OR2X2_176 ( .A(_3836_), .B(_3837_), .Y(_3838_) );
OR2X2 OR2X2_177 ( .A(_3838_), .B(_3835_), .Y(_3839_) );
OR2X2 OR2X2_178 ( .A(_3832_), .B(_3839_), .Y(_3840_) );
OR2X2 OR2X2_179 ( .A(_3825_), .B(_3840_), .Y(REG_A_15_) );
AND2X2 AND2X2_190 ( .A(_3369__bF_buf1), .B(REGs_REGS_4__16_), .Y(_3841_) );
AND2X2 AND2X2_191 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__16_), .Y(_3842_) );
OR2X2 OR2X2_180 ( .A(_3841_), .B(_3842_), .Y(_3843_) );
AND2X2 AND2X2_192 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__16_), .Y(_3844_) );
AND2X2 AND2X2_193 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__16_), .Y(_3845_) );
OR2X2 OR2X2_181 ( .A(_3845_), .B(_3844_), .Y(_3846_) );
OR2X2 OR2X2_182 ( .A(_3843_), .B(_3846_), .Y(_3847_) );
AND2X2 AND2X2_194 ( .A(_3386__bF_buf3), .B(gnd), .Y(_3848_) );
AND2X2 AND2X2_195 ( .A(_3388__bF_buf1), .B(REGs_REGS_3__16_), .Y(_3849_) );
AND2X2 AND2X2_196 ( .A(_3390__bF_buf1), .B(REGs_REGS_2__16_), .Y(_3850_) );
OR2X2 OR2X2_183 ( .A(_3849_), .B(_3850_), .Y(_3851_) );
OR2X2 OR2X2_184 ( .A(_3848_), .B(_3851_), .Y(_3852_) );
OR2X2 OR2X2_185 ( .A(_3852_), .B(_3847_), .Y(_3853_) );
AND2X2 AND2X2_197 ( .A(_2549_), .B(_3396__bF_buf3), .Y(_3854_) );
AND2X2 AND2X2_198 ( .A(_2553_), .B(_3398__bF_buf0), .Y(_3855_) );
OR2X2 OR2X2_186 ( .A(_3855_), .B(_3854_), .Y(_3856_) );
AND2X2 AND2X2_199 ( .A(_2558_), .B(_3401__bF_buf1), .Y(_3857_) );
AND2X2 AND2X2_200 ( .A(_2562_), .B(_3403__bF_buf4), .Y(_3858_) );
OR2X2 OR2X2_187 ( .A(_3858_), .B(_3857_), .Y(_3859_) );
OR2X2 OR2X2_188 ( .A(_3856_), .B(_3859_), .Y(_3860_) );
AND2X2 AND2X2_201 ( .A(_3409__bF_buf3), .B(_2568_), .Y(_3861_) );
AND2X2 AND2X2_202 ( .A(_3411__bF_buf3), .B(_2572_), .Y(_3862_) );
OR2X2 OR2X2_189 ( .A(_3861_), .B(_3862_), .Y(_3863_) );
AND2X2 AND2X2_203 ( .A(_2577_), .B(_3414__bF_buf1), .Y(_3864_) );
AND2X2 AND2X2_204 ( .A(_3416__bF_buf3), .B(_2581_), .Y(_3865_) );
OR2X2 OR2X2_190 ( .A(_3864_), .B(_3865_), .Y(_3866_) );
OR2X2 OR2X2_191 ( .A(_3866_), .B(_3863_), .Y(_3867_) );
OR2X2 OR2X2_192 ( .A(_3860_), .B(_3867_), .Y(_3868_) );
OR2X2 OR2X2_193 ( .A(_3853_), .B(_3868_), .Y(REG_A_16_) );
AND2X2 AND2X2_205 ( .A(_3369__bF_buf0), .B(REGs_REGS_4__17_), .Y(_3869_) );
AND2X2 AND2X2_206 ( .A(_3373__bF_buf2), .B(REGs_REGS_5__17_), .Y(_3870_) );
OR2X2 OR2X2_194 ( .A(_3869_), .B(_3870_), .Y(_3871_) );
AND2X2 AND2X2_207 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__17_), .Y(_3872_) );
AND2X2 AND2X2_208 ( .A(_3381__bF_buf0), .B(REGs_REGS_7__17_), .Y(_3873_) );
OR2X2 OR2X2_195 ( .A(_3873_), .B(_3872_), .Y(_3874_) );
OR2X2 OR2X2_196 ( .A(_3871_), .B(_3874_), .Y(_3875_) );
AND2X2 AND2X2_209 ( .A(_3386__bF_buf1), .B(gnd), .Y(_3876_) );
AND2X2 AND2X2_210 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__17_), .Y(_3877_) );
AND2X2 AND2X2_211 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__17_), .Y(_3878_) );
OR2X2 OR2X2_197 ( .A(_3877_), .B(_3878_), .Y(_3879_) );
OR2X2 OR2X2_198 ( .A(_3876_), .B(_3879_), .Y(_3880_) );
OR2X2 OR2X2_199 ( .A(_3880_), .B(_3875_), .Y(_3881_) );
AND2X2 AND2X2_212 ( .A(_2601_), .B(_3396__bF_buf2), .Y(_3882_) );
AND2X2 AND2X2_213 ( .A(_2605_), .B(_3398__bF_buf1), .Y(_3883_) );
OR2X2 OR2X2_200 ( .A(_3883_), .B(_3882_), .Y(_3884_) );
AND2X2 AND2X2_214 ( .A(_2610_), .B(_3401__bF_buf0), .Y(_3885_) );
AND2X2 AND2X2_215 ( .A(_2614_), .B(_3403__bF_buf3), .Y(_3886_) );
OR2X2 OR2X2_201 ( .A(_3886_), .B(_3885_), .Y(_3887_) );
OR2X2 OR2X2_202 ( .A(_3884_), .B(_3887_), .Y(_3888_) );
AND2X2 AND2X2_216 ( .A(_3409__bF_buf4), .B(_2620_), .Y(_3889_) );
AND2X2 AND2X2_217 ( .A(_3411__bF_buf2), .B(_2624_), .Y(_3890_) );
OR2X2 OR2X2_203 ( .A(_3889_), .B(_3890_), .Y(_3891_) );
AND2X2 AND2X2_218 ( .A(_2629_), .B(_3414__bF_buf4), .Y(_3892_) );
AND2X2 AND2X2_219 ( .A(_3416__bF_buf4), .B(_2633_), .Y(_3893_) );
OR2X2 OR2X2_204 ( .A(_3892_), .B(_3893_), .Y(_3894_) );
OR2X2 OR2X2_205 ( .A(_3894_), .B(_3891_), .Y(_3895_) );
OR2X2 OR2X2_206 ( .A(_3888_), .B(_3895_), .Y(_3896_) );
OR2X2 OR2X2_207 ( .A(_3881_), .B(_3896_), .Y(REG_A_17_) );
AND2X2 AND2X2_220 ( .A(_3369__bF_buf2), .B(REGs_REGS_4__18_), .Y(_3897_) );
AND2X2 AND2X2_221 ( .A(_3373__bF_buf2), .B(REGs_REGS_5__18_), .Y(_3898_) );
OR2X2 OR2X2_208 ( .A(_3897_), .B(_3898_), .Y(_3899_) );
AND2X2 AND2X2_222 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__18_), .Y(_3900_) );
AND2X2 AND2X2_223 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__18_), .Y(_3901_) );
OR2X2 OR2X2_209 ( .A(_3901_), .B(_3900_), .Y(_3902_) );
OR2X2 OR2X2_210 ( .A(_3899_), .B(_3902_), .Y(_3903_) );
AND2X2 AND2X2_224 ( .A(_3386__bF_buf0), .B(gnd), .Y(_3904_) );
AND2X2 AND2X2_225 ( .A(_3388__bF_buf2), .B(REGs_REGS_3__18_), .Y(_3905_) );
AND2X2 AND2X2_226 ( .A(_3390__bF_buf0), .B(REGs_REGS_2__18_), .Y(_3906_) );
OR2X2 OR2X2_211 ( .A(_3905_), .B(_3906_), .Y(_3907_) );
OR2X2 OR2X2_212 ( .A(_3904_), .B(_3907_), .Y(_3908_) );
OR2X2 OR2X2_213 ( .A(_3908_), .B(_3903_), .Y(_3909_) );
AND2X2 AND2X2_227 ( .A(_2653_), .B(_3396__bF_buf3), .Y(_3910_) );
AND2X2 AND2X2_228 ( .A(_2657_), .B(_3398__bF_buf4), .Y(_3911_) );
OR2X2 OR2X2_214 ( .A(_3911_), .B(_3910_), .Y(_3912_) );
AND2X2 AND2X2_229 ( .A(_2662_), .B(_3401__bF_buf4), .Y(_3913_) );
AND2X2 AND2X2_230 ( .A(_2666_), .B(_3403__bF_buf1), .Y(_3914_) );
OR2X2 OR2X2_215 ( .A(_3914_), .B(_3913_), .Y(_3915_) );
OR2X2 OR2X2_216 ( .A(_3912_), .B(_3915_), .Y(_3916_) );
AND2X2 AND2X2_231 ( .A(_3409__bF_buf3), .B(_2672_), .Y(_3917_) );
AND2X2 AND2X2_232 ( .A(_3411__bF_buf3), .B(_2676_), .Y(_3918_) );
OR2X2 OR2X2_217 ( .A(_3917_), .B(_3918_), .Y(_3919_) );
AND2X2 AND2X2_233 ( .A(_2681_), .B(_3414__bF_buf1), .Y(_3920_) );
AND2X2 AND2X2_234 ( .A(_3416__bF_buf3), .B(_2685_), .Y(_3921_) );
OR2X2 OR2X2_218 ( .A(_3920_), .B(_3921_), .Y(_3922_) );
OR2X2 OR2X2_219 ( .A(_3922_), .B(_3919_), .Y(_3923_) );
OR2X2 OR2X2_220 ( .A(_3916_), .B(_3923_), .Y(_3924_) );
OR2X2 OR2X2_221 ( .A(_3909_), .B(_3924_), .Y(REG_A_18_) );
AND2X2 AND2X2_235 ( .A(_3369__bF_buf0), .B(REGs_REGS_4__19_), .Y(_3925_) );
AND2X2 AND2X2_236 ( .A(_3373__bF_buf2), .B(REGs_REGS_5__19_), .Y(_3926_) );
OR2X2 OR2X2_222 ( .A(_3925_), .B(_3926_), .Y(_3927_) );
AND2X2 AND2X2_237 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__19_), .Y(_3928_) );
AND2X2 AND2X2_238 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__19_), .Y(_3929_) );
OR2X2 OR2X2_223 ( .A(_3929_), .B(_3928_), .Y(_3930_) );
OR2X2 OR2X2_224 ( .A(_3927_), .B(_3930_), .Y(_3931_) );
AND2X2 AND2X2_239 ( .A(_3386__bF_buf0), .B(gnd), .Y(_3932_) );
AND2X2 AND2X2_240 ( .A(_3388__bF_buf0), .B(REGs_REGS_3__19_), .Y(_3933_) );
AND2X2 AND2X2_241 ( .A(_3390__bF_buf2), .B(REGs_REGS_2__19_), .Y(_3934_) );
OR2X2 OR2X2_225 ( .A(_3933_), .B(_3934_), .Y(_3935_) );
OR2X2 OR2X2_226 ( .A(_3932_), .B(_3935_), .Y(_3936_) );
OR2X2 OR2X2_227 ( .A(_3936_), .B(_3931_), .Y(_3937_) );
AND2X2 AND2X2_242 ( .A(_2705_), .B(_3396__bF_buf4), .Y(_3938_) );
AND2X2 AND2X2_243 ( .A(_2709_), .B(_3398__bF_buf2), .Y(_3939_) );
OR2X2 OR2X2_228 ( .A(_3939_), .B(_3938_), .Y(_3940_) );
AND2X2 AND2X2_244 ( .A(_2714_), .B(_3401__bF_buf2), .Y(_3941_) );
AND2X2 AND2X2_245 ( .A(_2718_), .B(_3403__bF_buf0), .Y(_3942_) );
OR2X2 OR2X2_229 ( .A(_3942_), .B(_3941_), .Y(_3943_) );
OR2X2 OR2X2_230 ( .A(_3940_), .B(_3943_), .Y(_3944_) );
AND2X2 AND2X2_246 ( .A(_3409__bF_buf0), .B(_2724_), .Y(_3945_) );
AND2X2 AND2X2_247 ( .A(_3411__bF_buf4), .B(_2728_), .Y(_3946_) );
OR2X2 OR2X2_231 ( .A(_3945_), .B(_3946_), .Y(_3947_) );
AND2X2 AND2X2_248 ( .A(_2733_), .B(_3414__bF_buf0), .Y(_3948_) );
AND2X2 AND2X2_249 ( .A(_3416__bF_buf2), .B(_2737_), .Y(_3949_) );
OR2X2 OR2X2_232 ( .A(_3948_), .B(_3949_), .Y(_3950_) );
OR2X2 OR2X2_233 ( .A(_3950_), .B(_3947_), .Y(_3951_) );
OR2X2 OR2X2_234 ( .A(_3944_), .B(_3951_), .Y(_3952_) );
OR2X2 OR2X2_235 ( .A(_3937_), .B(_3952_), .Y(REG_A_19_) );
AND2X2 AND2X2_250 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__20_), .Y(_3953_) );
AND2X2 AND2X2_251 ( .A(_3373__bF_buf0), .B(REGs_REGS_5__20_), .Y(_3954_) );
OR2X2 OR2X2_236 ( .A(_3953_), .B(_3954_), .Y(_3955_) );
AND2X2 AND2X2_252 ( .A(_3378__bF_buf2), .B(REGs_REGS_6__20_), .Y(_3956_) );
AND2X2 AND2X2_253 ( .A(_3381__bF_buf2), .B(REGs_REGS_7__20_), .Y(_3957_) );
OR2X2 OR2X2_237 ( .A(_3957_), .B(_3956_), .Y(_3958_) );
OR2X2 OR2X2_238 ( .A(_3955_), .B(_3958_), .Y(_3959_) );
AND2X2 AND2X2_254 ( .A(_3386__bF_buf4), .B(gnd), .Y(_3960_) );
AND2X2 AND2X2_255 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__20_), .Y(_3961_) );
AND2X2 AND2X2_256 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__20_), .Y(_3962_) );
OR2X2 OR2X2_239 ( .A(_3961_), .B(_3962_), .Y(_3963_) );
OR2X2 OR2X2_240 ( .A(_3960_), .B(_3963_), .Y(_3964_) );
OR2X2 OR2X2_241 ( .A(_3964_), .B(_3959_), .Y(_3965_) );
AND2X2 AND2X2_257 ( .A(_2757_), .B(_3396__bF_buf2), .Y(_3966_) );
AND2X2 AND2X2_258 ( .A(_2761_), .B(_3398__bF_buf1), .Y(_3967_) );
OR2X2 OR2X2_242 ( .A(_3967_), .B(_3966_), .Y(_3968_) );
AND2X2 AND2X2_259 ( .A(_2766_), .B(_3401__bF_buf0), .Y(_3969_) );
AND2X2 AND2X2_260 ( .A(_2770_), .B(_3403__bF_buf3), .Y(_3970_) );
OR2X2 OR2X2_243 ( .A(_3970_), .B(_3969_), .Y(_3971_) );
OR2X2 OR2X2_244 ( .A(_3968_), .B(_3971_), .Y(_3972_) );
AND2X2 AND2X2_261 ( .A(_3409__bF_buf4), .B(_2776_), .Y(_3973_) );
AND2X2 AND2X2_262 ( .A(_3411__bF_buf2), .B(_2780_), .Y(_3974_) );
OR2X2 OR2X2_245 ( .A(_3973_), .B(_3974_), .Y(_3975_) );
AND2X2 AND2X2_263 ( .A(_2785_), .B(_3414__bF_buf4), .Y(_3976_) );
AND2X2 AND2X2_264 ( .A(_3416__bF_buf4), .B(_2789_), .Y(_3977_) );
OR2X2 OR2X2_246 ( .A(_3976_), .B(_3977_), .Y(_3978_) );
OR2X2 OR2X2_247 ( .A(_3978_), .B(_3975_), .Y(_3979_) );
OR2X2 OR2X2_248 ( .A(_3972_), .B(_3979_), .Y(_3980_) );
OR2X2 OR2X2_249 ( .A(_3965_), .B(_3980_), .Y(REG_A_20_) );
AND2X2 AND2X2_265 ( .A(_3369__bF_buf2), .B(REGs_REGS_4__21_), .Y(_3981_) );
AND2X2 AND2X2_266 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__21_), .Y(_3982_) );
OR2X2 OR2X2_250 ( .A(_3981_), .B(_3982_), .Y(_3983_) );
AND2X2 AND2X2_267 ( .A(_3378__bF_buf1), .B(REGs_REGS_6__21_), .Y(_3984_) );
AND2X2 AND2X2_268 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__21_), .Y(_3985_) );
OR2X2 OR2X2_251 ( .A(_3985_), .B(_3984_), .Y(_3986_) );
OR2X2 OR2X2_252 ( .A(_3983_), .B(_3986_), .Y(_3987_) );
AND2X2 AND2X2_269 ( .A(_3386__bF_buf0), .B(gnd), .Y(_3988_) );
AND2X2 AND2X2_270 ( .A(_3388__bF_buf2), .B(REGs_REGS_3__21_), .Y(_3989_) );
AND2X2 AND2X2_271 ( .A(_3390__bF_buf0), .B(REGs_REGS_2__21_), .Y(_3990_) );
OR2X2 OR2X2_253 ( .A(_3989_), .B(_3990_), .Y(_3991_) );
OR2X2 OR2X2_254 ( .A(_3988_), .B(_3991_), .Y(_3992_) );
OR2X2 OR2X2_255 ( .A(_3992_), .B(_3987_), .Y(_3993_) );
AND2X2 AND2X2_272 ( .A(_2809_), .B(_3396__bF_buf4), .Y(_3994_) );
AND2X2 AND2X2_273 ( .A(_2813_), .B(_3398__bF_buf2), .Y(_3995_) );
OR2X2 OR2X2_256 ( .A(_3995_), .B(_3994_), .Y(_3996_) );
AND2X2 AND2X2_274 ( .A(_2818_), .B(_3401__bF_buf4), .Y(_3997_) );
AND2X2 AND2X2_275 ( .A(_2822_), .B(_3403__bF_buf4), .Y(_3998_) );
OR2X2 OR2X2_257 ( .A(_3998_), .B(_3997_), .Y(_3999_) );
OR2X2 OR2X2_258 ( .A(_3996_), .B(_3999_), .Y(_4000_) );
AND2X2 AND2X2_276 ( .A(_3409__bF_buf2), .B(_2828_), .Y(_4001_) );
AND2X2 AND2X2_277 ( .A(_3411__bF_buf1), .B(_2832_), .Y(_4002_) );
OR2X2 OR2X2_259 ( .A(_4001_), .B(_4002_), .Y(_4003_) );
AND2X2 AND2X2_278 ( .A(_2837_), .B(_3414__bF_buf1), .Y(_4004_) );
AND2X2 AND2X2_279 ( .A(_3416__bF_buf3), .B(_2841_), .Y(_4005_) );
OR2X2 OR2X2_260 ( .A(_4004_), .B(_4005_), .Y(_4006_) );
OR2X2 OR2X2_261 ( .A(_4006_), .B(_4003_), .Y(_4007_) );
OR2X2 OR2X2_262 ( .A(_4000_), .B(_4007_), .Y(_4008_) );
OR2X2 OR2X2_263 ( .A(_3993_), .B(_4008_), .Y(REG_A_21_) );
AND2X2 AND2X2_280 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__22_), .Y(_4009_) );
AND2X2 AND2X2_281 ( .A(_3373__bF_buf1), .B(REGs_REGS_5__22_), .Y(_4010_) );
OR2X2 OR2X2_264 ( .A(_4009_), .B(_4010_), .Y(_4011_) );
AND2X2 AND2X2_282 ( .A(_3378__bF_buf0), .B(REGs_REGS_6__22_), .Y(_4012_) );
AND2X2 AND2X2_283 ( .A(_3381__bF_buf1), .B(REGs_REGS_7__22_), .Y(_4013_) );
OR2X2 OR2X2_265 ( .A(_4013_), .B(_4012_), .Y(_4014_) );
OR2X2 OR2X2_266 ( .A(_4011_), .B(_4014_), .Y(_4015_) );
AND2X2 AND2X2_284 ( .A(_3386__bF_buf4), .B(gnd), .Y(_4016_) );
AND2X2 AND2X2_285 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__22_), .Y(_4017_) );
AND2X2 AND2X2_286 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__22_), .Y(_4018_) );
OR2X2 OR2X2_267 ( .A(_4017_), .B(_4018_), .Y(_4019_) );
OR2X2 OR2X2_268 ( .A(_4016_), .B(_4019_), .Y(_4020_) );
OR2X2 OR2X2_269 ( .A(_4020_), .B(_4015_), .Y(_4021_) );
AND2X2 AND2X2_287 ( .A(_2861_), .B(_3396__bF_buf1), .Y(_4022_) );
AND2X2 AND2X2_288 ( .A(_2865_), .B(_3398__bF_buf3), .Y(_4023_) );
OR2X2 OR2X2_270 ( .A(_4023_), .B(_4022_), .Y(_4024_) );
AND2X2 AND2X2_289 ( .A(_2870_), .B(_3401__bF_buf3), .Y(_4025_) );
AND2X2 AND2X2_290 ( .A(_2874_), .B(_3403__bF_buf2), .Y(_4026_) );
OR2X2 OR2X2_271 ( .A(_4026_), .B(_4025_), .Y(_4027_) );
OR2X2 OR2X2_272 ( .A(_4024_), .B(_4027_), .Y(_4028_) );
AND2X2 AND2X2_291 ( .A(_3409__bF_buf1), .B(_2880_), .Y(_4029_) );
AND2X2 AND2X2_292 ( .A(_3411__bF_buf0), .B(_2884_), .Y(_4030_) );
OR2X2 OR2X2_273 ( .A(_4029_), .B(_4030_), .Y(_4031_) );
AND2X2 AND2X2_293 ( .A(_2889_), .B(_3414__bF_buf3), .Y(_4032_) );
AND2X2 AND2X2_294 ( .A(_3416__bF_buf0), .B(_2893_), .Y(_4033_) );
OR2X2 OR2X2_274 ( .A(_4032_), .B(_4033_), .Y(_4034_) );
OR2X2 OR2X2_275 ( .A(_4034_), .B(_4031_), .Y(_4035_) );
OR2X2 OR2X2_276 ( .A(_4028_), .B(_4035_), .Y(_4036_) );
OR2X2 OR2X2_277 ( .A(_4021_), .B(_4036_), .Y(REG_A_22_) );
AND2X2 AND2X2_295 ( .A(_3369__bF_buf1), .B(REGs_REGS_4__23_), .Y(_4037_) );
AND2X2 AND2X2_296 ( .A(_3373__bF_buf4), .B(REGs_REGS_5__23_), .Y(_4038_) );
OR2X2 OR2X2_278 ( .A(_4037_), .B(_4038_), .Y(_4039_) );
AND2X2 AND2X2_297 ( .A(_3378__bF_buf4), .B(REGs_REGS_6__23_), .Y(_4040_) );
AND2X2 AND2X2_298 ( .A(_3381__bF_buf4), .B(REGs_REGS_7__23_), .Y(_4041_) );
OR2X2 OR2X2_279 ( .A(_4041_), .B(_4040_), .Y(_4042_) );
OR2X2 OR2X2_280 ( .A(_4039_), .B(_4042_), .Y(_4043_) );
AND2X2 AND2X2_299 ( .A(_3386__bF_buf3), .B(gnd), .Y(_4044_) );
AND2X2 AND2X2_300 ( .A(_3388__bF_buf1), .B(REGs_REGS_3__23_), .Y(_4045_) );
AND2X2 AND2X2_301 ( .A(_3390__bF_buf1), .B(REGs_REGS_2__23_), .Y(_4046_) );
OR2X2 OR2X2_281 ( .A(_4045_), .B(_4046_), .Y(_4047_) );
OR2X2 OR2X2_282 ( .A(_4044_), .B(_4047_), .Y(_4048_) );
OR2X2 OR2X2_283 ( .A(_4048_), .B(_4043_), .Y(_4049_) );
AND2X2 AND2X2_302 ( .A(_2913_), .B(_3396__bF_buf0), .Y(_4050_) );
AND2X2 AND2X2_303 ( .A(_2917_), .B(_3398__bF_buf4), .Y(_4051_) );
OR2X2 OR2X2_284 ( .A(_4051_), .B(_4050_), .Y(_4052_) );
AND2X2 AND2X2_304 ( .A(_2922_), .B(_3401__bF_buf4), .Y(_4053_) );
AND2X2 AND2X2_305 ( .A(_2926_), .B(_3403__bF_buf1), .Y(_4054_) );
OR2X2 OR2X2_285 ( .A(_4054_), .B(_4053_), .Y(_4055_) );
OR2X2 OR2X2_286 ( .A(_4052_), .B(_4055_), .Y(_4056_) );
AND2X2 AND2X2_306 ( .A(_3409__bF_buf3), .B(_2932_), .Y(_4057_) );
AND2X2 AND2X2_307 ( .A(_3411__bF_buf3), .B(_2936_), .Y(_4058_) );
OR2X2 OR2X2_287 ( .A(_4057_), .B(_4058_), .Y(_4059_) );
AND2X2 AND2X2_308 ( .A(_2941_), .B(_3414__bF_buf2), .Y(_4060_) );
AND2X2 AND2X2_309 ( .A(_3416__bF_buf2), .B(_2945_), .Y(_4061_) );
OR2X2 OR2X2_288 ( .A(_4060_), .B(_4061_), .Y(_4062_) );
OR2X2 OR2X2_289 ( .A(_4062_), .B(_4059_), .Y(_4063_) );
OR2X2 OR2X2_290 ( .A(_4056_), .B(_4063_), .Y(_4064_) );
OR2X2 OR2X2_291 ( .A(_4049_), .B(_4064_), .Y(REG_A_23_) );
AND2X2 AND2X2_310 ( .A(_3369__bF_buf0), .B(REGs_REGS_4__24_), .Y(_4065_) );
AND2X2 AND2X2_311 ( .A(_3373__bF_buf2), .B(REGs_REGS_5__24_), .Y(_4066_) );
OR2X2 OR2X2_292 ( .A(_4065_), .B(_4066_), .Y(_4067_) );
AND2X2 AND2X2_312 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__24_), .Y(_4068_) );
AND2X2 AND2X2_313 ( .A(_3381__bF_buf0), .B(REGs_REGS_7__24_), .Y(_4069_) );
OR2X2 OR2X2_293 ( .A(_4069_), .B(_4068_), .Y(_4070_) );
OR2X2 OR2X2_294 ( .A(_4067_), .B(_4070_), .Y(_4071_) );
AND2X2 AND2X2_314 ( .A(_3386__bF_buf1), .B(gnd), .Y(_4072_) );
AND2X2 AND2X2_315 ( .A(_3388__bF_buf0), .B(REGs_REGS_3__24_), .Y(_4073_) );
AND2X2 AND2X2_316 ( .A(_3390__bF_buf2), .B(REGs_REGS_2__24_), .Y(_4074_) );
OR2X2 OR2X2_295 ( .A(_4073_), .B(_4074_), .Y(_4075_) );
OR2X2 OR2X2_296 ( .A(_4072_), .B(_4075_), .Y(_4076_) );
OR2X2 OR2X2_297 ( .A(_4076_), .B(_4071_), .Y(_4077_) );
AND2X2 AND2X2_317 ( .A(_2965_), .B(_3396__bF_buf4), .Y(_4078_) );
AND2X2 AND2X2_318 ( .A(_2969_), .B(_3398__bF_buf2), .Y(_4079_) );
OR2X2 OR2X2_298 ( .A(_4079_), .B(_4078_), .Y(_4080_) );
AND2X2 AND2X2_319 ( .A(_2974_), .B(_3401__bF_buf2), .Y(_4081_) );
AND2X2 AND2X2_320 ( .A(_2978_), .B(_3403__bF_buf0), .Y(_4082_) );
OR2X2 OR2X2_299 ( .A(_4082_), .B(_4081_), .Y(_4083_) );
OR2X2 OR2X2_300 ( .A(_4080_), .B(_4083_), .Y(_4084_) );
AND2X2 AND2X2_321 ( .A(_3409__bF_buf0), .B(_2984_), .Y(_4085_) );
AND2X2 AND2X2_322 ( .A(_3411__bF_buf4), .B(_2988_), .Y(_4086_) );
OR2X2 OR2X2_301 ( .A(_4085_), .B(_4086_), .Y(_4087_) );
AND2X2 AND2X2_323 ( .A(_2993_), .B(_3414__bF_buf0), .Y(_4088_) );
AND2X2 AND2X2_324 ( .A(_3416__bF_buf1), .B(_2997_), .Y(_4089_) );
OR2X2 OR2X2_302 ( .A(_4088_), .B(_4089_), .Y(_4090_) );
OR2X2 OR2X2_303 ( .A(_4090_), .B(_4087_), .Y(_4091_) );
OR2X2 OR2X2_304 ( .A(_4084_), .B(_4091_), .Y(_4092_) );
OR2X2 OR2X2_305 ( .A(_4077_), .B(_4092_), .Y(REG_A_24_) );
AND2X2 AND2X2_325 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__25_), .Y(_4093_) );
AND2X2 AND2X2_326 ( .A(_3373__bF_buf0), .B(REGs_REGS_5__25_), .Y(_4094_) );
OR2X2 OR2X2_306 ( .A(_4093_), .B(_4094_), .Y(_4095_) );
AND2X2 AND2X2_327 ( .A(_3378__bF_buf2), .B(REGs_REGS_6__25_), .Y(_4096_) );
AND2X2 AND2X2_328 ( .A(_3381__bF_buf2), .B(REGs_REGS_7__25_), .Y(_4097_) );
OR2X2 OR2X2_307 ( .A(_4097_), .B(_4096_), .Y(_4098_) );
OR2X2 OR2X2_308 ( .A(_4095_), .B(_4098_), .Y(_4099_) );
AND2X2 AND2X2_329 ( .A(_3386__bF_buf2), .B(gnd), .Y(_4100_) );
AND2X2 AND2X2_330 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__25_), .Y(_4101_) );
AND2X2 AND2X2_331 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__25_), .Y(_4102_) );
OR2X2 OR2X2_309 ( .A(_4101_), .B(_4102_), .Y(_4103_) );
OR2X2 OR2X2_310 ( .A(_4100_), .B(_4103_), .Y(_4104_) );
OR2X2 OR2X2_311 ( .A(_4104_), .B(_4099_), .Y(_4105_) );
AND2X2 AND2X2_332 ( .A(_3017_), .B(_3396__bF_buf4), .Y(_4106_) );
AND2X2 AND2X2_333 ( .A(_3021_), .B(_3398__bF_buf1), .Y(_4107_) );
OR2X2 OR2X2_312 ( .A(_4107_), .B(_4106_), .Y(_4108_) );
AND2X2 AND2X2_334 ( .A(_3026_), .B(_3401__bF_buf0), .Y(_4109_) );
AND2X2 AND2X2_335 ( .A(_3030_), .B(_3403__bF_buf3), .Y(_4110_) );
OR2X2 OR2X2_313 ( .A(_4110_), .B(_4109_), .Y(_4111_) );
OR2X2 OR2X2_314 ( .A(_4108_), .B(_4111_), .Y(_4112_) );
AND2X2 AND2X2_336 ( .A(_3409__bF_buf4), .B(_3036_), .Y(_4113_) );
AND2X2 AND2X2_337 ( .A(_3411__bF_buf2), .B(_3040_), .Y(_4114_) );
OR2X2 OR2X2_315 ( .A(_4113_), .B(_4114_), .Y(_4115_) );
AND2X2 AND2X2_338 ( .A(_3045_), .B(_3414__bF_buf4), .Y(_4116_) );
AND2X2 AND2X2_339 ( .A(_3416__bF_buf4), .B(_3049_), .Y(_4117_) );
OR2X2 OR2X2_316 ( .A(_4116_), .B(_4117_), .Y(_4118_) );
OR2X2 OR2X2_317 ( .A(_4118_), .B(_4115_), .Y(_4119_) );
OR2X2 OR2X2_318 ( .A(_4112_), .B(_4119_), .Y(_4120_) );
OR2X2 OR2X2_319 ( .A(_4105_), .B(_4120_), .Y(REG_A_25_) );
AND2X2 AND2X2_340 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__26_), .Y(_4121_) );
AND2X2 AND2X2_341 ( .A(_3373__bF_buf1), .B(REGs_REGS_5__26_), .Y(_4122_) );
OR2X2 OR2X2_320 ( .A(_4121_), .B(_4122_), .Y(_4123_) );
AND2X2 AND2X2_342 ( .A(_3378__bF_buf0), .B(REGs_REGS_6__26_), .Y(_4124_) );
AND2X2 AND2X2_343 ( .A(_3381__bF_buf1), .B(REGs_REGS_7__26_), .Y(_4125_) );
OR2X2 OR2X2_321 ( .A(_4125_), .B(_4124_), .Y(_4126_) );
OR2X2 OR2X2_322 ( .A(_4123_), .B(_4126_), .Y(_4127_) );
AND2X2 AND2X2_344 ( .A(_3386__bF_buf4), .B(gnd), .Y(_4128_) );
AND2X2 AND2X2_345 ( .A(_3388__bF_buf4), .B(REGs_REGS_3__26_), .Y(_4129_) );
AND2X2 AND2X2_346 ( .A(_3390__bF_buf4), .B(REGs_REGS_2__26_), .Y(_4130_) );
OR2X2 OR2X2_323 ( .A(_4129_), .B(_4130_), .Y(_4131_) );
OR2X2 OR2X2_324 ( .A(_4128_), .B(_4131_), .Y(_4132_) );
OR2X2 OR2X2_325 ( .A(_4132_), .B(_4127_), .Y(_4133_) );
AND2X2 AND2X2_347 ( .A(_3069_), .B(_3396__bF_buf1), .Y(_4134_) );
AND2X2 AND2X2_348 ( .A(_3073_), .B(_3398__bF_buf3), .Y(_4135_) );
OR2X2 OR2X2_326 ( .A(_4135_), .B(_4134_), .Y(_4136_) );
AND2X2 AND2X2_349 ( .A(_3078_), .B(_3401__bF_buf3), .Y(_4137_) );
AND2X2 AND2X2_350 ( .A(_3082_), .B(_3403__bF_buf3), .Y(_4138_) );
OR2X2 OR2X2_327 ( .A(_4138_), .B(_4137_), .Y(_4139_) );
OR2X2 OR2X2_328 ( .A(_4136_), .B(_4139_), .Y(_4140_) );
AND2X2 AND2X2_351 ( .A(_3409__bF_buf4), .B(_3088_), .Y(_4141_) );
AND2X2 AND2X2_352 ( .A(_3411__bF_buf0), .B(_3092_), .Y(_4142_) );
OR2X2 OR2X2_329 ( .A(_4141_), .B(_4142_), .Y(_4143_) );
AND2X2 AND2X2_353 ( .A(_3097_), .B(_3414__bF_buf3), .Y(_4144_) );
AND2X2 AND2X2_354 ( .A(_3416__bF_buf0), .B(_3101_), .Y(_4145_) );
OR2X2 OR2X2_330 ( .A(_4144_), .B(_4145_), .Y(_4146_) );
OR2X2 OR2X2_331 ( .A(_4146_), .B(_4143_), .Y(_4147_) );
OR2X2 OR2X2_332 ( .A(_4140_), .B(_4147_), .Y(_4148_) );
OR2X2 OR2X2_333 ( .A(_4133_), .B(_4148_), .Y(REG_A_26_) );
AND2X2 AND2X2_355 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__27_), .Y(_4149_) );
AND2X2 AND2X2_356 ( .A(_3373__bF_buf0), .B(REGs_REGS_5__27_), .Y(_4150_) );
OR2X2 OR2X2_334 ( .A(_4149_), .B(_4150_), .Y(_4151_) );
AND2X2 AND2X2_357 ( .A(_3378__bF_buf2), .B(REGs_REGS_6__27_), .Y(_4152_) );
AND2X2 AND2X2_358 ( .A(_3381__bF_buf2), .B(REGs_REGS_7__27_), .Y(_4153_) );
OR2X2 OR2X2_335 ( .A(_4153_), .B(_4152_), .Y(_4154_) );
OR2X2 OR2X2_336 ( .A(_4151_), .B(_4154_), .Y(_4155_) );
AND2X2 AND2X2_359 ( .A(_3386__bF_buf2), .B(gnd), .Y(_4156_) );
AND2X2 AND2X2_360 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__27_), .Y(_4157_) );
AND2X2 AND2X2_361 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__27_), .Y(_4158_) );
OR2X2 OR2X2_337 ( .A(_4157_), .B(_4158_), .Y(_4159_) );
OR2X2 OR2X2_338 ( .A(_4156_), .B(_4159_), .Y(_4160_) );
OR2X2 OR2X2_339 ( .A(_4160_), .B(_4155_), .Y(_4161_) );
AND2X2 AND2X2_362 ( .A(_3121_), .B(_3396__bF_buf2), .Y(_4162_) );
AND2X2 AND2X2_363 ( .A(_3125_), .B(_3398__bF_buf1), .Y(_4163_) );
OR2X2 OR2X2_340 ( .A(_4163_), .B(_4162_), .Y(_4164_) );
AND2X2 AND2X2_364 ( .A(_3130_), .B(_3401__bF_buf0), .Y(_4165_) );
AND2X2 AND2X2_365 ( .A(_3134_), .B(_3403__bF_buf3), .Y(_4166_) );
OR2X2 OR2X2_341 ( .A(_4166_), .B(_4165_), .Y(_4167_) );
OR2X2 OR2X2_342 ( .A(_4164_), .B(_4167_), .Y(_4168_) );
AND2X2 AND2X2_366 ( .A(_3409__bF_buf4), .B(_3140_), .Y(_4169_) );
AND2X2 AND2X2_367 ( .A(_3411__bF_buf2), .B(_3144_), .Y(_4170_) );
OR2X2 OR2X2_343 ( .A(_4169_), .B(_4170_), .Y(_4171_) );
AND2X2 AND2X2_368 ( .A(_3149_), .B(_3414__bF_buf4), .Y(_4172_) );
AND2X2 AND2X2_369 ( .A(_3416__bF_buf4), .B(_3153_), .Y(_4173_) );
OR2X2 OR2X2_344 ( .A(_4172_), .B(_4173_), .Y(_4174_) );
OR2X2 OR2X2_345 ( .A(_4174_), .B(_4171_), .Y(_4175_) );
OR2X2 OR2X2_346 ( .A(_4168_), .B(_4175_), .Y(_4176_) );
OR2X2 OR2X2_347 ( .A(_4161_), .B(_4176_), .Y(REG_A_27_) );
AND2X2 AND2X2_370 ( .A(_3369__bF_buf2), .B(REGs_REGS_4__28_), .Y(_4177_) );
AND2X2 AND2X2_371 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__28_), .Y(_4178_) );
OR2X2 OR2X2_348 ( .A(_4177_), .B(_4178_), .Y(_4179_) );
AND2X2 AND2X2_372 ( .A(_3378__bF_buf1), .B(REGs_REGS_6__28_), .Y(_4180_) );
AND2X2 AND2X2_373 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__28_), .Y(_4181_) );
OR2X2 OR2X2_349 ( .A(_4181_), .B(_4180_), .Y(_4182_) );
OR2X2 OR2X2_350 ( .A(_4179_), .B(_4182_), .Y(_4183_) );
AND2X2 AND2X2_374 ( .A(_3386__bF_buf0), .B(gnd), .Y(_4184_) );
AND2X2 AND2X2_375 ( .A(_3388__bF_buf2), .B(REGs_REGS_3__28_), .Y(_4185_) );
AND2X2 AND2X2_376 ( .A(_3390__bF_buf0), .B(REGs_REGS_2__28_), .Y(_4186_) );
OR2X2 OR2X2_351 ( .A(_4185_), .B(_4186_), .Y(_4187_) );
OR2X2 OR2X2_352 ( .A(_4184_), .B(_4187_), .Y(_4188_) );
OR2X2 OR2X2_353 ( .A(_4188_), .B(_4183_), .Y(_4189_) );
AND2X2 AND2X2_377 ( .A(_3173_), .B(_3396__bF_buf0), .Y(_4190_) );
AND2X2 AND2X2_378 ( .A(_3177_), .B(_3398__bF_buf4), .Y(_4191_) );
OR2X2 OR2X2_354 ( .A(_4191_), .B(_4190_), .Y(_4192_) );
AND2X2 AND2X2_379 ( .A(_3182_), .B(_3401__bF_buf4), .Y(_4193_) );
AND2X2 AND2X2_380 ( .A(_3186_), .B(_3403__bF_buf1), .Y(_4194_) );
OR2X2 OR2X2_355 ( .A(_4194_), .B(_4193_), .Y(_4195_) );
OR2X2 OR2X2_356 ( .A(_4192_), .B(_4195_), .Y(_4196_) );
AND2X2 AND2X2_381 ( .A(_3409__bF_buf2), .B(_3192_), .Y(_4197_) );
AND2X2 AND2X2_382 ( .A(_3411__bF_buf1), .B(_3196_), .Y(_4198_) );
OR2X2 OR2X2_357 ( .A(_4197_), .B(_4198_), .Y(_4199_) );
AND2X2 AND2X2_383 ( .A(_3201_), .B(_3414__bF_buf2), .Y(_4200_) );
AND2X2 AND2X2_384 ( .A(_3416__bF_buf2), .B(_3205_), .Y(_4201_) );
OR2X2 OR2X2_358 ( .A(_4200_), .B(_4201_), .Y(_4202_) );
OR2X2 OR2X2_359 ( .A(_4202_), .B(_4199_), .Y(_4203_) );
OR2X2 OR2X2_360 ( .A(_4196_), .B(_4203_), .Y(_4204_) );
OR2X2 OR2X2_361 ( .A(_4189_), .B(_4204_), .Y(REG_A_28_) );
AND2X2 AND2X2_385 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__29_), .Y(_4205_) );
AND2X2 AND2X2_386 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__29_), .Y(_4206_) );
OR2X2 OR2X2_362 ( .A(_4205_), .B(_4206_), .Y(_4207_) );
AND2X2 AND2X2_387 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__29_), .Y(_4208_) );
AND2X2 AND2X2_388 ( .A(_3381__bF_buf0), .B(REGs_REGS_7__29_), .Y(_4209_) );
OR2X2 OR2X2_363 ( .A(_4209_), .B(_4208_), .Y(_4210_) );
OR2X2 OR2X2_364 ( .A(_4207_), .B(_4210_), .Y(_4211_) );
AND2X2 AND2X2_389 ( .A(_3386__bF_buf2), .B(gnd), .Y(_4212_) );
AND2X2 AND2X2_390 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__29_), .Y(_4213_) );
AND2X2 AND2X2_391 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__29_), .Y(_4214_) );
OR2X2 OR2X2_365 ( .A(_4213_), .B(_4214_), .Y(_4215_) );
OR2X2 OR2X2_366 ( .A(_4212_), .B(_4215_), .Y(_4216_) );
OR2X2 OR2X2_367 ( .A(_4216_), .B(_4211_), .Y(_4217_) );
AND2X2 AND2X2_392 ( .A(_3225_), .B(_3396__bF_buf4), .Y(_4218_) );
AND2X2 AND2X2_393 ( .A(_3229_), .B(_3398__bF_buf2), .Y(_4219_) );
OR2X2 OR2X2_368 ( .A(_4219_), .B(_4218_), .Y(_4220_) );
AND2X2 AND2X2_394 ( .A(_3234_), .B(_3401__bF_buf2), .Y(_4221_) );
AND2X2 AND2X2_395 ( .A(_3238_), .B(_3403__bF_buf0), .Y(_4222_) );
OR2X2 OR2X2_369 ( .A(_4222_), .B(_4221_), .Y(_4223_) );
OR2X2 OR2X2_370 ( .A(_4220_), .B(_4223_), .Y(_4224_) );
AND2X2 AND2X2_396 ( .A(_3409__bF_buf0), .B(_3244_), .Y(_4225_) );
AND2X2 AND2X2_397 ( .A(_3411__bF_buf4), .B(_3248_), .Y(_4226_) );
OR2X2 OR2X2_371 ( .A(_4225_), .B(_4226_), .Y(_4227_) );
AND2X2 AND2X2_398 ( .A(_3253_), .B(_3414__bF_buf0), .Y(_4228_) );
AND2X2 AND2X2_399 ( .A(_3416__bF_buf1), .B(_3257_), .Y(_4229_) );
OR2X2 OR2X2_372 ( .A(_4228_), .B(_4229_), .Y(_4230_) );
OR2X2 OR2X2_373 ( .A(_4230_), .B(_4227_), .Y(_4231_) );
OR2X2 OR2X2_374 ( .A(_4224_), .B(_4231_), .Y(_4232_) );
OR2X2 OR2X2_375 ( .A(_4217_), .B(_4232_), .Y(REG_A_29_) );
AND2X2 AND2X2_400 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__30_), .Y(_4233_) );
AND2X2 AND2X2_401 ( .A(_3373__bF_buf0), .B(REGs_REGS_5__30_), .Y(_4234_) );
OR2X2 OR2X2_376 ( .A(_4233_), .B(_4234_), .Y(_4235_) );
AND2X2 AND2X2_402 ( .A(_3378__bF_buf2), .B(REGs_REGS_6__30_), .Y(_4236_) );
AND2X2 AND2X2_403 ( .A(_3381__bF_buf2), .B(REGs_REGS_7__30_), .Y(_4237_) );
OR2X2 OR2X2_377 ( .A(_4237_), .B(_4236_), .Y(_4238_) );
OR2X2 OR2X2_378 ( .A(_4235_), .B(_4238_), .Y(_4239_) );
AND2X2 AND2X2_404 ( .A(_3386__bF_buf2), .B(gnd), .Y(_4240_) );
AND2X2 AND2X2_405 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__30_), .Y(_4241_) );
AND2X2 AND2X2_406 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__30_), .Y(_4242_) );
OR2X2 OR2X2_379 ( .A(_4241_), .B(_4242_), .Y(_4243_) );
OR2X2 OR2X2_380 ( .A(_4240_), .B(_4243_), .Y(_4244_) );
OR2X2 OR2X2_381 ( .A(_4244_), .B(_4239_), .Y(_4245_) );
AND2X2 AND2X2_407 ( .A(_3277_), .B(_3396__bF_buf2), .Y(_4246_) );
AND2X2 AND2X2_408 ( .A(_3281_), .B(_3398__bF_buf1), .Y(_4247_) );
OR2X2 OR2X2_382 ( .A(_4247_), .B(_4246_), .Y(_4248_) );
AND2X2 AND2X2_409 ( .A(_3286_), .B(_3401__bF_buf0), .Y(_4249_) );
AND2X2 AND2X2_410 ( .A(_3290_), .B(_3403__bF_buf3), .Y(_4250_) );
OR2X2 OR2X2_383 ( .A(_4250_), .B(_4249_), .Y(_4251_) );
OR2X2 OR2X2_384 ( .A(_4248_), .B(_4251_), .Y(_4252_) );
AND2X2 AND2X2_411 ( .A(_3409__bF_buf4), .B(_3296_), .Y(_4253_) );
AND2X2 AND2X2_412 ( .A(_3411__bF_buf2), .B(_3300_), .Y(_4254_) );
OR2X2 OR2X2_385 ( .A(_4253_), .B(_4254_), .Y(_4255_) );
AND2X2 AND2X2_413 ( .A(_3305_), .B(_3414__bF_buf4), .Y(_4256_) );
AND2X2 AND2X2_414 ( .A(_3416__bF_buf4), .B(_3309_), .Y(_4257_) );
OR2X2 OR2X2_386 ( .A(_4256_), .B(_4257_), .Y(_4258_) );
OR2X2 OR2X2_387 ( .A(_4258_), .B(_4255_), .Y(_4259_) );
OR2X2 OR2X2_388 ( .A(_4252_), .B(_4259_), .Y(_4260_) );
OR2X2 OR2X2_389 ( .A(_4245_), .B(_4260_), .Y(REG_A_30_) );
AND2X2 AND2X2_415 ( .A(_3369__bF_buf0), .B(REGs_REGS_4__31_), .Y(_4261_) );
AND2X2 AND2X2_416 ( .A(_3373__bF_buf2), .B(REGs_REGS_5__31_), .Y(_4262_) );
OR2X2 OR2X2_390 ( .A(_4261_), .B(_4262_), .Y(_4263_) );
AND2X2 AND2X2_417 ( .A(_3378__bF_buf3), .B(REGs_REGS_6__31_), .Y(_4264_) );
AND2X2 AND2X2_418 ( .A(_3381__bF_buf3), .B(REGs_REGS_7__31_), .Y(_4265_) );
OR2X2 OR2X2_391 ( .A(_4265_), .B(_4264_), .Y(_4266_) );
OR2X2 OR2X2_392 ( .A(_4263_), .B(_4266_), .Y(_4267_) );
AND2X2 AND2X2_419 ( .A(_3386__bF_buf1), .B(gnd), .Y(_4268_) );
AND2X2 AND2X2_420 ( .A(_3388__bF_buf0), .B(REGs_REGS_3__31_), .Y(_4269_) );
AND2X2 AND2X2_421 ( .A(_3390__bF_buf2), .B(REGs_REGS_2__31_), .Y(_4270_) );
OR2X2 OR2X2_393 ( .A(_4269_), .B(_4270_), .Y(_4271_) );
OR2X2 OR2X2_394 ( .A(_4268_), .B(_4271_), .Y(_4272_) );
OR2X2 OR2X2_395 ( .A(_4272_), .B(_4267_), .Y(_4273_) );
AND2X2 AND2X2_422 ( .A(_3329_), .B(_3396__bF_buf0), .Y(_4274_) );
AND2X2 AND2X2_423 ( .A(_3333_), .B(_3398__bF_buf4), .Y(_4275_) );
OR2X2 OR2X2_396 ( .A(_4275_), .B(_4274_), .Y(_4276_) );
AND2X2 AND2X2_424 ( .A(_3338_), .B(_3401__bF_buf4), .Y(_4277_) );
AND2X2 AND2X2_425 ( .A(_3342_), .B(_3403__bF_buf1), .Y(_4278_) );
OR2X2 OR2X2_397 ( .A(_4278_), .B(_4277_), .Y(_4279_) );
OR2X2 OR2X2_398 ( .A(_4276_), .B(_4279_), .Y(_4280_) );
AND2X2 AND2X2_426 ( .A(_3409__bF_buf0), .B(_3348_), .Y(_4281_) );
AND2X2 AND2X2_427 ( .A(_3411__bF_buf4), .B(_3352_), .Y(_4282_) );
OR2X2 OR2X2_399 ( .A(_4281_), .B(_4282_), .Y(_4283_) );
AND2X2 AND2X2_428 ( .A(_3357_), .B(_3414__bF_buf0), .Y(_4284_) );
AND2X2 AND2X2_429 ( .A(_3416__bF_buf1), .B(_3361_), .Y(_4285_) );
OR2X2 OR2X2_400 ( .A(_4284_), .B(_4285_), .Y(_4286_) );
OR2X2 OR2X2_401 ( .A(_4286_), .B(_4283_), .Y(_4287_) );
OR2X2 OR2X2_402 ( .A(_4280_), .B(_4287_), .Y(_4288_) );
OR2X2 OR2X2_403 ( .A(_4273_), .B(_4288_), .Y(REG_A_31_) );
INVX1 INVX1_1 ( .A(REG_RFD_exec_pipe_1_), .Y(_4289_) );
NAND3X1 NAND3X1_1 ( .A(_4289_), .B(REG_RFD_exec_pipe_0_), .C(REG_RFD_exec_pipe_2_), .Y(_4290_) );
NOR2X1 NOR2X1_1 ( .A(_1569_), .B(_4290_), .Y(_4291_) );
NAND2X1 NAND2X1_1 ( .A(REGs_USR_REGS_5__0_), .B(_1573__bF_buf16), .Y(_4292_) );
MUX2X1 MUX2X1_1 ( .A(_1567__bF_buf0), .B(_4292_), .S(_4291__bF_buf0), .Y(_927_) );
NAND2X1 NAND2X1_2 ( .A(REGs_USR_REGS_5__1_), .B(_1573__bF_buf68), .Y(_4293_) );
MUX2X1 MUX2X1_2 ( .A(_1575__bF_buf1), .B(_4293_), .S(_4291__bF_buf2), .Y(_928_) );
NAND2X1 NAND2X1_3 ( .A(REGs_USR_REGS_5__2_), .B(_1573__bF_buf23), .Y(_4294_) );
MUX2X1 MUX2X1_3 ( .A(_1577__bF_buf2), .B(_4294_), .S(_4291__bF_buf1), .Y(_929_) );
NAND2X1 NAND2X1_4 ( .A(REGs_USR_REGS_5__3_), .B(_1573__bF_buf59), .Y(_4295_) );
MUX2X1 MUX2X1_4 ( .A(_1579__bF_buf0), .B(_4295_), .S(_4291__bF_buf1), .Y(_930_) );
NAND2X1 NAND2X1_5 ( .A(REGs_USR_REGS_5__4_), .B(_1573__bF_buf46), .Y(_4296_) );
MUX2X1 MUX2X1_5 ( .A(_1581__bF_buf3), .B(_4296_), .S(_4291__bF_buf4), .Y(_931_) );
NAND2X1 NAND2X1_6 ( .A(REGs_USR_REGS_5__5_), .B(_1573__bF_buf14), .Y(_4297_) );
MUX2X1 MUX2X1_6 ( .A(_1583__bF_buf2), .B(_4297_), .S(_4291__bF_buf3), .Y(_932_) );
NAND2X1 NAND2X1_7 ( .A(REGs_USR_REGS_5__6_), .B(_1573__bF_buf27), .Y(_4298_) );
MUX2X1 MUX2X1_7 ( .A(_1585__bF_buf1), .B(_4298_), .S(_4291__bF_buf4), .Y(_933_) );
NAND2X1 NAND2X1_8 ( .A(REGs_USR_REGS_5__7_), .B(_1573__bF_buf48), .Y(_4299_) );
MUX2X1 MUX2X1_8 ( .A(_1587__bF_buf2), .B(_4299_), .S(_4291__bF_buf4), .Y(_934_) );
NAND2X1 NAND2X1_9 ( .A(REGs_USR_REGS_5__8_), .B(_1573__bF_buf31), .Y(_4300_) );
MUX2X1 MUX2X1_9 ( .A(_1589__bF_buf0), .B(_4300_), .S(_4291__bF_buf3), .Y(_935_) );
NAND2X1 NAND2X1_10 ( .A(REGs_USR_REGS_5__9_), .B(_1573__bF_buf60), .Y(_4301_) );
MUX2X1 MUX2X1_10 ( .A(_1591__bF_buf3), .B(_4301_), .S(_4291__bF_buf3), .Y(_936_) );
NAND2X1 NAND2X1_11 ( .A(REGs_USR_REGS_5__10_), .B(_1573__bF_buf44), .Y(_4302_) );
MUX2X1 MUX2X1_11 ( .A(_1593__bF_buf2), .B(_4302_), .S(_4291__bF_buf3), .Y(_937_) );
NAND2X1 NAND2X1_12 ( .A(REGs_USR_REGS_5__11_), .B(_1573__bF_buf68), .Y(_4303_) );
MUX2X1 MUX2X1_12 ( .A(_1595__bF_buf0), .B(_4303_), .S(_4291__bF_buf2), .Y(_938_) );
NAND2X1 NAND2X1_13 ( .A(REGs_USR_REGS_5__12_), .B(_1573__bF_buf72), .Y(_4304_) );
MUX2X1 MUX2X1_13 ( .A(_1597__bF_buf3), .B(_4304_), .S(_4291__bF_buf4), .Y(_939_) );
NAND2X1 NAND2X1_14 ( .A(REGs_USR_REGS_5__13_), .B(_1573__bF_buf1), .Y(_4305_) );
MUX2X1 MUX2X1_14 ( .A(_1599__bF_buf3), .B(_4305_), .S(_4291__bF_buf0), .Y(_940_) );
NAND2X1 NAND2X1_15 ( .A(REGs_USR_REGS_5__14_), .B(_1573__bF_buf44), .Y(_4306_) );
MUX2X1 MUX2X1_15 ( .A(_1601__bF_buf2), .B(_4306_), .S(_4291__bF_buf3), .Y(_941_) );
NAND2X1 NAND2X1_16 ( .A(REGs_USR_REGS_5__15_), .B(_1573__bF_buf53), .Y(_4307_) );
MUX2X1 MUX2X1_16 ( .A(_1603__bF_buf0), .B(_4307_), .S(_4291__bF_buf2), .Y(_942_) );
NAND2X1 NAND2X1_17 ( .A(REGs_USR_REGS_5__16_), .B(_1573__bF_buf63), .Y(_4308_) );
MUX2X1 MUX2X1_17 ( .A(_1605__bF_buf3), .B(_4308_), .S(_4291__bF_buf2), .Y(_943_) );
NAND2X1 NAND2X1_18 ( .A(REGs_USR_REGS_5__17_), .B(_1573__bF_buf23), .Y(_4309_) );
MUX2X1 MUX2X1_18 ( .A(_1607__bF_buf3), .B(_4309_), .S(_4291__bF_buf1), .Y(_944_) );
NAND2X1 NAND2X1_19 ( .A(REGs_USR_REGS_5__18_), .B(_1573__bF_buf68), .Y(_4310_) );
MUX2X1 MUX2X1_19 ( .A(_1609__bF_buf2), .B(_4310_), .S(_4291__bF_buf2), .Y(_945_) );
NAND2X1 NAND2X1_20 ( .A(REGs_USR_REGS_5__19_), .B(_1573__bF_buf40), .Y(_4311_) );
MUX2X1 MUX2X1_20 ( .A(_1611__bF_buf1), .B(_4311_), .S(_4291__bF_buf0), .Y(_946_) );
NAND2X1 NAND2X1_21 ( .A(REGs_USR_REGS_5__20_), .B(_1573__bF_buf7), .Y(_4312_) );
MUX2X1 MUX2X1_21 ( .A(_1613__bF_buf0), .B(_4312_), .S(_4291__bF_buf1), .Y(_947_) );
NAND2X1 NAND2X1_22 ( .A(REGs_USR_REGS_5__21_), .B(_1573__bF_buf1), .Y(_4313_) );
MUX2X1 MUX2X1_22 ( .A(_1615__bF_buf3), .B(_4313_), .S(_4291__bF_buf0), .Y(_948_) );
NAND2X1 NAND2X1_23 ( .A(REGs_USR_REGS_5__22_), .B(_1573__bF_buf72), .Y(_4314_) );
MUX2X1 MUX2X1_23 ( .A(_1617__bF_buf2), .B(_4314_), .S(_4291__bF_buf4), .Y(_949_) );
NAND2X1 NAND2X1_24 ( .A(REGs_USR_REGS_5__23_), .B(_1573__bF_buf52), .Y(_4315_) );
MUX2X1 MUX2X1_24 ( .A(_1619__bF_buf3), .B(_4315_), .S(_4291__bF_buf3), .Y(_950_) );
NAND2X1 NAND2X1_25 ( .A(REGs_USR_REGS_5__24_), .B(_1573__bF_buf71), .Y(_4316_) );
MUX2X1 MUX2X1_25 ( .A(_1621__bF_buf0), .B(_4316_), .S(_4291__bF_buf1), .Y(_951_) );
NAND2X1 NAND2X1_26 ( .A(REGs_USR_REGS_5__25_), .B(_1573__bF_buf31), .Y(_4317_) );
MUX2X1 MUX2X1_26 ( .A(_1623__bF_buf0), .B(_4317_), .S(_4291__bF_buf3), .Y(_952_) );
NAND2X1 NAND2X1_27 ( .A(REGs_USR_REGS_5__26_), .B(_1573__bF_buf48), .Y(_4318_) );
MUX2X1 MUX2X1_27 ( .A(_1625__bF_buf0), .B(_4318_), .S(_4291__bF_buf4), .Y(_953_) );
NAND2X1 NAND2X1_28 ( .A(REGs_USR_REGS_5__27_), .B(_1573__bF_buf56), .Y(_4319_) );
MUX2X1 MUX2X1_28 ( .A(_1627__bF_buf2), .B(_4319_), .S(_4291__bF_buf4), .Y(_954_) );
NAND2X1 NAND2X1_29 ( .A(REGs_USR_REGS_5__28_), .B(_1573__bF_buf50), .Y(_4320_) );
MUX2X1 MUX2X1_29 ( .A(_1629__bF_buf2), .B(_4320_), .S(_4291__bF_buf0), .Y(_955_) );
NAND2X1 NAND2X1_30 ( .A(REGs_USR_REGS_5__29_), .B(_1573__bF_buf1), .Y(_4321_) );
MUX2X1 MUX2X1_30 ( .A(_1631__bF_buf0), .B(_4321_), .S(_4291__bF_buf0), .Y(_956_) );
NAND2X1 NAND2X1_31 ( .A(REGs_USR_REGS_5__30_), .B(_1573__bF_buf23), .Y(_4322_) );
MUX2X1 MUX2X1_31 ( .A(_1633__bF_buf3), .B(_4322_), .S(_4291__bF_buf1), .Y(_957_) );
NAND2X1 NAND2X1_32 ( .A(REGs_USR_REGS_5__31_), .B(_1573__bF_buf53), .Y(_4323_) );
MUX2X1 MUX2X1_32 ( .A(_1635__bF_buf2), .B(_4323_), .S(_4291__bF_buf2), .Y(_958_) );
NAND3X1 NAND3X1_2 ( .A(REG_RFD_exec_pipe_0_), .B(REG_RFD_exec_pipe_1_), .C(REG_RFD_exec_pipe_2_), .Y(_4324_) );
NOR2X1 NOR2X1_2 ( .A(_1569_), .B(_4324_), .Y(_4325_) );
NAND2X1 NAND2X1_33 ( .A(REGs_USR_REGS_7__0_), .B(_1573__bF_buf39), .Y(_4326_) );
MUX2X1 MUX2X1_33 ( .A(_1567__bF_buf0), .B(_4326_), .S(_4325__bF_buf1), .Y(_959_) );
NAND2X1 NAND2X1_34 ( .A(REGs_USR_REGS_7__1_), .B(_1573__bF_buf14), .Y(_4327_) );
MUX2X1 MUX2X1_34 ( .A(_1575__bF_buf1), .B(_4327_), .S(_4325__bF_buf4), .Y(_960_) );
NAND2X1 NAND2X1_35 ( .A(REGs_USR_REGS_7__2_), .B(_1573__bF_buf34), .Y(_4328_) );
MUX2X1 MUX2X1_35 ( .A(_1577__bF_buf0), .B(_4328_), .S(_4325__bF_buf1), .Y(_961_) );
NAND2X1 NAND2X1_36 ( .A(REGs_USR_REGS_7__3_), .B(_1573__bF_buf23), .Y(_4329_) );
MUX2X1 MUX2X1_36 ( .A(_1579__bF_buf0), .B(_4329_), .S(_4325__bF_buf1), .Y(_962_) );
NAND2X1 NAND2X1_37 ( .A(REGs_USR_REGS_7__4_), .B(_1573__bF_buf27), .Y(_4330_) );
MUX2X1 MUX2X1_37 ( .A(_1581__bF_buf2), .B(_4330_), .S(_4325__bF_buf2), .Y(_963_) );
NAND2X1 NAND2X1_38 ( .A(REGs_USR_REGS_7__5_), .B(_1573__bF_buf45), .Y(_4331_) );
MUX2X1 MUX2X1_38 ( .A(_1583__bF_buf1), .B(_4331_), .S(_4325__bF_buf0), .Y(_964_) );
NAND2X1 NAND2X1_39 ( .A(REGs_USR_REGS_7__6_), .B(_1573__bF_buf72), .Y(_4332_) );
MUX2X1 MUX2X1_39 ( .A(_1585__bF_buf1), .B(_4332_), .S(_4325__bF_buf2), .Y(_965_) );
NAND2X1 NAND2X1_40 ( .A(REGs_USR_REGS_7__7_), .B(_1573__bF_buf71), .Y(_4333_) );
MUX2X1 MUX2X1_40 ( .A(_1587__bF_buf1), .B(_4333_), .S(_4325__bF_buf3), .Y(_966_) );
NAND2X1 NAND2X1_41 ( .A(REGs_USR_REGS_7__8_), .B(_1573__bF_buf24), .Y(_4334_) );
MUX2X1 MUX2X1_41 ( .A(_1589__bF_buf1), .B(_4334_), .S(_4325__bF_buf1), .Y(_967_) );
NAND2X1 NAND2X1_42 ( .A(REGs_USR_REGS_7__9_), .B(_1573__bF_buf45), .Y(_4335_) );
MUX2X1 MUX2X1_42 ( .A(_1591__bF_buf1), .B(_4335_), .S(_4325__bF_buf0), .Y(_968_) );
NAND2X1 NAND2X1_43 ( .A(REGs_USR_REGS_7__10_), .B(_1573__bF_buf44), .Y(_4336_) );
MUX2X1 MUX2X1_43 ( .A(_1593__bF_buf2), .B(_4336_), .S(_4325__bF_buf4), .Y(_969_) );
NAND2X1 NAND2X1_44 ( .A(REGs_USR_REGS_7__11_), .B(_1573__bF_buf14), .Y(_4337_) );
MUX2X1 MUX2X1_44 ( .A(_1595__bF_buf3), .B(_4337_), .S(_4325__bF_buf4), .Y(_970_) );
NAND2X1 NAND2X1_45 ( .A(REGs_USR_REGS_7__12_), .B(_1573__bF_buf72), .Y(_4338_) );
MUX2X1 MUX2X1_45 ( .A(_1597__bF_buf1), .B(_4338_), .S(_4325__bF_buf2), .Y(_971_) );
NAND2X1 NAND2X1_46 ( .A(REGs_USR_REGS_7__13_), .B(_1573__bF_buf30), .Y(_4339_) );
MUX2X1 MUX2X1_46 ( .A(_1599__bF_buf3), .B(_4339_), .S(_4325__bF_buf3), .Y(_972_) );
NAND2X1 NAND2X1_47 ( .A(REGs_USR_REGS_7__14_), .B(_1573__bF_buf60), .Y(_4340_) );
MUX2X1 MUX2X1_47 ( .A(_1601__bF_buf2), .B(_4340_), .S(_4325__bF_buf4), .Y(_973_) );
NAND2X1 NAND2X1_48 ( .A(REGs_USR_REGS_7__15_), .B(_1573__bF_buf53), .Y(_4341_) );
MUX2X1 MUX2X1_48 ( .A(_1603__bF_buf0), .B(_4341_), .S(_4325__bF_buf4), .Y(_974_) );
NAND2X1 NAND2X1_49 ( .A(REGs_USR_REGS_7__16_), .B(_1573__bF_buf45), .Y(_4342_) );
MUX2X1 MUX2X1_49 ( .A(_1605__bF_buf0), .B(_4342_), .S(_4325__bF_buf0), .Y(_975_) );
NAND2X1 NAND2X1_50 ( .A(REGs_USR_REGS_7__17_), .B(_1573__bF_buf47), .Y(_4343_) );
MUX2X1 MUX2X1_50 ( .A(_1607__bF_buf3), .B(_4343_), .S(_4325__bF_buf1), .Y(_976_) );
NAND2X1 NAND2X1_51 ( .A(REGs_USR_REGS_7__18_), .B(_1573__bF_buf60), .Y(_4344_) );
MUX2X1 MUX2X1_51 ( .A(_1609__bF_buf2), .B(_4344_), .S(_4325__bF_buf4), .Y(_977_) );
NAND2X1 NAND2X1_52 ( .A(REGs_USR_REGS_7__19_), .B(_1573__bF_buf30), .Y(_4345_) );
MUX2X1 MUX2X1_52 ( .A(_1611__bF_buf2), .B(_4345_), .S(_4325__bF_buf3), .Y(_978_) );
NAND2X1 NAND2X1_53 ( .A(REGs_USR_REGS_7__20_), .B(_1573__bF_buf7), .Y(_4346_) );
MUX2X1 MUX2X1_53 ( .A(_1613__bF_buf0), .B(_4346_), .S(_4325__bF_buf3), .Y(_979_) );
NAND2X1 NAND2X1_54 ( .A(REGs_USR_REGS_7__21_), .B(_1573__bF_buf45), .Y(_4347_) );
MUX2X1 MUX2X1_54 ( .A(_1615__bF_buf0), .B(_4347_), .S(_4325__bF_buf0), .Y(_980_) );
NAND2X1 NAND2X1_55 ( .A(REGs_USR_REGS_7__22_), .B(_1573__bF_buf46), .Y(_4348_) );
MUX2X1 MUX2X1_55 ( .A(_1617__bF_buf2), .B(_4348_), .S(_4325__bF_buf2), .Y(_981_) );
NAND2X1 NAND2X1_56 ( .A(REGs_USR_REGS_7__23_), .B(_1573__bF_buf14), .Y(_4349_) );
MUX2X1 MUX2X1_56 ( .A(_1619__bF_buf3), .B(_4349_), .S(_4325__bF_buf4), .Y(_982_) );
NAND2X1 NAND2X1_57 ( .A(REGs_USR_REGS_7__24_), .B(_1573__bF_buf30), .Y(_4350_) );
MUX2X1 MUX2X1_57 ( .A(_1621__bF_buf1), .B(_4350_), .S(_4325__bF_buf3), .Y(_983_) );
NAND2X1 NAND2X1_58 ( .A(REGs_USR_REGS_7__25_), .B(_1573__bF_buf71), .Y(_4351_) );
MUX2X1 MUX2X1_58 ( .A(_1623__bF_buf3), .B(_4351_), .S(_4325__bF_buf3), .Y(_984_) );
NAND2X1 NAND2X1_59 ( .A(REGs_USR_REGS_7__26_), .B(_1573__bF_buf46), .Y(_4352_) );
MUX2X1 MUX2X1_59 ( .A(_1625__bF_buf0), .B(_4352_), .S(_4325__bF_buf2), .Y(_985_) );
NAND2X1 NAND2X1_60 ( .A(REGs_USR_REGS_7__27_), .B(_1573__bF_buf47), .Y(_4353_) );
MUX2X1 MUX2X1_60 ( .A(_1627__bF_buf1), .B(_4353_), .S(_4325__bF_buf2), .Y(_986_) );
NAND2X1 NAND2X1_61 ( .A(REGs_USR_REGS_7__28_), .B(_1573__bF_buf21), .Y(_4354_) );
MUX2X1 MUX2X1_61 ( .A(_1629__bF_buf0), .B(_4354_), .S(_4325__bF_buf0), .Y(_987_) );
NAND2X1 NAND2X1_62 ( .A(REGs_USR_REGS_7__29_), .B(_1573__bF_buf58), .Y(_4355_) );
MUX2X1 MUX2X1_62 ( .A(_1631__bF_buf3), .B(_4355_), .S(_4325__bF_buf1), .Y(_988_) );
NAND2X1 NAND2X1_63 ( .A(REGs_USR_REGS_7__30_), .B(_1573__bF_buf6), .Y(_4356_) );
MUX2X1 MUX2X1_63 ( .A(_1633__bF_buf2), .B(_4356_), .S(_4325__bF_buf3), .Y(_989_) );
NAND2X1 NAND2X1_64 ( .A(REGs_USR_REGS_7__31_), .B(_1573__bF_buf20), .Y(_4357_) );
MUX2X1 MUX2X1_64 ( .A(_1635__bF_buf2), .B(_4357_), .S(_4325__bF_buf0), .Y(_990_) );
NAND3X1 NAND3X1_3 ( .A(REG_RFD_exec_pipe_3_), .B(REG_Write_wb_pipe), .C(INTERRUPT_flag_bF_buf15_bF_buf3), .Y(_4358_) );
INVX1 INVX1_2 ( .A(REG_RFD_exec_pipe_2_), .Y(_4359_) );
NAND3X1 NAND3X1_4 ( .A(_1570_), .B(REG_RFD_exec_pipe_1_), .C(_4359_), .Y(_4360_) );
NOR2X1 NOR2X1_3 ( .A(_4360_), .B(_4358_), .Y(_4361_) );
NAND2X1 NAND2X1_65 ( .A(REGs_FIRQ_REGS_2__0_), .B(_1573__bF_buf59), .Y(_4362_) );
MUX2X1 MUX2X1_65 ( .A(_1567__bF_buf3), .B(_4362_), .S(_4361__bF_buf4), .Y(_991_) );
NAND2X1 NAND2X1_66 ( .A(REGs_FIRQ_REGS_2__1_), .B(_1573__bF_buf24), .Y(_4363_) );
MUX2X1 MUX2X1_66 ( .A(_1575__bF_buf2), .B(_4363_), .S(_4361__bF_buf1), .Y(_992_) );
NAND2X1 NAND2X1_67 ( .A(REGs_FIRQ_REGS_2__2_), .B(_1573__bF_buf55), .Y(_4364_) );
MUX2X1 MUX2X1_67 ( .A(_1577__bF_buf3), .B(_4364_), .S(_4361__bF_buf2), .Y(_993_) );
NAND2X1 NAND2X1_68 ( .A(REGs_FIRQ_REGS_2__3_), .B(_1573__bF_buf59), .Y(_4365_) );
MUX2X1 MUX2X1_68 ( .A(_1579__bF_buf1), .B(_4365_), .S(_4361__bF_buf4), .Y(_994_) );
NAND2X1 NAND2X1_69 ( .A(REGs_FIRQ_REGS_2__4_), .B(_1573__bF_buf37), .Y(_4366_) );
MUX2X1 MUX2X1_69 ( .A(_1581__bF_buf0), .B(_4366_), .S(_4361__bF_buf2), .Y(_995_) );
NAND2X1 NAND2X1_70 ( .A(REGs_FIRQ_REGS_2__5_), .B(_1573__bF_buf24), .Y(_4367_) );
MUX2X1 MUX2X1_70 ( .A(_1583__bF_buf0), .B(_4367_), .S(_4361__bF_buf1), .Y(_996_) );
NAND2X1 NAND2X1_71 ( .A(REGs_FIRQ_REGS_2__6_), .B(_1573__bF_buf69), .Y(_4368_) );
MUX2X1 MUX2X1_71 ( .A(_1585__bF_buf2), .B(_4368_), .S(_4361__bF_buf2), .Y(_997_) );
NAND2X1 NAND2X1_72 ( .A(REGs_FIRQ_REGS_2__7_), .B(_1573__bF_buf35), .Y(_4369_) );
MUX2X1 MUX2X1_72 ( .A(_1587__bF_buf0), .B(_4369_), .S(_4361__bF_buf3), .Y(_998_) );
NAND2X1 NAND2X1_73 ( .A(REGs_FIRQ_REGS_2__8_), .B(_1573__bF_buf54), .Y(_4370_) );
MUX2X1 MUX2X1_73 ( .A(_1589__bF_buf1), .B(_4370_), .S(_4361__bF_buf1), .Y(_999_) );
NAND2X1 NAND2X1_74 ( .A(REGs_FIRQ_REGS_2__9_), .B(_1573__bF_buf13), .Y(_4371_) );
MUX2X1 MUX2X1_74 ( .A(_1591__bF_buf0), .B(_4371_), .S(_4361__bF_buf0), .Y(_1000_) );
NAND2X1 NAND2X1_75 ( .A(REGs_FIRQ_REGS_2__10_), .B(_1573__bF_buf20), .Y(_4372_) );
MUX2X1 MUX2X1_75 ( .A(_1593__bF_buf3), .B(_4372_), .S(_4361__bF_buf0), .Y(_1001_) );
NAND2X1 NAND2X1_76 ( .A(REGs_FIRQ_REGS_2__11_), .B(_1573__bF_buf39), .Y(_4373_) );
MUX2X1 MUX2X1_76 ( .A(_1595__bF_buf1), .B(_4373_), .S(_4361__bF_buf4), .Y(_1002_) );
NAND2X1 NAND2X1_77 ( .A(REGs_FIRQ_REGS_2__12_), .B(_1573__bF_buf37), .Y(_4374_) );
MUX2X1 MUX2X1_77 ( .A(_1597__bF_buf2), .B(_4374_), .S(_4361__bF_buf2), .Y(_1003_) );
NAND2X1 NAND2X1_78 ( .A(REGs_FIRQ_REGS_2__13_), .B(_1573__bF_buf35), .Y(_4375_) );
MUX2X1 MUX2X1_78 ( .A(_1599__bF_buf1), .B(_4375_), .S(_4361__bF_buf3), .Y(_1004_) );
NAND2X1 NAND2X1_79 ( .A(REGs_FIRQ_REGS_2__14_), .B(_1573__bF_buf63), .Y(_4376_) );
MUX2X1 MUX2X1_79 ( .A(_1601__bF_buf1), .B(_4376_), .S(_4361__bF_buf0), .Y(_1005_) );
NAND2X1 NAND2X1_80 ( .A(REGs_FIRQ_REGS_2__15_), .B(_1573__bF_buf77), .Y(_4377_) );
MUX2X1 MUX2X1_80 ( .A(_1603__bF_buf1), .B(_4377_), .S(_4361__bF_buf0), .Y(_1006_) );
NAND2X1 NAND2X1_81 ( .A(REGs_FIRQ_REGS_2__16_), .B(_1573__bF_buf63), .Y(_4378_) );
MUX2X1 MUX2X1_81 ( .A(_1605__bF_buf3), .B(_4378_), .S(_4361__bF_buf0), .Y(_1007_) );
NAND2X1 NAND2X1_82 ( .A(REGs_FIRQ_REGS_2__17_), .B(_1573__bF_buf12), .Y(_4379_) );
MUX2X1 MUX2X1_82 ( .A(_1607__bF_buf2), .B(_4379_), .S(_4361__bF_buf3), .Y(_1008_) );
NAND2X1 NAND2X1_83 ( .A(REGs_FIRQ_REGS_2__18_), .B(_1573__bF_buf20), .Y(_4380_) );
MUX2X1 MUX2X1_83 ( .A(_1609__bF_buf3), .B(_4380_), .S(_4361__bF_buf0), .Y(_1009_) );
NAND2X1 NAND2X1_84 ( .A(REGs_FIRQ_REGS_2__19_), .B(_1573__bF_buf54), .Y(_4381_) );
MUX2X1 MUX2X1_84 ( .A(_1611__bF_buf0), .B(_4381_), .S(_4361__bF_buf1), .Y(_1010_) );
NAND2X1 NAND2X1_85 ( .A(REGs_FIRQ_REGS_2__20_), .B(_1573__bF_buf5), .Y(_4382_) );
MUX2X1 MUX2X1_85 ( .A(_1613__bF_buf3), .B(_4382_), .S(_4361__bF_buf3), .Y(_1011_) );
NAND2X1 NAND2X1_86 ( .A(REGs_FIRQ_REGS_2__21_), .B(_1573__bF_buf24), .Y(_4383_) );
MUX2X1 MUX2X1_86 ( .A(_1615__bF_buf2), .B(_4383_), .S(_4361__bF_buf1), .Y(_1012_) );
NAND2X1 NAND2X1_87 ( .A(REGs_FIRQ_REGS_2__22_), .B(_1573__bF_buf37), .Y(_4384_) );
MUX2X1 MUX2X1_87 ( .A(_1617__bF_buf1), .B(_4384_), .S(_4361__bF_buf2), .Y(_1013_) );
NAND2X1 NAND2X1_88 ( .A(REGs_FIRQ_REGS_2__23_), .B(_1573__bF_buf24), .Y(_4385_) );
MUX2X1 MUX2X1_88 ( .A(_1619__bF_buf1), .B(_4385_), .S(_4361__bF_buf1), .Y(_1014_) );
NAND2X1 NAND2X1_89 ( .A(REGs_FIRQ_REGS_2__24_), .B(_1573__bF_buf5), .Y(_4386_) );
MUX2X1 MUX2X1_89 ( .A(_1621__bF_buf0), .B(_4386_), .S(_4361__bF_buf3), .Y(_1015_) );
NAND2X1 NAND2X1_90 ( .A(REGs_FIRQ_REGS_2__25_), .B(_1573__bF_buf12), .Y(_4387_) );
MUX2X1 MUX2X1_90 ( .A(_1623__bF_buf1), .B(_4387_), .S(_4361__bF_buf3), .Y(_1016_) );
NAND2X1 NAND2X1_91 ( .A(REGs_FIRQ_REGS_2__26_), .B(_1573__bF_buf69), .Y(_4388_) );
MUX2X1 MUX2X1_91 ( .A(_1625__bF_buf3), .B(_4388_), .S(_4361__bF_buf2), .Y(_1017_) );
NAND2X1 NAND2X1_92 ( .A(REGs_FIRQ_REGS_2__27_), .B(_1573__bF_buf17), .Y(_4389_) );
MUX2X1 MUX2X1_92 ( .A(_1627__bF_buf3), .B(_4389_), .S(_4361__bF_buf3), .Y(_1018_) );
NAND2X1 NAND2X1_93 ( .A(REGs_FIRQ_REGS_2__28_), .B(_1573__bF_buf16), .Y(_4390_) );
MUX2X1 MUX2X1_93 ( .A(_1629__bF_buf1), .B(_4390_), .S(_4361__bF_buf4), .Y(_1019_) );
NAND2X1 NAND2X1_94 ( .A(REGs_FIRQ_REGS_2__29_), .B(_1573__bF_buf58), .Y(_4391_) );
MUX2X1 MUX2X1_94 ( .A(_1631__bF_buf3), .B(_4391_), .S(_4361__bF_buf4), .Y(_1020_) );
NAND2X1 NAND2X1_95 ( .A(REGs_FIRQ_REGS_2__30_), .B(_1573__bF_buf61), .Y(_4392_) );
MUX2X1 MUX2X1_95 ( .A(_1633__bF_buf2), .B(_4392_), .S(_4361__bF_buf4), .Y(_1021_) );
NAND2X1 NAND2X1_96 ( .A(REGs_FIRQ_REGS_2__31_), .B(_1573__bF_buf59), .Y(_4393_) );
MUX2X1 MUX2X1_96 ( .A(_1635__bF_buf3), .B(_4393_), .S(_4361__bF_buf4), .Y(_1022_) );
NAND3X1 NAND3X1_5 ( .A(_4359_), .B(REG_RFD_exec_pipe_0_), .C(REG_RFD_exec_pipe_1_), .Y(_4394_) );
NOR2X1 NOR2X1_4 ( .A(_4394_), .B(_4358_), .Y(_4395_) );
NAND2X1 NAND2X1_97 ( .A(REGs_FIRQ_REGS_3__0_), .B(_1573__bF_buf76), .Y(_4396_) );
MUX2X1 MUX2X1_97 ( .A(_1567__bF_buf2), .B(_4396_), .S(_4395__bF_buf3), .Y(_1023_) );
NAND2X1 NAND2X1_98 ( .A(REGs_FIRQ_REGS_3__1_), .B(_1573__bF_buf16), .Y(_4397_) );
MUX2X1 MUX2X1_98 ( .A(_1575__bF_buf2), .B(_4397_), .S(_4395__bF_buf0), .Y(_1024_) );
NAND2X1 NAND2X1_99 ( .A(REGs_FIRQ_REGS_3__2_), .B(_1573__bF_buf55), .Y(_4398_) );
MUX2X1 MUX2X1_99 ( .A(_1577__bF_buf3), .B(_4398_), .S(_4395__bF_buf4), .Y(_1025_) );
NAND2X1 NAND2X1_100 ( .A(REGs_FIRQ_REGS_3__3_), .B(_1573__bF_buf59), .Y(_4399_) );
MUX2X1 MUX2X1_100 ( .A(_1579__bF_buf1), .B(_4399_), .S(_4395__bF_buf0), .Y(_1026_) );
NAND2X1 NAND2X1_101 ( .A(REGs_FIRQ_REGS_3__4_), .B(_1573__bF_buf38), .Y(_4400_) );
MUX2X1 MUX2X1_101 ( .A(_1581__bF_buf0), .B(_4400_), .S(_4395__bF_buf4), .Y(_1027_) );
NAND2X1 NAND2X1_102 ( .A(REGs_FIRQ_REGS_3__5_), .B(_1573__bF_buf31), .Y(_4401_) );
MUX2X1 MUX2X1_102 ( .A(_1583__bF_buf2), .B(_4401_), .S(_4395__bF_buf2), .Y(_1028_) );
NAND2X1 NAND2X1_103 ( .A(REGs_FIRQ_REGS_3__6_), .B(_1573__bF_buf37), .Y(_4402_) );
MUX2X1 MUX2X1_103 ( .A(_1585__bF_buf2), .B(_4402_), .S(_4395__bF_buf4), .Y(_1029_) );
NAND2X1 NAND2X1_104 ( .A(REGs_FIRQ_REGS_3__7_), .B(_1573__bF_buf35), .Y(_4403_) );
MUX2X1 MUX2X1_104 ( .A(_1587__bF_buf0), .B(_4403_), .S(_4395__bF_buf3), .Y(_1030_) );
NAND2X1 NAND2X1_105 ( .A(REGs_FIRQ_REGS_3__8_), .B(_1573__bF_buf28), .Y(_4404_) );
MUX2X1 MUX2X1_105 ( .A(_1589__bF_buf1), .B(_4404_), .S(_4395__bF_buf1), .Y(_1031_) );
NAND2X1 NAND2X1_106 ( .A(REGs_FIRQ_REGS_3__9_), .B(_1573__bF_buf31), .Y(_4405_) );
MUX2X1 MUX2X1_106 ( .A(_1591__bF_buf3), .B(_4405_), .S(_4395__bF_buf2), .Y(_1032_) );
NAND2X1 NAND2X1_107 ( .A(REGs_FIRQ_REGS_3__10_), .B(_1573__bF_buf74), .Y(_4406_) );
MUX2X1 MUX2X1_107 ( .A(_1593__bF_buf1), .B(_4406_), .S(_4395__bF_buf2), .Y(_1033_) );
NAND2X1 NAND2X1_108 ( .A(REGs_FIRQ_REGS_3__11_), .B(_1573__bF_buf8), .Y(_4407_) );
MUX2X1 MUX2X1_108 ( .A(_1595__bF_buf0), .B(_4407_), .S(_4395__bF_buf2), .Y(_1034_) );
NAND2X1 NAND2X1_109 ( .A(REGs_FIRQ_REGS_3__12_), .B(_1573__bF_buf57), .Y(_4408_) );
MUX2X1 MUX2X1_109 ( .A(_1597__bF_buf3), .B(_4408_), .S(_4395__bF_buf4), .Y(_1035_) );
NAND2X1 NAND2X1_110 ( .A(REGs_FIRQ_REGS_3__13_), .B(_1573__bF_buf35), .Y(_4409_) );
MUX2X1 MUX2X1_110 ( .A(_1599__bF_buf1), .B(_4409_), .S(_4395__bF_buf3), .Y(_1036_) );
NAND2X1 NAND2X1_111 ( .A(REGs_FIRQ_REGS_3__14_), .B(_1573__bF_buf77), .Y(_4410_) );
MUX2X1 MUX2X1_111 ( .A(_1601__bF_buf1), .B(_4410_), .S(_4395__bF_buf1), .Y(_1037_) );
NAND2X1 NAND2X1_112 ( .A(REGs_FIRQ_REGS_3__15_), .B(_1573__bF_buf50), .Y(_4411_) );
MUX2X1 MUX2X1_112 ( .A(_1603__bF_buf1), .B(_4411_), .S(_4395__bF_buf1), .Y(_1038_) );
NAND2X1 NAND2X1_113 ( .A(REGs_FIRQ_REGS_3__16_), .B(_1573__bF_buf31), .Y(_4412_) );
MUX2X1 MUX2X1_113 ( .A(_1605__bF_buf1), .B(_4412_), .S(_4395__bF_buf2), .Y(_1039_) );
NAND2X1 NAND2X1_114 ( .A(REGs_FIRQ_REGS_3__17_), .B(_1573__bF_buf12), .Y(_4413_) );
MUX2X1 MUX2X1_114 ( .A(_1607__bF_buf2), .B(_4413_), .S(_4395__bF_buf3), .Y(_1040_) );
NAND2X1 NAND2X1_115 ( .A(REGs_FIRQ_REGS_3__18_), .B(_1573__bF_buf77), .Y(_4414_) );
MUX2X1 MUX2X1_115 ( .A(_1609__bF_buf3), .B(_4414_), .S(_4395__bF_buf1), .Y(_1041_) );
NAND2X1 NAND2X1_116 ( .A(REGs_FIRQ_REGS_3__19_), .B(_1573__bF_buf54), .Y(_4415_) );
MUX2X1 MUX2X1_116 ( .A(_1611__bF_buf0), .B(_4415_), .S(_4395__bF_buf0), .Y(_1042_) );
NAND2X1 NAND2X1_117 ( .A(REGs_FIRQ_REGS_3__20_), .B(_1573__bF_buf5), .Y(_4416_) );
MUX2X1 MUX2X1_117 ( .A(_1613__bF_buf3), .B(_4416_), .S(_4395__bF_buf3), .Y(_1043_) );
NAND2X1 NAND2X1_118 ( .A(REGs_FIRQ_REGS_3__21_), .B(_1573__bF_buf8), .Y(_4417_) );
MUX2X1 MUX2X1_118 ( .A(_1615__bF_buf3), .B(_4417_), .S(_4395__bF_buf2), .Y(_1044_) );
NAND2X1 NAND2X1_119 ( .A(REGs_FIRQ_REGS_3__22_), .B(_1573__bF_buf37), .Y(_4418_) );
MUX2X1 MUX2X1_119 ( .A(_1617__bF_buf1), .B(_4418_), .S(_4395__bF_buf4), .Y(_1045_) );
NAND2X1 NAND2X1_120 ( .A(REGs_FIRQ_REGS_3__23_), .B(_1573__bF_buf26), .Y(_4419_) );
MUX2X1 MUX2X1_120 ( .A(_1619__bF_buf1), .B(_4419_), .S(_4395__bF_buf1), .Y(_1046_) );
NAND2X1 NAND2X1_121 ( .A(REGs_FIRQ_REGS_3__24_), .B(_1573__bF_buf18), .Y(_4420_) );
MUX2X1 MUX2X1_121 ( .A(_1621__bF_buf3), .B(_4420_), .S(_4395__bF_buf0), .Y(_1047_) );
NAND2X1 NAND2X1_122 ( .A(REGs_FIRQ_REGS_3__25_), .B(_1573__bF_buf35), .Y(_4421_) );
MUX2X1 MUX2X1_122 ( .A(_1623__bF_buf1), .B(_4421_), .S(_4395__bF_buf3), .Y(_1048_) );
NAND2X1 NAND2X1_123 ( .A(REGs_FIRQ_REGS_3__26_), .B(_1573__bF_buf69), .Y(_4422_) );
MUX2X1 MUX2X1_123 ( .A(_1625__bF_buf3), .B(_4422_), .S(_4395__bF_buf4), .Y(_1049_) );
NAND2X1 NAND2X1_124 ( .A(REGs_FIRQ_REGS_3__27_), .B(_1573__bF_buf12), .Y(_4423_) );
MUX2X1 MUX2X1_124 ( .A(_1627__bF_buf3), .B(_4423_), .S(_4395__bF_buf3), .Y(_1050_) );
NAND2X1 NAND2X1_125 ( .A(REGs_FIRQ_REGS_3__28_), .B(_1573__bF_buf26), .Y(_4424_) );
MUX2X1 MUX2X1_125 ( .A(_1629__bF_buf2), .B(_4424_), .S(_4395__bF_buf1), .Y(_1051_) );
NAND2X1 NAND2X1_126 ( .A(REGs_FIRQ_REGS_3__29_), .B(_1573__bF_buf58), .Y(_4425_) );
MUX2X1 MUX2X1_126 ( .A(_1631__bF_buf3), .B(_4425_), .S(_4395__bF_buf0), .Y(_1052_) );
NAND2X1 NAND2X1_127 ( .A(REGs_FIRQ_REGS_3__30_), .B(_1573__bF_buf55), .Y(_4426_) );
MUX2X1 MUX2X1_127 ( .A(_1633__bF_buf0), .B(_4426_), .S(_4395__bF_buf4), .Y(_1053_) );
NAND2X1 NAND2X1_128 ( .A(REGs_FIRQ_REGS_3__31_), .B(_1573__bF_buf54), .Y(_4427_) );
MUX2X1 MUX2X1_128 ( .A(_1635__bF_buf0), .B(_4427_), .S(_4395__bF_buf0), .Y(_1054_) );
INVX1 INVX1_3 ( .A(_4358_), .Y(_4428_) );
NAND3X1 NAND3X1_6 ( .A(_4428_), .B(REG_RFD_exec_pipe_0_), .C(_1641_), .Y(_4429_) );
NAND2X1 NAND2X1_129 ( .A(REGs_FIRQ_REGS_1__0_), .B(_1573__bF_buf76), .Y(_4430_) );
MUX2X1 MUX2X1_129 ( .A(_4430_), .B(_1567__bF_buf2), .S(_4429__bF_buf4), .Y(_1055_) );
NAND2X1 NAND2X1_130 ( .A(REGs_FIRQ_REGS_1__1_), .B(_1573__bF_buf8), .Y(_4431_) );
MUX2X1 MUX2X1_130 ( .A(_4431_), .B(_1575__bF_buf0), .S(_4429__bF_buf3), .Y(_1056_) );
NAND2X1 NAND2X1_131 ( .A(REGs_FIRQ_REGS_1__2_), .B(_1573__bF_buf7), .Y(_4432_) );
MUX2X1 MUX2X1_131 ( .A(_4432_), .B(_1577__bF_buf3), .S(_4429__bF_buf1), .Y(_1057_) );
NAND2X1 NAND2X1_132 ( .A(REGs_FIRQ_REGS_1__3_), .B(_1573__bF_buf48), .Y(_4433_) );
MUX2X1 MUX2X1_132 ( .A(_4433_), .B(_1579__bF_buf3), .S(_4429__bF_buf0), .Y(_1058_) );
NAND2X1 NAND2X1_133 ( .A(REGs_FIRQ_REGS_1__4_), .B(_1573__bF_buf27), .Y(_4434_) );
MUX2X1 MUX2X1_133 ( .A(_4434_), .B(_1581__bF_buf2), .S(_4429__bF_buf0), .Y(_1059_) );
NAND2X1 NAND2X1_134 ( .A(REGs_FIRQ_REGS_1__5_), .B(_1573__bF_buf13), .Y(_4435_) );
MUX2X1 MUX2X1_134 ( .A(_4435_), .B(_1583__bF_buf0), .S(_4429__bF_buf2), .Y(_1060_) );
NAND2X1 NAND2X1_135 ( .A(REGs_FIRQ_REGS_1__6_), .B(_1573__bF_buf11), .Y(_4436_) );
MUX2X1 MUX2X1_135 ( .A(_4436_), .B(_1585__bF_buf0), .S(_4429__bF_buf0), .Y(_1061_) );
NAND2X1 NAND2X1_136 ( .A(REGs_FIRQ_REGS_1__7_), .B(_1573__bF_buf17), .Y(_4437_) );
MUX2X1 MUX2X1_136 ( .A(_4437_), .B(_1587__bF_buf1), .S(_4429__bF_buf4), .Y(_1062_) );
NAND2X1 NAND2X1_137 ( .A(REGs_FIRQ_REGS_1__8_), .B(_1573__bF_buf18), .Y(_4438_) );
MUX2X1 MUX2X1_137 ( .A(_4438_), .B(_1589__bF_buf2), .S(_4429__bF_buf1), .Y(_1063_) );
NAND2X1 NAND2X1_138 ( .A(REGs_FIRQ_REGS_1__9_), .B(_1573__bF_buf77), .Y(_4439_) );
MUX2X1 MUX2X1_138 ( .A(_4439_), .B(_1591__bF_buf0), .S(_4429__bF_buf2), .Y(_1064_) );
NAND2X1 NAND2X1_139 ( .A(REGs_FIRQ_REGS_1__10_), .B(_1573__bF_buf74), .Y(_4440_) );
MUX2X1 MUX2X1_139 ( .A(_4440_), .B(_1593__bF_buf1), .S(_4429__bF_buf3), .Y(_1065_) );
NAND2X1 NAND2X1_140 ( .A(REGs_FIRQ_REGS_1__11_), .B(_1573__bF_buf28), .Y(_4441_) );
MUX2X1 MUX2X1_140 ( .A(_4441_), .B(_1595__bF_buf0), .S(_4429__bF_buf3), .Y(_1066_) );
NAND2X1 NAND2X1_141 ( .A(REGs_FIRQ_REGS_1__12_), .B(_1573__bF_buf11), .Y(_4442_) );
MUX2X1 MUX2X1_141 ( .A(_4442_), .B(_1597__bF_buf2), .S(_4429__bF_buf0), .Y(_1067_) );
NAND2X1 NAND2X1_142 ( .A(REGs_FIRQ_REGS_1__13_), .B(_1573__bF_buf76), .Y(_4443_) );
MUX2X1 MUX2X1_142 ( .A(_4443_), .B(_1599__bF_buf1), .S(_4429__bF_buf4), .Y(_1068_) );
NAND2X1 NAND2X1_143 ( .A(REGs_FIRQ_REGS_1__14_), .B(_1573__bF_buf20), .Y(_4444_) );
MUX2X1 MUX2X1_143 ( .A(_4444_), .B(_1601__bF_buf0), .S(_4429__bF_buf2), .Y(_1069_) );
NAND2X1 NAND2X1_144 ( .A(REGs_FIRQ_REGS_1__15_), .B(_1573__bF_buf50), .Y(_4445_) );
MUX2X1 MUX2X1_144 ( .A(_4445_), .B(_1603__bF_buf0), .S(_4429__bF_buf3), .Y(_1070_) );
NAND2X1 NAND2X1_145 ( .A(REGs_FIRQ_REGS_1__16_), .B(_1573__bF_buf74), .Y(_4446_) );
MUX2X1 MUX2X1_145 ( .A(_4446_), .B(_1605__bF_buf3), .S(_4429__bF_buf3), .Y(_1071_) );
NAND2X1 NAND2X1_146 ( .A(REGs_FIRQ_REGS_1__17_), .B(_1573__bF_buf6), .Y(_4447_) );
MUX2X1 MUX2X1_146 ( .A(_4447_), .B(_1607__bF_buf1), .S(_4429__bF_buf1), .Y(_1072_) );
NAND2X1 NAND2X1_147 ( .A(REGs_FIRQ_REGS_1__18_), .B(_1573__bF_buf20), .Y(_4448_) );
MUX2X1 MUX2X1_147 ( .A(_4448_), .B(_1609__bF_buf0), .S(_4429__bF_buf2), .Y(_1073_) );
NAND2X1 NAND2X1_148 ( .A(REGs_FIRQ_REGS_1__19_), .B(_1573__bF_buf54), .Y(_4449_) );
MUX2X1 MUX2X1_148 ( .A(_4449_), .B(_1611__bF_buf0), .S(_4429__bF_buf2), .Y(_1074_) );
NAND2X1 NAND2X1_149 ( .A(REGs_FIRQ_REGS_1__20_), .B(_1573__bF_buf76), .Y(_4450_) );
MUX2X1 MUX2X1_149 ( .A(_4450_), .B(_1613__bF_buf3), .S(_4429__bF_buf4), .Y(_1075_) );
NAND2X1 NAND2X1_150 ( .A(REGs_FIRQ_REGS_1__21_), .B(_1573__bF_buf28), .Y(_4451_) );
MUX2X1 MUX2X1_150 ( .A(_4451_), .B(_1615__bF_buf2), .S(_4429__bF_buf3), .Y(_1076_) );
NAND2X1 NAND2X1_151 ( .A(REGs_FIRQ_REGS_1__22_), .B(_1573__bF_buf11), .Y(_4452_) );
MUX2X1 MUX2X1_151 ( .A(_4452_), .B(_1617__bF_buf3), .S(_4429__bF_buf0), .Y(_1077_) );
NAND2X1 NAND2X1_152 ( .A(REGs_FIRQ_REGS_1__23_), .B(_1573__bF_buf13), .Y(_4453_) );
MUX2X1 MUX2X1_152 ( .A(_4453_), .B(_1619__bF_buf0), .S(_4429__bF_buf2), .Y(_1078_) );
NAND2X1 NAND2X1_153 ( .A(REGs_FIRQ_REGS_1__24_), .B(_1573__bF_buf30), .Y(_4454_) );
MUX2X1 MUX2X1_153 ( .A(_4454_), .B(_1621__bF_buf1), .S(_4429__bF_buf1), .Y(_1079_) );
NAND2X1 NAND2X1_154 ( .A(REGs_FIRQ_REGS_1__25_), .B(_1573__bF_buf76), .Y(_4455_) );
MUX2X1 MUX2X1_154 ( .A(_4455_), .B(_1623__bF_buf3), .S(_4429__bF_buf4), .Y(_1080_) );
NAND2X1 NAND2X1_155 ( .A(REGs_FIRQ_REGS_1__26_), .B(_1573__bF_buf38), .Y(_4456_) );
MUX2X1 MUX2X1_155 ( .A(_4456_), .B(_1625__bF_buf2), .S(_4429__bF_buf0), .Y(_1081_) );
NAND2X1 NAND2X1_156 ( .A(REGs_FIRQ_REGS_1__27_), .B(_1573__bF_buf17), .Y(_4457_) );
MUX2X1 MUX2X1_156 ( .A(_4457_), .B(_1627__bF_buf3), .S(_4429__bF_buf4), .Y(_1082_) );
NAND2X1 NAND2X1_157 ( .A(REGs_FIRQ_REGS_1__28_), .B(_1573__bF_buf28), .Y(_4458_) );
MUX2X1 MUX2X1_157 ( .A(_4458_), .B(_1629__bF_buf1), .S(_4429__bF_buf3), .Y(_1083_) );
NAND2X1 NAND2X1_158 ( .A(REGs_FIRQ_REGS_1__29_), .B(_1573__bF_buf18), .Y(_4459_) );
MUX2X1 MUX2X1_158 ( .A(_4459_), .B(_1631__bF_buf1), .S(_4429__bF_buf1), .Y(_1084_) );
NAND2X1 NAND2X1_159 ( .A(REGs_FIRQ_REGS_1__30_), .B(_1573__bF_buf22), .Y(_4460_) );
MUX2X1 MUX2X1_159 ( .A(_4460_), .B(_1633__bF_buf0), .S(_4429__bF_buf4), .Y(_1085_) );
NAND2X1 NAND2X1_160 ( .A(REGs_FIRQ_REGS_1__31_), .B(_1573__bF_buf32), .Y(_4461_) );
MUX2X1 MUX2X1_160 ( .A(_4461_), .B(_1635__bF_buf3), .S(_4429__bF_buf1), .Y(_1086_) );
NAND3X1 NAND3X1_7 ( .A(_4428_), .B(_1570_), .C(_1641_), .Y(_4462_) );
NAND2X1 NAND2X1_161 ( .A(REGs_FIRQ_REGS_0__0_), .B(_1573__bF_buf30), .Y(_4463_) );
MUX2X1 MUX2X1_161 ( .A(_4463_), .B(_1567__bF_buf2), .S(_4462__bF_buf4), .Y(_1087_) );
NAND2X1 NAND2X1_162 ( .A(REGs_FIRQ_REGS_0__1_), .B(_1573__bF_buf25), .Y(_4464_) );
MUX2X1 MUX2X1_162 ( .A(_4464_), .B(_1575__bF_buf2), .S(_4462__bF_buf1), .Y(_1088_) );
NAND2X1 NAND2X1_163 ( .A(REGs_FIRQ_REGS_0__2_), .B(_1573__bF_buf61), .Y(_4465_) );
MUX2X1 MUX2X1_163 ( .A(_4465_), .B(_1577__bF_buf2), .S(_4462__bF_buf4), .Y(_1089_) );
NAND2X1 NAND2X1_164 ( .A(REGs_FIRQ_REGS_0__3_), .B(_1573__bF_buf47), .Y(_4466_) );
MUX2X1 MUX2X1_164 ( .A(_4466_), .B(_1579__bF_buf3), .S(_4462__bF_buf3), .Y(_1090_) );
NAND2X1 NAND2X1_165 ( .A(REGs_FIRQ_REGS_0__4_), .B(_1573__bF_buf3), .Y(_4467_) );
MUX2X1 MUX2X1_165 ( .A(_4467_), .B(_1581__bF_buf1), .S(_4462__bF_buf3), .Y(_1091_) );
NAND2X1 NAND2X1_166 ( .A(REGs_FIRQ_REGS_0__5_), .B(_1573__bF_buf24), .Y(_4468_) );
MUX2X1 MUX2X1_166 ( .A(_4468_), .B(_1583__bF_buf0), .S(_4462__bF_buf1), .Y(_1092_) );
NAND2X1 NAND2X1_167 ( .A(REGs_FIRQ_REGS_0__6_), .B(_1573__bF_buf66), .Y(_4469_) );
MUX2X1 MUX2X1_167 ( .A(_4469_), .B(_1585__bF_buf0), .S(_4462__bF_buf3), .Y(_1093_) );
NAND2X1 NAND2X1_168 ( .A(REGs_FIRQ_REGS_0__7_), .B(_1573__bF_buf69), .Y(_4470_) );
MUX2X1 MUX2X1_168 ( .A(_4470_), .B(_1587__bF_buf2), .S(_4462__bF_buf4), .Y(_1094_) );
NAND2X1 NAND2X1_169 ( .A(REGs_FIRQ_REGS_0__8_), .B(_1573__bF_buf40), .Y(_4471_) );
MUX2X1 MUX2X1_169 ( .A(_4471_), .B(_1589__bF_buf2), .S(_4462__bF_buf0), .Y(_1095_) );
NAND2X1 NAND2X1_170 ( .A(REGs_FIRQ_REGS_0__9_), .B(_1573__bF_buf74), .Y(_4472_) );
MUX2X1 MUX2X1_170 ( .A(_4472_), .B(_1591__bF_buf3), .S(_4462__bF_buf2), .Y(_1096_) );
NAND2X1 NAND2X1_171 ( .A(REGs_FIRQ_REGS_0__10_), .B(_1573__bF_buf68), .Y(_4473_) );
MUX2X1 MUX2X1_171 ( .A(_4473_), .B(_1593__bF_buf1), .S(_4462__bF_buf2), .Y(_1097_) );
NAND2X1 NAND2X1_172 ( .A(REGs_FIRQ_REGS_0__11_), .B(_1573__bF_buf39), .Y(_4474_) );
MUX2X1 MUX2X1_172 ( .A(_4474_), .B(_1595__bF_buf1), .S(_4462__bF_buf0), .Y(_1098_) );
NAND2X1 NAND2X1_173 ( .A(REGs_FIRQ_REGS_0__12_), .B(_1573__bF_buf3), .Y(_4475_) );
MUX2X1 MUX2X1_173 ( .A(_4475_), .B(_1597__bF_buf1), .S(_4462__bF_buf3), .Y(_1099_) );
NAND2X1 NAND2X1_174 ( .A(REGs_FIRQ_REGS_0__13_), .B(_1573__bF_buf32), .Y(_4476_) );
MUX2X1 MUX2X1_174 ( .A(_4476_), .B(_1599__bF_buf0), .S(_4462__bF_buf0), .Y(_1100_) );
NAND2X1 NAND2X1_175 ( .A(REGs_FIRQ_REGS_0__14_), .B(_1573__bF_buf77), .Y(_4477_) );
MUX2X1 MUX2X1_175 ( .A(_4477_), .B(_1601__bF_buf0), .S(_4462__bF_buf1), .Y(_1101_) );
NAND2X1 NAND2X1_176 ( .A(REGs_FIRQ_REGS_0__15_), .B(_1573__bF_buf50), .Y(_4478_) );
MUX2X1 MUX2X1_176 ( .A(_4478_), .B(_1603__bF_buf1), .S(_4462__bF_buf2), .Y(_1102_) );
NAND2X1 NAND2X1_177 ( .A(REGs_FIRQ_REGS_0__16_), .B(_1573__bF_buf74), .Y(_4479_) );
MUX2X1 MUX2X1_177 ( .A(_4479_), .B(_1605__bF_buf3), .S(_4462__bF_buf2), .Y(_1103_) );
NAND2X1 NAND2X1_178 ( .A(REGs_FIRQ_REGS_0__17_), .B(_1573__bF_buf57), .Y(_4480_) );
MUX2X1 MUX2X1_178 ( .A(_4480_), .B(_1607__bF_buf1), .S(_4462__bF_buf4), .Y(_1104_) );
NAND2X1 NAND2X1_179 ( .A(REGs_FIRQ_REGS_0__18_), .B(_1573__bF_buf13), .Y(_4481_) );
MUX2X1 MUX2X1_179 ( .A(_4481_), .B(_1609__bF_buf0), .S(_4462__bF_buf1), .Y(_1105_) );
NAND2X1 NAND2X1_180 ( .A(REGs_FIRQ_REGS_0__19_), .B(_1573__bF_buf40), .Y(_4482_) );
MUX2X1 MUX2X1_180 ( .A(_4482_), .B(_1611__bF_buf2), .S(_4462__bF_buf0), .Y(_1106_) );
NAND2X1 NAND2X1_181 ( .A(REGs_FIRQ_REGS_0__20_), .B(_1573__bF_buf48), .Y(_4483_) );
MUX2X1 MUX2X1_181 ( .A(_4483_), .B(_1613__bF_buf2), .S(_4462__bF_buf3), .Y(_1107_) );
NAND2X1 NAND2X1_182 ( .A(REGs_FIRQ_REGS_0__21_), .B(_1573__bF_buf8), .Y(_4484_) );
MUX2X1 MUX2X1_182 ( .A(_4484_), .B(_1615__bF_buf2), .S(_4462__bF_buf2), .Y(_1108_) );
NAND2X1 NAND2X1_183 ( .A(REGs_FIRQ_REGS_0__22_), .B(_1573__bF_buf11), .Y(_4485_) );
MUX2X1 MUX2X1_183 ( .A(_4485_), .B(_1617__bF_buf3), .S(_4462__bF_buf3), .Y(_1109_) );
NAND2X1 NAND2X1_184 ( .A(REGs_FIRQ_REGS_0__23_), .B(_1573__bF_buf68), .Y(_4486_) );
MUX2X1 MUX2X1_184 ( .A(_4486_), .B(_1619__bF_buf3), .S(_4462__bF_buf2), .Y(_1110_) );
NAND2X1 NAND2X1_185 ( .A(REGs_FIRQ_REGS_0__24_), .B(_1573__bF_buf32), .Y(_4487_) );
MUX2X1 MUX2X1_185 ( .A(_4487_), .B(_1621__bF_buf3), .S(_4462__bF_buf0), .Y(_1111_) );
NAND2X1 NAND2X1_186 ( .A(REGs_FIRQ_REGS_0__25_), .B(_1573__bF_buf76), .Y(_4488_) );
MUX2X1 MUX2X1_186 ( .A(_4488_), .B(_1623__bF_buf3), .S(_4462__bF_buf4), .Y(_1112_) );
NAND2X1 NAND2X1_187 ( .A(REGs_FIRQ_REGS_0__26_), .B(_1573__bF_buf69), .Y(_4489_) );
MUX2X1 MUX2X1_187 ( .A(_4489_), .B(_1625__bF_buf3), .S(_4462__bF_buf4), .Y(_1113_) );
NAND2X1 NAND2X1_188 ( .A(REGs_FIRQ_REGS_0__27_), .B(_1573__bF_buf57), .Y(_4490_) );
MUX2X1 MUX2X1_188 ( .A(_4490_), .B(_1627__bF_buf2), .S(_4462__bF_buf4), .Y(_1114_) );
NAND2X1 NAND2X1_189 ( .A(REGs_FIRQ_REGS_0__28_), .B(_1573__bF_buf13), .Y(_4491_) );
MUX2X1 MUX2X1_189 ( .A(_4491_), .B(_1629__bF_buf2), .S(_4462__bF_buf1), .Y(_1115_) );
NAND2X1 NAND2X1_190 ( .A(REGs_FIRQ_REGS_0__29_), .B(_1573__bF_buf58), .Y(_4492_) );
MUX2X1 MUX2X1_190 ( .A(_4492_), .B(_1631__bF_buf3), .S(_4462__bF_buf1), .Y(_1116_) );
NAND2X1 NAND2X1_191 ( .A(REGs_FIRQ_REGS_0__30_), .B(_1573__bF_buf56), .Y(_4493_) );
MUX2X1 MUX2X1_191 ( .A(_4493_), .B(_1633__bF_buf3), .S(_4462__bF_buf3), .Y(_1117_) );
NAND2X1 NAND2X1_192 ( .A(REGs_FIRQ_REGS_0__31_), .B(_1573__bF_buf18), .Y(_4494_) );
MUX2X1 MUX2X1_192 ( .A(_4494_), .B(_1635__bF_buf3), .S(_4462__bF_buf0), .Y(_1118_) );
NAND3X1 NAND3X1_8 ( .A(_1637_), .B(REG_Write_wb_pipe), .C(_1640_), .Y(_4495_) );
NOR2X1 NOR2X1_5 ( .A(_1571_), .B(_4495_), .Y(_4496_) );
NAND2X1 NAND2X1_193 ( .A(REGs_REGS_6__0_), .B(_1573__bF_buf2), .Y(_4497_) );
MUX2X1 MUX2X1_193 ( .A(_1567__bF_buf3), .B(_4497_), .S(_4496__bF_buf3), .Y(_1119_) );
NAND2X1 NAND2X1_194 ( .A(REGs_REGS_6__1_), .B(_1573__bF_buf2), .Y(_4498_) );
MUX2X1 MUX2X1_194 ( .A(_1575__bF_buf3), .B(_4498_), .S(_4496__bF_buf3), .Y(_1120_) );
NAND2X1 NAND2X1_195 ( .A(REGs_REGS_6__2_), .B(_1573__bF_buf36), .Y(_4499_) );
MUX2X1 MUX2X1_195 ( .A(_1577__bF_buf1), .B(_4499_), .S(_4496__bF_buf2), .Y(_1121_) );
NAND2X1 NAND2X1_196 ( .A(REGs_REGS_6__3_), .B(_1573__bF_buf36), .Y(_4500_) );
MUX2X1 MUX2X1_196 ( .A(_1579__bF_buf2), .B(_4500_), .S(_4496__bF_buf2), .Y(_1122_) );
NAND2X1 NAND2X1_197 ( .A(REGs_REGS_6__4_), .B(_1573__bF_buf15), .Y(_4501_) );
MUX2X1 MUX2X1_197 ( .A(_1581__bF_buf3), .B(_4501_), .S(_4496__bF_buf4), .Y(_1123_) );
NAND2X1 NAND2X1_198 ( .A(REGs_REGS_6__5_), .B(_1573__bF_buf2), .Y(_4502_) );
MUX2X1 MUX2X1_198 ( .A(_1583__bF_buf3), .B(_4502_), .S(_4496__bF_buf3), .Y(_1124_) );
NAND2X1 NAND2X1_199 ( .A(REGs_REGS_6__6_), .B(_1573__bF_buf15), .Y(_4503_) );
MUX2X1 MUX2X1_199 ( .A(_1585__bF_buf3), .B(_4503_), .S(_4496__bF_buf4), .Y(_1125_) );
NAND2X1 NAND2X1_200 ( .A(REGs_REGS_6__7_), .B(_1573__bF_buf66), .Y(_4504_) );
MUX2X1 MUX2X1_200 ( .A(_1587__bF_buf3), .B(_4504_), .S(_4496__bF_buf4), .Y(_1126_) );
NAND2X1 NAND2X1_201 ( .A(REGs_REGS_6__8_), .B(_1573__bF_buf25), .Y(_4505_) );
MUX2X1 MUX2X1_201 ( .A(_1589__bF_buf3), .B(_4505_), .S(_4496__bF_buf3), .Y(_1127_) );
NAND2X1 NAND2X1_202 ( .A(REGs_REGS_6__9_), .B(_1573__bF_buf29), .Y(_4506_) );
MUX2X1 MUX2X1_202 ( .A(_1591__bF_buf2), .B(_4506_), .S(_4496__bF_buf0), .Y(_1128_) );
NAND2X1 NAND2X1_203 ( .A(REGs_REGS_6__10_), .B(_1573__bF_buf62), .Y(_4507_) );
MUX2X1 MUX2X1_203 ( .A(_1593__bF_buf0), .B(_4507_), .S(_4496__bF_buf0), .Y(_1129_) );
NAND2X1 NAND2X1_204 ( .A(REGs_REGS_6__11_), .B(_1573__bF_buf73), .Y(_4508_) );
MUX2X1 MUX2X1_204 ( .A(_1595__bF_buf2), .B(_4508_), .S(_4496__bF_buf3), .Y(_1130_) );
NAND2X1 NAND2X1_205 ( .A(REGs_REGS_6__12_), .B(_1573__bF_buf66), .Y(_4509_) );
MUX2X1 MUX2X1_205 ( .A(_1597__bF_buf0), .B(_4509_), .S(_4496__bF_buf4), .Y(_1131_) );
NAND2X1 NAND2X1_206 ( .A(REGs_REGS_6__13_), .B(_1573__bF_buf51), .Y(_4510_) );
MUX2X1 MUX2X1_206 ( .A(_1599__bF_buf2), .B(_4510_), .S(_4496__bF_buf2), .Y(_1132_) );
NAND2X1 NAND2X1_207 ( .A(REGs_REGS_6__14_), .B(_1573__bF_buf9), .Y(_4511_) );
MUX2X1 MUX2X1_207 ( .A(_1601__bF_buf3), .B(_4511_), .S(_4496__bF_buf0), .Y(_1133_) );
NAND2X1 NAND2X1_208 ( .A(REGs_REGS_6__15_), .B(_1573__bF_buf62), .Y(_4512_) );
MUX2X1 MUX2X1_208 ( .A(_1603__bF_buf2), .B(_4512_), .S(_4496__bF_buf0), .Y(_1134_) );
NAND2X1 NAND2X1_209 ( .A(REGs_REGS_6__16_), .B(_1573__bF_buf62), .Y(_4513_) );
MUX2X1 MUX2X1_209 ( .A(_1605__bF_buf2), .B(_4513_), .S(_4496__bF_buf0), .Y(_1135_) );
NAND2X1 NAND2X1_210 ( .A(REGs_REGS_6__17_), .B(_1573__bF_buf42), .Y(_4514_) );
MUX2X1 MUX2X1_210 ( .A(_1607__bF_buf0), .B(_4514_), .S(_4496__bF_buf1), .Y(_1136_) );
NAND2X1 NAND2X1_211 ( .A(REGs_REGS_6__18_), .B(_1573__bF_buf49), .Y(_4515_) );
MUX2X1 MUX2X1_211 ( .A(_1609__bF_buf1), .B(_4515_), .S(_4496__bF_buf1), .Y(_1137_) );
NAND2X1 NAND2X1_212 ( .A(REGs_REGS_6__19_), .B(_1573__bF_buf42), .Y(_4516_) );
MUX2X1 MUX2X1_212 ( .A(_1611__bF_buf3), .B(_4516_), .S(_4496__bF_buf1), .Y(_1138_) );
NAND2X1 NAND2X1_213 ( .A(REGs_REGS_6__20_), .B(_1573__bF_buf15), .Y(_4517_) );
MUX2X1 MUX2X1_213 ( .A(_1613__bF_buf2), .B(_4517_), .S(_4496__bF_buf4), .Y(_1139_) );
NAND2X1 NAND2X1_214 ( .A(REGs_REGS_6__21_), .B(_1573__bF_buf2), .Y(_4518_) );
MUX2X1 MUX2X1_214 ( .A(_1615__bF_buf1), .B(_4518_), .S(_4496__bF_buf3), .Y(_1140_) );
NAND2X1 NAND2X1_215 ( .A(REGs_REGS_6__22_), .B(_1573__bF_buf67), .Y(_4519_) );
MUX2X1 MUX2X1_215 ( .A(_1617__bF_buf0), .B(_4519_), .S(_4496__bF_buf4), .Y(_1141_) );
NAND2X1 NAND2X1_216 ( .A(REGs_REGS_6__23_), .B(_1573__bF_buf9), .Y(_4520_) );
MUX2X1 MUX2X1_216 ( .A(_1619__bF_buf2), .B(_4520_), .S(_4496__bF_buf0), .Y(_1142_) );
NAND2X1 NAND2X1_217 ( .A(REGs_REGS_6__24_), .B(_1573__bF_buf33), .Y(_4521_) );
MUX2X1 MUX2X1_217 ( .A(_1621__bF_buf2), .B(_4521_), .S(_4496__bF_buf1), .Y(_1143_) );
NAND2X1 NAND2X1_218 ( .A(REGs_REGS_6__25_), .B(_1573__bF_buf19), .Y(_4522_) );
MUX2X1 MUX2X1_218 ( .A(_1623__bF_buf2), .B(_4522_), .S(_4496__bF_buf2), .Y(_1144_) );
NAND2X1 NAND2X1_219 ( .A(REGs_REGS_6__26_), .B(_1573__bF_buf15), .Y(_4523_) );
MUX2X1 MUX2X1_219 ( .A(_1625__bF_buf1), .B(_4523_), .S(_4496__bF_buf4), .Y(_1145_) );
NAND2X1 NAND2X1_220 ( .A(REGs_REGS_6__27_), .B(_1573__bF_buf19), .Y(_4524_) );
MUX2X1 MUX2X1_220 ( .A(_1627__bF_buf0), .B(_4524_), .S(_4496__bF_buf2), .Y(_1146_) );
NAND2X1 NAND2X1_221 ( .A(REGs_REGS_6__28_), .B(_1573__bF_buf73), .Y(_4525_) );
MUX2X1 MUX2X1_221 ( .A(_1629__bF_buf3), .B(_4525_), .S(_4496__bF_buf3), .Y(_1147_) );
NAND2X1 NAND2X1_222 ( .A(REGs_REGS_6__29_), .B(_1573__bF_buf42), .Y(_4526_) );
MUX2X1 MUX2X1_222 ( .A(_1631__bF_buf2), .B(_4526_), .S(_4496__bF_buf1), .Y(_1148_) );
NAND2X1 NAND2X1_223 ( .A(REGs_REGS_6__30_), .B(_1573__bF_buf19), .Y(_4527_) );
MUX2X1 MUX2X1_223 ( .A(_1633__bF_buf1), .B(_4527_), .S(_4496__bF_buf2), .Y(_1149_) );
NAND2X1 NAND2X1_224 ( .A(REGs_REGS_6__31_), .B(_1573__bF_buf49), .Y(_4528_) );
MUX2X1 MUX2X1_224 ( .A(_1635__bF_buf1), .B(_4528_), .S(_4496__bF_buf1), .Y(_1150_) );
NAND3X1 NAND3X1_9 ( .A(_1570_), .B(REG_RFD_exec_pipe_2_), .C(_4289_), .Y(_4529_) );
NOR2X1 NOR2X1_6 ( .A(_4529_), .B(_4495_), .Y(_4530_) );
NAND2X1 NAND2X1_225 ( .A(REGs_REGS_4__0_), .B(_1573__bF_buf34), .Y(_4531_) );
MUX2X1 MUX2X1_225 ( .A(_1567__bF_buf1), .B(_4531_), .S(_4530__bF_buf0), .Y(_1151_) );
NAND2X1 NAND2X1_226 ( .A(REGs_REGS_4__1_), .B(_1573__bF_buf73), .Y(_4532_) );
MUX2X1 MUX2X1_226 ( .A(_1575__bF_buf3), .B(_4532_), .S(_4530__bF_buf3), .Y(_1152_) );
NAND2X1 NAND2X1_227 ( .A(REGs_REGS_4__2_), .B(_1573__bF_buf34), .Y(_4533_) );
MUX2X1 MUX2X1_227 ( .A(_1577__bF_buf0), .B(_4533_), .S(_4530__bF_buf0), .Y(_1153_) );
NAND2X1 NAND2X1_228 ( .A(REGs_REGS_4__3_), .B(_1573__bF_buf36), .Y(_4534_) );
MUX2X1 MUX2X1_228 ( .A(_1579__bF_buf2), .B(_4534_), .S(_4530__bF_buf0), .Y(_1154_) );
NAND2X1 NAND2X1_229 ( .A(REGs_REGS_4__4_), .B(_1573__bF_buf66), .Y(_4535_) );
MUX2X1 MUX2X1_229 ( .A(_1581__bF_buf1), .B(_4535_), .S(_4530__bF_buf1), .Y(_1155_) );
NAND2X1 NAND2X1_230 ( .A(REGs_REGS_4__5_), .B(_1573__bF_buf73), .Y(_4536_) );
MUX2X1 MUX2X1_230 ( .A(_1583__bF_buf3), .B(_4536_), .S(_4530__bF_buf3), .Y(_1156_) );
NAND2X1 NAND2X1_231 ( .A(REGs_REGS_4__6_), .B(_1573__bF_buf67), .Y(_4537_) );
MUX2X1 MUX2X1_231 ( .A(_1585__bF_buf3), .B(_4537_), .S(_4530__bF_buf1), .Y(_1157_) );
NAND2X1 NAND2X1_232 ( .A(REGs_REGS_4__7_), .B(_1573__bF_buf67), .Y(_4538_) );
MUX2X1 MUX2X1_232 ( .A(_1587__bF_buf3), .B(_4538_), .S(_4530__bF_buf1), .Y(_1158_) );
NAND2X1 NAND2X1_233 ( .A(REGs_REGS_4__8_), .B(_1573__bF_buf25), .Y(_4539_) );
MUX2X1 MUX2X1_233 ( .A(_1589__bF_buf3), .B(_4539_), .S(_4530__bF_buf2), .Y(_1159_) );
NAND2X1 NAND2X1_234 ( .A(REGs_REGS_4__9_), .B(_1573__bF_buf29), .Y(_4540_) );
MUX2X1 MUX2X1_234 ( .A(_1591__bF_buf2), .B(_4540_), .S(_4530__bF_buf2), .Y(_1160_) );
NAND2X1 NAND2X1_235 ( .A(REGs_REGS_4__10_), .B(_1573__bF_buf62), .Y(_4541_) );
MUX2X1 MUX2X1_235 ( .A(_1593__bF_buf0), .B(_4541_), .S(_4530__bF_buf3), .Y(_1161_) );
NAND2X1 NAND2X1_236 ( .A(REGs_REGS_4__11_), .B(_1573__bF_buf73), .Y(_4542_) );
MUX2X1 MUX2X1_236 ( .A(_1595__bF_buf2), .B(_4542_), .S(_4530__bF_buf3), .Y(_1162_) );
NAND2X1 NAND2X1_237 ( .A(REGs_REGS_4__12_), .B(_1573__bF_buf66), .Y(_4543_) );
MUX2X1 MUX2X1_237 ( .A(_1597__bF_buf0), .B(_4543_), .S(_4530__bF_buf1), .Y(_1163_) );
NAND2X1 NAND2X1_238 ( .A(REGs_REGS_4__13_), .B(_1573__bF_buf10), .Y(_4544_) );
MUX2X1 MUX2X1_238 ( .A(_1599__bF_buf2), .B(_4544_), .S(_4530__bF_buf4), .Y(_1164_) );
NAND2X1 NAND2X1_239 ( .A(REGs_REGS_4__14_), .B(_1573__bF_buf9), .Y(_4545_) );
MUX2X1 MUX2X1_239 ( .A(_1601__bF_buf3), .B(_4545_), .S(_4530__bF_buf3), .Y(_1165_) );
NAND2X1 NAND2X1_240 ( .A(REGs_REGS_4__15_), .B(_1573__bF_buf64), .Y(_4546_) );
MUX2X1 MUX2X1_240 ( .A(_1603__bF_buf2), .B(_4546_), .S(_4530__bF_buf2), .Y(_1166_) );
NAND2X1 NAND2X1_241 ( .A(REGs_REGS_4__16_), .B(_1573__bF_buf62), .Y(_4547_) );
MUX2X1 MUX2X1_241 ( .A(_1605__bF_buf2), .B(_4547_), .S(_4530__bF_buf3), .Y(_1167_) );
NAND2X1 NAND2X1_242 ( .A(REGs_REGS_4__17_), .B(_1573__bF_buf33), .Y(_4548_) );
MUX2X1 MUX2X1_242 ( .A(_1607__bF_buf0), .B(_4548_), .S(_4530__bF_buf4), .Y(_1168_) );
NAND2X1 NAND2X1_243 ( .A(REGs_REGS_4__18_), .B(_1573__bF_buf29), .Y(_4549_) );
MUX2X1 MUX2X1_243 ( .A(_1609__bF_buf0), .B(_4549_), .S(_4530__bF_buf2), .Y(_1169_) );
NAND2X1 NAND2X1_244 ( .A(REGs_REGS_4__19_), .B(_1573__bF_buf33), .Y(_4550_) );
MUX2X1 MUX2X1_244 ( .A(_1611__bF_buf3), .B(_4550_), .S(_4530__bF_buf4), .Y(_1170_) );
NAND2X1 NAND2X1_245 ( .A(REGs_REGS_4__20_), .B(_1573__bF_buf36), .Y(_4551_) );
MUX2X1 MUX2X1_245 ( .A(_1613__bF_buf1), .B(_4551_), .S(_4530__bF_buf0), .Y(_1171_) );
NAND2X1 NAND2X1_246 ( .A(REGs_REGS_4__21_), .B(_1573__bF_buf25), .Y(_4552_) );
MUX2X1 MUX2X1_246 ( .A(_1615__bF_buf0), .B(_4552_), .S(_4530__bF_buf2), .Y(_1172_) );
NAND2X1 NAND2X1_247 ( .A(REGs_REGS_4__22_), .B(_1573__bF_buf67), .Y(_4553_) );
MUX2X1 MUX2X1_247 ( .A(_1617__bF_buf0), .B(_4553_), .S(_4530__bF_buf1), .Y(_1173_) );
NAND2X1 NAND2X1_248 ( .A(REGs_REGS_4__23_), .B(_1573__bF_buf64), .Y(_4554_) );
MUX2X1 MUX2X1_248 ( .A(_1619__bF_buf0), .B(_4554_), .S(_4530__bF_buf2), .Y(_1174_) );
NAND2X1 NAND2X1_249 ( .A(REGs_REGS_4__24_), .B(_1573__bF_buf33), .Y(_4555_) );
MUX2X1 MUX2X1_249 ( .A(_1621__bF_buf2), .B(_4555_), .S(_4530__bF_buf4), .Y(_1175_) );
NAND2X1 NAND2X1_250 ( .A(REGs_REGS_4__25_), .B(_1573__bF_buf51), .Y(_4556_) );
MUX2X1 MUX2X1_250 ( .A(_1623__bF_buf2), .B(_4556_), .S(_4530__bF_buf4), .Y(_1176_) );
NAND2X1 NAND2X1_251 ( .A(REGs_REGS_4__26_), .B(_1573__bF_buf15), .Y(_4557_) );
MUX2X1 MUX2X1_251 ( .A(_1625__bF_buf0), .B(_4557_), .S(_4530__bF_buf1), .Y(_1177_) );
NAND2X1 NAND2X1_252 ( .A(REGs_REGS_4__27_), .B(_1573__bF_buf51), .Y(_4558_) );
MUX2X1 MUX2X1_252 ( .A(_1627__bF_buf0), .B(_4558_), .S(_4530__bF_buf4), .Y(_1178_) );
NAND2X1 NAND2X1_253 ( .A(REGs_REGS_4__28_), .B(_1573__bF_buf29), .Y(_4559_) );
MUX2X1 MUX2X1_253 ( .A(_1629__bF_buf3), .B(_4559_), .S(_4530__bF_buf3), .Y(_1179_) );
NAND2X1 NAND2X1_254 ( .A(REGs_REGS_4__29_), .B(_1573__bF_buf36), .Y(_4560_) );
MUX2X1 MUX2X1_254 ( .A(_1631__bF_buf2), .B(_4560_), .S(_4530__bF_buf0), .Y(_1180_) );
NAND2X1 NAND2X1_255 ( .A(REGs_REGS_4__30_), .B(_1573__bF_buf34), .Y(_4561_) );
MUX2X1 MUX2X1_255 ( .A(_1633__bF_buf3), .B(_4561_), .S(_4530__bF_buf0), .Y(_1181_) );
NAND2X1 NAND2X1_256 ( .A(REGs_REGS_4__31_), .B(_1573__bF_buf33), .Y(_4562_) );
MUX2X1 MUX2X1_256 ( .A(_1635__bF_buf1), .B(_4562_), .S(_4530__bF_buf4), .Y(_1182_) );
NOR2X1 NOR2X1_7 ( .A(_4394_), .B(_4495_), .Y(_4563_) );
NAND2X1 NAND2X1_257 ( .A(REGs_REGS_3__0_), .B(_1573__bF_buf10), .Y(_4564_) );
MUX2X1 MUX2X1_257 ( .A(_1567__bF_buf1), .B(_4564_), .S(_4563__bF_buf1), .Y(_1183_) );
NAND2X1 NAND2X1_258 ( .A(REGs_REGS_3__1_), .B(_1573__bF_buf75), .Y(_4565_) );
MUX2X1 MUX2X1_258 ( .A(_1575__bF_buf3), .B(_4565_), .S(_4563__bF_buf1), .Y(_1184_) );
NAND2X1 NAND2X1_259 ( .A(REGs_REGS_3__2_), .B(_1573__bF_buf4), .Y(_4566_) );
MUX2X1 MUX2X1_259 ( .A(_1577__bF_buf1), .B(_4566_), .S(_4563__bF_buf3), .Y(_1185_) );
NAND2X1 NAND2X1_260 ( .A(REGs_REGS_3__3_), .B(_1573__bF_buf4), .Y(_4567_) );
MUX2X1 MUX2X1_260 ( .A(_1579__bF_buf2), .B(_4567_), .S(_4563__bF_buf3), .Y(_1186_) );
NAND2X1 NAND2X1_261 ( .A(REGs_REGS_3__4_), .B(_1573__bF_buf0), .Y(_4568_) );
MUX2X1 MUX2X1_261 ( .A(_1581__bF_buf3), .B(_4568_), .S(_4563__bF_buf2), .Y(_1187_) );
NAND2X1 NAND2X1_262 ( .A(REGs_REGS_3__5_), .B(_1573__bF_buf75), .Y(_4569_) );
MUX2X1 MUX2X1_262 ( .A(_1583__bF_buf3), .B(_4569_), .S(_4563__bF_buf0), .Y(_1188_) );
NAND2X1 NAND2X1_263 ( .A(REGs_REGS_3__6_), .B(_1573__bF_buf0), .Y(_4570_) );
MUX2X1 MUX2X1_263 ( .A(_1585__bF_buf3), .B(_4570_), .S(_4563__bF_buf2), .Y(_1189_) );
NAND2X1 NAND2X1_264 ( .A(REGs_REGS_3__7_), .B(_1573__bF_buf0), .Y(_4571_) );
MUX2X1 MUX2X1_264 ( .A(_1587__bF_buf3), .B(_4571_), .S(_4563__bF_buf2), .Y(_1190_) );
NAND2X1 NAND2X1_265 ( .A(REGs_REGS_3__8_), .B(_1573__bF_buf49), .Y(_4572_) );
MUX2X1 MUX2X1_265 ( .A(_1589__bF_buf1), .B(_4572_), .S(_4563__bF_buf4), .Y(_1191_) );
NAND2X1 NAND2X1_266 ( .A(REGs_REGS_3__9_), .B(_1573__bF_buf65), .Y(_4573_) );
MUX2X1 MUX2X1_266 ( .A(_1591__bF_buf2), .B(_4573_), .S(_4563__bF_buf4), .Y(_1192_) );
NAND2X1 NAND2X1_267 ( .A(REGs_REGS_3__10_), .B(_1573__bF_buf65), .Y(_4574_) );
MUX2X1 MUX2X1_267 ( .A(_1593__bF_buf0), .B(_4574_), .S(_4563__bF_buf0), .Y(_1193_) );
NAND2X1 NAND2X1_268 ( .A(REGs_REGS_3__11_), .B(_1573__bF_buf41), .Y(_4575_) );
MUX2X1 MUX2X1_268 ( .A(_1595__bF_buf2), .B(_4575_), .S(_4563__bF_buf4), .Y(_1194_) );
NAND2X1 NAND2X1_269 ( .A(REGs_REGS_3__12_), .B(_1573__bF_buf19), .Y(_4576_) );
MUX2X1 MUX2X1_269 ( .A(_1597__bF_buf3), .B(_4576_), .S(_4563__bF_buf2), .Y(_1195_) );
NAND2X1 NAND2X1_270 ( .A(REGs_REGS_3__13_), .B(_1573__bF_buf10), .Y(_4577_) );
MUX2X1 MUX2X1_270 ( .A(_1599__bF_buf2), .B(_4577_), .S(_4563__bF_buf1), .Y(_1196_) );
NAND2X1 NAND2X1_271 ( .A(REGs_REGS_3__14_), .B(_1573__bF_buf41), .Y(_4578_) );
MUX2X1 MUX2X1_271 ( .A(_1601__bF_buf0), .B(_4578_), .S(_4563__bF_buf4), .Y(_1197_) );
NAND2X1 NAND2X1_272 ( .A(REGs_REGS_3__15_), .B(_1573__bF_buf41), .Y(_4579_) );
MUX2X1 MUX2X1_272 ( .A(_1603__bF_buf2), .B(_4579_), .S(_4563__bF_buf4), .Y(_1198_) );
NAND2X1 NAND2X1_273 ( .A(REGs_REGS_3__16_), .B(_1573__bF_buf65), .Y(_4580_) );
MUX2X1 MUX2X1_273 ( .A(_1605__bF_buf2), .B(_4580_), .S(_4563__bF_buf0), .Y(_1199_) );
NAND2X1 NAND2X1_274 ( .A(REGs_REGS_3__17_), .B(_1573__bF_buf10), .Y(_4581_) );
MUX2X1 MUX2X1_274 ( .A(_1607__bF_buf0), .B(_4581_), .S(_4563__bF_buf1), .Y(_1200_) );
NAND2X1 NAND2X1_275 ( .A(REGs_REGS_3__18_), .B(_1573__bF_buf65), .Y(_4582_) );
MUX2X1 MUX2X1_275 ( .A(_1609__bF_buf1), .B(_4582_), .S(_4563__bF_buf0), .Y(_1201_) );
NAND2X1 NAND2X1_276 ( .A(REGs_REGS_3__19_), .B(_1573__bF_buf75), .Y(_4583_) );
MUX2X1 MUX2X1_276 ( .A(_1611__bF_buf3), .B(_4583_), .S(_4563__bF_buf0), .Y(_1202_) );
NAND2X1 NAND2X1_277 ( .A(REGs_REGS_3__20_), .B(_1573__bF_buf51), .Y(_4584_) );
MUX2X1 MUX2X1_277 ( .A(_1613__bF_buf1), .B(_4584_), .S(_4563__bF_buf3), .Y(_1203_) );
NAND2X1 NAND2X1_278 ( .A(REGs_REGS_3__21_), .B(_1573__bF_buf49), .Y(_4585_) );
MUX2X1 MUX2X1_278 ( .A(_1615__bF_buf1), .B(_4585_), .S(_4563__bF_buf4), .Y(_1204_) );
NAND2X1 NAND2X1_279 ( .A(REGs_REGS_3__22_), .B(_1573__bF_buf0), .Y(_4586_) );
MUX2X1 MUX2X1_279 ( .A(_1617__bF_buf2), .B(_4586_), .S(_4563__bF_buf2), .Y(_1205_) );
NAND2X1 NAND2X1_280 ( .A(REGs_REGS_3__23_), .B(_1573__bF_buf65), .Y(_4587_) );
MUX2X1 MUX2X1_280 ( .A(_1619__bF_buf0), .B(_4587_), .S(_4563__bF_buf0), .Y(_1206_) );
NAND2X1 NAND2X1_281 ( .A(REGs_REGS_3__24_), .B(_1573__bF_buf10), .Y(_4588_) );
MUX2X1 MUX2X1_281 ( .A(_1621__bF_buf2), .B(_4588_), .S(_4563__bF_buf1), .Y(_1207_) );
NAND2X1 NAND2X1_282 ( .A(REGs_REGS_3__25_), .B(_1573__bF_buf51), .Y(_4589_) );
MUX2X1 MUX2X1_282 ( .A(_1623__bF_buf2), .B(_4589_), .S(_4563__bF_buf3), .Y(_1208_) );
NAND2X1 NAND2X1_283 ( .A(REGs_REGS_3__26_), .B(_1573__bF_buf0), .Y(_4590_) );
MUX2X1 MUX2X1_283 ( .A(_1625__bF_buf1), .B(_4590_), .S(_4563__bF_buf2), .Y(_1209_) );
NAND2X1 NAND2X1_284 ( .A(REGs_REGS_3__27_), .B(_1573__bF_buf51), .Y(_4591_) );
MUX2X1 MUX2X1_284 ( .A(_1627__bF_buf0), .B(_4591_), .S(_4563__bF_buf3), .Y(_1210_) );
NAND2X1 NAND2X1_285 ( .A(REGs_REGS_3__28_), .B(_1573__bF_buf49), .Y(_4592_) );
MUX2X1 MUX2X1_285 ( .A(_1629__bF_buf3), .B(_4592_), .S(_4563__bF_buf4), .Y(_1211_) );
NAND2X1 NAND2X1_286 ( .A(REGs_REGS_3__29_), .B(_1573__bF_buf51), .Y(_4593_) );
MUX2X1 MUX2X1_286 ( .A(_1631__bF_buf2), .B(_4593_), .S(_4563__bF_buf3), .Y(_1212_) );
NAND2X1 NAND2X1_287 ( .A(REGs_REGS_3__30_), .B(_1573__bF_buf4), .Y(_4594_) );
MUX2X1 MUX2X1_287 ( .A(_1633__bF_buf1), .B(_4594_), .S(_4563__bF_buf3), .Y(_1213_) );
NAND2X1 NAND2X1_288 ( .A(REGs_REGS_3__31_), .B(_1573__bF_buf75), .Y(_4595_) );
MUX2X1 MUX2X1_288 ( .A(_1635__bF_buf1), .B(_4595_), .S(_4563__bF_buf1), .Y(_1214_) );
NOR2X1 NOR2X1_8 ( .A(_4529_), .B(_4358_), .Y(_4596_) );
NAND2X1 NAND2X1_289 ( .A(REGs_FIRQ_REGS_4__0_), .B(_1573__bF_buf54), .Y(_4597_) );
MUX2X1 MUX2X1_289 ( .A(_1567__bF_buf3), .B(_4597_), .S(_4596__bF_buf1), .Y(_1215_) );
NAND2X1 NAND2X1_290 ( .A(REGs_FIRQ_REGS_4__1_), .B(_1573__bF_buf53), .Y(_4598_) );
MUX2X1 MUX2X1_290 ( .A(_1575__bF_buf0), .B(_4598_), .S(_4596__bF_buf4), .Y(_1216_) );
NAND2X1 NAND2X1_291 ( .A(REGs_FIRQ_REGS_4__2_), .B(_1573__bF_buf58), .Y(_4599_) );
MUX2X1 MUX2X1_291 ( .A(_1577__bF_buf0), .B(_4599_), .S(_4596__bF_buf1), .Y(_1217_) );
NAND2X1 NAND2X1_292 ( .A(REGs_FIRQ_REGS_4__3_), .B(_1573__bF_buf23), .Y(_4600_) );
MUX2X1 MUX2X1_292 ( .A(_1579__bF_buf0), .B(_4600_), .S(_4596__bF_buf3), .Y(_1218_) );
NAND2X1 NAND2X1_293 ( .A(REGs_FIRQ_REGS_4__4_), .B(_1573__bF_buf66), .Y(_4601_) );
MUX2X1 MUX2X1_293 ( .A(_1581__bF_buf1), .B(_4601_), .S(_4596__bF_buf3), .Y(_1219_) );
NAND2X1 NAND2X1_294 ( .A(REGs_FIRQ_REGS_4__5_), .B(_1573__bF_buf44), .Y(_4602_) );
MUX2X1 MUX2X1_294 ( .A(_1583__bF_buf2), .B(_4602_), .S(_4596__bF_buf0), .Y(_1220_) );
NAND2X1 NAND2X1_295 ( .A(REGs_FIRQ_REGS_4__6_), .B(_1573__bF_buf38), .Y(_4603_) );
MUX2X1 MUX2X1_295 ( .A(_1585__bF_buf0), .B(_4603_), .S(_4596__bF_buf3), .Y(_1221_) );
NAND2X1 NAND2X1_296 ( .A(REGs_FIRQ_REGS_4__7_), .B(_1573__bF_buf5), .Y(_4604_) );
MUX2X1 MUX2X1_296 ( .A(_1587__bF_buf1), .B(_4604_), .S(_4596__bF_buf2), .Y(_1222_) );
NAND2X1 NAND2X1_297 ( .A(REGs_FIRQ_REGS_4__8_), .B(_1573__bF_buf74), .Y(_4605_) );
MUX2X1 MUX2X1_297 ( .A(_1589__bF_buf0), .B(_4605_), .S(_4596__bF_buf4), .Y(_1223_) );
NAND2X1 NAND2X1_298 ( .A(REGs_FIRQ_REGS_4__9_), .B(_1573__bF_buf60), .Y(_4606_) );
MUX2X1 MUX2X1_298 ( .A(_1591__bF_buf3), .B(_4606_), .S(_4596__bF_buf0), .Y(_1224_) );
NAND2X1 NAND2X1_299 ( .A(REGs_FIRQ_REGS_4__10_), .B(_1573__bF_buf70), .Y(_4607_) );
MUX2X1 MUX2X1_299 ( .A(_1593__bF_buf3), .B(_4607_), .S(_4596__bF_buf4), .Y(_1225_) );
NAND2X1 NAND2X1_300 ( .A(REGs_FIRQ_REGS_4__11_), .B(_1573__bF_buf63), .Y(_4608_) );
MUX2X1 MUX2X1_300 ( .A(_1595__bF_buf3), .B(_4608_), .S(_4596__bF_buf4), .Y(_1226_) );
NAND2X1 NAND2X1_301 ( .A(REGs_FIRQ_REGS_4__12_), .B(_1573__bF_buf3), .Y(_4609_) );
MUX2X1 MUX2X1_301 ( .A(_1597__bF_buf0), .B(_4609_), .S(_4596__bF_buf3), .Y(_1227_) );
NAND2X1 NAND2X1_302 ( .A(REGs_FIRQ_REGS_4__13_), .B(_1573__bF_buf40), .Y(_4610_) );
MUX2X1 MUX2X1_302 ( .A(_1599__bF_buf3), .B(_4610_), .S(_4596__bF_buf1), .Y(_1228_) );
NAND2X1 NAND2X1_303 ( .A(REGs_FIRQ_REGS_4__14_), .B(_1573__bF_buf60), .Y(_4611_) );
MUX2X1 MUX2X1_303 ( .A(_1601__bF_buf2), .B(_4611_), .S(_4596__bF_buf0), .Y(_1229_) );
NAND2X1 NAND2X1_304 ( .A(REGs_FIRQ_REGS_4__15_), .B(_1573__bF_buf14), .Y(_4612_) );
MUX2X1 MUX2X1_304 ( .A(_1603__bF_buf3), .B(_4612_), .S(_4596__bF_buf4), .Y(_1230_) );
NAND2X1 NAND2X1_305 ( .A(REGs_FIRQ_REGS_4__16_), .B(_1573__bF_buf52), .Y(_4613_) );
MUX2X1 MUX2X1_305 ( .A(_1605__bF_buf1), .B(_4613_), .S(_4596__bF_buf0), .Y(_1231_) );
NAND2X1 NAND2X1_306 ( .A(REGs_FIRQ_REGS_4__17_), .B(_1573__bF_buf6), .Y(_4614_) );
MUX2X1 MUX2X1_306 ( .A(_1607__bF_buf1), .B(_4614_), .S(_4596__bF_buf2), .Y(_1232_) );
NAND2X1 NAND2X1_307 ( .A(REGs_FIRQ_REGS_4__18_), .B(_1573__bF_buf52), .Y(_4615_) );
MUX2X1 MUX2X1_307 ( .A(_1609__bF_buf2), .B(_4615_), .S(_4596__bF_buf0), .Y(_1233_) );
NAND2X1 NAND2X1_308 ( .A(REGs_FIRQ_REGS_4__19_), .B(_1573__bF_buf40), .Y(_4616_) );
MUX2X1 MUX2X1_308 ( .A(_1611__bF_buf1), .B(_4616_), .S(_4596__bF_buf1), .Y(_1234_) );
NAND2X1 NAND2X1_309 ( .A(REGs_FIRQ_REGS_4__20_), .B(_1573__bF_buf5), .Y(_4617_) );
MUX2X1 MUX2X1_309 ( .A(_1613__bF_buf3), .B(_4617_), .S(_4596__bF_buf2), .Y(_1235_) );
NAND2X1 NAND2X1_310 ( .A(REGs_FIRQ_REGS_4__21_), .B(_1573__bF_buf28), .Y(_4618_) );
MUX2X1 MUX2X1_310 ( .A(_1615__bF_buf3), .B(_4618_), .S(_4596__bF_buf1), .Y(_1236_) );
NAND2X1 NAND2X1_311 ( .A(REGs_FIRQ_REGS_4__22_), .B(_1573__bF_buf3), .Y(_4619_) );
MUX2X1 MUX2X1_311 ( .A(_1617__bF_buf0), .B(_4619_), .S(_4596__bF_buf3), .Y(_1237_) );
NAND2X1 NAND2X1_312 ( .A(REGs_FIRQ_REGS_4__23_), .B(_1573__bF_buf52), .Y(_4620_) );
MUX2X1 MUX2X1_312 ( .A(_1619__bF_buf3), .B(_4620_), .S(_4596__bF_buf0), .Y(_1238_) );
NAND2X1 NAND2X1_313 ( .A(REGs_FIRQ_REGS_4__24_), .B(_1573__bF_buf71), .Y(_4621_) );
MUX2X1 MUX2X1_313 ( .A(_1621__bF_buf0), .B(_4621_), .S(_4596__bF_buf2), .Y(_1239_) );
NAND2X1 NAND2X1_314 ( .A(REGs_FIRQ_REGS_4__25_), .B(_1573__bF_buf71), .Y(_4622_) );
MUX2X1 MUX2X1_314 ( .A(_1623__bF_buf3), .B(_4622_), .S(_4596__bF_buf2), .Y(_1240_) );
NAND2X1 NAND2X1_315 ( .A(REGs_FIRQ_REGS_4__26_), .B(_1573__bF_buf55), .Y(_4623_) );
MUX2X1 MUX2X1_315 ( .A(_1625__bF_buf2), .B(_4623_), .S(_4596__bF_buf2), .Y(_1241_) );
NAND2X1 NAND2X1_316 ( .A(REGs_FIRQ_REGS_4__27_), .B(_1573__bF_buf56), .Y(_4624_) );
MUX2X1 MUX2X1_316 ( .A(_1627__bF_buf1), .B(_4624_), .S(_4596__bF_buf3), .Y(_1242_) );
NAND2X1 NAND2X1_317 ( .A(REGs_FIRQ_REGS_4__28_), .B(_1573__bF_buf20), .Y(_4625_) );
MUX2X1 MUX2X1_317 ( .A(_1629__bF_buf2), .B(_4625_), .S(_4596__bF_buf4), .Y(_1243_) );
NAND2X1 NAND2X1_318 ( .A(REGs_FIRQ_REGS_4__29_), .B(_1573__bF_buf39), .Y(_4626_) );
MUX2X1 MUX2X1_318 ( .A(_1631__bF_buf1), .B(_4626_), .S(_4596__bF_buf1), .Y(_1244_) );
NAND2X1 NAND2X1_319 ( .A(REGs_FIRQ_REGS_4__30_), .B(_1573__bF_buf56), .Y(_4627_) );
MUX2X1 MUX2X1_319 ( .A(_1633__bF_buf3), .B(_4627_), .S(_4596__bF_buf3), .Y(_1245_) );
NAND2X1 NAND2X1_320 ( .A(REGs_FIRQ_REGS_4__31_), .B(_1573__bF_buf63), .Y(_4628_) );
MUX2X1 MUX2X1_320 ( .A(_1635__bF_buf2), .B(_4628_), .S(_4596__bF_buf4), .Y(_1246_) );
NAND3X1 NAND3X1_10 ( .A(_1639_), .B(REG_RFD_exec_pipe_0_), .C(_1641_), .Y(_4629_) );
NAND2X1 NAND2X1_321 ( .A(REGs_USR_REGS_1__0_), .B(_1573__bF_buf76), .Y(_4630_) );
MUX2X1 MUX2X1_321 ( .A(_4630_), .B(_1567__bF_buf2), .S(_4629__bF_buf0), .Y(_1247_) );
NAND2X1 NAND2X1_322 ( .A(REGs_USR_REGS_1__1_), .B(_1573__bF_buf50), .Y(_4631_) );
MUX2X1 MUX2X1_322 ( .A(_4631_), .B(_1575__bF_buf0), .S(_4629__bF_buf2), .Y(_1248_) );
NAND2X1 NAND2X1_323 ( .A(REGs_USR_REGS_1__2_), .B(_1573__bF_buf61), .Y(_4632_) );
MUX2X1 MUX2X1_323 ( .A(_4632_), .B(_1577__bF_buf3), .S(_4629__bF_buf4), .Y(_1249_) );
NAND2X1 NAND2X1_324 ( .A(REGs_USR_REGS_1__3_), .B(_1573__bF_buf48), .Y(_4633_) );
MUX2X1 MUX2X1_324 ( .A(_4633_), .B(_1579__bF_buf3), .S(_4629__bF_buf3), .Y(_1250_) );
NAND2X1 NAND2X1_325 ( .A(REGs_USR_REGS_1__4_), .B(_1573__bF_buf38), .Y(_4634_) );
MUX2X1 MUX2X1_325 ( .A(_4634_), .B(_1581__bF_buf0), .S(_4629__bF_buf3), .Y(_1251_) );
NAND2X1 NAND2X1_326 ( .A(REGs_USR_REGS_1__5_), .B(_1573__bF_buf50), .Y(_4635_) );
MUX2X1 MUX2X1_326 ( .A(_4635_), .B(_1583__bF_buf2), .S(_4629__bF_buf1), .Y(_1252_) );
NAND2X1 NAND2X1_327 ( .A(REGs_USR_REGS_1__6_), .B(_1573__bF_buf11), .Y(_4636_) );
MUX2X1 MUX2X1_327 ( .A(_4636_), .B(_1585__bF_buf2), .S(_4629__bF_buf3), .Y(_1253_) );
NAND2X1 NAND2X1_328 ( .A(REGs_USR_REGS_1__7_), .B(_1573__bF_buf12), .Y(_4637_) );
MUX2X1 MUX2X1_328 ( .A(_4637_), .B(_1587__bF_buf0), .S(_4629__bF_buf0), .Y(_1254_) );
NAND2X1 NAND2X1_329 ( .A(REGs_USR_REGS_1__8_), .B(_1573__bF_buf40), .Y(_4638_) );
MUX2X1 MUX2X1_329 ( .A(_4638_), .B(_1589__bF_buf2), .S(_4629__bF_buf4), .Y(_1255_) );
NAND2X1 NAND2X1_330 ( .A(REGs_USR_REGS_1__9_), .B(_1573__bF_buf13), .Y(_4639_) );
MUX2X1 MUX2X1_330 ( .A(_4639_), .B(_1591__bF_buf0), .S(_4629__bF_buf1), .Y(_1256_) );
NAND2X1 NAND2X1_331 ( .A(REGs_USR_REGS_1__10_), .B(_1573__bF_buf74), .Y(_4640_) );
MUX2X1 MUX2X1_331 ( .A(_4640_), .B(_1593__bF_buf1), .S(_4629__bF_buf2), .Y(_1257_) );
NAND2X1 NAND2X1_332 ( .A(REGs_USR_REGS_1__11_), .B(_1573__bF_buf8), .Y(_4641_) );
MUX2X1 MUX2X1_332 ( .A(_4641_), .B(_1595__bF_buf0), .S(_4629__bF_buf2), .Y(_1258_) );
NAND2X1 NAND2X1_333 ( .A(REGs_USR_REGS_1__12_), .B(_1573__bF_buf37), .Y(_4642_) );
MUX2X1 MUX2X1_333 ( .A(_4642_), .B(_1597__bF_buf2), .S(_4629__bF_buf3), .Y(_1259_) );
NAND2X1 NAND2X1_334 ( .A(REGs_USR_REGS_1__13_), .B(_1573__bF_buf32), .Y(_4643_) );
MUX2X1 MUX2X1_334 ( .A(_4643_), .B(_1599__bF_buf0), .S(_4629__bF_buf4), .Y(_1260_) );
NAND2X1 NAND2X1_335 ( .A(REGs_USR_REGS_1__14_), .B(_1573__bF_buf20), .Y(_4644_) );
MUX2X1 MUX2X1_335 ( .A(_4644_), .B(_1601__bF_buf1), .S(_4629__bF_buf1), .Y(_1261_) );
NAND2X1 NAND2X1_336 ( .A(REGs_USR_REGS_1__15_), .B(_1573__bF_buf50), .Y(_4645_) );
MUX2X1 MUX2X1_336 ( .A(_4645_), .B(_1603__bF_buf0), .S(_4629__bF_buf2), .Y(_1262_) );
NAND2X1 NAND2X1_337 ( .A(REGs_USR_REGS_1__16_), .B(_1573__bF_buf77), .Y(_4646_) );
MUX2X1 MUX2X1_337 ( .A(_4646_), .B(_1605__bF_buf3), .S(_4629__bF_buf1), .Y(_1263_) );
NAND2X1 NAND2X1_338 ( .A(REGs_USR_REGS_1__17_), .B(_1573__bF_buf12), .Y(_4647_) );
MUX2X1 MUX2X1_338 ( .A(_4647_), .B(_1607__bF_buf2), .S(_4629__bF_buf0), .Y(_1264_) );
NAND2X1 NAND2X1_339 ( .A(REGs_USR_REGS_1__18_), .B(_1573__bF_buf20), .Y(_4648_) );
MUX2X1 MUX2X1_339 ( .A(_4648_), .B(_1609__bF_buf3), .S(_4629__bF_buf1), .Y(_1265_) );
NAND2X1 NAND2X1_340 ( .A(REGs_USR_REGS_1__19_), .B(_1573__bF_buf16), .Y(_4649_) );
MUX2X1 MUX2X1_340 ( .A(_4649_), .B(_1611__bF_buf1), .S(_4629__bF_buf4), .Y(_1266_) );
NAND2X1 NAND2X1_341 ( .A(REGs_USR_REGS_1__20_), .B(_1573__bF_buf22), .Y(_4650_) );
MUX2X1 MUX2X1_341 ( .A(_4650_), .B(_1613__bF_buf2), .S(_4629__bF_buf3), .Y(_1267_) );
NAND2X1 NAND2X1_342 ( .A(REGs_USR_REGS_1__21_), .B(_1573__bF_buf28), .Y(_4651_) );
MUX2X1 MUX2X1_342 ( .A(_4651_), .B(_1615__bF_buf2), .S(_4629__bF_buf2), .Y(_1268_) );
NAND2X1 NAND2X1_343 ( .A(REGs_USR_REGS_1__22_), .B(_1573__bF_buf11), .Y(_4652_) );
MUX2X1 MUX2X1_343 ( .A(_4652_), .B(_1617__bF_buf1), .S(_4629__bF_buf3), .Y(_1269_) );
NAND2X1 NAND2X1_344 ( .A(REGs_USR_REGS_1__23_), .B(_1573__bF_buf77), .Y(_4653_) );
MUX2X1 MUX2X1_344 ( .A(_4653_), .B(_1619__bF_buf1), .S(_4629__bF_buf1), .Y(_1270_) );
NAND2X1 NAND2X1_345 ( .A(REGs_USR_REGS_1__24_), .B(_1573__bF_buf71), .Y(_4654_) );
MUX2X1 MUX2X1_345 ( .A(_4654_), .B(_1621__bF_buf0), .S(_4629__bF_buf4), .Y(_1271_) );
NAND2X1 NAND2X1_346 ( .A(REGs_USR_REGS_1__25_), .B(_1573__bF_buf17), .Y(_4655_) );
MUX2X1 MUX2X1_346 ( .A(_4655_), .B(_1623__bF_buf1), .S(_4629__bF_buf0), .Y(_1272_) );
NAND2X1 NAND2X1_347 ( .A(REGs_USR_REGS_1__26_), .B(_1573__bF_buf38), .Y(_4656_) );
MUX2X1 MUX2X1_347 ( .A(_4656_), .B(_1625__bF_buf2), .S(_4629__bF_buf3), .Y(_1273_) );
NAND2X1 NAND2X1_348 ( .A(REGs_USR_REGS_1__27_), .B(_1573__bF_buf17), .Y(_4657_) );
MUX2X1 MUX2X1_348 ( .A(_4657_), .B(_1627__bF_buf3), .S(_4629__bF_buf0), .Y(_1274_) );
NAND2X1 NAND2X1_349 ( .A(REGs_USR_REGS_1__28_), .B(_1573__bF_buf28), .Y(_4658_) );
MUX2X1 MUX2X1_349 ( .A(_4658_), .B(_1629__bF_buf1), .S(_4629__bF_buf2), .Y(_1275_) );
NAND2X1 NAND2X1_350 ( .A(REGs_USR_REGS_1__29_), .B(_1573__bF_buf39), .Y(_4659_) );
MUX2X1 MUX2X1_350 ( .A(_4659_), .B(_1631__bF_buf1), .S(_4629__bF_buf4), .Y(_1276_) );
NAND2X1 NAND2X1_351 ( .A(REGs_USR_REGS_1__30_), .B(_1573__bF_buf22), .Y(_4660_) );
MUX2X1 MUX2X1_351 ( .A(_4660_), .B(_1633__bF_buf2), .S(_4629__bF_buf0), .Y(_1277_) );
NAND2X1 NAND2X1_352 ( .A(REGs_USR_REGS_1__31_), .B(_1573__bF_buf32), .Y(_4661_) );
MUX2X1 MUX2X1_352 ( .A(_4661_), .B(_1635__bF_buf3), .S(_4629__bF_buf4), .Y(_1278_) );
NOR2X1 NOR2X1_9 ( .A(_4360_), .B(_4495_), .Y(_4662_) );
NAND2X1 NAND2X1_353 ( .A(REGs_REGS_2__0_), .B(_1573__bF_buf10), .Y(_4663_) );
MUX2X1 MUX2X1_353 ( .A(_1567__bF_buf1), .B(_4663_), .S(_4662__bF_buf2), .Y(_1279_) );
NAND2X1 NAND2X1_354 ( .A(REGs_REGS_2__1_), .B(_1573__bF_buf75), .Y(_4664_) );
MUX2X1 MUX2X1_354 ( .A(_1575__bF_buf3), .B(_4664_), .S(_4662__bF_buf2), .Y(_1280_) );
NAND2X1 NAND2X1_355 ( .A(REGs_REGS_2__2_), .B(_1573__bF_buf4), .Y(_4665_) );
MUX2X1 MUX2X1_355 ( .A(_1577__bF_buf1), .B(_4665_), .S(_4662__bF_buf4), .Y(_1281_) );
NAND2X1 NAND2X1_356 ( .A(REGs_REGS_2__3_), .B(_1573__bF_buf4), .Y(_4666_) );
MUX2X1 MUX2X1_356 ( .A(_1579__bF_buf2), .B(_4666_), .S(_4662__bF_buf4), .Y(_1282_) );
NAND2X1 NAND2X1_357 ( .A(REGs_REGS_2__4_), .B(_1573__bF_buf0), .Y(_4667_) );
MUX2X1 MUX2X1_357 ( .A(_1581__bF_buf3), .B(_4667_), .S(_4662__bF_buf1), .Y(_1283_) );
NAND2X1 NAND2X1_358 ( .A(REGs_REGS_2__5_), .B(_1573__bF_buf75), .Y(_4668_) );
MUX2X1 MUX2X1_358 ( .A(_1583__bF_buf3), .B(_4668_), .S(_4662__bF_buf0), .Y(_1284_) );
NAND2X1 NAND2X1_359 ( .A(REGs_REGS_2__6_), .B(_1573__bF_buf0), .Y(_4669_) );
MUX2X1 MUX2X1_359 ( .A(_1585__bF_buf3), .B(_4669_), .S(_4662__bF_buf1), .Y(_1285_) );
NAND2X1 NAND2X1_360 ( .A(REGs_REGS_2__7_), .B(_1573__bF_buf0), .Y(_4670_) );
MUX2X1 MUX2X1_360 ( .A(_1587__bF_buf3), .B(_4670_), .S(_4662__bF_buf1), .Y(_1286_) );
NAND2X1 NAND2X1_361 ( .A(REGs_REGS_2__8_), .B(_1573__bF_buf49), .Y(_4671_) );
MUX2X1 MUX2X1_361 ( .A(_1589__bF_buf1), .B(_4671_), .S(_4662__bF_buf3), .Y(_1287_) );
NAND2X1 NAND2X1_362 ( .A(REGs_REGS_2__9_), .B(_1573__bF_buf41), .Y(_4672_) );
MUX2X1 MUX2X1_362 ( .A(_1591__bF_buf2), .B(_4672_), .S(_4662__bF_buf3), .Y(_1288_) );
NAND2X1 NAND2X1_363 ( .A(REGs_REGS_2__10_), .B(_1573__bF_buf65), .Y(_4673_) );
MUX2X1 MUX2X1_363 ( .A(_1593__bF_buf0), .B(_4673_), .S(_4662__bF_buf0), .Y(_1289_) );
NAND2X1 NAND2X1_364 ( .A(REGs_REGS_2__11_), .B(_1573__bF_buf41), .Y(_4674_) );
MUX2X1 MUX2X1_364 ( .A(_1595__bF_buf2), .B(_4674_), .S(_4662__bF_buf3), .Y(_1290_) );
NAND2X1 NAND2X1_365 ( .A(REGs_REGS_2__12_), .B(_1573__bF_buf19), .Y(_4675_) );
MUX2X1 MUX2X1_365 ( .A(_1597__bF_buf3), .B(_4675_), .S(_4662__bF_buf1), .Y(_1291_) );
NAND2X1 NAND2X1_366 ( .A(REGs_REGS_2__13_), .B(_1573__bF_buf10), .Y(_4676_) );
MUX2X1 MUX2X1_366 ( .A(_1599__bF_buf2), .B(_4676_), .S(_4662__bF_buf2), .Y(_1292_) );
NAND2X1 NAND2X1_367 ( .A(REGs_REGS_2__14_), .B(_1573__bF_buf41), .Y(_4677_) );
MUX2X1 MUX2X1_367 ( .A(_1601__bF_buf0), .B(_4677_), .S(_4662__bF_buf3), .Y(_1293_) );
NAND2X1 NAND2X1_368 ( .A(REGs_REGS_2__15_), .B(_1573__bF_buf41), .Y(_4678_) );
MUX2X1 MUX2X1_368 ( .A(_1603__bF_buf2), .B(_4678_), .S(_4662__bF_buf3), .Y(_1294_) );
NAND2X1 NAND2X1_369 ( .A(REGs_REGS_2__16_), .B(_1573__bF_buf65), .Y(_4679_) );
MUX2X1 MUX2X1_369 ( .A(_1605__bF_buf2), .B(_4679_), .S(_4662__bF_buf0), .Y(_1295_) );
NAND2X1 NAND2X1_370 ( .A(REGs_REGS_2__17_), .B(_1573__bF_buf10), .Y(_4680_) );
MUX2X1 MUX2X1_370 ( .A(_1607__bF_buf0), .B(_4680_), .S(_4662__bF_buf2), .Y(_1296_) );
NAND2X1 NAND2X1_371 ( .A(REGs_REGS_2__18_), .B(_1573__bF_buf65), .Y(_4681_) );
MUX2X1 MUX2X1_371 ( .A(_1609__bF_buf1), .B(_4681_), .S(_4662__bF_buf0), .Y(_1297_) );
NAND2X1 NAND2X1_372 ( .A(REGs_REGS_2__19_), .B(_1573__bF_buf75), .Y(_4682_) );
MUX2X1 MUX2X1_372 ( .A(_1611__bF_buf3), .B(_4682_), .S(_4662__bF_buf0), .Y(_1298_) );
NAND2X1 NAND2X1_373 ( .A(REGs_REGS_2__20_), .B(_1573__bF_buf51), .Y(_4683_) );
MUX2X1 MUX2X1_373 ( .A(_1613__bF_buf1), .B(_4683_), .S(_4662__bF_buf4), .Y(_1299_) );
NAND2X1 NAND2X1_374 ( .A(REGs_REGS_2__21_), .B(_1573__bF_buf41), .Y(_4684_) );
MUX2X1 MUX2X1_374 ( .A(_1615__bF_buf1), .B(_4684_), .S(_4662__bF_buf3), .Y(_1300_) );
NAND2X1 NAND2X1_375 ( .A(REGs_REGS_2__22_), .B(_1573__bF_buf19), .Y(_4685_) );
MUX2X1 MUX2X1_375 ( .A(_1617__bF_buf2), .B(_4685_), .S(_4662__bF_buf1), .Y(_1301_) );
NAND2X1 NAND2X1_376 ( .A(REGs_REGS_2__23_), .B(_1573__bF_buf65), .Y(_4686_) );
MUX2X1 MUX2X1_376 ( .A(_1619__bF_buf0), .B(_4686_), .S(_4662__bF_buf0), .Y(_1302_) );
NAND2X1 NAND2X1_377 ( .A(REGs_REGS_2__24_), .B(_1573__bF_buf10), .Y(_4687_) );
MUX2X1 MUX2X1_377 ( .A(_1621__bF_buf2), .B(_4687_), .S(_4662__bF_buf2), .Y(_1303_) );
NAND2X1 NAND2X1_378 ( .A(REGs_REGS_2__25_), .B(_1573__bF_buf4), .Y(_4688_) );
MUX2X1 MUX2X1_378 ( .A(_1623__bF_buf2), .B(_4688_), .S(_4662__bF_buf4), .Y(_1304_) );
NAND2X1 NAND2X1_379 ( .A(REGs_REGS_2__26_), .B(_1573__bF_buf19), .Y(_4689_) );
MUX2X1 MUX2X1_379 ( .A(_1625__bF_buf1), .B(_4689_), .S(_4662__bF_buf1), .Y(_1305_) );
NAND2X1 NAND2X1_380 ( .A(REGs_REGS_2__27_), .B(_1573__bF_buf4), .Y(_4690_) );
MUX2X1 MUX2X1_380 ( .A(_1627__bF_buf0), .B(_4690_), .S(_4662__bF_buf4), .Y(_1306_) );
NAND2X1 NAND2X1_381 ( .A(REGs_REGS_2__28_), .B(_1573__bF_buf49), .Y(_4691_) );
MUX2X1 MUX2X1_381 ( .A(_1629__bF_buf3), .B(_4691_), .S(_4662__bF_buf3), .Y(_1307_) );
NAND2X1 NAND2X1_382 ( .A(REGs_REGS_2__29_), .B(_1573__bF_buf51), .Y(_4692_) );
MUX2X1 MUX2X1_382 ( .A(_1631__bF_buf2), .B(_4692_), .S(_4662__bF_buf4), .Y(_1308_) );
NAND2X1 NAND2X1_383 ( .A(REGs_REGS_2__30_), .B(_1573__bF_buf4), .Y(_4693_) );
MUX2X1 MUX2X1_383 ( .A(_1633__bF_buf1), .B(_4693_), .S(_4662__bF_buf4), .Y(_1309_) );
NAND2X1 NAND2X1_384 ( .A(REGs_REGS_2__31_), .B(_1573__bF_buf75), .Y(_4694_) );
MUX2X1 MUX2X1_384 ( .A(_1635__bF_buf1), .B(_4694_), .S(_4662__bF_buf2), .Y(_1310_) );
NOR2X1 NOR2X1_10 ( .A(_4290_), .B(_4358_), .Y(_4695_) );
NAND2X1 NAND2X1_385 ( .A(REGs_FIRQ_REGS_5__0_), .B(_1573__bF_buf40), .Y(_4696_) );
MUX2X1 MUX2X1_385 ( .A(_1567__bF_buf0), .B(_4696_), .S(_4695__bF_buf3), .Y(_1311_) );
NAND2X1 NAND2X1_386 ( .A(REGs_FIRQ_REGS_5__1_), .B(_1573__bF_buf14), .Y(_4697_) );
MUX2X1 MUX2X1_386 ( .A(_1575__bF_buf1), .B(_4697_), .S(_4695__bF_buf0), .Y(_1312_) );
NAND2X1 NAND2X1_387 ( .A(REGs_FIRQ_REGS_5__2_), .B(_1573__bF_buf23), .Y(_4698_) );
MUX2X1 MUX2X1_387 ( .A(_1577__bF_buf2), .B(_4698_), .S(_4695__bF_buf2), .Y(_1313_) );
NAND2X1 NAND2X1_388 ( .A(REGs_FIRQ_REGS_5__3_), .B(_1573__bF_buf59), .Y(_4699_) );
MUX2X1 MUX2X1_388 ( .A(_1579__bF_buf1), .B(_4699_), .S(_4695__bF_buf2), .Y(_1314_) );
NAND2X1 NAND2X1_389 ( .A(REGs_FIRQ_REGS_5__4_), .B(_1573__bF_buf27), .Y(_4700_) );
MUX2X1 MUX2X1_389 ( .A(_1581__bF_buf2), .B(_4700_), .S(_4695__bF_buf1), .Y(_1315_) );
NAND2X1 NAND2X1_390 ( .A(REGs_FIRQ_REGS_5__5_), .B(_1573__bF_buf78), .Y(_4701_) );
MUX2X1 MUX2X1_390 ( .A(_1583__bF_buf1), .B(_4701_), .S(_4695__bF_buf4), .Y(_1316_) );
NAND2X1 NAND2X1_391 ( .A(REGs_FIRQ_REGS_5__6_), .B(_1573__bF_buf72), .Y(_4702_) );
MUX2X1 MUX2X1_391 ( .A(_1585__bF_buf1), .B(_4702_), .S(_4695__bF_buf1), .Y(_1317_) );
NAND2X1 NAND2X1_392 ( .A(REGs_FIRQ_REGS_5__7_), .B(_1573__bF_buf56), .Y(_4703_) );
MUX2X1 MUX2X1_392 ( .A(_1587__bF_buf2), .B(_4703_), .S(_4695__bF_buf2), .Y(_1318_) );
NAND2X1 NAND2X1_393 ( .A(REGs_FIRQ_REGS_5__8_), .B(_1573__bF_buf68), .Y(_4704_) );
MUX2X1 MUX2X1_393 ( .A(_1589__bF_buf0), .B(_4704_), .S(_4695__bF_buf0), .Y(_1319_) );
NAND2X1 NAND2X1_394 ( .A(REGs_FIRQ_REGS_5__9_), .B(_1573__bF_buf78), .Y(_4705_) );
MUX2X1 MUX2X1_394 ( .A(_1591__bF_buf1), .B(_4705_), .S(_4695__bF_buf4), .Y(_1320_) );
NAND2X1 NAND2X1_395 ( .A(REGs_FIRQ_REGS_5__10_), .B(_1573__bF_buf44), .Y(_4706_) );
MUX2X1 MUX2X1_395 ( .A(_1593__bF_buf2), .B(_4706_), .S(_4695__bF_buf4), .Y(_1321_) );
NAND2X1 NAND2X1_396 ( .A(REGs_FIRQ_REGS_5__11_), .B(_1573__bF_buf68), .Y(_4707_) );
MUX2X1 MUX2X1_396 ( .A(_1595__bF_buf0), .B(_4707_), .S(_4695__bF_buf0), .Y(_1322_) );
NAND2X1 NAND2X1_397 ( .A(REGs_FIRQ_REGS_5__12_), .B(_1573__bF_buf72), .Y(_4708_) );
MUX2X1 MUX2X1_397 ( .A(_1597__bF_buf1), .B(_4708_), .S(_4695__bF_buf1), .Y(_1323_) );
NAND2X1 NAND2X1_398 ( .A(REGs_FIRQ_REGS_5__13_), .B(_1573__bF_buf1), .Y(_4709_) );
MUX2X1 MUX2X1_398 ( .A(_1599__bF_buf3), .B(_4709_), .S(_4695__bF_buf3), .Y(_1324_) );
NAND2X1 NAND2X1_399 ( .A(REGs_FIRQ_REGS_5__14_), .B(_1573__bF_buf44), .Y(_4710_) );
MUX2X1 MUX2X1_399 ( .A(_1601__bF_buf2), .B(_4710_), .S(_4695__bF_buf0), .Y(_1325_) );
NAND2X1 NAND2X1_400 ( .A(REGs_FIRQ_REGS_5__15_), .B(_1573__bF_buf53), .Y(_4711_) );
MUX2X1 MUX2X1_400 ( .A(_1603__bF_buf3), .B(_4711_), .S(_4695__bF_buf4), .Y(_1326_) );
NAND2X1 NAND2X1_401 ( .A(REGs_FIRQ_REGS_5__16_), .B(_1573__bF_buf70), .Y(_4712_) );
MUX2X1 MUX2X1_401 ( .A(_1605__bF_buf0), .B(_4712_), .S(_4695__bF_buf4), .Y(_1327_) );
NAND2X1 NAND2X1_402 ( .A(REGs_FIRQ_REGS_5__17_), .B(_1573__bF_buf23), .Y(_4713_) );
MUX2X1 MUX2X1_402 ( .A(_1607__bF_buf3), .B(_4713_), .S(_4695__bF_buf2), .Y(_1328_) );
NAND2X1 NAND2X1_403 ( .A(REGs_FIRQ_REGS_5__18_), .B(_1573__bF_buf52), .Y(_4714_) );
MUX2X1 MUX2X1_403 ( .A(_1609__bF_buf2), .B(_4714_), .S(_4695__bF_buf0), .Y(_1329_) );
NAND2X1 NAND2X1_404 ( .A(REGs_FIRQ_REGS_5__19_), .B(_1573__bF_buf43), .Y(_4715_) );
MUX2X1 MUX2X1_404 ( .A(_1611__bF_buf2), .B(_4715_), .S(_4695__bF_buf3), .Y(_1330_) );
NAND2X1 NAND2X1_405 ( .A(REGs_FIRQ_REGS_5__20_), .B(_1573__bF_buf56), .Y(_4716_) );
MUX2X1 MUX2X1_405 ( .A(_1613__bF_buf1), .B(_4716_), .S(_4695__bF_buf2), .Y(_1331_) );
NAND2X1 NAND2X1_406 ( .A(REGs_FIRQ_REGS_5__21_), .B(_1573__bF_buf1), .Y(_4717_) );
MUX2X1 MUX2X1_406 ( .A(_1615__bF_buf3), .B(_4717_), .S(_4695__bF_buf3), .Y(_1332_) );
NAND2X1 NAND2X1_407 ( .A(REGs_FIRQ_REGS_5__22_), .B(_1573__bF_buf46), .Y(_4718_) );
MUX2X1 MUX2X1_407 ( .A(_1617__bF_buf2), .B(_4718_), .S(_4695__bF_buf1), .Y(_1333_) );
NAND2X1 NAND2X1_408 ( .A(REGs_FIRQ_REGS_5__23_), .B(_1573__bF_buf60), .Y(_4719_) );
MUX2X1 MUX2X1_408 ( .A(_1619__bF_buf3), .B(_4719_), .S(_4695__bF_buf0), .Y(_1334_) );
NAND2X1 NAND2X1_409 ( .A(REGs_FIRQ_REGS_5__24_), .B(_1573__bF_buf43), .Y(_4720_) );
MUX2X1 MUX2X1_409 ( .A(_1621__bF_buf1), .B(_4720_), .S(_4695__bF_buf3), .Y(_1335_) );
NAND2X1 NAND2X1_410 ( .A(REGs_FIRQ_REGS_5__25_), .B(_1573__bF_buf1), .Y(_4721_) );
MUX2X1 MUX2X1_410 ( .A(_1623__bF_buf0), .B(_4721_), .S(_4695__bF_buf3), .Y(_1336_) );
NAND2X1 NAND2X1_411 ( .A(REGs_FIRQ_REGS_5__26_), .B(_1573__bF_buf46), .Y(_4722_) );
MUX2X1 MUX2X1_411 ( .A(_1625__bF_buf0), .B(_4722_), .S(_4695__bF_buf1), .Y(_1337_) );
NAND2X1 NAND2X1_412 ( .A(REGs_FIRQ_REGS_5__27_), .B(_1573__bF_buf46), .Y(_4723_) );
MUX2X1 MUX2X1_412 ( .A(_1627__bF_buf1), .B(_4723_), .S(_4695__bF_buf1), .Y(_1338_) );
NAND2X1 NAND2X1_413 ( .A(REGs_FIRQ_REGS_5__28_), .B(_1573__bF_buf53), .Y(_4724_) );
MUX2X1 MUX2X1_413 ( .A(_1629__bF_buf2), .B(_4724_), .S(_4695__bF_buf4), .Y(_1339_) );
NAND2X1 NAND2X1_414 ( .A(REGs_FIRQ_REGS_5__29_), .B(_1573__bF_buf1), .Y(_4725_) );
MUX2X1 MUX2X1_414 ( .A(_1631__bF_buf0), .B(_4725_), .S(_4695__bF_buf3), .Y(_1340_) );
NAND2X1 NAND2X1_415 ( .A(REGs_FIRQ_REGS_5__30_), .B(_1573__bF_buf23), .Y(_4726_) );
MUX2X1 MUX2X1_415 ( .A(_1633__bF_buf3), .B(_4726_), .S(_4695__bF_buf2), .Y(_1341_) );
NAND2X1 NAND2X1_416 ( .A(REGs_FIRQ_REGS_5__31_), .B(_1573__bF_buf70), .Y(_4727_) );
MUX2X1 MUX2X1_416 ( .A(_1635__bF_buf2), .B(_4727_), .S(_4695__bF_buf4), .Y(_1342_) );
NOR2X1 NOR2X1_11 ( .A(_1571_), .B(_4358_), .Y(_4728_) );
NAND2X1 NAND2X1_417 ( .A(REGs_FIRQ_REGS_6__0_), .B(_1573__bF_buf59), .Y(_4729_) );
MUX2X1 MUX2X1_417 ( .A(_1567__bF_buf3), .B(_4729_), .S(_4728__bF_buf0), .Y(_1343_) );
NAND2X1 NAND2X1_418 ( .A(REGs_FIRQ_REGS_6__1_), .B(_1573__bF_buf53), .Y(_4730_) );
MUX2X1 MUX2X1_418 ( .A(_1575__bF_buf0), .B(_4730_), .S(_4728__bF_buf4), .Y(_1344_) );
NAND2X1 NAND2X1_419 ( .A(REGs_FIRQ_REGS_6__2_), .B(_1573__bF_buf61), .Y(_4731_) );
MUX2X1 MUX2X1_419 ( .A(_1577__bF_buf2), .B(_4731_), .S(_4728__bF_buf0), .Y(_1345_) );
NAND2X1 NAND2X1_420 ( .A(REGs_FIRQ_REGS_6__3_), .B(_1573__bF_buf61), .Y(_4732_) );
MUX2X1 MUX2X1_420 ( .A(_1579__bF_buf0), .B(_4732_), .S(_4728__bF_buf0), .Y(_1346_) );
NAND2X1 NAND2X1_421 ( .A(REGs_FIRQ_REGS_6__4_), .B(_1573__bF_buf27), .Y(_4733_) );
MUX2X1 MUX2X1_421 ( .A(_1581__bF_buf2), .B(_4733_), .S(_4728__bF_buf2), .Y(_1347_) );
NAND2X1 NAND2X1_422 ( .A(REGs_FIRQ_REGS_6__5_), .B(_1573__bF_buf45), .Y(_4734_) );
MUX2X1 MUX2X1_422 ( .A(_1583__bF_buf1), .B(_4734_), .S(_4728__bF_buf1), .Y(_1348_) );
NAND2X1 NAND2X1_423 ( .A(REGs_FIRQ_REGS_6__6_), .B(_1573__bF_buf38), .Y(_4735_) );
MUX2X1 MUX2X1_423 ( .A(_1585__bF_buf1), .B(_4735_), .S(_4728__bF_buf2), .Y(_1349_) );
NAND2X1 NAND2X1_424 ( .A(REGs_FIRQ_REGS_6__7_), .B(_1573__bF_buf55), .Y(_4736_) );
MUX2X1 MUX2X1_424 ( .A(_1587__bF_buf2), .B(_4736_), .S(_4728__bF_buf2), .Y(_1350_) );
NAND2X1 NAND2X1_425 ( .A(REGs_FIRQ_REGS_6__8_), .B(_1573__bF_buf74), .Y(_4737_) );
MUX2X1 MUX2X1_425 ( .A(_1589__bF_buf0), .B(_4737_), .S(_4728__bF_buf4), .Y(_1351_) );
NAND2X1 NAND2X1_426 ( .A(REGs_FIRQ_REGS_6__9_), .B(_1573__bF_buf45), .Y(_4738_) );
MUX2X1 MUX2X1_426 ( .A(_1591__bF_buf1), .B(_4738_), .S(_4728__bF_buf4), .Y(_1352_) );
NAND2X1 NAND2X1_427 ( .A(REGs_FIRQ_REGS_6__10_), .B(_1573__bF_buf9), .Y(_4739_) );
MUX2X1 MUX2X1_427 ( .A(_1593__bF_buf3), .B(_4739_), .S(_4728__bF_buf1), .Y(_1353_) );
NAND2X1 NAND2X1_428 ( .A(REGs_FIRQ_REGS_6__11_), .B(_1573__bF_buf78), .Y(_4740_) );
MUX2X1 MUX2X1_428 ( .A(_1595__bF_buf3), .B(_4740_), .S(_4728__bF_buf4), .Y(_1354_) );
NAND2X1 NAND2X1_429 ( .A(REGs_FIRQ_REGS_6__12_), .B(_1573__bF_buf22), .Y(_4741_) );
MUX2X1 MUX2X1_429 ( .A(_1597__bF_buf3), .B(_4741_), .S(_4728__bF_buf3), .Y(_1355_) );
NAND2X1 NAND2X1_430 ( .A(REGs_FIRQ_REGS_6__13_), .B(_1573__bF_buf32), .Y(_4742_) );
MUX2X1 MUX2X1_430 ( .A(_1599__bF_buf0), .B(_4742_), .S(_4728__bF_buf3), .Y(_1356_) );
NAND2X1 NAND2X1_431 ( .A(REGs_FIRQ_REGS_6__14_), .B(_1573__bF_buf9), .Y(_4743_) );
MUX2X1 MUX2X1_431 ( .A(_1601__bF_buf3), .B(_4743_), .S(_4728__bF_buf1), .Y(_1357_) );
NAND2X1 NAND2X1_432 ( .A(REGs_FIRQ_REGS_6__15_), .B(_1573__bF_buf44), .Y(_4744_) );
MUX2X1 MUX2X1_432 ( .A(_1603__bF_buf3), .B(_4744_), .S(_4728__bF_buf4), .Y(_1358_) );
NAND2X1 NAND2X1_433 ( .A(REGs_FIRQ_REGS_6__16_), .B(_1573__bF_buf45), .Y(_4745_) );
MUX2X1 MUX2X1_433 ( .A(_1605__bF_buf0), .B(_4745_), .S(_4728__bF_buf4), .Y(_1359_) );
NAND2X1 NAND2X1_434 ( .A(REGs_FIRQ_REGS_6__17_), .B(_1573__bF_buf61), .Y(_4746_) );
MUX2X1 MUX2X1_434 ( .A(_1607__bF_buf3), .B(_4746_), .S(_4728__bF_buf0), .Y(_1360_) );
NAND2X1 NAND2X1_435 ( .A(REGs_FIRQ_REGS_6__18_), .B(_1573__bF_buf70), .Y(_4747_) );
MUX2X1 MUX2X1_435 ( .A(_1609__bF_buf3), .B(_4747_), .S(_4728__bF_buf4), .Y(_1361_) );
NAND2X1 NAND2X1_436 ( .A(REGs_FIRQ_REGS_6__19_), .B(_1573__bF_buf43), .Y(_4748_) );
MUX2X1 MUX2X1_436 ( .A(_1611__bF_buf2), .B(_4748_), .S(_4728__bF_buf3), .Y(_1362_) );
NAND2X1 NAND2X1_437 ( .A(REGs_FIRQ_REGS_6__20_), .B(_1573__bF_buf32), .Y(_4749_) );
MUX2X1 MUX2X1_437 ( .A(_1613__bF_buf0), .B(_4749_), .S(_4728__bF_buf0), .Y(_1363_) );
NAND2X1 NAND2X1_438 ( .A(REGs_FIRQ_REGS_6__21_), .B(_1573__bF_buf64), .Y(_4750_) );
MUX2X1 MUX2X1_438 ( .A(_1615__bF_buf0), .B(_4750_), .S(_4728__bF_buf1), .Y(_1364_) );
NAND2X1 NAND2X1_439 ( .A(REGs_FIRQ_REGS_6__22_), .B(_1573__bF_buf27), .Y(_4751_) );
MUX2X1 MUX2X1_439 ( .A(_1617__bF_buf3), .B(_4751_), .S(_4728__bF_buf2), .Y(_1365_) );
NAND2X1 NAND2X1_440 ( .A(REGs_FIRQ_REGS_6__23_), .B(_1573__bF_buf64), .Y(_4752_) );
MUX2X1 MUX2X1_440 ( .A(_1619__bF_buf2), .B(_4752_), .S(_4728__bF_buf1), .Y(_1366_) );
NAND2X1 NAND2X1_441 ( .A(REGs_FIRQ_REGS_6__24_), .B(_1573__bF_buf43), .Y(_4753_) );
MUX2X1 MUX2X1_441 ( .A(_1621__bF_buf1), .B(_4753_), .S(_4728__bF_buf3), .Y(_1367_) );
NAND2X1 NAND2X1_442 ( .A(REGs_FIRQ_REGS_6__25_), .B(_1573__bF_buf71), .Y(_4754_) );
MUX2X1 MUX2X1_442 ( .A(_1623__bF_buf0), .B(_4754_), .S(_4728__bF_buf3), .Y(_1368_) );
NAND2X1 NAND2X1_443 ( .A(REGs_FIRQ_REGS_6__26_), .B(_1573__bF_buf48), .Y(_4755_) );
MUX2X1 MUX2X1_443 ( .A(_1625__bF_buf0), .B(_4755_), .S(_4728__bF_buf2), .Y(_1369_) );
NAND2X1 NAND2X1_444 ( .A(REGs_FIRQ_REGS_6__27_), .B(_1573__bF_buf48), .Y(_4756_) );
MUX2X1 MUX2X1_444 ( .A(_1627__bF_buf2), .B(_4756_), .S(_4728__bF_buf2), .Y(_1370_) );
NAND2X1 NAND2X1_445 ( .A(REGs_FIRQ_REGS_6__28_), .B(_1573__bF_buf21), .Y(_4757_) );
MUX2X1 MUX2X1_445 ( .A(_1629__bF_buf0), .B(_4757_), .S(_4728__bF_buf1), .Y(_1371_) );
NAND2X1 NAND2X1_446 ( .A(REGs_FIRQ_REGS_6__29_), .B(_1573__bF_buf30), .Y(_4758_) );
MUX2X1 MUX2X1_446 ( .A(_1631__bF_buf0), .B(_4758_), .S(_4728__bF_buf3), .Y(_1372_) );
NAND2X1 NAND2X1_447 ( .A(REGs_FIRQ_REGS_6__30_), .B(_1573__bF_buf22), .Y(_4759_) );
MUX2X1 MUX2X1_447 ( .A(_1633__bF_buf0), .B(_4759_), .S(_4728__bF_buf3), .Y(_1373_) );
NAND2X1 NAND2X1_448 ( .A(REGs_FIRQ_REGS_6__31_), .B(_1573__bF_buf58), .Y(_4760_) );
MUX2X1 MUX2X1_448 ( .A(_1635__bF_buf0), .B(_4760_), .S(_4728__bF_buf0), .Y(_1374_) );
NOR2X1 NOR2X1_12 ( .A(_4529_), .B(_1569_), .Y(_4761_) );
NAND2X1 NAND2X1_449 ( .A(REGs_USR_REGS_4__0_), .B(_1573__bF_buf54), .Y(_4762_) );
MUX2X1 MUX2X1_449 ( .A(_1567__bF_buf3), .B(_4762_), .S(_4761__bF_buf0), .Y(_1375_) );
NAND2X1 NAND2X1_450 ( .A(REGs_USR_REGS_4__1_), .B(_1573__bF_buf52), .Y(_4763_) );
MUX2X1 MUX2X1_450 ( .A(_1575__bF_buf1), .B(_4763_), .S(_4761__bF_buf1), .Y(_1376_) );
NAND2X1 NAND2X1_451 ( .A(REGs_USR_REGS_4__2_), .B(_1573__bF_buf34), .Y(_4764_) );
MUX2X1 MUX2X1_451 ( .A(_1577__bF_buf0), .B(_4764_), .S(_4761__bF_buf4), .Y(_1377_) );
NAND2X1 NAND2X1_452 ( .A(REGs_USR_REGS_4__3_), .B(_1573__bF_buf23), .Y(_4765_) );
MUX2X1 MUX2X1_452 ( .A(_1579__bF_buf0), .B(_4765_), .S(_4761__bF_buf4), .Y(_1378_) );
NAND2X1 NAND2X1_453 ( .A(REGs_USR_REGS_4__4_), .B(_1573__bF_buf27), .Y(_4766_) );
MUX2X1 MUX2X1_453 ( .A(_1581__bF_buf2), .B(_4766_), .S(_4761__bF_buf4), .Y(_1379_) );
NAND2X1 NAND2X1_454 ( .A(REGs_USR_REGS_4__5_), .B(_1573__bF_buf14), .Y(_4767_) );
MUX2X1 MUX2X1_454 ( .A(_1583__bF_buf2), .B(_4767_), .S(_4761__bF_buf2), .Y(_1380_) );
NAND2X1 NAND2X1_455 ( .A(REGs_USR_REGS_4__6_), .B(_1573__bF_buf38), .Y(_4768_) );
MUX2X1 MUX2X1_455 ( .A(_1585__bF_buf0), .B(_4768_), .S(_4761__bF_buf4), .Y(_1381_) );
NAND2X1 NAND2X1_456 ( .A(REGs_USR_REGS_4__7_), .B(_1573__bF_buf5), .Y(_4769_) );
MUX2X1 MUX2X1_456 ( .A(_1587__bF_buf1), .B(_4769_), .S(_4761__bF_buf3), .Y(_1382_) );
NAND2X1 NAND2X1_457 ( .A(REGs_USR_REGS_4__8_), .B(_1573__bF_buf26), .Y(_4770_) );
MUX2X1 MUX2X1_457 ( .A(_1589__bF_buf3), .B(_4770_), .S(_4761__bF_buf0), .Y(_1383_) );
NAND2X1 NAND2X1_458 ( .A(REGs_USR_REGS_4__9_), .B(_1573__bF_buf60), .Y(_4771_) );
MUX2X1 MUX2X1_458 ( .A(_1591__bF_buf3), .B(_4771_), .S(_4761__bF_buf1), .Y(_1384_) );
NAND2X1 NAND2X1_459 ( .A(REGs_USR_REGS_4__10_), .B(_1573__bF_buf70), .Y(_4772_) );
MUX2X1 MUX2X1_459 ( .A(_1593__bF_buf3), .B(_4772_), .S(_4761__bF_buf2), .Y(_1385_) );
NAND2X1 NAND2X1_460 ( .A(REGs_USR_REGS_4__11_), .B(_1573__bF_buf53), .Y(_4773_) );
MUX2X1 MUX2X1_460 ( .A(_1595__bF_buf3), .B(_4773_), .S(_4761__bF_buf2), .Y(_1386_) );
NAND2X1 NAND2X1_461 ( .A(REGs_USR_REGS_4__12_), .B(_1573__bF_buf3), .Y(_4774_) );
MUX2X1 MUX2X1_461 ( .A(_1597__bF_buf1), .B(_4774_), .S(_4761__bF_buf4), .Y(_1387_) );
NAND2X1 NAND2X1_462 ( .A(REGs_USR_REGS_4__13_), .B(_1573__bF_buf1), .Y(_4775_) );
MUX2X1 MUX2X1_462 ( .A(_1599__bF_buf3), .B(_4775_), .S(_4761__bF_buf0), .Y(_1388_) );
NAND2X1 NAND2X1_463 ( .A(REGs_USR_REGS_4__14_), .B(_1573__bF_buf60), .Y(_4776_) );
MUX2X1 MUX2X1_463 ( .A(_1601__bF_buf2), .B(_4776_), .S(_4761__bF_buf1), .Y(_1389_) );
NAND2X1 NAND2X1_464 ( .A(REGs_USR_REGS_4__15_), .B(_1573__bF_buf63), .Y(_4777_) );
MUX2X1 MUX2X1_464 ( .A(_1603__bF_buf3), .B(_4777_), .S(_4761__bF_buf2), .Y(_1390_) );
NAND2X1 NAND2X1_465 ( .A(REGs_USR_REGS_4__16_), .B(_1573__bF_buf52), .Y(_4778_) );
MUX2X1 MUX2X1_465 ( .A(_1605__bF_buf1), .B(_4778_), .S(_4761__bF_buf1), .Y(_1391_) );
NAND2X1 NAND2X1_466 ( .A(REGs_USR_REGS_4__17_), .B(_1573__bF_buf6), .Y(_4779_) );
MUX2X1 MUX2X1_466 ( .A(_1607__bF_buf1), .B(_4779_), .S(_4761__bF_buf3), .Y(_1392_) );
NAND2X1 NAND2X1_467 ( .A(REGs_USR_REGS_4__18_), .B(_1573__bF_buf52), .Y(_4780_) );
MUX2X1 MUX2X1_467 ( .A(_1609__bF_buf2), .B(_4780_), .S(_4761__bF_buf1), .Y(_1393_) );
NAND2X1 NAND2X1_468 ( .A(REGs_USR_REGS_4__19_), .B(_1573__bF_buf16), .Y(_4781_) );
MUX2X1 MUX2X1_468 ( .A(_1611__bF_buf1), .B(_4781_), .S(_4761__bF_buf0), .Y(_1394_) );
NAND2X1 NAND2X1_469 ( .A(REGs_USR_REGS_4__20_), .B(_1573__bF_buf5), .Y(_4782_) );
MUX2X1 MUX2X1_469 ( .A(_1613__bF_buf3), .B(_4782_), .S(_4761__bF_buf3), .Y(_1395_) );
NAND2X1 NAND2X1_470 ( .A(REGs_USR_REGS_4__21_), .B(_1573__bF_buf26), .Y(_4783_) );
MUX2X1 MUX2X1_470 ( .A(_1615__bF_buf2), .B(_4783_), .S(_4761__bF_buf0), .Y(_1396_) );
NAND2X1 NAND2X1_471 ( .A(REGs_USR_REGS_4__22_), .B(_1573__bF_buf38), .Y(_4784_) );
MUX2X1 MUX2X1_471 ( .A(_1617__bF_buf3), .B(_4784_), .S(_4761__bF_buf4), .Y(_1397_) );
NAND2X1 NAND2X1_472 ( .A(REGs_USR_REGS_4__23_), .B(_1573__bF_buf52), .Y(_4785_) );
MUX2X1 MUX2X1_472 ( .A(_1619__bF_buf3), .B(_4785_), .S(_4761__bF_buf1), .Y(_1398_) );
NAND2X1 NAND2X1_473 ( .A(REGs_USR_REGS_4__24_), .B(_1573__bF_buf71), .Y(_4786_) );
MUX2X1 MUX2X1_473 ( .A(_1621__bF_buf0), .B(_4786_), .S(_4761__bF_buf3), .Y(_1399_) );
NAND2X1 NAND2X1_474 ( .A(REGs_USR_REGS_4__25_), .B(_1573__bF_buf71), .Y(_4787_) );
MUX2X1 MUX2X1_474 ( .A(_1623__bF_buf3), .B(_4787_), .S(_4761__bF_buf3), .Y(_1400_) );
NAND2X1 NAND2X1_475 ( .A(REGs_USR_REGS_4__26_), .B(_1573__bF_buf38), .Y(_4788_) );
MUX2X1 MUX2X1_475 ( .A(_1625__bF_buf2), .B(_4788_), .S(_4761__bF_buf4), .Y(_1401_) );
NAND2X1 NAND2X1_476 ( .A(REGs_USR_REGS_4__27_), .B(_1573__bF_buf22), .Y(_4789_) );
MUX2X1 MUX2X1_476 ( .A(_1627__bF_buf2), .B(_4789_), .S(_4761__bF_buf3), .Y(_1402_) );
NAND2X1 NAND2X1_477 ( .A(REGs_USR_REGS_4__28_), .B(_1573__bF_buf70), .Y(_4790_) );
MUX2X1 MUX2X1_477 ( .A(_1629__bF_buf0), .B(_4790_), .S(_4761__bF_buf2), .Y(_1403_) );
NAND2X1 NAND2X1_478 ( .A(REGs_USR_REGS_4__29_), .B(_1573__bF_buf39), .Y(_4791_) );
MUX2X1 MUX2X1_478 ( .A(_1631__bF_buf1), .B(_4791_), .S(_4761__bF_buf0), .Y(_1404_) );
NAND2X1 NAND2X1_479 ( .A(REGs_USR_REGS_4__30_), .B(_1573__bF_buf7), .Y(_4792_) );
MUX2X1 MUX2X1_479 ( .A(_1633__bF_buf2), .B(_4792_), .S(_4761__bF_buf3), .Y(_1405_) );
NAND2X1 NAND2X1_480 ( .A(REGs_USR_REGS_4__31_), .B(_1573__bF_buf70), .Y(_4793_) );
MUX2X1 MUX2X1_480 ( .A(_1635__bF_buf2), .B(_4793_), .S(_4761__bF_buf2), .Y(_1406_) );
NOR2X1 NOR2X1_13 ( .A(_4324_), .B(_4358_), .Y(_4794_) );
NAND2X1 NAND2X1_481 ( .A(REGs_FIRQ_REGS_7__0_), .B(_1573__bF_buf40), .Y(_4795_) );
MUX2X1 MUX2X1_481 ( .A(_1567__bF_buf0), .B(_4795_), .S(_4794__bF_buf1), .Y(_1407_) );
NAND2X1 NAND2X1_482 ( .A(REGs_FIRQ_REGS_7__1_), .B(_1573__bF_buf14), .Y(_4796_) );
MUX2X1 MUX2X1_482 ( .A(_1575__bF_buf1), .B(_4796_), .S(_4794__bF_buf4), .Y(_1408_) );
NAND2X1 NAND2X1_483 ( .A(REGs_FIRQ_REGS_7__2_), .B(_1573__bF_buf34), .Y(_4797_) );
MUX2X1 MUX2X1_483 ( .A(_1577__bF_buf0), .B(_4797_), .S(_4794__bF_buf3), .Y(_1409_) );
NAND2X1 NAND2X1_484 ( .A(REGs_FIRQ_REGS_7__3_), .B(_1573__bF_buf47), .Y(_4798_) );
MUX2X1 MUX2X1_484 ( .A(_1579__bF_buf3), .B(_4798_), .S(_4794__bF_buf2), .Y(_1410_) );
NAND2X1 NAND2X1_485 ( .A(REGs_FIRQ_REGS_7__4_), .B(_1573__bF_buf72), .Y(_4799_) );
MUX2X1 MUX2X1_485 ( .A(_1581__bF_buf3), .B(_4799_), .S(_4794__bF_buf2), .Y(_1411_) );
NAND2X1 NAND2X1_486 ( .A(REGs_FIRQ_REGS_7__5_), .B(_1573__bF_buf78), .Y(_4800_) );
MUX2X1 MUX2X1_486 ( .A(_1583__bF_buf1), .B(_4800_), .S(_4794__bF_buf4), .Y(_1412_) );
NAND2X1 NAND2X1_487 ( .A(REGs_FIRQ_REGS_7__6_), .B(_1573__bF_buf72), .Y(_4801_) );
MUX2X1 MUX2X1_487 ( .A(_1585__bF_buf1), .B(_4801_), .S(_4794__bF_buf2), .Y(_1413_) );
NAND2X1 NAND2X1_488 ( .A(REGs_FIRQ_REGS_7__7_), .B(_1573__bF_buf7), .Y(_4802_) );
MUX2X1 MUX2X1_488 ( .A(_1587__bF_buf2), .B(_4802_), .S(_4794__bF_buf3), .Y(_1414_) );
NAND2X1 NAND2X1_489 ( .A(REGs_FIRQ_REGS_7__8_), .B(_1573__bF_buf64), .Y(_4803_) );
MUX2X1 MUX2X1_489 ( .A(_1589__bF_buf3), .B(_4803_), .S(_4794__bF_buf0), .Y(_1415_) );
NAND2X1 NAND2X1_490 ( .A(REGs_FIRQ_REGS_7__9_), .B(_1573__bF_buf21), .Y(_4804_) );
MUX2X1 MUX2X1_490 ( .A(_1591__bF_buf1), .B(_4804_), .S(_4794__bF_buf0), .Y(_1416_) );
NAND2X1 NAND2X1_491 ( .A(REGs_FIRQ_REGS_7__10_), .B(_1573__bF_buf44), .Y(_4805_) );
MUX2X1 MUX2X1_491 ( .A(_1593__bF_buf2), .B(_4805_), .S(_4794__bF_buf4), .Y(_1417_) );
NAND2X1 NAND2X1_492 ( .A(REGs_FIRQ_REGS_7__11_), .B(_1573__bF_buf14), .Y(_4806_) );
MUX2X1 MUX2X1_492 ( .A(_1595__bF_buf3), .B(_4806_), .S(_4794__bF_buf4), .Y(_1418_) );
NAND2X1 NAND2X1_493 ( .A(REGs_FIRQ_REGS_7__12_), .B(_1573__bF_buf72), .Y(_4807_) );
MUX2X1 MUX2X1_493 ( .A(_1597__bF_buf1), .B(_4807_), .S(_4794__bF_buf2), .Y(_1419_) );
NAND2X1 NAND2X1_494 ( .A(REGs_FIRQ_REGS_7__13_), .B(_1573__bF_buf43), .Y(_4808_) );
MUX2X1 MUX2X1_494 ( .A(_1599__bF_buf3), .B(_4808_), .S(_4794__bF_buf1), .Y(_1420_) );
NAND2X1 NAND2X1_495 ( .A(REGs_FIRQ_REGS_7__14_), .B(_1573__bF_buf60), .Y(_4809_) );
MUX2X1 MUX2X1_495 ( .A(_1601__bF_buf2), .B(_4809_), .S(_4794__bF_buf4), .Y(_1421_) );
NAND2X1 NAND2X1_496 ( .A(REGs_FIRQ_REGS_7__15_), .B(_1573__bF_buf78), .Y(_4810_) );
MUX2X1 MUX2X1_496 ( .A(_1603__bF_buf3), .B(_4810_), .S(_4794__bF_buf4), .Y(_1422_) );
NAND2X1 NAND2X1_497 ( .A(REGs_FIRQ_REGS_7__16_), .B(_1573__bF_buf45), .Y(_4811_) );
MUX2X1 MUX2X1_497 ( .A(_1605__bF_buf0), .B(_4811_), .S(_4794__bF_buf0), .Y(_1423_) );
NAND2X1 NAND2X1_498 ( .A(REGs_FIRQ_REGS_7__17_), .B(_1573__bF_buf47), .Y(_4812_) );
MUX2X1 MUX2X1_498 ( .A(_1607__bF_buf3), .B(_4812_), .S(_4794__bF_buf3), .Y(_1424_) );
NAND2X1 NAND2X1_499 ( .A(REGs_FIRQ_REGS_7__18_), .B(_1573__bF_buf44), .Y(_4813_) );
MUX2X1 MUX2X1_499 ( .A(_1609__bF_buf2), .B(_4813_), .S(_4794__bF_buf4), .Y(_1425_) );
NAND2X1 NAND2X1_500 ( .A(REGs_FIRQ_REGS_7__19_), .B(_1573__bF_buf43), .Y(_4814_) );
MUX2X1 MUX2X1_500 ( .A(_1611__bF_buf2), .B(_4814_), .S(_4794__bF_buf1), .Y(_1426_) );
NAND2X1 NAND2X1_501 ( .A(REGs_FIRQ_REGS_7__20_), .B(_1573__bF_buf7), .Y(_4815_) );
MUX2X1 MUX2X1_501 ( .A(_1613__bF_buf0), .B(_4815_), .S(_4794__bF_buf3), .Y(_1427_) );
NAND2X1 NAND2X1_502 ( .A(REGs_FIRQ_REGS_7__21_), .B(_1573__bF_buf64), .Y(_4816_) );
MUX2X1 MUX2X1_502 ( .A(_1615__bF_buf0), .B(_4816_), .S(_4794__bF_buf0), .Y(_1428_) );
NAND2X1 NAND2X1_503 ( .A(REGs_FIRQ_REGS_7__22_), .B(_1573__bF_buf46), .Y(_4817_) );
MUX2X1 MUX2X1_503 ( .A(_1617__bF_buf2), .B(_4817_), .S(_4794__bF_buf2), .Y(_1429_) );
NAND2X1 NAND2X1_504 ( .A(REGs_FIRQ_REGS_7__23_), .B(_1573__bF_buf21), .Y(_4818_) );
MUX2X1 MUX2X1_504 ( .A(_1619__bF_buf2), .B(_4818_), .S(_4794__bF_buf0), .Y(_1430_) );
NAND2X1 NAND2X1_505 ( .A(REGs_FIRQ_REGS_7__24_), .B(_1573__bF_buf43), .Y(_4819_) );
MUX2X1 MUX2X1_505 ( .A(_1621__bF_buf1), .B(_4819_), .S(_4794__bF_buf1), .Y(_1431_) );
NAND2X1 NAND2X1_506 ( .A(REGs_FIRQ_REGS_7__25_), .B(_1573__bF_buf30), .Y(_4820_) );
MUX2X1 MUX2X1_506 ( .A(_1623__bF_buf0), .B(_4820_), .S(_4794__bF_buf1), .Y(_1432_) );
NAND2X1 NAND2X1_507 ( .A(REGs_FIRQ_REGS_7__26_), .B(_1573__bF_buf55), .Y(_4821_) );
MUX2X1 MUX2X1_507 ( .A(_1625__bF_buf2), .B(_4821_), .S(_4794__bF_buf3), .Y(_1433_) );
NAND2X1 NAND2X1_508 ( .A(REGs_FIRQ_REGS_7__27_), .B(_1573__bF_buf46), .Y(_4822_) );
MUX2X1 MUX2X1_508 ( .A(_1627__bF_buf1), .B(_4822_), .S(_4794__bF_buf3), .Y(_1434_) );
NAND2X1 NAND2X1_509 ( .A(REGs_FIRQ_REGS_7__28_), .B(_1573__bF_buf21), .Y(_4823_) );
MUX2X1 MUX2X1_509 ( .A(_1629__bF_buf0), .B(_4823_), .S(_4794__bF_buf0), .Y(_1435_) );
NAND2X1 NAND2X1_510 ( .A(REGs_FIRQ_REGS_7__29_), .B(_1573__bF_buf43), .Y(_4824_) );
MUX2X1 MUX2X1_510 ( .A(_1631__bF_buf0), .B(_4824_), .S(_4794__bF_buf1), .Y(_1436_) );
NAND2X1 NAND2X1_511 ( .A(REGs_FIRQ_REGS_7__30_), .B(_1573__bF_buf7), .Y(_4825_) );
MUX2X1 MUX2X1_511 ( .A(_1633__bF_buf2), .B(_4825_), .S(_4794__bF_buf3), .Y(_1437_) );
NAND2X1 NAND2X1_512 ( .A(REGs_FIRQ_REGS_7__31_), .B(_1573__bF_buf24), .Y(_4826_) );
MUX2X1 MUX2X1_512 ( .A(_1635__bF_buf0), .B(_4826_), .S(_4794__bF_buf2), .Y(_1438_) );
NOR2X1 NOR2X1_14 ( .A(_1569_), .B(_4394_), .Y(_4827_) );
NAND2X1 NAND2X1_513 ( .A(REGs_USR_REGS_3__0_), .B(_1573__bF_buf76), .Y(_4828_) );
MUX2X1 MUX2X1_513 ( .A(_1567__bF_buf2), .B(_4828_), .S(_4827__bF_buf2), .Y(_1439_) );
NAND2X1 NAND2X1_514 ( .A(REGs_USR_REGS_3__1_), .B(_1573__bF_buf26), .Y(_4829_) );
MUX2X1 MUX2X1_514 ( .A(_1575__bF_buf2), .B(_4829_), .S(_4827__bF_buf0), .Y(_1440_) );
NAND2X1 NAND2X1_515 ( .A(REGs_USR_REGS_3__2_), .B(_1573__bF_buf61), .Y(_4830_) );
MUX2X1 MUX2X1_515 ( .A(_1577__bF_buf2), .B(_4830_), .S(_4827__bF_buf3), .Y(_1441_) );
NAND2X1 NAND2X1_516 ( .A(REGs_USR_REGS_3__3_), .B(_1573__bF_buf59), .Y(_4831_) );
MUX2X1 MUX2X1_516 ( .A(_1579__bF_buf1), .B(_4831_), .S(_4827__bF_buf3), .Y(_1442_) );
NAND2X1 NAND2X1_517 ( .A(REGs_USR_REGS_3__4_), .B(_1573__bF_buf11), .Y(_4832_) );
MUX2X1 MUX2X1_517 ( .A(_1581__bF_buf0), .B(_4832_), .S(_4827__bF_buf2), .Y(_1443_) );
NAND2X1 NAND2X1_518 ( .A(REGs_USR_REGS_3__5_), .B(_1573__bF_buf8), .Y(_4833_) );
MUX2X1 MUX2X1_518 ( .A(_1583__bF_buf2), .B(_4833_), .S(_4827__bF_buf4), .Y(_1444_) );
NAND2X1 NAND2X1_519 ( .A(REGs_USR_REGS_3__6_), .B(_1573__bF_buf37), .Y(_4834_) );
MUX2X1 MUX2X1_519 ( .A(_1585__bF_buf2), .B(_4834_), .S(_4827__bF_buf2), .Y(_1445_) );
NAND2X1 NAND2X1_520 ( .A(REGs_USR_REGS_3__7_), .B(_1573__bF_buf35), .Y(_4835_) );
MUX2X1 MUX2X1_520 ( .A(_1587__bF_buf0), .B(_4835_), .S(_4827__bF_buf1), .Y(_1446_) );
NAND2X1 NAND2X1_521 ( .A(REGs_USR_REGS_3__8_), .B(_1573__bF_buf28), .Y(_4836_) );
MUX2X1 MUX2X1_521 ( .A(_1589__bF_buf2), .B(_4836_), .S(_4827__bF_buf4), .Y(_1447_) );
NAND2X1 NAND2X1_522 ( .A(REGs_USR_REGS_3__9_), .B(_1573__bF_buf13), .Y(_4837_) );
MUX2X1 MUX2X1_522 ( .A(_1591__bF_buf0), .B(_4837_), .S(_4827__bF_buf0), .Y(_1448_) );
NAND2X1 NAND2X1_523 ( .A(REGs_USR_REGS_3__10_), .B(_1573__bF_buf68), .Y(_4838_) );
MUX2X1 MUX2X1_523 ( .A(_1593__bF_buf2), .B(_4838_), .S(_4827__bF_buf4), .Y(_1449_) );
NAND2X1 NAND2X1_524 ( .A(REGs_USR_REGS_3__11_), .B(_1573__bF_buf28), .Y(_4839_) );
MUX2X1 MUX2X1_524 ( .A(_1595__bF_buf1), .B(_4839_), .S(_4827__bF_buf4), .Y(_1450_) );
NAND2X1 NAND2X1_525 ( .A(REGs_USR_REGS_3__12_), .B(_1573__bF_buf57), .Y(_4840_) );
MUX2X1 MUX2X1_525 ( .A(_1597__bF_buf2), .B(_4840_), .S(_4827__bF_buf2), .Y(_1451_) );
NAND2X1 NAND2X1_526 ( .A(REGs_USR_REGS_3__13_), .B(_1573__bF_buf35), .Y(_4841_) );
MUX2X1 MUX2X1_526 ( .A(_1599__bF_buf1), .B(_4841_), .S(_4827__bF_buf1), .Y(_1452_) );
NAND2X1 NAND2X1_527 ( .A(REGs_USR_REGS_3__14_), .B(_1573__bF_buf77), .Y(_4842_) );
MUX2X1 MUX2X1_527 ( .A(_1601__bF_buf1), .B(_4842_), .S(_4827__bF_buf0), .Y(_1453_) );
NAND2X1 NAND2X1_528 ( .A(REGs_USR_REGS_3__15_), .B(_1573__bF_buf50), .Y(_4843_) );
MUX2X1 MUX2X1_528 ( .A(_1603__bF_buf1), .B(_4843_), .S(_4827__bF_buf0), .Y(_1454_) );
NAND2X1 NAND2X1_529 ( .A(REGs_USR_REGS_3__16_), .B(_1573__bF_buf68), .Y(_4844_) );
MUX2X1 MUX2X1_529 ( .A(_1605__bF_buf1), .B(_4844_), .S(_4827__bF_buf4), .Y(_1455_) );
NAND2X1 NAND2X1_530 ( .A(REGs_USR_REGS_3__17_), .B(_1573__bF_buf12), .Y(_4845_) );
MUX2X1 MUX2X1_530 ( .A(_1607__bF_buf2), .B(_4845_), .S(_4827__bF_buf1), .Y(_1456_) );
NAND2X1 NAND2X1_531 ( .A(REGs_USR_REGS_3__18_), .B(_1573__bF_buf25), .Y(_4846_) );
MUX2X1 MUX2X1_531 ( .A(_1609__bF_buf0), .B(_4846_), .S(_4827__bF_buf0), .Y(_1457_) );
NAND2X1 NAND2X1_532 ( .A(REGs_USR_REGS_3__19_), .B(_1573__bF_buf54), .Y(_4847_) );
MUX2X1 MUX2X1_532 ( .A(_1611__bF_buf0), .B(_4847_), .S(_4827__bF_buf3), .Y(_1458_) );
NAND2X1 NAND2X1_533 ( .A(REGs_USR_REGS_3__20_), .B(_1573__bF_buf5), .Y(_4848_) );
MUX2X1 MUX2X1_533 ( .A(_1613__bF_buf3), .B(_4848_), .S(_4827__bF_buf1), .Y(_1459_) );
NAND2X1 NAND2X1_534 ( .A(REGs_USR_REGS_3__21_), .B(_1573__bF_buf8), .Y(_4849_) );
MUX2X1 MUX2X1_534 ( .A(_1615__bF_buf3), .B(_4849_), .S(_4827__bF_buf4), .Y(_1460_) );
NAND2X1 NAND2X1_535 ( .A(REGs_USR_REGS_3__22_), .B(_1573__bF_buf11), .Y(_4850_) );
MUX2X1 MUX2X1_535 ( .A(_1617__bF_buf1), .B(_4850_), .S(_4827__bF_buf2), .Y(_1461_) );
NAND2X1 NAND2X1_536 ( .A(REGs_USR_REGS_3__23_), .B(_1573__bF_buf26), .Y(_4851_) );
MUX2X1 MUX2X1_536 ( .A(_1619__bF_buf1), .B(_4851_), .S(_4827__bF_buf0), .Y(_1462_) );
NAND2X1 NAND2X1_537 ( .A(REGs_USR_REGS_3__24_), .B(_1573__bF_buf18), .Y(_4852_) );
MUX2X1 MUX2X1_537 ( .A(_1621__bF_buf3), .B(_4852_), .S(_4827__bF_buf3), .Y(_1463_) );
NAND2X1 NAND2X1_538 ( .A(REGs_USR_REGS_3__25_), .B(_1573__bF_buf35), .Y(_4853_) );
MUX2X1 MUX2X1_538 ( .A(_1623__bF_buf1), .B(_4853_), .S(_4827__bF_buf1), .Y(_1464_) );
NAND2X1 NAND2X1_539 ( .A(REGs_USR_REGS_3__26_), .B(_1573__bF_buf69), .Y(_4854_) );
MUX2X1 MUX2X1_539 ( .A(_1625__bF_buf3), .B(_4854_), .S(_4827__bF_buf2), .Y(_1465_) );
NAND2X1 NAND2X1_540 ( .A(REGs_USR_REGS_3__27_), .B(_1573__bF_buf12), .Y(_4855_) );
MUX2X1 MUX2X1_540 ( .A(_1627__bF_buf3), .B(_4855_), .S(_4827__bF_buf1), .Y(_1466_) );
NAND2X1 NAND2X1_541 ( .A(REGs_USR_REGS_3__28_), .B(_1573__bF_buf8), .Y(_4856_) );
MUX2X1 MUX2X1_541 ( .A(_1629__bF_buf2), .B(_4856_), .S(_4827__bF_buf4), .Y(_1467_) );
NAND2X1 NAND2X1_542 ( .A(REGs_USR_REGS_3__29_), .B(_1573__bF_buf58), .Y(_4857_) );
MUX2X1 MUX2X1_542 ( .A(_1631__bF_buf3), .B(_4857_), .S(_4827__bF_buf3), .Y(_1468_) );
NAND2X1 NAND2X1_543 ( .A(REGs_USR_REGS_3__30_), .B(_1573__bF_buf61), .Y(_4858_) );
MUX2X1 MUX2X1_543 ( .A(_1633__bF_buf2), .B(_4858_), .S(_4827__bF_buf3), .Y(_1469_) );
NAND2X1 NAND2X1_544 ( .A(REGs_USR_REGS_3__31_), .B(_1573__bF_buf54), .Y(_4859_) );
MUX2X1 MUX2X1_544 ( .A(_1635__bF_buf0), .B(_4859_), .S(_4827__bF_buf3), .Y(_1470_) );
NOR2X1 NOR2X1_15 ( .A(_4360_), .B(_1569_), .Y(_4860_) );
NAND2X1 NAND2X1_545 ( .A(REGs_USR_REGS_2__0_), .B(_1573__bF_buf58), .Y(_4861_) );
MUX2X1 MUX2X1_545 ( .A(_1567__bF_buf3), .B(_4861_), .S(_4860__bF_buf0), .Y(_1471_) );
NAND2X1 NAND2X1_546 ( .A(REGs_USR_REGS_2__1_), .B(_1573__bF_buf16), .Y(_4862_) );
MUX2X1 MUX2X1_546 ( .A(_1575__bF_buf2), .B(_4862_), .S(_4860__bF_buf0), .Y(_1472_) );
NAND2X1 NAND2X1_547 ( .A(REGs_USR_REGS_2__2_), .B(_1573__bF_buf22), .Y(_4863_) );
MUX2X1 MUX2X1_547 ( .A(_1577__bF_buf3), .B(_4863_), .S(_4860__bF_buf3), .Y(_1473_) );
NAND2X1 NAND2X1_548 ( .A(REGs_USR_REGS_2__3_), .B(_1573__bF_buf18), .Y(_4864_) );
MUX2X1 MUX2X1_548 ( .A(_1579__bF_buf1), .B(_4864_), .S(_4860__bF_buf1), .Y(_1474_) );
NAND2X1 NAND2X1_549 ( .A(REGs_USR_REGS_2__4_), .B(_1573__bF_buf37), .Y(_4865_) );
MUX2X1 MUX2X1_549 ( .A(_1581__bF_buf0), .B(_4865_), .S(_4860__bF_buf3), .Y(_1475_) );
NAND2X1 NAND2X1_550 ( .A(REGs_USR_REGS_2__5_), .B(_1573__bF_buf13), .Y(_4866_) );
MUX2X1 MUX2X1_550 ( .A(_1583__bF_buf0), .B(_4866_), .S(_4860__bF_buf0), .Y(_1476_) );
NAND2X1 NAND2X1_551 ( .A(REGs_USR_REGS_2__6_), .B(_1573__bF_buf69), .Y(_4867_) );
MUX2X1 MUX2X1_551 ( .A(_1585__bF_buf2), .B(_4867_), .S(_4860__bF_buf3), .Y(_1477_) );
NAND2X1 NAND2X1_552 ( .A(REGs_USR_REGS_2__7_), .B(_1573__bF_buf17), .Y(_4868_) );
MUX2X1 MUX2X1_552 ( .A(_1587__bF_buf0), .B(_4868_), .S(_4860__bF_buf2), .Y(_1478_) );
NAND2X1 NAND2X1_553 ( .A(REGs_USR_REGS_2__8_), .B(_1573__bF_buf16), .Y(_4869_) );
MUX2X1 MUX2X1_553 ( .A(_1589__bF_buf2), .B(_4869_), .S(_4860__bF_buf1), .Y(_1479_) );
NAND2X1 NAND2X1_554 ( .A(REGs_USR_REGS_2__9_), .B(_1573__bF_buf13), .Y(_4870_) );
MUX2X1 MUX2X1_554 ( .A(_1591__bF_buf0), .B(_4870_), .S(_4860__bF_buf0), .Y(_1480_) );
NAND2X1 NAND2X1_555 ( .A(REGs_USR_REGS_2__10_), .B(_1573__bF_buf63), .Y(_4871_) );
MUX2X1 MUX2X1_555 ( .A(_1593__bF_buf2), .B(_4871_), .S(_4860__bF_buf4), .Y(_1481_) );
NAND2X1 NAND2X1_556 ( .A(REGs_USR_REGS_2__11_), .B(_1573__bF_buf39), .Y(_4872_) );
MUX2X1 MUX2X1_556 ( .A(_1595__bF_buf1), .B(_4872_), .S(_4860__bF_buf1), .Y(_1482_) );
NAND2X1 NAND2X1_557 ( .A(REGs_USR_REGS_2__12_), .B(_1573__bF_buf57), .Y(_4873_) );
MUX2X1 MUX2X1_557 ( .A(_1597__bF_buf2), .B(_4873_), .S(_4860__bF_buf3), .Y(_1483_) );
NAND2X1 NAND2X1_558 ( .A(REGs_USR_REGS_2__13_), .B(_1573__bF_buf35), .Y(_4874_) );
MUX2X1 MUX2X1_558 ( .A(_1599__bF_buf1), .B(_4874_), .S(_4860__bF_buf2), .Y(_1484_) );
NAND2X1 NAND2X1_559 ( .A(REGs_USR_REGS_2__14_), .B(_1573__bF_buf63), .Y(_4875_) );
MUX2X1 MUX2X1_559 ( .A(_1601__bF_buf1), .B(_4875_), .S(_4860__bF_buf4), .Y(_1485_) );
NAND2X1 NAND2X1_560 ( .A(REGs_USR_REGS_2__15_), .B(_1573__bF_buf50), .Y(_4876_) );
MUX2X1 MUX2X1_560 ( .A(_1603__bF_buf1), .B(_4876_), .S(_4860__bF_buf4), .Y(_1486_) );
NAND2X1 NAND2X1_561 ( .A(REGs_USR_REGS_2__16_), .B(_1573__bF_buf63), .Y(_4877_) );
MUX2X1 MUX2X1_561 ( .A(_1605__bF_buf3), .B(_4877_), .S(_4860__bF_buf4), .Y(_1487_) );
NAND2X1 NAND2X1_562 ( .A(REGs_USR_REGS_2__17_), .B(_1573__bF_buf12), .Y(_4878_) );
MUX2X1 MUX2X1_562 ( .A(_1607__bF_buf2), .B(_4878_), .S(_4860__bF_buf2), .Y(_1488_) );
NAND2X1 NAND2X1_563 ( .A(REGs_USR_REGS_2__18_), .B(_1573__bF_buf20), .Y(_4879_) );
MUX2X1 MUX2X1_563 ( .A(_1609__bF_buf3), .B(_4879_), .S(_4860__bF_buf4), .Y(_1489_) );
NAND2X1 NAND2X1_564 ( .A(REGs_USR_REGS_2__19_), .B(_1573__bF_buf24), .Y(_4880_) );
MUX2X1 MUX2X1_564 ( .A(_1611__bF_buf0), .B(_4880_), .S(_4860__bF_buf0), .Y(_1490_) );
NAND2X1 NAND2X1_565 ( .A(REGs_USR_REGS_2__20_), .B(_1573__bF_buf22), .Y(_4881_) );
MUX2X1 MUX2X1_565 ( .A(_1613__bF_buf2), .B(_4881_), .S(_4860__bF_buf3), .Y(_1491_) );
NAND2X1 NAND2X1_566 ( .A(REGs_USR_REGS_2__21_), .B(_1573__bF_buf26), .Y(_4882_) );
MUX2X1 MUX2X1_566 ( .A(_1615__bF_buf2), .B(_4882_), .S(_4860__bF_buf4), .Y(_1492_) );
NAND2X1 NAND2X1_567 ( .A(REGs_USR_REGS_2__22_), .B(_1573__bF_buf37), .Y(_4883_) );
MUX2X1 MUX2X1_567 ( .A(_1617__bF_buf1), .B(_4883_), .S(_4860__bF_buf3), .Y(_1493_) );
NAND2X1 NAND2X1_568 ( .A(REGs_USR_REGS_2__23_), .B(_1573__bF_buf26), .Y(_4884_) );
MUX2X1 MUX2X1_568 ( .A(_1619__bF_buf1), .B(_4884_), .S(_4860__bF_buf0), .Y(_1494_) );
NAND2X1 NAND2X1_569 ( .A(REGs_USR_REGS_2__24_), .B(_1573__bF_buf18), .Y(_4885_) );
MUX2X1 MUX2X1_569 ( .A(_1621__bF_buf3), .B(_4885_), .S(_4860__bF_buf1), .Y(_1495_) );
NAND2X1 NAND2X1_570 ( .A(REGs_USR_REGS_2__25_), .B(_1573__bF_buf17), .Y(_4886_) );
MUX2X1 MUX2X1_570 ( .A(_1623__bF_buf1), .B(_4886_), .S(_4860__bF_buf2), .Y(_1496_) );
NAND2X1 NAND2X1_571 ( .A(REGs_USR_REGS_2__26_), .B(_1573__bF_buf69), .Y(_4887_) );
MUX2X1 MUX2X1_571 ( .A(_1625__bF_buf3), .B(_4887_), .S(_4860__bF_buf2), .Y(_1497_) );
NAND2X1 NAND2X1_572 ( .A(REGs_USR_REGS_2__27_), .B(_1573__bF_buf17), .Y(_4888_) );
MUX2X1 MUX2X1_572 ( .A(_1627__bF_buf3), .B(_4888_), .S(_4860__bF_buf2), .Y(_1498_) );
NAND2X1 NAND2X1_573 ( .A(REGs_USR_REGS_2__28_), .B(_1573__bF_buf16), .Y(_4889_) );
MUX2X1 MUX2X1_573 ( .A(_1629__bF_buf1), .B(_4889_), .S(_4860__bF_buf4), .Y(_1499_) );
NAND2X1 NAND2X1_574 ( .A(REGs_USR_REGS_2__29_), .B(_1573__bF_buf39), .Y(_4890_) );
MUX2X1 MUX2X1_574 ( .A(_1631__bF_buf1), .B(_4890_), .S(_4860__bF_buf1), .Y(_1500_) );
NAND2X1 NAND2X1_575 ( .A(REGs_USR_REGS_2__30_), .B(_1573__bF_buf22), .Y(_4891_) );
MUX2X1 MUX2X1_575 ( .A(_1633__bF_buf0), .B(_4891_), .S(_4860__bF_buf3), .Y(_1501_) );
NAND2X1 NAND2X1_576 ( .A(REGs_USR_REGS_2__31_), .B(_1573__bF_buf59), .Y(_4892_) );
MUX2X1 MUX2X1_576 ( .A(_1635__bF_buf3), .B(_4892_), .S(_4860__bF_buf1), .Y(_1502_) );
NOR2X1 NOR2X1_16 ( .A(_4495_), .B(_4324_), .Y(_4893_) );
NAND2X1 NAND2X1_577 ( .A(REGs_REGS_7__0_), .B(_1573__bF_buf42), .Y(_4894_) );
MUX2X1 MUX2X1_577 ( .A(_1567__bF_buf1), .B(_4894_), .S(_4893__bF_buf3), .Y(_1503_) );
NAND2X1 NAND2X1_578 ( .A(REGs_REGS_7__1_), .B(_1573__bF_buf42), .Y(_4895_) );
MUX2X1 MUX2X1_578 ( .A(_1575__bF_buf3), .B(_4895_), .S(_4893__bF_buf3), .Y(_1504_) );
NAND2X1 NAND2X1_579 ( .A(REGs_REGS_7__2_), .B(_1573__bF_buf36), .Y(_4896_) );
MUX2X1 MUX2X1_579 ( .A(_1577__bF_buf1), .B(_4896_), .S(_4893__bF_buf0), .Y(_1505_) );
NAND2X1 NAND2X1_580 ( .A(REGs_REGS_7__3_), .B(_1573__bF_buf19), .Y(_4897_) );
MUX2X1 MUX2X1_580 ( .A(_1579__bF_buf2), .B(_4897_), .S(_4893__bF_buf0), .Y(_1506_) );
NAND2X1 NAND2X1_581 ( .A(REGs_REGS_7__4_), .B(_1573__bF_buf15), .Y(_4898_) );
MUX2X1 MUX2X1_581 ( .A(_1581__bF_buf3), .B(_4898_), .S(_4893__bF_buf2), .Y(_1507_) );
NAND2X1 NAND2X1_582 ( .A(REGs_REGS_7__5_), .B(_1573__bF_buf2), .Y(_4899_) );
MUX2X1 MUX2X1_582 ( .A(_1583__bF_buf3), .B(_4899_), .S(_4893__bF_buf4), .Y(_1508_) );
NAND2X1 NAND2X1_583 ( .A(REGs_REGS_7__6_), .B(_1573__bF_buf15), .Y(_4900_) );
MUX2X1 MUX2X1_583 ( .A(_1585__bF_buf3), .B(_4900_), .S(_4893__bF_buf2), .Y(_1509_) );
NAND2X1 NAND2X1_584 ( .A(REGs_REGS_7__7_), .B(_1573__bF_buf66), .Y(_4901_) );
MUX2X1 MUX2X1_584 ( .A(_1587__bF_buf3), .B(_4901_), .S(_4893__bF_buf2), .Y(_1510_) );
NAND2X1 NAND2X1_585 ( .A(REGs_REGS_7__8_), .B(_1573__bF_buf25), .Y(_4902_) );
MUX2X1 MUX2X1_585 ( .A(_1589__bF_buf3), .B(_4902_), .S(_4893__bF_buf1), .Y(_1511_) );
NAND2X1 NAND2X1_586 ( .A(REGs_REGS_7__9_), .B(_1573__bF_buf29), .Y(_4903_) );
MUX2X1 MUX2X1_586 ( .A(_1591__bF_buf2), .B(_4903_), .S(_4893__bF_buf1), .Y(_1512_) );
NAND2X1 NAND2X1_587 ( .A(REGs_REGS_7__10_), .B(_1573__bF_buf9), .Y(_4904_) );
MUX2X1 MUX2X1_587 ( .A(_1593__bF_buf3), .B(_4904_), .S(_4893__bF_buf1), .Y(_1513_) );
NAND2X1 NAND2X1_588 ( .A(REGs_REGS_7__11_), .B(_1573__bF_buf73), .Y(_4905_) );
MUX2X1 MUX2X1_588 ( .A(_1595__bF_buf2), .B(_4905_), .S(_4893__bF_buf4), .Y(_1514_) );
NAND2X1 NAND2X1_589 ( .A(REGs_REGS_7__12_), .B(_1573__bF_buf66), .Y(_4906_) );
MUX2X1 MUX2X1_589 ( .A(_1597__bF_buf0), .B(_4906_), .S(_4893__bF_buf2), .Y(_1515_) );
NAND2X1 NAND2X1_590 ( .A(REGs_REGS_7__13_), .B(_1573__bF_buf36), .Y(_4907_) );
MUX2X1 MUX2X1_590 ( .A(_1599__bF_buf2), .B(_4907_), .S(_4893__bF_buf3), .Y(_1516_) );
NAND2X1 NAND2X1_591 ( .A(REGs_REGS_7__14_), .B(_1573__bF_buf62), .Y(_4908_) );
MUX2X1 MUX2X1_591 ( .A(_1601__bF_buf3), .B(_4908_), .S(_4893__bF_buf1), .Y(_1517_) );
NAND2X1 NAND2X1_592 ( .A(REGs_REGS_7__15_), .B(_1573__bF_buf62), .Y(_4909_) );
MUX2X1 MUX2X1_592 ( .A(_1603__bF_buf2), .B(_4909_), .S(_4893__bF_buf1), .Y(_1518_) );
NAND2X1 NAND2X1_593 ( .A(REGs_REGS_7__16_), .B(_1573__bF_buf41), .Y(_4910_) );
MUX2X1 MUX2X1_593 ( .A(_1605__bF_buf2), .B(_4910_), .S(_4893__bF_buf4), .Y(_1519_) );
NAND2X1 NAND2X1_594 ( .A(REGs_REGS_7__17_), .B(_1573__bF_buf36), .Y(_4911_) );
MUX2X1 MUX2X1_594 ( .A(_1607__bF_buf3), .B(_4911_), .S(_4893__bF_buf3), .Y(_1520_) );
NAND2X1 NAND2X1_595 ( .A(REGs_REGS_7__18_), .B(_1573__bF_buf73), .Y(_4912_) );
MUX2X1 MUX2X1_595 ( .A(_1609__bF_buf1), .B(_4912_), .S(_4893__bF_buf4), .Y(_1521_) );
NAND2X1 NAND2X1_596 ( .A(REGs_REGS_7__19_), .B(_1573__bF_buf49), .Y(_4913_) );
MUX2X1 MUX2X1_596 ( .A(_1611__bF_buf3), .B(_4913_), .S(_4893__bF_buf4), .Y(_1522_) );
NAND2X1 NAND2X1_597 ( .A(REGs_REGS_7__20_), .B(_1573__bF_buf15), .Y(_4914_) );
MUX2X1 MUX2X1_597 ( .A(_1613__bF_buf2), .B(_4914_), .S(_4893__bF_buf0), .Y(_1523_) );
NAND2X1 NAND2X1_598 ( .A(REGs_REGS_7__21_), .B(_1573__bF_buf2), .Y(_4915_) );
MUX2X1 MUX2X1_598 ( .A(_1615__bF_buf1), .B(_4915_), .S(_4893__bF_buf4), .Y(_1524_) );
NAND2X1 NAND2X1_599 ( .A(REGs_REGS_7__22_), .B(_1573__bF_buf67), .Y(_4916_) );
MUX2X1 MUX2X1_599 ( .A(_1617__bF_buf0), .B(_4916_), .S(_4893__bF_buf2), .Y(_1525_) );
NAND2X1 NAND2X1_600 ( .A(REGs_REGS_7__23_), .B(_1573__bF_buf9), .Y(_4917_) );
MUX2X1 MUX2X1_600 ( .A(_1619__bF_buf2), .B(_4917_), .S(_4893__bF_buf1), .Y(_1526_) );
NAND2X1 NAND2X1_601 ( .A(REGs_REGS_7__24_), .B(_1573__bF_buf33), .Y(_4918_) );
MUX2X1 MUX2X1_601 ( .A(_1621__bF_buf2), .B(_4918_), .S(_4893__bF_buf3), .Y(_1527_) );
NAND2X1 NAND2X1_602 ( .A(REGs_REGS_7__25_), .B(_1573__bF_buf47), .Y(_4919_) );
MUX2X1 MUX2X1_602 ( .A(_1623__bF_buf2), .B(_4919_), .S(_4893__bF_buf0), .Y(_1528_) );
NAND2X1 NAND2X1_603 ( .A(REGs_REGS_7__26_), .B(_1573__bF_buf46), .Y(_4920_) );
MUX2X1 MUX2X1_603 ( .A(_1625__bF_buf1), .B(_4920_), .S(_4893__bF_buf2), .Y(_1529_) );
NAND2X1 NAND2X1_604 ( .A(REGs_REGS_7__27_), .B(_1573__bF_buf19), .Y(_4921_) );
MUX2X1 MUX2X1_604 ( .A(_1627__bF_buf0), .B(_4921_), .S(_4893__bF_buf0), .Y(_1530_) );
NAND2X1 NAND2X1_605 ( .A(REGs_REGS_7__28_), .B(_1573__bF_buf73), .Y(_4922_) );
MUX2X1 MUX2X1_605 ( .A(_1629__bF_buf3), .B(_4922_), .S(_4893__bF_buf4), .Y(_1531_) );
NAND2X1 NAND2X1_606 ( .A(REGs_REGS_7__29_), .B(_1573__bF_buf42), .Y(_4923_) );
MUX2X1 MUX2X1_606 ( .A(_1631__bF_buf2), .B(_4923_), .S(_4893__bF_buf3), .Y(_1532_) );
NAND2X1 NAND2X1_607 ( .A(REGs_REGS_7__30_), .B(_1573__bF_buf36), .Y(_4924_) );
MUX2X1 MUX2X1_607 ( .A(_1633__bF_buf1), .B(_4924_), .S(_4893__bF_buf0), .Y(_1533_) );
NAND2X1 NAND2X1_608 ( .A(REGs_REGS_7__31_), .B(_1573__bF_buf2), .Y(_4925_) );
MUX2X1 MUX2X1_608 ( .A(_1635__bF_buf0), .B(_4925_), .S(_4893__bF_buf3), .Y(_1534_) );
NOR2X1 NOR2X1_17 ( .A(_4290_), .B(_4495_), .Y(_4926_) );
NAND2X1 NAND2X1_609 ( .A(REGs_REGS_5__0_), .B(_1573__bF_buf42), .Y(_4927_) );
MUX2X1 MUX2X1_609 ( .A(_1567__bF_buf1), .B(_4927_), .S(_4926__bF_buf3), .Y(_1535_) );
NAND2X1 NAND2X1_610 ( .A(REGs_REGS_5__1_), .B(_1573__bF_buf42), .Y(_4928_) );
MUX2X1 MUX2X1_610 ( .A(_1575__bF_buf3), .B(_4928_), .S(_4926__bF_buf3), .Y(_1536_) );
NAND2X1 NAND2X1_611 ( .A(REGs_REGS_5__2_), .B(_1573__bF_buf34), .Y(_4929_) );
MUX2X1 MUX2X1_611 ( .A(_1577__bF_buf1), .B(_4929_), .S(_4926__bF_buf1), .Y(_1537_) );
NAND2X1 NAND2X1_612 ( .A(REGs_REGS_5__3_), .B(_1573__bF_buf47), .Y(_4930_) );
MUX2X1 MUX2X1_612 ( .A(_1579__bF_buf2), .B(_4930_), .S(_4926__bF_buf1), .Y(_1538_) );
NAND2X1 NAND2X1_613 ( .A(REGs_REGS_5__4_), .B(_1573__bF_buf67), .Y(_4931_) );
MUX2X1 MUX2X1_613 ( .A(_1581__bF_buf1), .B(_4931_), .S(_4926__bF_buf0), .Y(_1539_) );
NAND2X1 NAND2X1_614 ( .A(REGs_REGS_5__5_), .B(_1573__bF_buf73), .Y(_4932_) );
MUX2X1 MUX2X1_614 ( .A(_1583__bF_buf3), .B(_4932_), .S(_4926__bF_buf3), .Y(_1540_) );
NAND2X1 NAND2X1_615 ( .A(REGs_REGS_5__6_), .B(_1573__bF_buf67), .Y(_4933_) );
MUX2X1 MUX2X1_615 ( .A(_1585__bF_buf3), .B(_4933_), .S(_4926__bF_buf0), .Y(_1541_) );
NAND2X1 NAND2X1_616 ( .A(REGs_REGS_5__7_), .B(_1573__bF_buf67), .Y(_4934_) );
MUX2X1 MUX2X1_616 ( .A(_1587__bF_buf3), .B(_4934_), .S(_4926__bF_buf0), .Y(_1542_) );
NAND2X1 NAND2X1_617 ( .A(REGs_REGS_5__8_), .B(_1573__bF_buf25), .Y(_4935_) );
MUX2X1 MUX2X1_617 ( .A(_1589__bF_buf3), .B(_4935_), .S(_4926__bF_buf4), .Y(_1543_) );
NAND2X1 NAND2X1_618 ( .A(REGs_REGS_5__9_), .B(_1573__bF_buf29), .Y(_4936_) );
MUX2X1 MUX2X1_618 ( .A(_1591__bF_buf2), .B(_4936_), .S(_4926__bF_buf4), .Y(_1544_) );
NAND2X1 NAND2X1_619 ( .A(REGs_REGS_5__10_), .B(_1573__bF_buf62), .Y(_4937_) );
MUX2X1 MUX2X1_619 ( .A(_1593__bF_buf0), .B(_4937_), .S(_4926__bF_buf4), .Y(_1545_) );
NAND2X1 NAND2X1_620 ( .A(REGs_REGS_5__11_), .B(_1573__bF_buf29), .Y(_4938_) );
MUX2X1 MUX2X1_620 ( .A(_1595__bF_buf2), .B(_4938_), .S(_4926__bF_buf3), .Y(_1546_) );
NAND2X1 NAND2X1_621 ( .A(REGs_REGS_5__12_), .B(_1573__bF_buf66), .Y(_4939_) );
MUX2X1 MUX2X1_621 ( .A(_1597__bF_buf0), .B(_4939_), .S(_4926__bF_buf0), .Y(_1547_) );
NAND2X1 NAND2X1_622 ( .A(REGs_REGS_5__13_), .B(_1573__bF_buf33), .Y(_4940_) );
MUX2X1 MUX2X1_622 ( .A(_1599__bF_buf2), .B(_4940_), .S(_4926__bF_buf2), .Y(_1548_) );
NAND2X1 NAND2X1_623 ( .A(REGs_REGS_5__14_), .B(_1573__bF_buf9), .Y(_4941_) );
MUX2X1 MUX2X1_623 ( .A(_1601__bF_buf3), .B(_4941_), .S(_4926__bF_buf4), .Y(_1549_) );
NAND2X1 NAND2X1_624 ( .A(REGs_REGS_5__15_), .B(_1573__bF_buf64), .Y(_4942_) );
MUX2X1 MUX2X1_624 ( .A(_1603__bF_buf2), .B(_4942_), .S(_4926__bF_buf4), .Y(_1550_) );
NAND2X1 NAND2X1_625 ( .A(REGs_REGS_5__16_), .B(_1573__bF_buf62), .Y(_4943_) );
MUX2X1 MUX2X1_625 ( .A(_1605__bF_buf2), .B(_4943_), .S(_4926__bF_buf4), .Y(_1551_) );
NAND2X1 NAND2X1_626 ( .A(REGs_REGS_5__17_), .B(_1573__bF_buf33), .Y(_4944_) );
MUX2X1 MUX2X1_626 ( .A(_1607__bF_buf0), .B(_4944_), .S(_4926__bF_buf2), .Y(_1552_) );
NAND2X1 NAND2X1_627 ( .A(REGs_REGS_5__18_), .B(_1573__bF_buf49), .Y(_4945_) );
MUX2X1 MUX2X1_627 ( .A(_1609__bF_buf1), .B(_4945_), .S(_4926__bF_buf2), .Y(_1553_) );
NAND2X1 NAND2X1_628 ( .A(REGs_REGS_5__19_), .B(_1573__bF_buf42), .Y(_4946_) );
MUX2X1 MUX2X1_628 ( .A(_1611__bF_buf3), .B(_4946_), .S(_4926__bF_buf2), .Y(_1554_) );
NAND2X1 NAND2X1_629 ( .A(REGs_REGS_5__20_), .B(_1573__bF_buf34), .Y(_4947_) );
MUX2X1 MUX2X1_629 ( .A(_1613__bF_buf1), .B(_4947_), .S(_4926__bF_buf1), .Y(_1555_) );
NAND2X1 NAND2X1_630 ( .A(REGs_REGS_5__21_), .B(_1573__bF_buf29), .Y(_4948_) );
MUX2X1 MUX2X1_630 ( .A(_1615__bF_buf1), .B(_4948_), .S(_4926__bF_buf3), .Y(_1556_) );
NAND2X1 NAND2X1_631 ( .A(REGs_REGS_5__22_), .B(_1573__bF_buf67), .Y(_4949_) );
MUX2X1 MUX2X1_631 ( .A(_1617__bF_buf0), .B(_4949_), .S(_4926__bF_buf0), .Y(_1557_) );
NAND2X1 NAND2X1_632 ( .A(REGs_REGS_5__23_), .B(_1573__bF_buf64), .Y(_4950_) );
MUX2X1 MUX2X1_632 ( .A(_1619__bF_buf2), .B(_4950_), .S(_4926__bF_buf4), .Y(_1558_) );
NAND2X1 NAND2X1_633 ( .A(REGs_REGS_5__24_), .B(_1573__bF_buf33), .Y(_4951_) );
MUX2X1 MUX2X1_633 ( .A(_1621__bF_buf2), .B(_4951_), .S(_4926__bF_buf2), .Y(_1559_) );
NAND2X1 NAND2X1_634 ( .A(REGs_REGS_5__25_), .B(_1573__bF_buf47), .Y(_4952_) );
MUX2X1 MUX2X1_634 ( .A(_1623__bF_buf2), .B(_4952_), .S(_4926__bF_buf1), .Y(_1560_) );
NAND2X1 NAND2X1_635 ( .A(REGs_REGS_5__26_), .B(_1573__bF_buf15), .Y(_4953_) );
MUX2X1 MUX2X1_635 ( .A(_1625__bF_buf1), .B(_4953_), .S(_4926__bF_buf0), .Y(_1561_) );
NAND2X1 NAND2X1_636 ( .A(REGs_REGS_5__27_), .B(_1573__bF_buf47), .Y(_4954_) );
MUX2X1 MUX2X1_636 ( .A(_1627__bF_buf1), .B(_4954_), .S(_4926__bF_buf1), .Y(_1562_) );
NAND2X1 NAND2X1_637 ( .A(REGs_REGS_5__28_), .B(_1573__bF_buf29), .Y(_4955_) );
MUX2X1 MUX2X1_637 ( .A(_1629__bF_buf3), .B(_4955_), .S(_4926__bF_buf3), .Y(_1563_) );
NAND2X1 NAND2X1_638 ( .A(REGs_REGS_5__29_), .B(_1573__bF_buf2), .Y(_4956_) );
MUX2X1 MUX2X1_638 ( .A(_1631__bF_buf2), .B(_4956_), .S(_4926__bF_buf3), .Y(_1564_) );
NAND2X1 NAND2X1_639 ( .A(REGs_REGS_5__30_), .B(_1573__bF_buf34), .Y(_4957_) );
MUX2X1 MUX2X1_639 ( .A(_1633__bF_buf1), .B(_4957_), .S(_4926__bF_buf1), .Y(_1565_) );
NAND2X1 NAND2X1_640 ( .A(REGs_REGS_5__31_), .B(_1573__bF_buf75), .Y(_4958_) );
MUX2X1 MUX2X1_640 ( .A(_1635__bF_buf1), .B(_4958_), .S(_4926__bF_buf2), .Y(_1566_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf50), .D(_1023_), .Q(REGs_FIRQ_REGS_3__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf9), .D(_1024_), .Q(REGs_FIRQ_REGS_3__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf56), .D(_1025_), .Q(REGs_FIRQ_REGS_3__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf58), .D(_1026_), .Q(REGs_FIRQ_REGS_3__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf49), .D(_1027_), .Q(REGs_FIRQ_REGS_3__4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf76), .D(_1028_), .Q(REGs_FIRQ_REGS_3__5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf45), .D(_1029_), .Q(REGs_FIRQ_REGS_3__6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf30), .D(_1030_), .Q(REGs_FIRQ_REGS_3__7_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf9), .D(_1031_), .Q(REGs_FIRQ_REGS_3__8_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf62), .D(_1032_), .Q(REGs_FIRQ_REGS_3__9_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf26), .D(_1033_), .Q(REGs_FIRQ_REGS_3__10_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf54), .D(_1034_), .Q(REGs_FIRQ_REGS_3__11_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf38), .D(_1035_), .Q(REGs_FIRQ_REGS_3__12_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf30), .D(_1036_), .Q(REGs_FIRQ_REGS_3__13_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf59), .D(_1037_), .Q(REGs_FIRQ_REGS_3__14_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf10), .D(_1038_), .Q(REGs_FIRQ_REGS_3__15_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf62), .D(_1039_), .Q(REGs_FIRQ_REGS_3__16_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf30), .D(_1040_), .Q(REGs_FIRQ_REGS_3__17_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf59), .D(_1041_), .Q(REGs_FIRQ_REGS_3__18_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf70), .D(_1042_), .Q(REGs_FIRQ_REGS_3__19_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf31), .D(_1043_), .Q(REGs_FIRQ_REGS_3__20_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf76), .D(_1044_), .Q(REGs_FIRQ_REGS_3__21_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf45), .D(_1045_), .Q(REGs_FIRQ_REGS_3__22_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf66), .D(_1046_), .Q(REGs_FIRQ_REGS_3__23_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf12), .D(_1047_), .Q(REGs_FIRQ_REGS_3__24_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf30), .D(_1048_), .Q(REGs_FIRQ_REGS_3__25_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf29), .D(_1049_), .Q(REGs_FIRQ_REGS_3__26_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf30), .D(_1050_), .Q(REGs_FIRQ_REGS_3__27_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf10), .D(_1051_), .Q(REGs_FIRQ_REGS_3__28_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf58), .D(_1052_), .Q(REGs_FIRQ_REGS_3__29_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf56), .D(_1053_), .Q(REGs_FIRQ_REGS_3__30_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf4), .D(_1054_), .Q(REGs_FIRQ_REGS_3__31_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf70), .D(_1343_), .Q(REGs_FIRQ_REGS_6__0_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf47), .D(_1344_), .Q(REGs_FIRQ_REGS_6__1_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf7), .D(_1345_), .Q(REGs_FIRQ_REGS_6__2_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf7), .D(_1346_), .Q(REGs_FIRQ_REGS_6__3_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf86), .D(_1347_), .Q(REGs_FIRQ_REGS_6__4_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf78), .D(_1348_), .Q(REGs_FIRQ_REGS_6__5_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf49), .D(_1349_), .Q(REGs_FIRQ_REGS_6__6_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf18), .D(_1350_), .Q(REGs_FIRQ_REGS_6__7_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf15), .D(_1351_), .Q(REGs_FIRQ_REGS_6__8_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf78), .D(_1352_), .Q(REGs_FIRQ_REGS_6__9_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf0), .D(_1353_), .Q(REGs_FIRQ_REGS_6__10_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf20), .D(_1354_), .Q(REGs_FIRQ_REGS_6__11_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf50), .D(_1355_), .Q(REGs_FIRQ_REGS_6__12_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf79), .D(_1356_), .Q(REGs_FIRQ_REGS_6__13_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf0), .D(_1357_), .Q(REGs_FIRQ_REGS_6__14_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf20), .D(_1358_), .Q(REGs_FIRQ_REGS_6__15_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf78), .D(_1359_), .Q(REGs_FIRQ_REGS_6__16_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf7), .D(_1360_), .Q(REGs_FIRQ_REGS_6__17_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf32), .D(_1361_), .Q(REGs_FIRQ_REGS_6__18_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf52), .D(_1362_), .Q(REGs_FIRQ_REGS_6__19_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf2), .D(_1363_), .Q(REGs_FIRQ_REGS_6__20_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf35), .D(_1364_), .Q(REGs_FIRQ_REGS_6__21_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf88), .D(_1365_), .Q(REGs_FIRQ_REGS_6__22_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf35), .D(_1366_), .Q(REGs_FIRQ_REGS_6__23_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf11), .D(_1367_), .Q(REGs_FIRQ_REGS_6__24_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf13), .D(_1368_), .Q(REGs_FIRQ_REGS_6__25_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf18), .D(_1369_), .Q(REGs_FIRQ_REGS_6__26_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf18), .D(_1370_), .Q(REGs_FIRQ_REGS_6__27_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf78), .D(_1371_), .Q(REGs_FIRQ_REGS_6__28_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf79), .D(_1372_), .Q(REGs_FIRQ_REGS_6__29_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf50), .D(_1373_), .Q(REGs_FIRQ_REGS_6__30_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf82), .D(_1374_), .Q(REGs_FIRQ_REGS_6__31_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf50), .D(_1055_), .Q(REGs_FIRQ_REGS_1__0_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf76), .D(_1056_), .Q(REGs_FIRQ_REGS_1__1_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf24), .D(_1057_), .Q(REGs_FIRQ_REGS_1__2_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf18), .D(_1058_), .Q(REGs_FIRQ_REGS_1__3_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf88), .D(_1059_), .Q(REGs_FIRQ_REGS_1__4_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf66), .D(_1060_), .Q(REGs_FIRQ_REGS_1__5_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf49), .D(_1061_), .Q(REGs_FIRQ_REGS_1__6_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf80), .D(_1062_), .Q(REGs_FIRQ_REGS_1__7_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf34), .D(_1063_), .Q(REGs_FIRQ_REGS_1__8_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf42), .D(_1064_), .Q(REGs_FIRQ_REGS_1__9_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf26), .D(_1065_), .Q(REGs_FIRQ_REGS_1__10_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf54), .D(_1066_), .Q(REGs_FIRQ_REGS_1__11_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf49), .D(_1067_), .Q(REGs_FIRQ_REGS_1__12_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf80), .D(_1068_), .Q(REGs_FIRQ_REGS_1__13_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf42), .D(_1069_), .Q(REGs_FIRQ_REGS_1__14_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf62), .D(_1070_), .Q(REGs_FIRQ_REGS_1__15_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf15), .D(_1071_), .Q(REGs_FIRQ_REGS_1__16_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf13), .D(_1072_), .Q(REGs_FIRQ_REGS_1__17_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf42), .D(_1073_), .Q(REGs_FIRQ_REGS_1__18_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf70), .D(_1074_), .Q(REGs_FIRQ_REGS_1__19_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf50), .D(_1075_), .Q(REGs_FIRQ_REGS_1__20_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf54), .D(_1076_), .Q(REGs_FIRQ_REGS_1__21_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf49), .D(_1077_), .Q(REGs_FIRQ_REGS_1__22_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf41), .D(_1078_), .Q(REGs_FIRQ_REGS_1__23_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf79), .D(_1079_), .Q(REGs_FIRQ_REGS_1__24_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf80), .D(_1080_), .Q(REGs_FIRQ_REGS_1__25_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf49), .D(_1081_), .Q(REGs_FIRQ_REGS_1__26_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf80), .D(_1082_), .Q(REGs_FIRQ_REGS_1__27_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf54), .D(_1083_), .Q(REGs_FIRQ_REGS_1__28_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf34), .D(_1084_), .Q(REGs_FIRQ_REGS_1__29_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf50), .D(_1085_), .Q(REGs_FIRQ_REGS_1__30_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf2), .D(_1086_), .Q(REGs_FIRQ_REGS_1__31_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf58), .D(_991_), .Q(REGs_FIRQ_REGS_2__0_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf66), .D(_992_), .Q(REGs_FIRQ_REGS_2__1_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf56), .D(_993_), .Q(REGs_FIRQ_REGS_2__2_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf58), .D(_994_), .Q(REGs_FIRQ_REGS_2__3_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf45), .D(_995_), .Q(REGs_FIRQ_REGS_2__4_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf4), .D(_996_), .Q(REGs_FIRQ_REGS_2__5_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf23), .D(_997_), .Q(REGs_FIRQ_REGS_2__6_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf1), .D(_998_), .Q(REGs_FIRQ_REGS_2__7_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf70), .D(_999_), .Q(REGs_FIRQ_REGS_2__8_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf41), .D(_1000_), .Q(REGs_FIRQ_REGS_2__9_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf25), .D(_1001_), .Q(REGs_FIRQ_REGS_2__10_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf44), .D(_1002_), .Q(REGs_FIRQ_REGS_2__11_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf23), .D(_1003_), .Q(REGs_FIRQ_REGS_2__12_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf1), .D(_1004_), .Q(REGs_FIRQ_REGS_2__13_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf32), .D(_1005_), .Q(REGs_FIRQ_REGS_2__14_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf59), .D(_1006_), .Q(REGs_FIRQ_REGS_2__15_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf15), .D(_1007_), .Q(REGs_FIRQ_REGS_2__16_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf1), .D(_1008_), .Q(REGs_FIRQ_REGS_2__17_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf42), .D(_1009_), .Q(REGs_FIRQ_REGS_2__18_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf70), .D(_1010_), .Q(REGs_FIRQ_REGS_2__19_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf80), .D(_1011_), .Q(REGs_FIRQ_REGS_2__20_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf66), .D(_1012_), .Q(REGs_FIRQ_REGS_2__21_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf23), .D(_1013_), .Q(REGs_FIRQ_REGS_2__22_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf66), .D(_1014_), .Q(REGs_FIRQ_REGS_2__23_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf31), .D(_1015_), .Q(REGs_FIRQ_REGS_2__24_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf1), .D(_1016_), .Q(REGs_FIRQ_REGS_2__25_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf23), .D(_1017_), .Q(REGs_FIRQ_REGS_2__26_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf29), .D(_1018_), .Q(REGs_FIRQ_REGS_2__27_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf9), .D(_1019_), .Q(REGs_FIRQ_REGS_2__28_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf82), .D(_1020_), .Q(REGs_FIRQ_REGS_2__29_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf2), .D(_1021_), .Q(REGs_FIRQ_REGS_2__30_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf58), .D(_1022_), .Q(REGs_FIRQ_REGS_2__31_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf60), .D(_1183_), .Q(REGs_REGS_3__0_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf64), .D(_1184_), .Q(REGs_REGS_3__1_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf63), .D(_1185_), .Q(REGs_REGS_3__2_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf61), .D(_1186_), .Q(REGs_REGS_3__3_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf48), .D(_1187_), .Q(REGs_REGS_3__4_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf64), .D(_1188_), .Q(REGs_REGS_3__5_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf48), .D(_1189_), .Q(REGs_REGS_3__6_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf57), .D(_1190_), .Q(REGs_REGS_3__7_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf81), .D(_1191_), .Q(REGs_REGS_3__8_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf77), .D(_1192_), .Q(REGs_REGS_3__9_) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf51), .D(_1193_), .Q(REGs_REGS_3__10_) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf64), .D(_1194_), .Q(REGs_REGS_3__11_) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf48), .D(_1195_), .Q(REGs_REGS_3__12_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf60), .D(_1196_), .Q(REGs_REGS_3__13_) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf77), .D(_1197_), .Q(REGs_REGS_3__14_) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf19), .D(_1198_), .Q(REGs_REGS_3__15_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf51), .D(_1199_), .Q(REGs_REGS_3__16_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf63), .D(_1200_), .Q(REGs_REGS_3__17_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf51), .D(_1201_), .Q(REGs_REGS_3__18_) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf64), .D(_1202_), .Q(REGs_REGS_3__19_) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf43), .D(_1203_), .Q(REGs_REGS_3__20_) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf87), .D(_1204_), .Q(REGs_REGS_3__21_) );
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf48), .D(_1205_), .Q(REGs_REGS_3__22_) );
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf77), .D(_1206_), .Q(REGs_REGS_3__23_) );
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf60), .D(_1207_), .Q(REGs_REGS_3__24_) );
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf63), .D(_1208_), .Q(REGs_REGS_3__25_) );
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf48), .D(_1209_), .Q(REGs_REGS_3__26_) );
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf43), .D(_1210_), .Q(REGs_REGS_3__27_) );
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf81), .D(_1211_), .Q(REGs_REGS_3__28_) );
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf63), .D(_1212_), .Q(REGs_REGS_3__29_) );
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf43), .D(_1213_), .Q(REGs_REGS_3__30_) );
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf64), .D(_1214_), .Q(REGs_REGS_3__31_) );
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf39), .D(_1151_), .Q(REGs_REGS_4__0_) );
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf46), .D(_1152_), .Q(REGs_REGS_4__1_) );
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf39), .D(_1153_), .Q(REGs_REGS_4__2_) );
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf16), .D(_1154_), .Q(REGs_REGS_4__3_) );
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf22), .D(_1155_), .Q(REGs_REGS_4__4_) );
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf55), .D(_1156_), .Q(REGs_REGS_4__5_) );
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf68), .D(_1157_), .Q(REGs_REGS_4__6_) );
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf68), .D(_1158_), .Q(REGs_REGS_4__7_) );
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf55), .D(_1159_), .Q(REGs_REGS_4__8_) );
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf85), .D(_1160_), .Q(REGs_REGS_4__9_) );
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf69), .D(_1161_), .Q(REGs_REGS_4__10_) );
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf87), .D(_1162_), .Q(REGs_REGS_4__11_) );
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf22), .D(_1163_), .Q(REGs_REGS_4__12_) );
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf63), .D(_1164_), .Q(REGs_REGS_4__13_) );
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf6), .D(_1165_), .Q(REGs_REGS_4__14_) );
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf85), .D(_1166_), .Q(REGs_REGS_4__15_) );
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf87), .D(_1167_), .Q(REGs_REGS_4__16_) );
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf27), .D(_1168_), .Q(REGs_REGS_4__17_) );
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf69), .D(_1169_), .Q(REGs_REGS_4__18_) );
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf27), .D(_1170_), .Q(REGs_REGS_4__19_) );
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf33), .D(_1171_), .Q(REGs_REGS_4__20_) );
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf55), .D(_1172_), .Q(REGs_REGS_4__21_) );
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf57), .D(_1173_), .Q(REGs_REGS_4__22_) );
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf85), .D(_1174_), .Q(REGs_REGS_4__23_) );
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf27), .D(_1175_), .Q(REGs_REGS_4__24_) );
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf63), .D(_1176_), .Q(REGs_REGS_4__25_) );
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf84), .D(_1177_), .Q(REGs_REGS_4__26_) );
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf16), .D(_1178_), .Q(REGs_REGS_4__27_) );
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf55), .D(_1179_), .Q(REGs_REGS_4__28_) );
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf39), .D(_1180_), .Q(REGs_REGS_4__29_) );
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf71), .D(_1181_), .Q(REGs_REGS_4__30_) );
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf27), .D(_1182_), .Q(REGs_REGS_4__31_) );
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf39), .D(_1535_), .Q(REGs_REGS_5__0_) );
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf46), .D(_1536_), .Q(REGs_REGS_5__1_) );
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf39), .D(_1537_), .Q(REGs_REGS_5__2_) );
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf33), .D(_1538_), .Q(REGs_REGS_5__3_) );
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf68), .D(_1539_), .Q(REGs_REGS_5__4_) );
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf55), .D(_1540_), .Q(REGs_REGS_5__5_) );
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf68), .D(_1541_), .Q(REGs_REGS_5__6_) );
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf36), .D(_1542_), .Q(REGs_REGS_5__7_) );
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf85), .D(_1543_), .Q(REGs_REGS_5__8_) );
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf85), .D(_1544_), .Q(REGs_REGS_5__9_) );
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf6), .D(_1545_), .Q(REGs_REGS_5__10_) );
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf69), .D(_1546_), .Q(REGs_REGS_5__11_) );
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf68), .D(_1547_), .Q(REGs_REGS_5__12_) );
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf27), .D(_1548_), .Q(REGs_REGS_5__13_) );
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf0), .D(_1549_), .Q(REGs_REGS_5__14_) );
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf35), .D(_1550_), .Q(REGs_REGS_5__15_) );
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf69), .D(_1551_), .Q(REGs_REGS_5__16_) );
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf63), .D(_1552_), .Q(REGs_REGS_5__17_) );
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf64), .D(_1553_), .Q(REGs_REGS_5__18_) );
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf46), .D(_1554_), .Q(REGs_REGS_5__19_) );
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf71), .D(_1555_), .Q(REGs_REGS_5__20_) );
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf55), .D(_1556_), .Q(REGs_REGS_5__21_) );
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf57), .D(_1557_), .Q(REGs_REGS_5__22_) );
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf35), .D(_1558_), .Q(REGs_REGS_5__23_) );
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf27), .D(_1559_), .Q(REGs_REGS_5__24_) );
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf33), .D(_1560_), .Q(REGs_REGS_5__25_) );
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf37), .D(_1561_), .Q(REGs_REGS_5__26_) );
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf33), .D(_1562_), .Q(REGs_REGS_5__27_) );
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf55), .D(_1563_), .Q(REGs_REGS_5__28_) );
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf46), .D(_1564_), .Q(REGs_REGS_5__29_) );
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf39), .D(_1565_), .Q(REGs_REGS_5__30_) );
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf27), .D(_1566_), .Q(REGs_REGS_5__31_) );
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf82), .D(_1119_), .Q(REGs_REGS_6__0_) );
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf46), .D(_1120_), .Q(REGs_REGS_6__1_) );
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf16), .D(_1121_), .Q(REGs_REGS_6__2_) );
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf16), .D(_1122_), .Q(REGs_REGS_6__3_) );
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf68), .D(_1123_), .Q(REGs_REGS_6__4_) );
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf55), .D(_1124_), .Q(REGs_REGS_6__5_) );
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf37), .D(_1125_), .Q(REGs_REGS_6__6_) );
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf68), .D(_1126_), .Q(REGs_REGS_6__7_) );
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf41), .D(_1127_), .Q(REGs_REGS_6__8_) );
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf85), .D(_1128_), .Q(REGs_REGS_6__9_) );
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf53), .D(_1129_), .Q(REGs_REGS_6__10_) );
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf55), .D(_1130_), .Q(REGs_REGS_6__11_) );
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf22), .D(_1131_), .Q(REGs_REGS_6__12_) );
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf16), .D(_1132_), .Q(REGs_REGS_6__13_) );
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf6), .D(_1133_), .Q(REGs_REGS_6__14_) );
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf69), .D(_1134_), .Q(REGs_REGS_6__15_) );
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf69), .D(_1135_), .Q(REGs_REGS_6__16_) );
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf16), .D(_1136_), .Q(REGs_REGS_6__17_) );
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf81), .D(_1137_), .Q(REGs_REGS_6__18_) );
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf46), .D(_1138_), .Q(REGs_REGS_6__19_) );
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf37), .D(_1139_), .Q(REGs_REGS_6__20_) );
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf4), .D(_1140_), .Q(REGs_REGS_6__21_) );
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf68), .D(_1141_), .Q(REGs_REGS_6__22_) );
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf0), .D(_1142_), .Q(REGs_REGS_6__23_) );
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf27), .D(_1143_), .Q(REGs_REGS_6__24_) );
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf48), .D(_1144_), .Q(REGs_REGS_6__25_) );
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf37), .D(_1145_), .Q(REGs_REGS_6__26_) );
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf43), .D(_1146_), .Q(REGs_REGS_6__27_) );
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf46), .D(_1147_), .Q(REGs_REGS_6__28_) );
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf16), .D(_1148_), .Q(REGs_REGS_6__29_) );
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf33), .D(_1149_), .Q(REGs_REGS_6__30_) );
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf81), .D(_1150_), .Q(REGs_REGS_6__31_) );
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf39), .D(_1503_), .Q(REGs_REGS_7__0_) );
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf46), .D(_1504_), .Q(REGs_REGS_7__1_) );
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf39), .D(_1505_), .Q(REGs_REGS_7__2_) );
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf33), .D(_1506_), .Q(REGs_REGS_7__3_) );
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf84), .D(_1507_), .Q(REGs_REGS_7__4_) );
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf55), .D(_1508_), .Q(REGs_REGS_7__5_) );
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf68), .D(_1509_), .Q(REGs_REGS_7__6_) );
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf68), .D(_1510_), .Q(REGs_REGS_7__7_) );
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf85), .D(_1511_), .Q(REGs_REGS_7__8_) );
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf69), .D(_1512_), .Q(REGs_REGS_7__9_) );
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf6), .D(_1513_), .Q(REGs_REGS_7__10_) );
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf81), .D(_1514_), .Q(REGs_REGS_7__11_) );
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf84), .D(_1515_), .Q(REGs_REGS_7__12_) );
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf63), .D(_1516_), .Q(REGs_REGS_7__13_) );
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf6), .D(_1517_), .Q(REGs_REGS_7__14_) );
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf69), .D(_1518_), .Q(REGs_REGS_7__15_) );
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf87), .D(_1519_), .Q(REGs_REGS_7__16_) );
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf16), .D(_1520_), .Q(REGs_REGS_7__17_) );
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf81), .D(_1521_), .Q(REGs_REGS_7__18_) );
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf81), .D(_1522_), .Q(REGs_REGS_7__19_) );
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf37), .D(_1523_), .Q(REGs_REGS_7__20_) );
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf4), .D(_1524_), .Q(REGs_REGS_7__21_) );
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf57), .D(_1525_), .Q(REGs_REGS_7__22_) );
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf0), .D(_1526_), .Q(REGs_REGS_7__23_) );
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf46), .D(_1527_), .Q(REGs_REGS_7__24_) );
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf33), .D(_1528_), .Q(REGs_REGS_7__25_) );
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf37), .D(_1529_), .Q(REGs_REGS_7__26_) );
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf33), .D(_1530_), .Q(REGs_REGS_7__27_) );
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf81), .D(_1531_), .Q(REGs_REGS_7__28_) );
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf16), .D(_1532_), .Q(REGs_REGS_7__29_) );
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf39), .D(_1533_), .Q(REGs_REGS_7__30_) );
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf82), .D(_1534_), .Q(REGs_REGS_7__31_) );
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf34), .D(_1407_), .Q(REGs_FIRQ_REGS_7__0_) );
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf73), .D(_1408_), .Q(REGs_FIRQ_REGS_7__1_) );
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf82), .D(_1409_), .Q(REGs_FIRQ_REGS_7__2_) );
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf33), .D(_1410_), .Q(REGs_FIRQ_REGS_7__3_) );
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf86), .D(_1411_), .Q(REGs_FIRQ_REGS_7__4_) );
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf20), .D(_1412_), .Q(REGs_FIRQ_REGS_7__5_) );
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf84), .D(_1413_), .Q(REGs_FIRQ_REGS_7__6_) );
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf24), .D(_1414_), .Q(REGs_FIRQ_REGS_7__7_) );
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf85), .D(_1415_), .Q(REGs_FIRQ_REGS_7__8_) );
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf78), .D(_1416_), .Q(REGs_FIRQ_REGS_7__9_) );
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf75), .D(_1417_), .Q(REGs_FIRQ_REGS_7__10_) );
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf20), .D(_1418_), .Q(REGs_FIRQ_REGS_7__11_) );
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf84), .D(_1419_), .Q(REGs_FIRQ_REGS_7__12_) );
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf11), .D(_1420_), .Q(REGs_FIRQ_REGS_7__13_) );
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf75), .D(_1421_), .Q(REGs_FIRQ_REGS_7__14_) );
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf20), .D(_1422_), .Q(REGs_FIRQ_REGS_7__15_) );
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf25), .D(_1423_), .Q(REGs_FIRQ_REGS_7__16_) );
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf67), .D(_1424_), .Q(REGs_FIRQ_REGS_7__17_) );
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf75), .D(_1425_), .Q(REGs_FIRQ_REGS_7__18_) );
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf11), .D(_1426_), .Q(REGs_FIRQ_REGS_7__19_) );
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf2), .D(_1427_), .Q(REGs_FIRQ_REGS_7__20_) );
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf35), .D(_1428_), .Q(REGs_FIRQ_REGS_7__21_) );
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf74), .D(_1429_), .Q(REGs_FIRQ_REGS_7__22_) );
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf0), .D(_1430_), .Q(REGs_FIRQ_REGS_7__23_) );
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf11), .D(_1431_), .Q(REGs_FIRQ_REGS_7__24_) );
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf79), .D(_1432_), .Q(REGs_FIRQ_REGS_7__25_) );
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf56), .D(_1433_), .Q(REGs_FIRQ_REGS_7__26_) );
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf74), .D(_1434_), .Q(REGs_FIRQ_REGS_7__27_) );
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf0), .D(_1435_), .Q(REGs_FIRQ_REGS_7__28_) );
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf11), .D(_1436_), .Q(REGs_FIRQ_REGS_7__29_) );
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf24), .D(_1437_), .Q(REGs_FIRQ_REGS_7__30_) );
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf4), .D(_1438_), .Q(REGs_FIRQ_REGS_7__31_) );
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf60), .D(_1279_), .Q(REGs_REGS_2__0_) );
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf64), .D(_1280_), .Q(REGs_REGS_2__1_) );
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf61), .D(_1281_), .Q(REGs_REGS_2__2_) );
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf61), .D(_1282_), .Q(REGs_REGS_2__3_) );
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf48), .D(_1283_), .Q(REGs_REGS_2__4_) );
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf64), .D(_1284_), .Q(REGs_REGS_2__5_) );
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf57), .D(_1285_), .Q(REGs_REGS_2__6_) );
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf57), .D(_1286_), .Q(REGs_REGS_2__7_) );
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf81), .D(_1287_), .Q(REGs_REGS_2__8_) );
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf87), .D(_1288_), .Q(REGs_REGS_2__9_) );
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf51), .D(_1289_), .Q(REGs_REGS_2__10_) );
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf87), .D(_1290_), .Q(REGs_REGS_2__11_) );
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf43), .D(_1291_), .Q(REGs_REGS_2__12_) );
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf60), .D(_1292_), .Q(REGs_REGS_2__13_) );
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf77), .D(_1293_), .Q(REGs_REGS_2__14_) );
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf19), .D(_1294_), .Q(REGs_REGS_2__15_) );
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf51), .D(_1295_), .Q(REGs_REGS_2__16_) );
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf60), .D(_1296_), .Q(REGs_REGS_2__17_) );
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf51), .D(_1297_), .Q(REGs_REGS_2__18_) );
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf64), .D(_1298_), .Q(REGs_REGS_2__19_) );
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf43), .D(_1299_), .Q(REGs_REGS_2__20_) );
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf87), .D(_1300_), .Q(REGs_REGS_2__21_) );
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf48), .D(_1301_), .Q(REGs_REGS_2__22_) );
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf51), .D(_1302_), .Q(REGs_REGS_2__23_) );
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf60), .D(_1303_), .Q(REGs_REGS_2__24_) );
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf63), .D(_1304_), .Q(REGs_REGS_2__25_) );
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf48), .D(_1305_), .Q(REGs_REGS_2__26_) );
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf43), .D(_1306_), .Q(REGs_REGS_2__27_) );
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf64), .D(_1307_), .Q(REGs_REGS_2__28_) );
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf63), .D(_1308_), .Q(REGs_REGS_2__29_) );
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf43), .D(_1309_), .Q(REGs_REGS_2__30_) );
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf60), .D(_1310_), .Q(REGs_REGS_2__31_) );
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf83), .D(_895_), .Q(REGs_USR_REGS_0__0_) );
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf41), .D(_896_), .Q(REGs_USR_REGS_0__1_) );
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf24), .D(_897_), .Q(REGs_USR_REGS_0__2_) );
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf67), .D(_898_), .Q(REGs_USR_REGS_0__3_) );
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf88), .D(_899_), .Q(REGs_USR_REGS_0__4_) );
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf41), .D(_900_), .Q(REGs_USR_REGS_0__5_) );
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf22), .D(_901_), .Q(REGs_USR_REGS_0__6_) );
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf29), .D(_902_), .Q(REGs_USR_REGS_0__7_) );
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf34), .D(_903_), .Q(REGs_USR_REGS_0__8_) );
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf62), .D(_904_), .Q(REGs_USR_REGS_0__9_) );
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf26), .D(_905_), .Q(REGs_USR_REGS_0__10_) );
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf34), .D(_906_), .Q(REGs_USR_REGS_0__11_) );
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf88), .D(_907_), .Q(REGs_USR_REGS_0__12_) );
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf79), .D(_908_), .Q(REGs_USR_REGS_0__13_) );
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf42), .D(_909_), .Q(REGs_USR_REGS_0__14_) );
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf15), .D(_910_), .Q(REGs_USR_REGS_0__15_) );
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf62), .D(_911_), .Q(REGs_USR_REGS_0__16_) );
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf38), .D(_912_), .Q(REGs_USR_REGS_0__17_) );
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf42), .D(_913_), .Q(REGs_USR_REGS_0__18_) );
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf11), .D(_914_), .Q(REGs_USR_REGS_0__19_) );
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf74), .D(_915_), .Q(REGs_USR_REGS_0__20_) );
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf76), .D(_916_), .Q(REGs_USR_REGS_0__21_) );
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf88), .D(_917_), .Q(REGs_USR_REGS_0__22_) );
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf42), .D(_918_), .Q(REGs_USR_REGS_0__23_) );
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf79), .D(_919_), .Q(REGs_USR_REGS_0__24_) );
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf38), .D(_920_), .Q(REGs_USR_REGS_0__25_) );
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf29), .D(_921_), .Q(REGs_USR_REGS_0__26_) );
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf38), .D(_922_), .Q(REGs_USR_REGS_0__27_) );
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf10), .D(_923_), .Q(REGs_USR_REGS_0__28_) );
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf82), .D(_924_), .Q(REGs_USR_REGS_0__29_) );
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf67), .D(_925_), .Q(REGs_USR_REGS_0__30_) );
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf2), .D(_926_), .Q(REGs_USR_REGS_0__31_) );
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf83), .D(_1087_), .Q(REGs_FIRQ_REGS_0__0_) );
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf41), .D(_1088_), .Q(REGs_FIRQ_REGS_0__1_) );
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf2), .D(_1089_), .Q(REGs_FIRQ_REGS_0__2_) );
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf37), .D(_1090_), .Q(REGs_FIRQ_REGS_0__3_) );
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf22), .D(_1091_), .Q(REGs_FIRQ_REGS_0__4_) );
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf4), .D(_1092_), .Q(REGs_FIRQ_REGS_0__5_) );
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf22), .D(_1093_), .Q(REGs_FIRQ_REGS_0__6_) );
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf29), .D(_1094_), .Q(REGs_FIRQ_REGS_0__7_) );
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf34), .D(_1095_), .Q(REGs_FIRQ_REGS_0__8_) );
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf26), .D(_1096_), .Q(REGs_FIRQ_REGS_0__9_) );
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf26), .D(_1097_), .Q(REGs_FIRQ_REGS_0__10_) );
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf12), .D(_1098_), .Q(REGs_FIRQ_REGS_0__11_) );
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf22), .D(_1099_), .Q(REGs_FIRQ_REGS_0__12_) );
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf83), .D(_1100_), .Q(REGs_FIRQ_REGS_0__13_) );
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf59), .D(_1101_), .Q(REGs_FIRQ_REGS_0__14_) );
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf10), .D(_1102_), .Q(REGs_FIRQ_REGS_0__15_) );
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf10), .D(_1103_), .Q(REGs_FIRQ_REGS_0__16_) );
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf29), .D(_1104_), .Q(REGs_FIRQ_REGS_0__17_) );
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf42), .D(_1105_), .Q(REGs_FIRQ_REGS_0__18_) );
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf34), .D(_1106_), .Q(REGs_FIRQ_REGS_0__19_) );
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf74), .D(_1107_), .Q(REGs_FIRQ_REGS_0__20_) );
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf54), .D(_1108_), .Q(REGs_FIRQ_REGS_0__21_) );
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf88), .D(_1109_), .Q(REGs_FIRQ_REGS_0__22_) );
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf26), .D(_1110_), .Q(REGs_FIRQ_REGS_0__23_) );
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf79), .D(_1111_), .Q(REGs_FIRQ_REGS_0__24_) );
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf38), .D(_1112_), .Q(REGs_FIRQ_REGS_0__25_) );
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf38), .D(_1113_), .Q(REGs_FIRQ_REGS_0__26_) );
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf38), .D(_1114_), .Q(REGs_FIRQ_REGS_0__27_) );
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf66), .D(_1115_), .Q(REGs_FIRQ_REGS_0__28_) );
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf82), .D(_1116_), .Q(REGs_FIRQ_REGS_0__29_) );
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf67), .D(_1117_), .Q(REGs_FIRQ_REGS_0__30_) );
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf2), .D(_1118_), .Q(REGs_FIRQ_REGS_0__31_) );
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf44), .D(_1311_), .Q(REGs_FIRQ_REGS_5__0_) );
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf47), .D(_1312_), .Q(REGs_FIRQ_REGS_5__1_) );
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf67), .D(_1313_), .Q(REGs_FIRQ_REGS_5__2_) );
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf58), .D(_1314_), .Q(REGs_FIRQ_REGS_5__3_) );
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf86), .D(_1315_), .Q(REGs_FIRQ_REGS_5__4_) );
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf20), .D(_1316_), .Q(REGs_FIRQ_REGS_5__5_) );
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf86), .D(_1317_), .Q(REGs_FIRQ_REGS_5__6_) );
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf67), .D(_1318_), .Q(REGs_FIRQ_REGS_5__7_) );
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf62), .D(_1319_), .Q(REGs_FIRQ_REGS_5__8_) );
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf3), .D(_1320_), .Q(REGs_FIRQ_REGS_5__9_) );
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf73), .D(_1321_), .Q(REGs_FIRQ_REGS_5__10_) );
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf26), .D(_1322_), .Q(REGs_FIRQ_REGS_5__11_) );
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf86), .D(_1323_), .Q(REGs_FIRQ_REGS_5__12_) );
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf52), .D(_1324_), .Q(REGs_FIRQ_REGS_5__13_) );
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf73), .D(_1325_), .Q(REGs_FIRQ_REGS_5__14_) );
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf47), .D(_1326_), .Q(REGs_FIRQ_REGS_5__15_) );
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf3), .D(_1327_), .Q(REGs_FIRQ_REGS_5__16_) );
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf71), .D(_1328_), .Q(REGs_FIRQ_REGS_5__17_) );
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf14), .D(_1329_), .Q(REGs_FIRQ_REGS_5__18_) );
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf11), .D(_1330_), .Q(REGs_FIRQ_REGS_5__19_) );
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf67), .D(_1331_), .Q(REGs_FIRQ_REGS_5__20_) );
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf52), .D(_1332_), .Q(REGs_FIRQ_REGS_5__21_) );
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf74), .D(_1333_), .Q(REGs_FIRQ_REGS_5__22_) );
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf75), .D(_1334_), .Q(REGs_FIRQ_REGS_5__23_) );
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf11), .D(_1335_), .Q(REGs_FIRQ_REGS_5__24_) );
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf52), .D(_1336_), .Q(REGs_FIRQ_REGS_5__25_) );
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf74), .D(_1337_), .Q(REGs_FIRQ_REGS_5__26_) );
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf74), .D(_1338_), .Q(REGs_FIRQ_REGS_5__27_) );
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf15), .D(_1339_), .Q(REGs_FIRQ_REGS_5__28_) );
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf52), .D(_1340_), .Q(REGs_FIRQ_REGS_5__29_) );
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf71), .D(_1341_), .Q(REGs_FIRQ_REGS_5__30_) );
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf3), .D(_1342_), .Q(REGs_FIRQ_REGS_5__31_) );
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf80), .D(_1247_), .Q(REGs_USR_REGS_1__0_) );
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf10), .D(_1248_), .Q(REGs_USR_REGS_1__1_) );
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf2), .D(_1249_), .Q(REGs_USR_REGS_1__2_) );
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf18), .D(_1250_), .Q(REGs_USR_REGS_1__3_) );
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf49), .D(_1251_), .Q(REGs_USR_REGS_1__4_) );
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf10), .D(_1252_), .Q(REGs_USR_REGS_1__5_) );
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf49), .D(_1253_), .Q(REGs_USR_REGS_1__6_) );
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf1), .D(_1254_), .Q(REGs_USR_REGS_1__7_) );
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf44), .D(_1255_), .Q(REGs_USR_REGS_1__8_) );
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf41), .D(_1256_), .Q(REGs_USR_REGS_1__9_) );
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf62), .D(_1257_), .Q(REGs_USR_REGS_1__10_) );
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf76), .D(_1258_), .Q(REGs_USR_REGS_1__11_) );
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf45), .D(_1259_), .Q(REGs_USR_REGS_1__12_) );
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf83), .D(_1260_), .Q(REGs_USR_REGS_1__13_) );
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf59), .D(_1261_), .Q(REGs_USR_REGS_1__14_) );
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf76), .D(_1262_), .Q(REGs_USR_REGS_1__15_) );
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf10), .D(_1263_), .Q(REGs_USR_REGS_1__16_) );
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf80), .D(_1264_), .Q(REGs_USR_REGS_1__17_) );
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf42), .D(_1265_), .Q(REGs_USR_REGS_1__18_) );
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf44), .D(_1266_), .Q(REGs_USR_REGS_1__19_) );
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf50), .D(_1267_), .Q(REGs_USR_REGS_1__20_) );
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf54), .D(_1268_), .Q(REGs_USR_REGS_1__21_) );
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf49), .D(_1269_), .Q(REGs_USR_REGS_1__22_) );
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf59), .D(_1270_), .Q(REGs_USR_REGS_1__23_) );
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf13), .D(_1271_), .Q(REGs_USR_REGS_1__24_) );
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf80), .D(_1272_), .Q(REGs_USR_REGS_1__25_) );
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf45), .D(_1273_), .Q(REGs_USR_REGS_1__26_) );
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf29), .D(_1274_), .Q(REGs_USR_REGS_1__27_) );
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf54), .D(_1275_), .Q(REGs_USR_REGS_1__28_) );
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf34), .D(_1276_), .Q(REGs_USR_REGS_1__29_) );
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf24), .D(_1277_), .Q(REGs_USR_REGS_1__30_) );
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf2), .D(_1278_), .Q(REGs_USR_REGS_1__31_) );
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf82), .D(_1471_), .Q(REGs_USR_REGS_2__0_) );
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf9), .D(_1472_), .Q(REGs_USR_REGS_2__1_) );
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf24), .D(_1473_), .Q(REGs_USR_REGS_2__2_) );
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf12), .D(_1474_), .Q(REGs_USR_REGS_2__3_) );
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf23), .D(_1475_), .Q(REGs_USR_REGS_2__4_) );
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf41), .D(_1476_), .Q(REGs_USR_REGS_2__5_) );
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf23), .D(_1477_), .Q(REGs_USR_REGS_2__6_) );
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf1), .D(_1478_), .Q(REGs_USR_REGS_2__7_) );
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf44), .D(_1479_), .Q(REGs_USR_REGS_2__8_) );
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf41), .D(_1480_), .Q(REGs_USR_REGS_2__9_) );
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf15), .D(_1481_), .Q(REGs_USR_REGS_2__10_) );
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf70), .D(_1482_), .Q(REGs_USR_REGS_2__11_) );
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf38), .D(_1483_), .Q(REGs_USR_REGS_2__12_) );
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf1), .D(_1484_), .Q(REGs_USR_REGS_2__13_) );
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf32), .D(_1485_), .Q(REGs_USR_REGS_2__14_) );
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf59), .D(_1486_), .Q(REGs_USR_REGS_2__15_) );
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf32), .D(_1487_), .Q(REGs_USR_REGS_2__16_) );
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf80), .D(_1488_), .Q(REGs_USR_REGS_2__17_) );
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf25), .D(_1489_), .Q(REGs_USR_REGS_2__18_) );
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf4), .D(_1490_), .Q(REGs_USR_REGS_2__19_) );
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf50), .D(_1491_), .Q(REGs_USR_REGS_2__20_) );
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf66), .D(_1492_), .Q(REGs_USR_REGS_2__21_) );
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf45), .D(_1493_), .Q(REGs_USR_REGS_2__22_) );
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf66), .D(_1494_), .Q(REGs_USR_REGS_2__23_) );
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf12), .D(_1495_), .Q(REGs_USR_REGS_2__24_) );
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf1), .D(_1496_), .Q(REGs_USR_REGS_2__25_) );
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf23), .D(_1497_), .Q(REGs_USR_REGS_2__26_) );
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf29), .D(_1498_), .Q(REGs_USR_REGS_2__27_) );
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf9), .D(_1499_), .Q(REGs_USR_REGS_2__28_) );
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf12), .D(_1500_), .Q(REGs_USR_REGS_2__29_) );
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf50), .D(_1501_), .Q(REGs_USR_REGS_2__30_) );
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf58), .D(_1502_), .Q(REGs_USR_REGS_2__31_) );
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf50), .D(_1439_), .Q(REGs_USR_REGS_3__0_) );
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf9), .D(_1440_), .Q(REGs_USR_REGS_3__1_) );
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf7), .D(_1441_), .Q(REGs_USR_REGS_3__2_) );
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf58), .D(_1442_), .Q(REGs_USR_REGS_3__3_) );
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf45), .D(_1443_), .Q(REGs_USR_REGS_3__4_) );
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf76), .D(_1444_), .Q(REGs_USR_REGS_3__5_) );
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf45), .D(_1445_), .Q(REGs_USR_REGS_3__6_) );
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf30), .D(_1446_), .Q(REGs_USR_REGS_3__7_) );
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf54), .D(_1447_), .Q(REGs_USR_REGS_3__8_) );
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf59), .D(_1448_), .Q(REGs_USR_REGS_3__9_) );
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf26), .D(_1449_), .Q(REGs_USR_REGS_3__10_) );
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf9), .D(_1450_), .Q(REGs_USR_REGS_3__11_) );
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf23), .D(_1451_), .Q(REGs_USR_REGS_3__12_) );
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf30), .D(_1452_), .Q(REGs_USR_REGS_3__13_) );
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf59), .D(_1453_), .Q(REGs_USR_REGS_3__14_) );
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf59), .D(_1454_), .Q(REGs_USR_REGS_3__15_) );
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf62), .D(_1455_), .Q(REGs_USR_REGS_3__16_) );
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf1), .D(_1456_), .Q(REGs_USR_REGS_3__17_) );
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf85), .D(_1457_), .Q(REGs_USR_REGS_3__18_) );
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf70), .D(_1458_), .Q(REGs_USR_REGS_3__19_) );
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf80), .D(_1459_), .Q(REGs_USR_REGS_3__20_) );
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf76), .D(_1460_), .Q(REGs_USR_REGS_3__21_) );
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf45), .D(_1461_), .Q(REGs_USR_REGS_3__22_) );
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf66), .D(_1462_), .Q(REGs_USR_REGS_3__23_) );
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf12), .D(_1463_), .Q(REGs_USR_REGS_3__24_) );
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf30), .D(_1464_), .Q(REGs_USR_REGS_3__25_) );
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf29), .D(_1465_), .Q(REGs_USR_REGS_3__26_) );
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf30), .D(_1466_), .Q(REGs_USR_REGS_3__27_) );
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf10), .D(_1467_), .Q(REGs_USR_REGS_3__28_) );
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf82), .D(_1468_), .Q(REGs_USR_REGS_3__29_) );
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf7), .D(_1469_), .Q(REGs_USR_REGS_3__30_) );
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf70), .D(_1470_), .Q(REGs_USR_REGS_3__31_) );
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf70), .D(_1375_), .Q(REGs_USR_REGS_4__0_) );
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf47), .D(_1376_), .Q(REGs_USR_REGS_4__1_) );
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf71), .D(_1377_), .Q(REGs_USR_REGS_4__2_) );
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf7), .D(_1378_), .Q(REGs_USR_REGS_4__3_) );
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf86), .D(_1379_), .Q(REGs_USR_REGS_4__4_) );
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf73), .D(_1380_), .Q(REGs_USR_REGS_4__5_) );
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf88), .D(_1381_), .Q(REGs_USR_REGS_4__6_) );
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf13), .D(_1382_), .Q(REGs_USR_REGS_4__7_) );
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf66), .D(_1383_), .Q(REGs_USR_REGS_4__8_) );
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf14), .D(_1384_), .Q(REGs_USR_REGS_4__9_) );
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf3), .D(_1385_), .Q(REGs_USR_REGS_4__10_) );
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf32), .D(_1386_), .Q(REGs_USR_REGS_4__11_) );
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf88), .D(_1387_), .Q(REGs_USR_REGS_4__12_) );
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf52), .D(_1388_), .Q(REGs_USR_REGS_4__13_) );
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf75), .D(_1389_), .Q(REGs_USR_REGS_4__14_) );
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf32), .D(_1390_), .Q(REGs_USR_REGS_4__15_) );
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf14), .D(_1391_), .Q(REGs_USR_REGS_4__16_) );
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf83), .D(_1392_), .Q(REGs_USR_REGS_4__17_) );
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf14), .D(_1393_), .Q(REGs_USR_REGS_4__18_) );
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf9), .D(_1394_), .Q(REGs_USR_REGS_4__19_) );
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf13), .D(_1395_), .Q(REGs_USR_REGS_4__20_) );
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf54), .D(_1396_), .Q(REGs_USR_REGS_4__21_) );
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf88), .D(_1397_), .Q(REGs_USR_REGS_4__22_) );
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf14), .D(_1398_), .Q(REGs_USR_REGS_4__23_) );
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf5), .D(_1399_), .Q(REGs_USR_REGS_4__24_) );
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf5), .D(_1400_), .Q(REGs_USR_REGS_4__25_) );
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf49), .D(_1401_), .Q(REGs_USR_REGS_4__26_) );
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf56), .D(_1402_), .Q(REGs_USR_REGS_4__27_) );
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf25), .D(_1403_), .Q(REGs_USR_REGS_4__28_) );
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf34), .D(_1404_), .Q(REGs_USR_REGS_4__29_) );
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf24), .D(_1405_), .Q(REGs_USR_REGS_4__30_) );
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf32), .D(_1406_), .Q(REGs_USR_REGS_4__31_) );
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf44), .D(_927_), .Q(REGs_USR_REGS_5__0_) );
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf47), .D(_928_), .Q(REGs_USR_REGS_5__1_) );
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf67), .D(_929_), .Q(REGs_USR_REGS_5__2_) );
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf58), .D(_930_), .Q(REGs_USR_REGS_5__3_) );
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf84), .D(_931_), .Q(REGs_USR_REGS_5__4_) );
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf73), .D(_932_), .Q(REGs_USR_REGS_5__5_) );
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf86), .D(_933_), .Q(REGs_USR_REGS_5__6_) );
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf18), .D(_934_), .Q(REGs_USR_REGS_5__7_) );
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf62), .D(_935_), .Q(REGs_USR_REGS_5__8_) );
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf75), .D(_936_), .Q(REGs_USR_REGS_5__9_) );
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf73), .D(_937_), .Q(REGs_USR_REGS_5__10_) );
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf26), .D(_938_), .Q(REGs_USR_REGS_5__11_) );
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf84), .D(_939_), .Q(REGs_USR_REGS_5__12_) );
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf52), .D(_940_), .Q(REGs_USR_REGS_5__13_) );
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf73), .D(_941_), .Q(REGs_USR_REGS_5__14_) );
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf47), .D(_942_), .Q(REGs_USR_REGS_5__15_) );
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf20), .D(_943_), .Q(REGs_USR_REGS_5__16_) );
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf71), .D(_944_), .Q(REGs_USR_REGS_5__17_) );
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf47), .D(_945_), .Q(REGs_USR_REGS_5__18_) );
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf44), .D(_946_), .Q(REGs_USR_REGS_5__19_) );
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf7), .D(_947_), .Q(REGs_USR_REGS_5__20_) );
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf52), .D(_948_), .Q(REGs_USR_REGS_5__21_) );
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf84), .D(_949_), .Q(REGs_USR_REGS_5__22_) );
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf14), .D(_950_), .Q(REGs_USR_REGS_5__23_) );
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf5), .D(_951_), .Q(REGs_USR_REGS_5__24_) );
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf62), .D(_952_), .Q(REGs_USR_REGS_5__25_) );
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf74), .D(_953_), .Q(REGs_USR_REGS_5__26_) );
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf18), .D(_954_), .Q(REGs_USR_REGS_5__27_) );
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf76), .D(_955_), .Q(REGs_USR_REGS_5__28_) );
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf52), .D(_956_), .Q(REGs_USR_REGS_5__29_) );
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf71), .D(_957_), .Q(REGs_USR_REGS_5__30_) );
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf20), .D(_958_), .Q(REGs_USR_REGS_5__31_) );
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf12), .D(_863_), .Q(REGs_USR_REGS_6__0_) );
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf15), .D(_864_), .Q(REGs_USR_REGS_6__1_) );
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf7), .D(_865_), .Q(REGs_USR_REGS_6__2_) );
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf67), .D(_866_), .Q(REGs_USR_REGS_6__3_) );
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf18), .D(_867_), .Q(REGs_USR_REGS_6__4_) );
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf3), .D(_868_), .Q(REGs_USR_REGS_6__5_) );
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf23), .D(_869_), .Q(REGs_USR_REGS_6__6_) );
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf18), .D(_870_), .Q(REGs_USR_REGS_6__7_) );
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf76), .D(_871_), .Q(REGs_USR_REGS_6__8_) );
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf3), .D(_872_), .Q(REGs_USR_REGS_6__9_) );
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf78), .D(_873_), .Q(REGs_USR_REGS_6__10_) );
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf3), .D(_874_), .Q(REGs_USR_REGS_6__11_) );
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf38), .D(_875_), .Q(REGs_USR_REGS_6__12_) );
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf83), .D(_876_), .Q(REGs_USR_REGS_6__13_) );
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf0), .D(_877_), .Q(REGs_USR_REGS_6__14_) );
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf3), .D(_878_), .Q(REGs_USR_REGS_6__15_) );
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf78), .D(_879_), .Q(REGs_USR_REGS_6__16_) );
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf83), .D(_880_), .Q(REGs_USR_REGS_6__17_) );
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf25), .D(_881_), .Q(REGs_USR_REGS_6__18_) );
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf9), .D(_882_), .Q(REGs_USR_REGS_6__19_) );
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf24), .D(_883_), .Q(REGs_USR_REGS_6__20_) );
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf35), .D(_884_), .Q(REGs_USR_REGS_6__21_) );
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf86), .D(_885_), .Q(REGs_USR_REGS_6__22_) );
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf35), .D(_886_), .Q(REGs_USR_REGS_6__23_) );
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf11), .D(_887_), .Q(REGs_USR_REGS_6__24_) );
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf83), .D(_888_), .Q(REGs_USR_REGS_6__25_) );
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf56), .D(_889_), .Q(REGs_USR_REGS_6__26_) );
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf56), .D(_890_), .Q(REGs_USR_REGS_6__27_) );
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf78), .D(_891_), .Q(REGs_USR_REGS_6__28_) );
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf12), .D(_892_), .Q(REGs_USR_REGS_6__29_) );
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf56), .D(_893_), .Q(REGs_USR_REGS_6__30_) );
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf25), .D(_894_), .Q(REGs_USR_REGS_6__31_) );
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf12), .D(_959_), .Q(REGs_USR_REGS_7__0_) );
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf73), .D(_960_), .Q(REGs_USR_REGS_7__1_) );
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf82), .D(_961_), .Q(REGs_USR_REGS_7__2_) );
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf71), .D(_962_), .Q(REGs_USR_REGS_7__3_) );
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf86), .D(_963_), .Q(REGs_USR_REGS_7__4_) );
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf78), .D(_964_), .Q(REGs_USR_REGS_7__5_) );
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf86), .D(_965_), .Q(REGs_USR_REGS_7__6_) );
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf13), .D(_966_), .Q(REGs_USR_REGS_7__7_) );
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf4), .D(_967_), .Q(REGs_USR_REGS_7__8_) );
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf78), .D(_968_), .Q(REGs_USR_REGS_7__9_) );
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf73), .D(_969_), .Q(REGs_USR_REGS_7__10_) );
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf47), .D(_970_), .Q(REGs_USR_REGS_7__11_) );
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf84), .D(_971_), .Q(REGs_USR_REGS_7__12_) );
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf79), .D(_972_), .Q(REGs_USR_REGS_7__13_) );
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf75), .D(_973_), .Q(REGs_USR_REGS_7__14_) );
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf47), .D(_974_), .Q(REGs_USR_REGS_7__15_) );
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf25), .D(_975_), .Q(REGs_USR_REGS_7__16_) );
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf71), .D(_976_), .Q(REGs_USR_REGS_7__17_) );
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf75), .D(_977_), .Q(REGs_USR_REGS_7__18_) );
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf79), .D(_978_), .Q(REGs_USR_REGS_7__19_) );
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf24), .D(_979_), .Q(REGs_USR_REGS_7__20_) );
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf35), .D(_980_), .Q(REGs_USR_REGS_7__21_) );
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf74), .D(_981_), .Q(REGs_USR_REGS_7__22_) );
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf47), .D(_982_), .Q(REGs_USR_REGS_7__23_) );
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf79), .D(_983_), .Q(REGs_USR_REGS_7__24_) );
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf13), .D(_984_), .Q(REGs_USR_REGS_7__25_) );
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf37), .D(_985_), .Q(REGs_USR_REGS_7__26_) );
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf37), .D(_986_), .Q(REGs_USR_REGS_7__27_) );
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf35), .D(_987_), .Q(REGs_USR_REGS_7__28_) );
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf4), .D(_988_), .Q(REGs_USR_REGS_7__29_) );
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf83), .D(_989_), .Q(REGs_USR_REGS_7__30_) );
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf25), .D(_990_), .Q(REGs_USR_REGS_7__31_) );
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf70), .D(_1215_), .Q(REGs_FIRQ_REGS_4__0_) );
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf15), .D(_1216_), .Q(REGs_FIRQ_REGS_4__1_) );
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf58), .D(_1217_), .Q(REGs_FIRQ_REGS_4__2_) );
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf71), .D(_1218_), .Q(REGs_FIRQ_REGS_4__3_) );
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf22), .D(_1219_), .Q(REGs_FIRQ_REGS_4__4_) );
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf73), .D(_1220_), .Q(REGs_FIRQ_REGS_4__5_) );
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf88), .D(_1221_), .Q(REGs_FIRQ_REGS_4__6_) );
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf13), .D(_1222_), .Q(REGs_FIRQ_REGS_4__7_) );
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf15), .D(_1223_), .Q(REGs_FIRQ_REGS_4__8_) );
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf75), .D(_1224_), .Q(REGs_FIRQ_REGS_4__9_) );
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf3), .D(_1225_), .Q(REGs_FIRQ_REGS_4__10_) );
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf32), .D(_1226_), .Q(REGs_FIRQ_REGS_4__11_) );
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf84), .D(_1227_), .Q(REGs_FIRQ_REGS_4__12_) );
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf52), .D(_1228_), .Q(REGs_FIRQ_REGS_4__13_) );
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf75), .D(_1229_), .Q(REGs_FIRQ_REGS_4__14_) );
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf20), .D(_1230_), .Q(REGs_FIRQ_REGS_4__15_) );
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf14), .D(_1231_), .Q(REGs_FIRQ_REGS_4__16_) );
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf83), .D(_1232_), .Q(REGs_FIRQ_REGS_4__17_) );
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf14), .D(_1233_), .Q(REGs_FIRQ_REGS_4__18_) );
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf44), .D(_1234_), .Q(REGs_FIRQ_REGS_4__19_) );
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf31), .D(_1235_), .Q(REGs_FIRQ_REGS_4__20_) );
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf54), .D(_1236_), .Q(REGs_FIRQ_REGS_4__21_) );
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf22), .D(_1237_), .Q(REGs_FIRQ_REGS_4__22_) );
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf14), .D(_1238_), .Q(REGs_FIRQ_REGS_4__23_) );
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf31), .D(_1239_), .Q(REGs_FIRQ_REGS_4__24_) );
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf5), .D(_1240_), .Q(REGs_FIRQ_REGS_4__25_) );
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf56), .D(_1241_), .Q(REGs_FIRQ_REGS_4__26_) );
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf74), .D(_1242_), .Q(REGs_FIRQ_REGS_4__27_) );
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf25), .D(_1243_), .Q(REGs_FIRQ_REGS_4__28_) );
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf44), .D(_1244_), .Q(REGs_FIRQ_REGS_4__29_) );
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf67), .D(_1245_), .Q(REGs_FIRQ_REGS_4__30_) );
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf32), .D(_1246_), .Q(REGs_FIRQ_REGS_4__31_) );
INVX2 INVX2_1 ( .A(ULA_B_3_bF_buf7), .Y(_5289_) );
OR2X2 OR2X2_404 ( .A(ULA_B_0_bF_buf3), .B(ULA_B_1_bF_buf1), .Y(_5300_) );
OR2X2 OR2X2_405 ( .A(ULA_B_2_bF_buf1), .B(_5300_), .Y(_5310_) );
NAND2X1 NAND2X1_641 ( .A(ULA_cin_bF_buf2), .B(_5310_), .Y(_5321_) );
XOR2X1 XOR2X1_1 ( .A(_5289__bF_buf5), .B(_5321_), .Y(_5332_) );
AND2X2 AND2X2_430 ( .A(_5300_), .B(ULA_cin_bF_buf2), .Y(_5342_) );
XNOR2X1 XNOR2X1_1 ( .A(ULA_B_2_bF_buf0), .B(_5342_), .Y(_5353_) );
MUX2X1 MUX2X1_641 ( .A(ULA_A_25_), .B(ULA_A_24_), .S(ULA_B_0_bF_buf2), .Y(_5364_) );
OR2X2 OR2X2_406 ( .A(ULA_cin_bF_buf2), .B(ULA_B_1_bF_buf2), .Y(_5374_) );
INVX1 INVX1_4 ( .A(_5374_), .Y(_5385_) );
XNOR2X1 XNOR2X1_2 ( .A(ULA_B_0_bF_buf7), .B(ULA_B_1_bF_buf3), .Y(_5396_) );
AND2X2 AND2X2_431 ( .A(_5396_), .B(ULA_cin_bF_buf2), .Y(_5406_) );
OR2X2 OR2X2_407 ( .A(_5385_), .B(_5406_), .Y(_5417_) );
AND2X2 AND2X2_432 ( .A(_5417__bF_buf2), .B(_5364_), .Y(_5428_) );
INVX2 INVX2_2 ( .A(ULA_cin_bF_buf1), .Y(_5438_) );
XOR2X1 XOR2X1_2 ( .A(ULA_B_0_bF_buf7), .B(ULA_B_1_bF_buf3), .Y(_5449_) );
OR2X2 OR2X2_408 ( .A(_5438__bF_buf3), .B(_5449_), .Y(_5460_) );
AND2X2 AND2X2_433 ( .A(_5460_), .B(_5374_), .Y(_5470_) );
MUX2X1 MUX2X1_642 ( .A(ULA_A_27_), .B(ULA_A_26_), .S(ULA_B_0_bF_buf2), .Y(_5481_) );
AND2X2 AND2X2_434 ( .A(_5470__bF_buf3), .B(_5481_), .Y(_5492_) );
OR2X2 OR2X2_409 ( .A(_5428_), .B(_5492_), .Y(_5502_) );
AND2X2 AND2X2_435 ( .A(_5502_), .B(_5353__bF_buf3), .Y(_5513_) );
XOR2X1 XOR2X1_3 ( .A(ULA_B_2_bF_buf0), .B(_5342_), .Y(_5524_) );
MUX2X1 MUX2X1_643 ( .A(ULA_A_31_), .B(ULA_A_30_), .S(ULA_B_0_bF_buf6), .Y(_5534_) );
AND2X2 AND2X2_436 ( .A(_5470__bF_buf3), .B(_5534_), .Y(_5545_) );
MUX2X1 MUX2X1_644 ( .A(ULA_A_29_), .B(ULA_A_28_), .S(ULA_B_0_bF_buf4), .Y(_5556_) );
AND2X2 AND2X2_437 ( .A(_5417__bF_buf2), .B(_5556_), .Y(_5566_) );
OR2X2 OR2X2_410 ( .A(_5566_), .B(_5545_), .Y(_5577_) );
AND2X2 AND2X2_438 ( .A(_5577_), .B(_5524__bF_buf3), .Y(_5588_) );
OR2X2 OR2X2_411 ( .A(_5513_), .B(_5588_), .Y(_5598_) );
AND2X2 AND2X2_439 ( .A(_5598_), .B(_5332__bF_buf0), .Y(_5609_) );
XOR2X1 XOR2X1_4 ( .A(ULA_B_3_bF_buf5), .B(_5321_), .Y(_5620_) );
MUX2X1 MUX2X1_645 ( .A(ULA_A_21_), .B(ULA_A_20_), .S(ULA_B_0_bF_buf2), .Y(_5630_) );
AND2X2 AND2X2_440 ( .A(_5417__bF_buf3), .B(_5630_), .Y(_5641_) );
MUX2X1 MUX2X1_646 ( .A(ULA_A_23_), .B(ULA_A_22_), .S(ULA_B_0_bF_buf2), .Y(_5652_) );
AND2X2 AND2X2_441 ( .A(_5470__bF_buf3), .B(_5652_), .Y(_5657_) );
OR2X2 OR2X2_412 ( .A(_5641_), .B(_5657_), .Y(_5658_) );
AND2X2 AND2X2_442 ( .A(_5658_), .B(_5524__bF_buf0), .Y(_5659_) );
MUX2X1 MUX2X1_647 ( .A(ULA_A_17_), .B(ULA_A_16_), .S(ULA_B_0_bF_buf7), .Y(_5660_) );
AND2X2 AND2X2_443 ( .A(_5417__bF_buf3), .B(_5660_), .Y(_5661_) );
MUX2X1 MUX2X1_648 ( .A(ULA_A_19_), .B(ULA_A_18_), .S(ULA_B_0_bF_buf2), .Y(_5662_) );
AND2X2 AND2X2_444 ( .A(_5470__bF_buf0), .B(_5662_), .Y(_5663_) );
OR2X2 OR2X2_413 ( .A(_5661_), .B(_5663_), .Y(_5664_) );
AND2X2 AND2X2_445 ( .A(_5664_), .B(_5353__bF_buf1), .Y(_5665_) );
OR2X2 OR2X2_414 ( .A(_5659_), .B(_5665_), .Y(_5666_) );
AND2X2 AND2X2_446 ( .A(_5666_), .B(_5620__bF_buf0), .Y(_5667_) );
OR2X2 OR2X2_415 ( .A(_5609_), .B(_5667_), .Y(_5668_) );
INVX1 INVX1_5 ( .A(ULA_B_4_bF_buf2), .Y(_5669_) );
OR2X2 OR2X2_416 ( .A(ULA_B_3_bF_buf0), .B(_5310_), .Y(_5670_) );
AND2X2 AND2X2_447 ( .A(_5670_), .B(ULA_cin_bF_buf2), .Y(_5671_) );
XOR2X1 XOR2X1_5 ( .A(_5669__bF_buf3), .B(_5671_), .Y(_5672_) );
INVX1 INVX1_6 ( .A(CORE_ULA_ctrl_2_), .Y(_5673_) );
INVX1 INVX1_7 ( .A(CORE_ULA_ctrl_1_), .Y(_5674_) );
NAND3X1 NAND3X1_11 ( .A(_5673_), .B(CORE_ULA_ctrl_3_), .C(_5674_), .Y(_5675_) );
AND2X2 AND2X2_448 ( .A(CORE_ULA_ctrl_2_), .B(CORE_ULA_ctrl_1_), .Y(_5676_) );
NAND2X1 NAND2X1_642 ( .A(CORE_ULA_ctrl_3_), .B(_5676_), .Y(_5677_) );
AND2X2 AND2X2_449 ( .A(_5675_), .B(_5677_), .Y(_5678_) );
OR2X2 OR2X2_417 ( .A(_5672_), .B(_5678_), .Y(_5679_) );
OR2X2 OR2X2_418 ( .A(_5679_), .B(_5668_), .Y(_5680_) );
INVX2 INVX2_3 ( .A(ULA_B_2_bF_buf3), .Y(_5681_) );
INVX2 INVX2_4 ( .A(ULA_B_1_bF_buf2), .Y(_5682_) );
AND2X2 AND2X2_450 ( .A(_5660_), .B(_5682__bF_buf1), .Y(_5683_) );
AND2X2 AND2X2_451 ( .A(_5662_), .B(ULA_B_1_bF_buf2), .Y(_5684_) );
OR2X2 OR2X2_419 ( .A(_5683_), .B(_5684_), .Y(_5685_) );
AND2X2 AND2X2_452 ( .A(_5685_), .B(_5681__bF_buf5), .Y(_5686_) );
AND2X2 AND2X2_453 ( .A(_5630_), .B(_5682__bF_buf3), .Y(_5687_) );
AND2X2 AND2X2_454 ( .A(_5652_), .B(ULA_B_1_bF_buf3), .Y(_5688_) );
OR2X2 OR2X2_420 ( .A(_5687_), .B(_5688_), .Y(_5689_) );
AND2X2 AND2X2_455 ( .A(_5689_), .B(ULA_B_2_bF_buf1), .Y(_5690_) );
OR2X2 OR2X2_421 ( .A(_5686_), .B(_5690_), .Y(_5691_) );
AND2X2 AND2X2_456 ( .A(_5691_), .B(_5289__bF_buf3), .Y(_5692_) );
AND2X2 AND2X2_457 ( .A(_5556_), .B(_5682__bF_buf1), .Y(_5693_) );
AND2X2 AND2X2_458 ( .A(_5534_), .B(ULA_B_1_bF_buf0), .Y(_5694_) );
OR2X2 OR2X2_422 ( .A(_5693_), .B(_5694_), .Y(_5695_) );
AND2X2 AND2X2_459 ( .A(_5695_), .B(ULA_B_2_bF_buf1), .Y(_5696_) );
AND2X2 AND2X2_460 ( .A(_5481_), .B(ULA_B_1_bF_buf3), .Y(_5697_) );
AND2X2 AND2X2_461 ( .A(_5364_), .B(_5682__bF_buf3), .Y(_5698_) );
OR2X2 OR2X2_423 ( .A(_5697_), .B(_5698_), .Y(_5699_) );
AND2X2 AND2X2_462 ( .A(_5699_), .B(_5681__bF_buf3), .Y(_5700_) );
OR2X2 OR2X2_424 ( .A(_5696_), .B(_5700_), .Y(_5701_) );
AND2X2 AND2X2_463 ( .A(_5701_), .B(ULA_B_3_bF_buf4), .Y(_5702_) );
OR2X2 OR2X2_425 ( .A(_5692_), .B(_5702_), .Y(_5703_) );
INVX1 INVX1_8 ( .A(CORE_ULA_ctrl_3_), .Y(_5704_) );
NOR3X1 NOR3X1_1 ( .A(_5704_), .B(CORE_ULA_ctrl_2_), .C(_5674_), .Y(_5705_) );
NAND2X1 NAND2X1_643 ( .A(ULA_B_4_bF_buf1), .B(_5705_), .Y(_5706_) );
OR2X2 OR2X2_426 ( .A(_5706_), .B(_5703_), .Y(_5707_) );
MUX2X1 MUX2X1_649 ( .A(ULA_A_9_), .B(ULA_A_8_), .S(ULA_B_0_bF_buf0), .Y(_5708_) );
AND2X2 AND2X2_464 ( .A(_5708_), .B(_5682__bF_buf4), .Y(_5709_) );
MUX2X1 MUX2X1_650 ( .A(ULA_A_11_), .B(ULA_A_10_), .S(ULA_B_0_bF_buf0), .Y(_5710_) );
AND2X2 AND2X2_465 ( .A(_5710_), .B(ULA_B_1_bF_buf2), .Y(_5711_) );
OR2X2 OR2X2_427 ( .A(_5709_), .B(_5711_), .Y(_5712_) );
AND2X2 AND2X2_466 ( .A(_5712_), .B(_5681__bF_buf5), .Y(_5713_) );
MUX2X1 MUX2X1_651 ( .A(ULA_A_13_), .B(ULA_A_12_), .S(ULA_B_0_bF_buf0), .Y(_5714_) );
AND2X2 AND2X2_467 ( .A(_5714_), .B(_5682__bF_buf4), .Y(_5715_) );
MUX2X1 MUX2X1_652 ( .A(ULA_A_15_), .B(ULA_A_14_), .S(ULA_B_0_bF_buf7), .Y(_5716_) );
AND2X2 AND2X2_468 ( .A(_5716_), .B(ULA_B_1_bF_buf2), .Y(_5717_) );
OR2X2 OR2X2_428 ( .A(_5715_), .B(_5717_), .Y(_5718_) );
AND2X2 AND2X2_469 ( .A(_5718_), .B(ULA_B_2_bF_buf0), .Y(_5719_) );
OR2X2 OR2X2_429 ( .A(_5713_), .B(_5719_), .Y(_5720_) );
AND2X2 AND2X2_470 ( .A(_5720_), .B(ULA_B_3_bF_buf0), .Y(_5721_) );
MUX2X1 MUX2X1_653 ( .A(ULA_A_3_), .B(ULA_A_2_), .S(ULA_B_0_bF_buf5), .Y(_5722_) );
MUX2X1 MUX2X1_654 ( .A(ULA_A_1_), .B(ULA_A_0_), .S(ULA_B_0_bF_buf5), .Y(_5723_) );
MUX2X1 MUX2X1_655 ( .A(_5723_), .B(_5722_), .S(_5682__bF_buf4), .Y(_5724_) );
MUX2X1 MUX2X1_656 ( .A(ULA_A_7_), .B(ULA_A_6_), .S(ULA_B_0_bF_buf7), .Y(_5725_) );
MUX2X1 MUX2X1_657 ( .A(ULA_A_5_), .B(ULA_A_4_), .S(ULA_B_0_bF_buf0), .Y(_5726_) );
MUX2X1 MUX2X1_658 ( .A(_5726_), .B(_5725_), .S(_5682__bF_buf4), .Y(_5727_) );
MUX2X1 MUX2X1_659 ( .A(_5727_), .B(_5724_), .S(ULA_B_2_bF_buf0), .Y(_5728_) );
AND2X2 AND2X2_471 ( .A(_5728_), .B(_5289__bF_buf5), .Y(_5729_) );
NAND2X1 NAND2X1_644 ( .A(_5669__bF_buf0), .B(_5705_), .Y(_5730_) );
OR2X2 OR2X2_430 ( .A(_5730__bF_buf1), .B(_5729_), .Y(_5731_) );
OR2X2 OR2X2_431 ( .A(_5721_), .B(_5731_), .Y(_5732_) );
OR2X2 OR2X2_432 ( .A(ULA_A_0_), .B(ULA_B_0_bF_buf6), .Y(_5733_) );
NOR3X1 NOR3X1_2 ( .A(_5673_), .B(CORE_ULA_ctrl_3_), .C(CORE_ULA_ctrl_1_), .Y(_5734_) );
AND2X2 AND2X2_472 ( .A(_5704_), .B(_5676_), .Y(_5735_) );
NAND2X1 NAND2X1_645 ( .A(ULA_A_0_), .B(ULA_B_0_bF_buf6), .Y(_5736_) );
AND2X2 AND2X2_473 ( .A(_5735__bF_buf4), .B(_5736_), .Y(_5737_) );
OAI21X1 OAI21X1_1 ( .A(_5737_), .B(_5734__bF_buf2), .C(_5733_), .Y(_5738_) );
NAND3X1 NAND3X1_12 ( .A(_5704_), .B(_5673_), .C(_5674_), .Y(_5739_) );
NOR3X1 NOR3X1_3 ( .A(_5674_), .B(CORE_ULA_ctrl_3_), .C(CORE_ULA_ctrl_2_), .Y(_5740_) );
XOR2X1 XOR2X1_6 ( .A(_5438__bF_buf2), .B(_5736_), .Y(_5741_) );
NAND2X1 NAND2X1_646 ( .A(_5741_), .B(_5740__bF_buf3), .Y(_5742_) );
AND2X2 AND2X2_474 ( .A(_5742_), .B(_5739__bF_buf2), .Y(_5743_) );
AND2X2 AND2X2_475 ( .A(_5743_), .B(_5738_), .Y(_5744_) );
INVX1 INVX1_9 ( .A(_5670_), .Y(_5745_) );
NAND3X1 NAND3X1_13 ( .A(_5674_), .B(CORE_ULA_ctrl_3_), .C(CORE_ULA_ctrl_2_), .Y(_5746_) );
NOR2X1 NOR2X1_18 ( .A(_5746_), .B(ULA_B_4_bF_buf3), .Y(_5747_) );
NAND3X1 NAND3X1_14 ( .A(_5747_), .B(ULA_A_0_), .C(_5745_), .Y(_5748_) );
AND2X2 AND2X2_476 ( .A(_5748_), .B(_5744_), .Y(_5749_) );
AND2X2 AND2X2_477 ( .A(_5732_), .B(_5749_), .Y(_5750_) );
AND2X2 AND2X2_478 ( .A(_5750_), .B(_5707_), .Y(_5751_) );
MUX2X1 MUX2X1_660 ( .A(_5714_), .B(_5716_), .S(_5417__bF_buf5), .Y(_5752_) );
MUX2X1 MUX2X1_661 ( .A(_5708_), .B(_5710_), .S(_5417__bF_buf5), .Y(_5753_) );
MUX2X1 MUX2X1_662 ( .A(_5753_), .B(_5752_), .S(_5353__bF_buf0), .Y(_5754_) );
AND2X2 AND2X2_479 ( .A(_5754_), .B(_5332__bF_buf3), .Y(_5755_) );
MUX2X1 MUX2X1_663 ( .A(_5723_), .B(_5722_), .S(_5417__bF_buf1), .Y(_5756_) );
MUX2X1 MUX2X1_664 ( .A(_5726_), .B(_5725_), .S(_5417__bF_buf1), .Y(_5757_) );
MUX2X1 MUX2X1_665 ( .A(_5757_), .B(_5756_), .S(_5524__bF_buf2), .Y(_5758_) );
AND2X2 AND2X2_480 ( .A(_5758_), .B(_5620__bF_buf3), .Y(_5759_) );
XOR2X1 XOR2X1_7 ( .A(ULA_B_4_bF_buf2), .B(_5671_), .Y(_5760_) );
OR2X2 OR2X2_433 ( .A(_5760_), .B(_5678_), .Y(_5761_) );
OR2X2 OR2X2_434 ( .A(_5761_), .B(_5759_), .Y(_5762_) );
OR2X2 OR2X2_435 ( .A(_5755_), .B(_5762_), .Y(_5763_) );
AND2X2 AND2X2_481 ( .A(_5751_), .B(_5763_), .Y(_5764_) );
AND2X2 AND2X2_482 ( .A(_5764_), .B(_5680_), .Y(_5765_) );
NOR2X1 NOR2X1_19 ( .A(_5739__bF_buf1), .B(ULA_OUT_0__0_), .Y(_5766_) );
OR2X2 OR2X2_436 ( .A(_5766_), .B(_5765_), .Y(_5767_) );
INVX1 INVX1_10 ( .A(_5767_), .Y(ULA_ULA_OUT_0_) );
NOR2X1 NOR2X1_20 ( .A(_5739__bF_buf5), .B(ULA_OUT_0__1_), .Y(_5768_) );
MUX2X1 MUX2X1_666 ( .A(ULA_A_18_), .B(ULA_A_17_), .S(ULA_B_0_bF_buf3), .Y(_5769_) );
AND2X2 AND2X2_483 ( .A(_5769_), .B(_5682__bF_buf2), .Y(_5770_) );
MUX2X1 MUX2X1_667 ( .A(ULA_A_20_), .B(ULA_A_19_), .S(ULA_B_0_bF_buf1), .Y(_5771_) );
AND2X2 AND2X2_484 ( .A(_5771_), .B(ULA_B_1_bF_buf6), .Y(_5772_) );
OR2X2 OR2X2_437 ( .A(_5770_), .B(_5772_), .Y(_5773_) );
AND2X2 AND2X2_485 ( .A(_5773_), .B(_5681__bF_buf4), .Y(_5774_) );
MUX2X1 MUX2X1_668 ( .A(ULA_A_22_), .B(ULA_A_21_), .S(ULA_B_0_bF_buf7), .Y(_5775_) );
AND2X2 AND2X2_486 ( .A(_5775_), .B(_5682__bF_buf5), .Y(_5776_) );
MUX2X1 MUX2X1_669 ( .A(ULA_A_24_), .B(ULA_A_23_), .S(ULA_B_0_bF_buf7), .Y(_5777_) );
AND2X2 AND2X2_487 ( .A(_5777_), .B(ULA_B_1_bF_buf5), .Y(_5778_) );
OR2X2 OR2X2_438 ( .A(_5776_), .B(_5778_), .Y(_5779_) );
AND2X2 AND2X2_488 ( .A(_5779_), .B(ULA_B_2_bF_buf3), .Y(_5780_) );
OR2X2 OR2X2_439 ( .A(_5774_), .B(_5780_), .Y(_5781_) );
AND2X2 AND2X2_489 ( .A(_5781_), .B(_5289__bF_buf1), .Y(_5782_) );
MUX2X1 MUX2X1_670 ( .A(ULA_A_26_), .B(ULA_A_25_), .S(ULA_B_0_bF_buf7), .Y(_5783_) );
AND2X2 AND2X2_490 ( .A(_5783_), .B(_5682__bF_buf5), .Y(_5784_) );
MUX2X1 MUX2X1_671 ( .A(ULA_A_28_), .B(ULA_A_27_), .S(ULA_B_0_bF_buf5), .Y(_5785_) );
AND2X2 AND2X2_491 ( .A(_5785_), .B(ULA_B_1_bF_buf5), .Y(_5786_) );
OR2X2 OR2X2_440 ( .A(_5784_), .B(_5786_), .Y(_5787_) );
AND2X2 AND2X2_492 ( .A(_5787_), .B(_5681__bF_buf2), .Y(_5788_) );
INVX1 INVX1_11 ( .A(ULA_B_0_bF_buf6), .Y(_5789_) );
NAND3X1 NAND3X1_15 ( .A(_5789_), .B(ULA_B_1_bF_buf4), .C(ULA_A_31_), .Y(_5790_) );
MUX2X1 MUX2X1_672 ( .A(ULA_A_30_), .B(ULA_A_29_), .S(ULA_B_0_bF_buf1), .Y(_5791_) );
OR2X2 OR2X2_441 ( .A(ULA_B_1_bF_buf1), .B(_5791_), .Y(_5792_) );
AND2X2 AND2X2_493 ( .A(_5790_), .B(_5792_), .Y(_5793_) );
AND2X2 AND2X2_494 ( .A(_5793_), .B(ULA_B_2_bF_buf4), .Y(_5794_) );
OR2X2 OR2X2_442 ( .A(_5788_), .B(_5794_), .Y(_5795_) );
AND2X2 AND2X2_495 ( .A(_5795_), .B(ULA_B_3_bF_buf3), .Y(_5796_) );
OR2X2 OR2X2_443 ( .A(_5782_), .B(_5796_), .Y(_5797_) );
AND2X2 AND2X2_496 ( .A(_5797_), .B(ULA_B_4_bF_buf0), .Y(_5798_) );
NAND3X1 NAND3X1_16 ( .A(_5673_), .B(CORE_ULA_ctrl_3_), .C(CORE_ULA_ctrl_1_), .Y(_5799_) );
MUX2X1 MUX2X1_673 ( .A(ULA_A_2_), .B(ULA_A_1_), .S(ULA_B_0_bF_buf1), .Y(_5800_) );
OR2X2 OR2X2_444 ( .A(ULA_B_1_bF_buf5), .B(_5800_), .Y(_5801_) );
MUX2X1 MUX2X1_674 ( .A(ULA_A_4_), .B(ULA_A_3_), .S(ULA_B_0_bF_buf0), .Y(_5802_) );
OR2X2 OR2X2_445 ( .A(_5682__bF_buf2), .B(_5802_), .Y(_5803_) );
AND2X2 AND2X2_497 ( .A(_5803_), .B(_5681__bF_buf4), .Y(_5804_) );
AND2X2 AND2X2_498 ( .A(_5804_), .B(_5801_), .Y(_5805_) );
MUX2X1 MUX2X1_675 ( .A(ULA_A_6_), .B(ULA_A_5_), .S(ULA_B_0_bF_buf0), .Y(_5806_) );
AND2X2 AND2X2_499 ( .A(_5806_), .B(_5682__bF_buf2), .Y(_5807_) );
MUX2X1 MUX2X1_676 ( .A(ULA_A_8_), .B(ULA_A_7_), .S(ULA_B_0_bF_buf0), .Y(_5808_) );
AND2X2 AND2X2_500 ( .A(_5808_), .B(ULA_B_1_bF_buf6), .Y(_5809_) );
OR2X2 OR2X2_446 ( .A(_5807_), .B(_5809_), .Y(_5810_) );
AND2X2 AND2X2_501 ( .A(_5810_), .B(ULA_B_2_bF_buf3), .Y(_5811_) );
OR2X2 OR2X2_447 ( .A(_5805_), .B(_5811_), .Y(_5812_) );
AND2X2 AND2X2_502 ( .A(_5812_), .B(_5289__bF_buf0), .Y(_5813_) );
MUX2X1 MUX2X1_677 ( .A(ULA_A_10_), .B(ULA_A_9_), .S(ULA_B_0_bF_buf0), .Y(_5814_) );
AND2X2 AND2X2_503 ( .A(_5814_), .B(_5682__bF_buf2), .Y(_5815_) );
MUX2X1 MUX2X1_678 ( .A(ULA_A_12_), .B(ULA_A_11_), .S(ULA_B_0_bF_buf3), .Y(_5816_) );
AND2X2 AND2X2_504 ( .A(_5816_), .B(ULA_B_1_bF_buf6), .Y(_5817_) );
OR2X2 OR2X2_448 ( .A(_5815_), .B(_5817_), .Y(_5818_) );
AND2X2 AND2X2_505 ( .A(_5818_), .B(_5681__bF_buf4), .Y(_5819_) );
MUX2X1 MUX2X1_679 ( .A(ULA_A_14_), .B(ULA_A_13_), .S(ULA_B_0_bF_buf3), .Y(_5820_) );
AND2X2 AND2X2_506 ( .A(_5820_), .B(_5682__bF_buf2), .Y(_5821_) );
MUX2X1 MUX2X1_680 ( .A(ULA_A_16_), .B(ULA_A_15_), .S(ULA_B_0_bF_buf3), .Y(_5822_) );
AND2X2 AND2X2_507 ( .A(_5822_), .B(ULA_B_1_bF_buf6), .Y(_5823_) );
OR2X2 OR2X2_449 ( .A(_5821_), .B(_5823_), .Y(_5824_) );
AND2X2 AND2X2_508 ( .A(_5824_), .B(ULA_B_2_bF_buf3), .Y(_5825_) );
OR2X2 OR2X2_450 ( .A(_5819_), .B(_5825_), .Y(_5826_) );
AND2X2 AND2X2_509 ( .A(_5826_), .B(ULA_B_3_bF_buf7), .Y(_5827_) );
OR2X2 OR2X2_451 ( .A(_5813_), .B(_5827_), .Y(_5828_) );
AND2X2 AND2X2_510 ( .A(_5828_), .B(_5669__bF_buf2), .Y(_5829_) );
OR2X2 OR2X2_452 ( .A(_5799_), .B(_5829_), .Y(_5830_) );
OR2X2 OR2X2_453 ( .A(_5798_), .B(_5830_), .Y(_5831_) );
NOR2X1 NOR2X1_21 ( .A(ULA_A_1_), .B(ULA_B_1_bF_buf7), .Y(_5832_) );
NAND2X1 NAND2X1_647 ( .A(ULA_A_1_), .B(ULA_B_1_bF_buf7), .Y(_5833_) );
AOI21X1 AOI21X1_1 ( .A(_5833_), .B(_5735__bF_buf2), .C(_5734__bF_buf4), .Y(_5834_) );
OR2X2 OR2X2_454 ( .A(_5832_), .B(_5834_), .Y(_5835_) );
NAND2X1 NAND2X1_648 ( .A(_5438__bF_buf3), .B(_5833_), .Y(_5836_) );
NAND3X1 NAND3X1_17 ( .A(ULA_A_1_), .B(ULA_cin_bF_buf3), .C(ULA_B_1_bF_buf7), .Y(_5837_) );
NAND3X1 NAND3X1_18 ( .A(_5836_), .B(_5740__bF_buf2), .C(_5837_), .Y(_5838_) );
AND2X2 AND2X2_511 ( .A(_5838_), .B(_5739__bF_buf5), .Y(_5839_) );
AND2X2 AND2X2_512 ( .A(_5835_), .B(_5839_), .Y(_5840_) );
MUX2X1 MUX2X1_681 ( .A(ULA_A_0_), .B(ULA_A_1_), .S(ULA_B_0_bF_buf1), .Y(_5841_) );
OR2X2 OR2X2_455 ( .A(ULA_B_1_bF_buf4), .B(_5841_), .Y(_5842_) );
OR2X2 OR2X2_456 ( .A(ULA_B_2_bF_buf6), .B(_5842_), .Y(_5843_) );
INVX1 INVX1_12 ( .A(_5843_), .Y(_5844_) );
NAND2X1 NAND2X1_649 ( .A(CORE_ULA_ctrl_3_), .B(CORE_ULA_ctrl_2_), .Y(_5845_) );
NOR2X1 NOR2X1_22 ( .A(_5845_), .B(ULA_B_4_bF_buf1), .Y(_5846_) );
NAND3X1 NAND3X1_19 ( .A(_5844_), .B(_5289__bF_buf3), .C(_5846_), .Y(_5847_) );
AND2X2 AND2X2_513 ( .A(_5840_), .B(_5847_), .Y(_5848_) );
AND2X2 AND2X2_514 ( .A(_5831_), .B(_5848_), .Y(_5849_) );
OR2X2 OR2X2_457 ( .A(_5791_), .B(_5470__bF_buf1), .Y(_5850_) );
AND2X2 AND2X2_515 ( .A(_5850_), .B(_5790_), .Y(_5851_) );
AND2X2 AND2X2_516 ( .A(_5851_), .B(_5524__bF_buf2), .Y(_5852_) );
AND2X2 AND2X2_517 ( .A(_5417__bF_buf1), .B(_5783_), .Y(_5853_) );
AND2X2 AND2X2_518 ( .A(_5470__bF_buf1), .B(_5785_), .Y(_5854_) );
OR2X2 OR2X2_458 ( .A(_5853_), .B(_5854_), .Y(_5855_) );
AND2X2 AND2X2_519 ( .A(_5855_), .B(_5353__bF_buf0), .Y(_5856_) );
OR2X2 OR2X2_459 ( .A(_5852_), .B(_5856_), .Y(_5857_) );
AND2X2 AND2X2_520 ( .A(_5857_), .B(_5332__bF_buf2), .Y(_5858_) );
MUX2X1 MUX2X1_682 ( .A(_5775_), .B(_5777_), .S(_5417__bF_buf5), .Y(_5859_) );
MUX2X1 MUX2X1_683 ( .A(_5769_), .B(_5771_), .S(_5417__bF_buf4), .Y(_5860_) );
MUX2X1 MUX2X1_684 ( .A(_5860_), .B(_5859_), .S(_5353__bF_buf4), .Y(_5861_) );
AND2X2 AND2X2_521 ( .A(_5861_), .B(_5620__bF_buf2), .Y(_5862_) );
OR2X2 OR2X2_460 ( .A(_5858_), .B(_5862_), .Y(_5863_) );
OR2X2 OR2X2_461 ( .A(_5679_), .B(_5863_), .Y(_5864_) );
AND2X2 AND2X2_522 ( .A(_5417__bF_buf1), .B(_5806_), .Y(_5865_) );
AND2X2 AND2X2_523 ( .A(_5470__bF_buf1), .B(_5808_), .Y(_5866_) );
OR2X2 OR2X2_462 ( .A(_5865_), .B(_5866_), .Y(_5867_) );
OR2X2 OR2X2_463 ( .A(_5353__bF_buf4), .B(_5867_), .Y(_5868_) );
AND2X2 AND2X2_524 ( .A(_5470__bF_buf1), .B(_5802_), .Y(_5869_) );
AND2X2 AND2X2_525 ( .A(_5417__bF_buf4), .B(_5800_), .Y(_5870_) );
OR2X2 OR2X2_464 ( .A(_5524__bF_buf2), .B(_5870_), .Y(_5871_) );
OR2X2 OR2X2_465 ( .A(_5869_), .B(_5871_), .Y(_5872_) );
AND2X2 AND2X2_526 ( .A(_5872_), .B(_5620__bF_buf1), .Y(_5873_) );
AND2X2 AND2X2_527 ( .A(_5873_), .B(_5868_), .Y(_5874_) );
AND2X2 AND2X2_528 ( .A(_5417__bF_buf0), .B(_5820_), .Y(_5875_) );
AND2X2 AND2X2_529 ( .A(_5470__bF_buf2), .B(_5822_), .Y(_5876_) );
OR2X2 OR2X2_466 ( .A(_5875_), .B(_5876_), .Y(_5877_) );
AND2X2 AND2X2_530 ( .A(_5877_), .B(_5524__bF_buf1), .Y(_5878_) );
AND2X2 AND2X2_531 ( .A(_5417__bF_buf4), .B(_5814_), .Y(_5879_) );
AND2X2 AND2X2_532 ( .A(_5470__bF_buf2), .B(_5816_), .Y(_5880_) );
OR2X2 OR2X2_467 ( .A(_5879_), .B(_5880_), .Y(_5881_) );
AND2X2 AND2X2_533 ( .A(_5881_), .B(_5353__bF_buf4), .Y(_5882_) );
OR2X2 OR2X2_468 ( .A(_5878_), .B(_5882_), .Y(_5883_) );
AND2X2 AND2X2_534 ( .A(_5883_), .B(_5332__bF_buf2), .Y(_5884_) );
OR2X2 OR2X2_469 ( .A(_5874_), .B(_5884_), .Y(_5885_) );
OR2X2 OR2X2_470 ( .A(_5761_), .B(_5885_), .Y(_5886_) );
AND2X2 AND2X2_535 ( .A(_5864_), .B(_5886_), .Y(_5887_) );
AND2X2 AND2X2_536 ( .A(_5887_), .B(_5849_), .Y(_5888_) );
OR2X2 OR2X2_471 ( .A(_5768_), .B(_5888_), .Y(_5889_) );
INVX1 INVX1_13 ( .A(_5889_), .Y(ULA_ULA_OUT_1_) );
NOR2X1 NOR2X1_23 ( .A(_5739__bF_buf5), .B(ULA_OUT_0__2_), .Y(_5890_) );
AND2X2 AND2X2_537 ( .A(_5710_), .B(_5682__bF_buf4), .Y(_5891_) );
AND2X2 AND2X2_538 ( .A(_5714_), .B(ULA_B_1_bF_buf2), .Y(_5892_) );
OR2X2 OR2X2_472 ( .A(_5891_), .B(_5892_), .Y(_5893_) );
AND2X2 AND2X2_539 ( .A(_5893_), .B(_5681__bF_buf5), .Y(_5894_) );
AND2X2 AND2X2_540 ( .A(_5716_), .B(_5682__bF_buf1), .Y(_5895_) );
AND2X2 AND2X2_541 ( .A(_5660_), .B(ULA_B_1_bF_buf2), .Y(_5896_) );
OR2X2 OR2X2_473 ( .A(_5895_), .B(_5896_), .Y(_5897_) );
AND2X2 AND2X2_542 ( .A(_5897_), .B(ULA_B_2_bF_buf0), .Y(_5898_) );
OR2X2 OR2X2_474 ( .A(_5894_), .B(_5898_), .Y(_5899_) );
AND2X2 AND2X2_543 ( .A(_5899_), .B(ULA_B_3_bF_buf5), .Y(_5900_) );
AND2X2 AND2X2_544 ( .A(_5722_), .B(_5682__bF_buf4), .Y(_5901_) );
AND2X2 AND2X2_545 ( .A(_5726_), .B(ULA_B_1_bF_buf5), .Y(_5902_) );
OR2X2 OR2X2_475 ( .A(_5901_), .B(_5902_), .Y(_5903_) );
AND2X2 AND2X2_546 ( .A(_5903_), .B(_5681__bF_buf5), .Y(_5904_) );
AND2X2 AND2X2_547 ( .A(_5708_), .B(ULA_B_1_bF_buf2), .Y(_5905_) );
AND2X2 AND2X2_548 ( .A(_5725_), .B(_5682__bF_buf4), .Y(_5906_) );
OR2X2 OR2X2_476 ( .A(_5905_), .B(_5906_), .Y(_5907_) );
AND2X2 AND2X2_549 ( .A(_5907_), .B(ULA_B_2_bF_buf0), .Y(_5908_) );
OR2X2 OR2X2_477 ( .A(_5904_), .B(_5908_), .Y(_5909_) );
AND2X2 AND2X2_550 ( .A(_5909_), .B(_5289__bF_buf5), .Y(_5910_) );
OR2X2 OR2X2_478 ( .A(_5730__bF_buf1), .B(_5910_), .Y(_5911_) );
OR2X2 OR2X2_479 ( .A(_5900_), .B(_5911_), .Y(_5912_) );
AND2X2 AND2X2_551 ( .A(_5662_), .B(_5682__bF_buf1), .Y(_5913_) );
AND2X2 AND2X2_552 ( .A(_5630_), .B(ULA_B_1_bF_buf2), .Y(_5914_) );
OR2X2 OR2X2_480 ( .A(_5913_), .B(_5914_), .Y(_5915_) );
AND2X2 AND2X2_553 ( .A(_5915_), .B(_5681__bF_buf6), .Y(_5916_) );
AND2X2 AND2X2_554 ( .A(_5364_), .B(ULA_B_1_bF_buf3), .Y(_5917_) );
AND2X2 AND2X2_555 ( .A(_5652_), .B(_5682__bF_buf3), .Y(_5918_) );
OR2X2 OR2X2_481 ( .A(_5917_), .B(_5918_), .Y(_5919_) );
AND2X2 AND2X2_556 ( .A(_5919_), .B(ULA_B_2_bF_buf5), .Y(_5920_) );
OR2X2 OR2X2_482 ( .A(_5916_), .B(_5920_), .Y(_5921_) );
AND2X2 AND2X2_557 ( .A(_5921_), .B(_5289__bF_buf2), .Y(_5922_) );
OR2X2 OR2X2_483 ( .A(ULA_B_1_bF_buf0), .B(_5534_), .Y(_5923_) );
AND2X2 AND2X2_558 ( .A(_5923_), .B(ULA_B_2_bF_buf5), .Y(_5924_) );
AND2X2 AND2X2_559 ( .A(_5556_), .B(ULA_B_1_bF_buf0), .Y(_5925_) );
AND2X2 AND2X2_560 ( .A(_5481_), .B(_5682__bF_buf3), .Y(_5926_) );
OR2X2 OR2X2_484 ( .A(_5925_), .B(_5926_), .Y(_5927_) );
AND2X2 AND2X2_561 ( .A(_5927_), .B(_5681__bF_buf6), .Y(_5928_) );
OR2X2 OR2X2_485 ( .A(_5924_), .B(_5928_), .Y(_5929_) );
AND2X2 AND2X2_562 ( .A(_5929_), .B(ULA_B_3_bF_buf4), .Y(_5930_) );
OR2X2 OR2X2_486 ( .A(_5930_), .B(_5922_), .Y(_5931_) );
OR2X2 OR2X2_487 ( .A(_5706_), .B(_5931_), .Y(_5932_) );
NAND3X1 NAND3X1_20 ( .A(_5704_), .B(CORE_ULA_ctrl_2_), .C(_5674_), .Y(_5933_) );
OR2X2 OR2X2_488 ( .A(ULA_A_2_), .B(ULA_B_2_bF_buf6), .Y(_5934_) );
INVX1 INVX1_14 ( .A(_5934_), .Y(_5935_) );
OR2X2 OR2X2_489 ( .A(_5935_), .B(_5933_), .Y(_5936_) );
NAND2X1 NAND2X1_650 ( .A(ULA_A_2_), .B(ULA_B_2_bF_buf6), .Y(_5937_) );
NAND3X1 NAND3X1_21 ( .A(_5735__bF_buf4), .B(_5934_), .C(_5937_), .Y(_5938_) );
AND2X2 AND2X2_563 ( .A(_5938_), .B(_5936_), .Y(_5939_) );
NAND3X1 NAND3X1_22 ( .A(_5704_), .B(CORE_ULA_ctrl_1_), .C(_5673_), .Y(_5940_) );
XOR2X1 XOR2X1_8 ( .A(ULA_cin_bF_buf6), .B(_5937_), .Y(_5941_) );
OR2X2 OR2X2_490 ( .A(_5941_), .B(_5940_), .Y(_5942_) );
AND2X2 AND2X2_564 ( .A(_5942_), .B(_5739__bF_buf2), .Y(_5943_) );
AND2X2 AND2X2_565 ( .A(_5939_), .B(_5943_), .Y(_5944_) );
INVX1 INVX1_15 ( .A(_5846_), .Y(_5945_) );
MUX2X1 MUX2X1_685 ( .A(ULA_A_1_), .B(ULA_A_2_), .S(ULA_B_0_bF_buf5), .Y(_5946_) );
OR2X2 OR2X2_491 ( .A(ULA_B_1_bF_buf0), .B(_5946_), .Y(_5947_) );
NAND3X1 NAND3X1_23 ( .A(_5789_), .B(ULA_A_0_), .C(ULA_B_1_bF_buf0), .Y(_5948_) );
AND2X2 AND2X2_566 ( .A(_5948_), .B(_5947_), .Y(_5949_) );
OR2X2 OR2X2_492 ( .A(ULA_B_2_bF_buf5), .B(_5949_), .Y(_5950_) );
OR2X2 OR2X2_493 ( .A(ULA_B_3_bF_buf6), .B(_5950_), .Y(_5951_) );
OR2X2 OR2X2_494 ( .A(_5945__bF_buf3), .B(_5951_), .Y(_5952_) );
AND2X2 AND2X2_567 ( .A(_5952_), .B(_5944_), .Y(_5953_) );
AND2X2 AND2X2_568 ( .A(_5932_), .B(_5953_), .Y(_5954_) );
AND2X2 AND2X2_569 ( .A(_5954_), .B(_5912_), .Y(_5955_) );
OR2X2 OR2X2_495 ( .A(_5534_), .B(_5470__bF_buf3), .Y(_5956_) );
AND2X2 AND2X2_570 ( .A(_5956_), .B(_5524__bF_buf3), .Y(_5957_) );
AND2X2 AND2X2_571 ( .A(_5417__bF_buf2), .B(_5481_), .Y(_5958_) );
AND2X2 AND2X2_572 ( .A(_5470__bF_buf3), .B(_5556_), .Y(_5959_) );
OR2X2 OR2X2_496 ( .A(_5958_), .B(_5959_), .Y(_5960_) );
AND2X2 AND2X2_573 ( .A(_5960_), .B(_5353__bF_buf3), .Y(_5961_) );
OR2X2 OR2X2_497 ( .A(_5957_), .B(_5961_), .Y(_5962_) );
AND2X2 AND2X2_574 ( .A(_5962_), .B(_5332__bF_buf0), .Y(_5963_) );
AND2X2 AND2X2_575 ( .A(_5417__bF_buf2), .B(_5652_), .Y(_5964_) );
AND2X2 AND2X2_576 ( .A(_5470__bF_buf3), .B(_5364_), .Y(_5965_) );
OR2X2 OR2X2_498 ( .A(_5964_), .B(_5965_), .Y(_5966_) );
AND2X2 AND2X2_577 ( .A(_5966_), .B(_5524__bF_buf3), .Y(_5967_) );
AND2X2 AND2X2_578 ( .A(_5417__bF_buf3), .B(_5662_), .Y(_5968_) );
AND2X2 AND2X2_579 ( .A(_5470__bF_buf0), .B(_5630_), .Y(_5969_) );
OR2X2 OR2X2_499 ( .A(_5968_), .B(_5969_), .Y(_5970_) );
AND2X2 AND2X2_580 ( .A(_5970_), .B(_5353__bF_buf3), .Y(_5971_) );
OR2X2 OR2X2_500 ( .A(_5967_), .B(_5971_), .Y(_5972_) );
AND2X2 AND2X2_581 ( .A(_5972_), .B(_5620__bF_buf0), .Y(_5973_) );
OR2X2 OR2X2_501 ( .A(_5963_), .B(_5973_), .Y(_5974_) );
OR2X2 OR2X2_502 ( .A(_5679_), .B(_5974_), .Y(_5975_) );
AND2X2 AND2X2_582 ( .A(_5470__bF_buf1), .B(_5726_), .Y(_5976_) );
AND2X2 AND2X2_583 ( .A(_5417__bF_buf5), .B(_5722_), .Y(_5977_) );
OR2X2 OR2X2_503 ( .A(_5524__bF_buf0), .B(_5977_), .Y(_5978_) );
OR2X2 OR2X2_504 ( .A(_5976_), .B(_5978_), .Y(_5979_) );
AND2X2 AND2X2_584 ( .A(_5417__bF_buf2), .B(_5725_), .Y(_5980_) );
AND2X2 AND2X2_585 ( .A(_5470__bF_buf0), .B(_5708_), .Y(_5981_) );
OR2X2 OR2X2_505 ( .A(_5980_), .B(_5981_), .Y(_5982_) );
OR2X2 OR2X2_506 ( .A(_5353__bF_buf1), .B(_5982_), .Y(_5983_) );
AND2X2 AND2X2_586 ( .A(_5983_), .B(_5979_), .Y(_5984_) );
OR2X2 OR2X2_507 ( .A(_5332__bF_buf3), .B(_5984_), .Y(_5985_) );
AND2X2 AND2X2_587 ( .A(_5417__bF_buf3), .B(_5716_), .Y(_5986_) );
AND2X2 AND2X2_588 ( .A(_5470__bF_buf0), .B(_5660_), .Y(_5987_) );
OR2X2 OR2X2_508 ( .A(_5986_), .B(_5987_), .Y(_5988_) );
AND2X2 AND2X2_589 ( .A(_5988_), .B(_5524__bF_buf0), .Y(_5989_) );
AND2X2 AND2X2_590 ( .A(_5417__bF_buf5), .B(_5710_), .Y(_5990_) );
AND2X2 AND2X2_591 ( .A(_5470__bF_buf0), .B(_5714_), .Y(_5991_) );
OR2X2 OR2X2_509 ( .A(_5990_), .B(_5991_), .Y(_5992_) );
AND2X2 AND2X2_592 ( .A(_5992_), .B(_5353__bF_buf1), .Y(_5993_) );
OR2X2 OR2X2_510 ( .A(_5989_), .B(_5993_), .Y(_5994_) );
OR2X2 OR2X2_511 ( .A(_5620__bF_buf0), .B(_5994_), .Y(_5995_) );
AND2X2 AND2X2_593 ( .A(_5985_), .B(_5995_), .Y(_5996_) );
OR2X2 OR2X2_512 ( .A(_5761_), .B(_5996_), .Y(_5997_) );
AND2X2 AND2X2_594 ( .A(_5997_), .B(_5975_), .Y(_5998_) );
AND2X2 AND2X2_595 ( .A(_5998_), .B(_5955_), .Y(_5999_) );
OR2X2 OR2X2_513 ( .A(_5890_), .B(_5999_), .Y(_6000_) );
INVX1 INVX1_16 ( .A(_6000_), .Y(ULA_ULA_OUT_2_) );
NOR2X1 NOR2X1_24 ( .A(_5739__bF_buf1), .B(ULA_OUT_0__3_), .Y(_6001_) );
NOR2X1 NOR2X1_25 ( .A(ULA_B_0_bF_buf1), .B(ULA_B_1_bF_buf4), .Y(_6002_) );
NAND3X1 NAND3X1_24 ( .A(_6002_), .B(ULA_B_2_bF_buf1), .C(ULA_A_31_), .Y(_6003_) );
AND2X2 AND2X2_596 ( .A(_5417__bF_buf1), .B(_5785_), .Y(_6004_) );
AND2X2 AND2X2_597 ( .A(_5470__bF_buf1), .B(_5791_), .Y(_6005_) );
OR2X2 OR2X2_514 ( .A(_6004_), .B(_6005_), .Y(_6006_) );
OR2X2 OR2X2_515 ( .A(_5524__bF_buf2), .B(_6006_), .Y(_6007_) );
AND2X2 AND2X2_598 ( .A(_6007_), .B(_6003_), .Y(_6008_) );
AND2X2 AND2X2_599 ( .A(_6008_), .B(_5332__bF_buf1), .Y(_6009_) );
AND2X2 AND2X2_600 ( .A(_5417__bF_buf0), .B(_5777_), .Y(_6010_) );
AND2X2 AND2X2_601 ( .A(_5470__bF_buf2), .B(_5783_), .Y(_6011_) );
OR2X2 OR2X2_516 ( .A(_6010_), .B(_6011_), .Y(_6012_) );
AND2X2 AND2X2_602 ( .A(_6012_), .B(_5524__bF_buf1), .Y(_6013_) );
AND2X2 AND2X2_603 ( .A(_5417__bF_buf4), .B(_5771_), .Y(_6014_) );
AND2X2 AND2X2_604 ( .A(_5470__bF_buf2), .B(_5775_), .Y(_6015_) );
OR2X2 OR2X2_517 ( .A(_6014_), .B(_6015_), .Y(_6016_) );
AND2X2 AND2X2_605 ( .A(_6016_), .B(_5353__bF_buf2), .Y(_6017_) );
OR2X2 OR2X2_518 ( .A(_6013_), .B(_6017_), .Y(_6018_) );
AND2X2 AND2X2_606 ( .A(_6018_), .B(_5620__bF_buf2), .Y(_6019_) );
OR2X2 OR2X2_519 ( .A(_6009_), .B(_6019_), .Y(_6020_) );
OR2X2 OR2X2_520 ( .A(_5679_), .B(_6020_), .Y(_6021_) );
AND2X2 AND2X2_607 ( .A(_5841_), .B(ULA_B_1_bF_buf4), .Y(_6022_) );
MUX2X1 MUX2X1_686 ( .A(ULA_A_2_), .B(ULA_A_3_), .S(ULA_B_0_bF_buf1), .Y(_6023_) );
AND2X2 AND2X2_608 ( .A(_6023_), .B(_5682__bF_buf6), .Y(_6024_) );
OR2X2 OR2X2_521 ( .A(_6022_), .B(_6024_), .Y(_6025_) );
NOR3X1 NOR3X1_4 ( .A(_6025_), .B(ULA_B_2_bF_buf6), .C(ULA_B_3_bF_buf0), .Y(_6026_) );
NAND2X1 NAND2X1_651 ( .A(_5846_), .B(_6026_), .Y(_6027_) );
NOR2X1 NOR2X1_26 ( .A(ULA_A_3_), .B(ULA_B_3_bF_buf6), .Y(_6028_) );
NAND2X1 NAND2X1_652 ( .A(ULA_A_3_), .B(ULA_B_3_bF_buf6), .Y(_6029_) );
AOI21X1 AOI21X1_2 ( .A(_6029_), .B(_5735__bF_buf2), .C(_5734__bF_buf4), .Y(_6030_) );
OR2X2 OR2X2_522 ( .A(_6028_), .B(_6030_), .Y(_6031_) );
NAND3X1 NAND3X1_25 ( .A(ULA_cin_bF_buf3), .B(ULA_A_3_), .C(ULA_B_3_bF_buf6), .Y(_6032_) );
NAND2X1 NAND2X1_653 ( .A(_5438__bF_buf3), .B(_6029_), .Y(_6033_) );
NAND3X1 NAND3X1_26 ( .A(_6033_), .B(_5740__bF_buf2), .C(_6032_), .Y(_6034_) );
AND2X2 AND2X2_609 ( .A(_6034_), .B(_5739__bF_buf1), .Y(_6035_) );
AND2X2 AND2X2_610 ( .A(_6031_), .B(_6035_), .Y(_6036_) );
AND2X2 AND2X2_611 ( .A(_6027_), .B(_6036_), .Y(_6037_) );
AND2X2 AND2X2_612 ( .A(_6037_), .B(_6021_), .Y(_6038_) );
AND2X2 AND2X2_613 ( .A(_5771_), .B(_5682__bF_buf2), .Y(_6039_) );
AND2X2 AND2X2_614 ( .A(_5775_), .B(ULA_B_1_bF_buf5), .Y(_6040_) );
OR2X2 OR2X2_523 ( .A(_6039_), .B(_6040_), .Y(_6041_) );
AND2X2 AND2X2_615 ( .A(_6041_), .B(_5681__bF_buf2), .Y(_6042_) );
AND2X2 AND2X2_616 ( .A(_5777_), .B(_5682__bF_buf5), .Y(_6043_) );
AND2X2 AND2X2_617 ( .A(_5783_), .B(ULA_B_1_bF_buf5), .Y(_6044_) );
OR2X2 OR2X2_524 ( .A(_6043_), .B(_6044_), .Y(_6045_) );
AND2X2 AND2X2_618 ( .A(_6045_), .B(ULA_B_2_bF_buf2), .Y(_6046_) );
OR2X2 OR2X2_525 ( .A(_6042_), .B(_6046_), .Y(_6047_) );
AND2X2 AND2X2_619 ( .A(_6047_), .B(_5289__bF_buf0), .Y(_6048_) );
AND2X2 AND2X2_620 ( .A(_5785_), .B(_5682__bF_buf5), .Y(_6049_) );
AND2X2 AND2X2_621 ( .A(_5791_), .B(ULA_B_1_bF_buf1), .Y(_6050_) );
OR2X2 OR2X2_526 ( .A(_6049_), .B(_6050_), .Y(_6051_) );
OR2X2 OR2X2_527 ( .A(ULA_B_2_bF_buf6), .B(_6051_), .Y(_6052_) );
AND2X2 AND2X2_622 ( .A(_6052_), .B(_6003_), .Y(_6053_) );
AND2X2 AND2X2_623 ( .A(_6053_), .B(ULA_B_3_bF_buf1), .Y(_6054_) );
OR2X2 OR2X2_528 ( .A(_6048_), .B(_6054_), .Y(_6055_) );
AND2X2 AND2X2_624 ( .A(_6055_), .B(ULA_B_4_bF_buf2), .Y(_6056_) );
OR2X2 OR2X2_529 ( .A(ULA_B_1_bF_buf6), .B(_5802_), .Y(_6057_) );
OR2X2 OR2X2_530 ( .A(_5682__bF_buf2), .B(_5806_), .Y(_6058_) );
AND2X2 AND2X2_625 ( .A(_6058_), .B(_5681__bF_buf4), .Y(_6059_) );
AND2X2 AND2X2_626 ( .A(_6059_), .B(_6057_), .Y(_6060_) );
AND2X2 AND2X2_627 ( .A(_5808_), .B(_5682__bF_buf2), .Y(_6061_) );
AND2X2 AND2X2_628 ( .A(_5814_), .B(ULA_B_1_bF_buf6), .Y(_6062_) );
OR2X2 OR2X2_531 ( .A(_6061_), .B(_6062_), .Y(_6063_) );
AND2X2 AND2X2_629 ( .A(_6063_), .B(ULA_B_2_bF_buf3), .Y(_6064_) );
OR2X2 OR2X2_532 ( .A(_6060_), .B(_6064_), .Y(_6065_) );
AND2X2 AND2X2_630 ( .A(_6065_), .B(_5289__bF_buf5), .Y(_6066_) );
AND2X2 AND2X2_631 ( .A(_5816_), .B(_5682__bF_buf2), .Y(_6067_) );
AND2X2 AND2X2_632 ( .A(_5820_), .B(ULA_B_1_bF_buf6), .Y(_6068_) );
OR2X2 OR2X2_533 ( .A(_6067_), .B(_6068_), .Y(_6069_) );
AND2X2 AND2X2_633 ( .A(_6069_), .B(_5681__bF_buf4), .Y(_6070_) );
AND2X2 AND2X2_634 ( .A(_5822_), .B(_5682__bF_buf4), .Y(_6071_) );
AND2X2 AND2X2_635 ( .A(_5769_), .B(ULA_B_1_bF_buf6), .Y(_6072_) );
OR2X2 OR2X2_534 ( .A(_6071_), .B(_6072_), .Y(_6073_) );
AND2X2 AND2X2_636 ( .A(_6073_), .B(ULA_B_2_bF_buf2), .Y(_6074_) );
OR2X2 OR2X2_535 ( .A(_6070_), .B(_6074_), .Y(_6075_) );
AND2X2 AND2X2_637 ( .A(_6075_), .B(ULA_B_3_bF_buf7), .Y(_6076_) );
OR2X2 OR2X2_536 ( .A(_6066_), .B(_6076_), .Y(_6077_) );
AND2X2 AND2X2_638 ( .A(_6077_), .B(_5669__bF_buf2), .Y(_6078_) );
OR2X2 OR2X2_537 ( .A(_5799_), .B(_6078_), .Y(_6079_) );
OR2X2 OR2X2_538 ( .A(_6056_), .B(_6079_), .Y(_6080_) );
MUX2X1 MUX2X1_687 ( .A(_5822_), .B(_5769_), .S(_5417__bF_buf4), .Y(_6081_) );
MUX2X1 MUX2X1_688 ( .A(_5816_), .B(_5820_), .S(_5417__bF_buf0), .Y(_6082_) );
MUX2X1 MUX2X1_689 ( .A(_6082_), .B(_6081_), .S(_5353__bF_buf2), .Y(_6083_) );
OR2X2 OR2X2_539 ( .A(_5620__bF_buf2), .B(_6083_), .Y(_6084_) );
MUX2X1 MUX2X1_690 ( .A(_5808_), .B(_5814_), .S(_5417__bF_buf0), .Y(_6085_) );
MUX2X1 MUX2X1_691 ( .A(_5802_), .B(_5806_), .S(_5417__bF_buf0), .Y(_6086_) );
MUX2X1 MUX2X1_692 ( .A(_6086_), .B(_6085_), .S(_5353__bF_buf2), .Y(_6087_) );
OR2X2 OR2X2_540 ( .A(_5332__bF_buf1), .B(_6087_), .Y(_6088_) );
AND2X2 AND2X2_639 ( .A(_6084_), .B(_6088_), .Y(_6089_) );
OR2X2 OR2X2_541 ( .A(_5761_), .B(_6089_), .Y(_6090_) );
AND2X2 AND2X2_640 ( .A(_6090_), .B(_6080_), .Y(_6091_) );
AND2X2 AND2X2_641 ( .A(_6091_), .B(_6038_), .Y(_6092_) );
OR2X2 OR2X2_542 ( .A(_6001_), .B(_6092_), .Y(_6093_) );
INVX1 INVX1_17 ( .A(_6093_), .Y(ULA_ULA_OUT_3_) );
NOR2X1 NOR2X1_27 ( .A(_5739__bF_buf1), .B(ULA_OUT_0__4_), .Y(_6094_) );
OR2X2 OR2X2_543 ( .A(_5524__bF_buf3), .B(_5577_), .Y(_6095_) );
AND2X2 AND2X2_642 ( .A(_6095_), .B(_5332__bF_buf0), .Y(_6096_) );
AND2X2 AND2X2_643 ( .A(_5502_), .B(_5524__bF_buf3), .Y(_6097_) );
AND2X2 AND2X2_644 ( .A(_5658_), .B(_5353__bF_buf1), .Y(_6098_) );
OR2X2 OR2X2_544 ( .A(_6097_), .B(_6098_), .Y(_6099_) );
AND2X2 AND2X2_645 ( .A(_6099_), .B(_5620__bF_buf3), .Y(_6100_) );
OR2X2 OR2X2_545 ( .A(_6096_), .B(_6100_), .Y(_6101_) );
OR2X2 OR2X2_546 ( .A(_5679_), .B(_6101_), .Y(_6102_) );
AOI21X1 AOI21X1_3 ( .A(ULA_A_0_), .B(_6002_), .C(_5681__bF_buf3), .Y(_6103_) );
AND2X2 AND2X2_646 ( .A(_5946_), .B(ULA_B_1_bF_buf0), .Y(_6104_) );
MUX2X1 MUX2X1_693 ( .A(ULA_A_3_), .B(ULA_A_4_), .S(ULA_B_0_bF_buf6), .Y(_6105_) );
AND2X2 AND2X2_647 ( .A(_6105_), .B(_5682__bF_buf1), .Y(_6106_) );
OR2X2 OR2X2_547 ( .A(_6104_), .B(_6106_), .Y(_6107_) );
AND2X2 AND2X2_648 ( .A(_6107_), .B(_5681__bF_buf6), .Y(_6108_) );
OR2X2 OR2X2_548 ( .A(_6103_), .B(_6108_), .Y(_6109_) );
OR2X2 OR2X2_549 ( .A(ULA_B_3_bF_buf4), .B(_6109_), .Y(_6110_) );
OR2X2 OR2X2_550 ( .A(_5945__bF_buf3), .B(_6110_), .Y(_6111_) );
OR2X2 OR2X2_551 ( .A(ULA_A_4_), .B(ULA_B_4_bF_buf3), .Y(_6112_) );
NAND2X1 NAND2X1_654 ( .A(ULA_A_4_), .B(ULA_B_4_bF_buf3), .Y(_6113_) );
AND2X2 AND2X2_649 ( .A(_5735__bF_buf4), .B(_6113_), .Y(_6114_) );
OAI21X1 OAI21X1_2 ( .A(_6114_), .B(_5734__bF_buf2), .C(_6112_), .Y(_6115_) );
XOR2X1 XOR2X1_9 ( .A(ULA_cin_bF_buf6), .B(_6113_), .Y(_6116_) );
OR2X2 OR2X2_552 ( .A(_6116_), .B(_5940_), .Y(_6117_) );
AND2X2 AND2X2_650 ( .A(_6117_), .B(_5739__bF_buf2), .Y(_6118_) );
AND2X2 AND2X2_651 ( .A(_6115_), .B(_6118_), .Y(_6119_) );
AND2X2 AND2X2_652 ( .A(_6111_), .B(_6119_), .Y(_6120_) );
AND2X2 AND2X2_653 ( .A(_5725_), .B(ULA_B_1_bF_buf6), .Y(_6121_) );
AND2X2 AND2X2_654 ( .A(_5726_), .B(_5682__bF_buf4), .Y(_6122_) );
OR2X2 OR2X2_553 ( .A(_6121_), .B(_6122_), .Y(_6123_) );
OR2X2 OR2X2_554 ( .A(ULA_B_2_bF_buf0), .B(_6123_), .Y(_6124_) );
OR2X2 OR2X2_555 ( .A(_5681__bF_buf5), .B(_5712_), .Y(_6125_) );
AND2X2 AND2X2_655 ( .A(_6124_), .B(_6125_), .Y(_6126_) );
AND2X2 AND2X2_656 ( .A(_6126_), .B(_5289__bF_buf5), .Y(_6127_) );
AND2X2 AND2X2_657 ( .A(_5718_), .B(_5681__bF_buf5), .Y(_6128_) );
AND2X2 AND2X2_658 ( .A(_5685_), .B(ULA_B_2_bF_buf0), .Y(_6129_) );
OR2X2 OR2X2_556 ( .A(_6128_), .B(_6129_), .Y(_6130_) );
AND2X2 AND2X2_659 ( .A(_6130_), .B(ULA_B_3_bF_buf5), .Y(_6131_) );
OR2X2 OR2X2_557 ( .A(_6131_), .B(_6127_), .Y(_6132_) );
OR2X2 OR2X2_558 ( .A(_5730__bF_buf2), .B(_6132_), .Y(_6133_) );
AND2X2 AND2X2_660 ( .A(_6133_), .B(_6120_), .Y(_6134_) );
AND2X2 AND2X2_661 ( .A(_5664_), .B(_5524__bF_buf0), .Y(_6135_) );
AND2X2 AND2X2_662 ( .A(_5417__bF_buf5), .B(_5714_), .Y(_6136_) );
AND2X2 AND2X2_663 ( .A(_5470__bF_buf0), .B(_5716_), .Y(_6137_) );
OR2X2 OR2X2_559 ( .A(_6136_), .B(_6137_), .Y(_6138_) );
AND2X2 AND2X2_664 ( .A(_6138_), .B(_5353__bF_buf0), .Y(_6139_) );
OR2X2 OR2X2_560 ( .A(_6135_), .B(_6139_), .Y(_6140_) );
OR2X2 OR2X2_561 ( .A(_5620__bF_buf3), .B(_5761_), .Y(_6141_) );
OR2X2 OR2X2_562 ( .A(_6141_), .B(_6140_), .Y(_6142_) );
MUX2X1 MUX2X1_694 ( .A(_5757_), .B(_5753_), .S(_5353__bF_buf0), .Y(_6143_) );
OR2X2 OR2X2_563 ( .A(_5332__bF_buf3), .B(_5761_), .Y(_6144_) );
OR2X2 OR2X2_564 ( .A(_6144_), .B(_6143_), .Y(_6145_) );
OR2X2 OR2X2_565 ( .A(ULA_B_2_bF_buf1), .B(_5695_), .Y(_6146_) );
OR2X2 OR2X2_566 ( .A(_5289__bF_buf3), .B(_6146_), .Y(_6147_) );
AND2X2 AND2X2_665 ( .A(_5689_), .B(_5681__bF_buf3), .Y(_6148_) );
AND2X2 AND2X2_666 ( .A(_5699_), .B(ULA_B_2_bF_buf1), .Y(_6149_) );
OR2X2 OR2X2_567 ( .A(_6148_), .B(_6149_), .Y(_6150_) );
OR2X2 OR2X2_568 ( .A(ULA_B_3_bF_buf5), .B(_6150_), .Y(_6151_) );
AND2X2 AND2X2_667 ( .A(_6151_), .B(_6147_), .Y(_6152_) );
OR2X2 OR2X2_569 ( .A(_5706_), .B(_6152_), .Y(_6153_) );
AND2X2 AND2X2_668 ( .A(_6145_), .B(_6153_), .Y(_6154_) );
AND2X2 AND2X2_669 ( .A(_6154_), .B(_6142_), .Y(_6155_) );
AND2X2 AND2X2_670 ( .A(_6155_), .B(_6134_), .Y(_6156_) );
AND2X2 AND2X2_671 ( .A(_6156_), .B(_6102_), .Y(_6157_) );
OR2X2 OR2X2_570 ( .A(_6094_), .B(_6157_), .Y(_6158_) );
INVX1 INVX1_18 ( .A(_6158_), .Y(ULA_ULA_OUT_4_) );
AND2X2 AND2X2_672 ( .A(_5417__bF_buf4), .B(_5769_), .Y(_6159_) );
AND2X2 AND2X2_673 ( .A(_5470__bF_buf2), .B(_5771_), .Y(_6160_) );
OR2X2 OR2X2_571 ( .A(_6159_), .B(_6160_), .Y(_6161_) );
AND2X2 AND2X2_674 ( .A(_6161_), .B(_5524__bF_buf1), .Y(_6162_) );
AND2X2 AND2X2_675 ( .A(_5877_), .B(_5353__bF_buf4), .Y(_6163_) );
OR2X2 OR2X2_572 ( .A(_6162_), .B(_6163_), .Y(_6164_) );
INVX1 INVX1_19 ( .A(_6164_), .Y(_6165_) );
MUX2X1 MUX2X1_695 ( .A(_5881_), .B(_5867_), .S(_5524__bF_buf1), .Y(_6166_) );
MUX2X1 MUX2X1_696 ( .A(_6165_), .B(_6166_), .S(_5332__bF_buf2), .Y(_6167_) );
AND2X2 AND2X2_676 ( .A(_6167_), .B(_5672_), .Y(_6168_) );
AOI21X1 AOI21X1_4 ( .A(_5790_), .B(_5850_), .C(_5524__bF_buf2), .Y(_6169_) );
NOR2X1 NOR2X1_28 ( .A(_6169_), .B(_5620__bF_buf1), .Y(_6170_) );
MUX2X1 MUX2X1_697 ( .A(_5783_), .B(_5785_), .S(_5417__bF_buf1), .Y(_6171_) );
MUX2X1 MUX2X1_698 ( .A(_5859_), .B(_6171_), .S(_5353__bF_buf0), .Y(_6172_) );
AND2X2 AND2X2_677 ( .A(_6172_), .B(_5620__bF_buf1), .Y(_6173_) );
OR2X2 OR2X2_573 ( .A(_6173_), .B(_6170_), .Y(_6174_) );
AND2X2 AND2X2_678 ( .A(_6174_), .B(_5760_), .Y(_6175_) );
OR2X2 OR2X2_574 ( .A(_5678_), .B(_6175_), .Y(_6176_) );
OR2X2 OR2X2_575 ( .A(_6176_), .B(_6168_), .Y(_6177_) );
INVX1 INVX1_20 ( .A(_5845_), .Y(_6178_) );
AND2X2 AND2X2_679 ( .A(_5842_), .B(ULA_B_2_bF_buf6), .Y(_6179_) );
AND2X2 AND2X2_680 ( .A(_6023_), .B(ULA_B_1_bF_buf4), .Y(_6180_) );
MUX2X1 MUX2X1_699 ( .A(ULA_A_4_), .B(ULA_A_5_), .S(ULA_B_0_bF_buf1), .Y(_6181_) );
AND2X2 AND2X2_681 ( .A(_6181_), .B(_5682__bF_buf6), .Y(_6182_) );
OR2X2 OR2X2_576 ( .A(_6180_), .B(_6182_), .Y(_6183_) );
AND2X2 AND2X2_682 ( .A(_6183_), .B(_5681__bF_buf1), .Y(_6184_) );
NOR3X1 NOR3X1_5 ( .A(_6184_), .B(ULA_B_3_bF_buf1), .C(_6179_), .Y(_6185_) );
NAND3X1 NAND3X1_27 ( .A(_6185_), .B(_5669__bF_buf1), .C(_6178_), .Y(_6186_) );
NOR2X1 NOR2X1_29 ( .A(ULA_A_5_), .B(ULA_B_5_), .Y(_6187_) );
NAND2X1 NAND2X1_655 ( .A(ULA_A_5_), .B(ULA_B_5_), .Y(_6188_) );
AOI21X1 AOI21X1_5 ( .A(_6188_), .B(_5735__bF_buf2), .C(_5734__bF_buf4), .Y(_6189_) );
OR2X2 OR2X2_577 ( .A(_6187_), .B(_6189_), .Y(_6190_) );
NAND3X1 NAND3X1_28 ( .A(ULA_cin_bF_buf3), .B(ULA_A_5_), .C(ULA_B_5_), .Y(_6191_) );
NAND2X1 NAND2X1_656 ( .A(_5438__bF_buf3), .B(_6188_), .Y(_6192_) );
NAND3X1 NAND3X1_29 ( .A(_6192_), .B(_5740__bF_buf2), .C(_6191_), .Y(_6193_) );
AND2X2 AND2X2_683 ( .A(_6193_), .B(_5739__bF_buf1), .Y(_6194_) );
AND2X2 AND2X2_684 ( .A(_6190_), .B(_6194_), .Y(_6195_) );
AND2X2 AND2X2_685 ( .A(_6186_), .B(_6195_), .Y(_6196_) );
AND2X2 AND2X2_686 ( .A(_5779_), .B(_5681__bF_buf4), .Y(_6197_) );
AND2X2 AND2X2_687 ( .A(_5787_), .B(ULA_B_2_bF_buf2), .Y(_6198_) );
OR2X2 OR2X2_578 ( .A(_6197_), .B(_6198_), .Y(_6199_) );
AND2X2 AND2X2_688 ( .A(_6199_), .B(_5289__bF_buf1), .Y(_6200_) );
OR2X2 OR2X2_579 ( .A(ULA_B_2_bF_buf4), .B(_5793_), .Y(_6201_) );
AND2X2 AND2X2_689 ( .A(_6201_), .B(ULA_B_3_bF_buf3), .Y(_6202_) );
OR2X2 OR2X2_580 ( .A(_6202_), .B(_6200_), .Y(_6203_) );
OR2X2 OR2X2_581 ( .A(_5706_), .B(_6203_), .Y(_6204_) );
NAND2X1 NAND2X1_657 ( .A(_5681__bF_buf4), .B(_5810_), .Y(_6205_) );
NAND2X1 NAND2X1_658 ( .A(ULA_B_2_bF_buf3), .B(_5818_), .Y(_6206_) );
NAND3X1 NAND3X1_30 ( .A(_6205_), .B(_5289__bF_buf5), .C(_6206_), .Y(_6207_) );
AND2X2 AND2X2_690 ( .A(_5824_), .B(_5681__bF_buf4), .Y(_6208_) );
AND2X2 AND2X2_691 ( .A(_5773_), .B(ULA_B_2_bF_buf3), .Y(_6209_) );
OR2X2 OR2X2_582 ( .A(_6208_), .B(_6209_), .Y(_6210_) );
OR2X2 OR2X2_583 ( .A(_5289__bF_buf0), .B(_6210_), .Y(_6211_) );
AND2X2 AND2X2_692 ( .A(_6207_), .B(_6211_), .Y(_6212_) );
OR2X2 OR2X2_584 ( .A(_5730__bF_buf1), .B(_6212_), .Y(_6213_) );
AND2X2 AND2X2_693 ( .A(_6213_), .B(_6204_), .Y(_6214_) );
AND2X2 AND2X2_694 ( .A(_6214_), .B(_6196_), .Y(_6215_) );
AND2X2 AND2X2_695 ( .A(_6177_), .B(_6215_), .Y(_6216_) );
NOR2X1 NOR2X1_30 ( .A(_5739__bF_buf1), .B(ULA_OUT_0__5_), .Y(_6217_) );
OR2X2 OR2X2_585 ( .A(_6217_), .B(_6216_), .Y(_6218_) );
INVX1 INVX1_21 ( .A(_6218_), .Y(ULA_ULA_OUT_5_) );
NOR2X1 NOR2X1_31 ( .A(_5739__bF_buf1), .B(ULA_OUT_0__6_), .Y(_6219_) );
INVX1 INVX1_22 ( .A(_5534_), .Y(_6220_) );
NAND3X1 NAND3X1_31 ( .A(_6220_), .B(_5353__bF_buf3), .C(_5417__bF_buf2), .Y(_6221_) );
AND2X2 AND2X2_696 ( .A(_6221_), .B(_5332__bF_buf0), .Y(_6222_) );
AND2X2 AND2X2_697 ( .A(_5960_), .B(_5524__bF_buf3), .Y(_6223_) );
AND2X2 AND2X2_698 ( .A(_5966_), .B(_5353__bF_buf3), .Y(_6224_) );
OR2X2 OR2X2_586 ( .A(_6223_), .B(_6224_), .Y(_6225_) );
AND2X2 AND2X2_699 ( .A(_6225_), .B(_5620__bF_buf0), .Y(_6226_) );
OR2X2 OR2X2_587 ( .A(_6222_), .B(_6226_), .Y(_6227_) );
OR2X2 OR2X2_588 ( .A(_5679_), .B(_6227_), .Y(_6228_) );
AND2X2 AND2X2_700 ( .A(_5949_), .B(ULA_B_2_bF_buf5), .Y(_6229_) );
AND2X2 AND2X2_701 ( .A(_6105_), .B(ULA_B_1_bF_buf0), .Y(_6230_) );
MUX2X1 MUX2X1_700 ( .A(ULA_A_5_), .B(ULA_A_6_), .S(ULA_B_0_bF_buf4), .Y(_6231_) );
AND2X2 AND2X2_702 ( .A(_6231_), .B(_5682__bF_buf1), .Y(_6232_) );
OR2X2 OR2X2_589 ( .A(_6230_), .B(_6232_), .Y(_6233_) );
AND2X2 AND2X2_703 ( .A(_6233_), .B(_5681__bF_buf6), .Y(_6234_) );
OR2X2 OR2X2_590 ( .A(_6234_), .B(_6229_), .Y(_6235_) );
OR2X2 OR2X2_591 ( .A(ULA_B_3_bF_buf6), .B(_6235_), .Y(_6236_) );
OR2X2 OR2X2_592 ( .A(_5945__bF_buf2), .B(_6236_), .Y(_6237_) );
OR2X2 OR2X2_593 ( .A(ULA_A_6_), .B(ULA_B_6_), .Y(_6238_) );
NAND2X1 NAND2X1_659 ( .A(ULA_A_6_), .B(ULA_B_6_), .Y(_6239_) );
AND2X2 AND2X2_704 ( .A(_5735__bF_buf2), .B(_6239_), .Y(_6240_) );
OAI21X1 OAI21X1_3 ( .A(_6240_), .B(_5734__bF_buf4), .C(_6238_), .Y(_6241_) );
NOR2X1 NOR2X1_32 ( .A(_6239_), .B(_5438__bF_buf3), .Y(_6242_) );
AOI21X1 AOI21X1_6 ( .A(ULA_A_6_), .B(ULA_B_6_), .C(ULA_cin_bF_buf3), .Y(_6243_) );
OR2X2 OR2X2_594 ( .A(_6243_), .B(_5940_), .Y(_6244_) );
OR2X2 OR2X2_595 ( .A(_6242_), .B(_6244_), .Y(_6245_) );
AND2X2 AND2X2_705 ( .A(_6245_), .B(_5739__bF_buf5), .Y(_6246_) );
AND2X2 AND2X2_706 ( .A(_6241_), .B(_6246_), .Y(_6247_) );
AND2X2 AND2X2_707 ( .A(_6237_), .B(_6247_), .Y(_6248_) );
NOR2X1 NOR2X1_33 ( .A(_5678_), .B(_5760_), .Y(_6249_) );
MUX2X1 MUX2X1_701 ( .A(_5992_), .B(_5982_), .S(_5524__bF_buf0), .Y(_6250_) );
NAND3X1 NAND3X1_32 ( .A(_6250_), .B(_5620__bF_buf3), .C(_6249_), .Y(_6251_) );
AND2X2 AND2X2_708 ( .A(_6251_), .B(_6248_), .Y(_6252_) );
NOR2X1 NOR2X1_34 ( .A(_5799_), .B(ULA_B_4_bF_buf1), .Y(_6253_) );
MUX2X1 MUX2X1_702 ( .A(_5907_), .B(_5893_), .S(_5681__bF_buf5), .Y(_6254_) );
OR2X2 OR2X2_596 ( .A(ULA_B_3_bF_buf5), .B(_6254_), .Y(_6255_) );
AND2X2 AND2X2_709 ( .A(_5897_), .B(_5681__bF_buf5), .Y(_6256_) );
AND2X2 AND2X2_710 ( .A(_5915_), .B(ULA_B_2_bF_buf5), .Y(_6257_) );
OR2X2 OR2X2_597 ( .A(_6256_), .B(_6257_), .Y(_6258_) );
NAND2X1 NAND2X1_660 ( .A(ULA_B_3_bF_buf5), .B(_6258_), .Y(_6259_) );
NAND3X1 NAND3X1_33 ( .A(_6259_), .B(_6253_), .C(_6255_), .Y(_6260_) );
NAND3X1 NAND3X1_34 ( .A(_6220_), .B(_5682__bF_buf1), .C(_5681__bF_buf6), .Y(_6261_) );
AND2X2 AND2X2_711 ( .A(_6261_), .B(ULA_B_3_bF_buf2), .Y(_6262_) );
AND2X2 AND2X2_712 ( .A(_5927_), .B(ULA_B_2_bF_buf5), .Y(_6263_) );
AND2X2 AND2X2_713 ( .A(_5919_), .B(_5681__bF_buf6), .Y(_6264_) );
OR2X2 OR2X2_598 ( .A(_6263_), .B(_6264_), .Y(_6265_) );
AND2X2 AND2X2_714 ( .A(_6265_), .B(_5289__bF_buf2), .Y(_6266_) );
OR2X2 OR2X2_599 ( .A(_6266_), .B(_6262_), .Y(_6267_) );
OR2X2 OR2X2_600 ( .A(_5706_), .B(_6267_), .Y(_6268_) );
MUX2X1 MUX2X1_703 ( .A(_5662_), .B(_5630_), .S(_5417__bF_buf3), .Y(_6269_) );
MUX2X1 MUX2X1_704 ( .A(_5716_), .B(_5660_), .S(_5417__bF_buf3), .Y(_6270_) );
MUX2X1 MUX2X1_705 ( .A(_6270_), .B(_6269_), .S(_5353__bF_buf1), .Y(_6271_) );
OR2X2 OR2X2_601 ( .A(_6141_), .B(_6271_), .Y(_6272_) );
AND2X2 AND2X2_715 ( .A(_6272_), .B(_6268_), .Y(_6273_) );
AND2X2 AND2X2_716 ( .A(_6260_), .B(_6273_), .Y(_6274_) );
AND2X2 AND2X2_717 ( .A(_6274_), .B(_6252_), .Y(_6275_) );
AND2X2 AND2X2_718 ( .A(_6275_), .B(_6228_), .Y(_6276_) );
OR2X2 OR2X2_602 ( .A(_6219_), .B(_6276_), .Y(_6277_) );
INVX1 INVX1_23 ( .A(_6277_), .Y(ULA_ULA_OUT_6_) );
NOR2X1 NOR2X1_35 ( .A(_5739__bF_buf5), .B(ULA_OUT_0__7_), .Y(_6278_) );
INVX1 INVX1_24 ( .A(_5310_), .Y(_6279_) );
NAND3X1 NAND3X1_35 ( .A(_6279_), .B(ULA_B_3_bF_buf0), .C(ULA_A_31_), .Y(_6280_) );
AND2X2 AND2X2_719 ( .A(_6012_), .B(_5353__bF_buf4), .Y(_6281_) );
AND2X2 AND2X2_720 ( .A(_6006_), .B(_5524__bF_buf2), .Y(_6282_) );
OR2X2 OR2X2_603 ( .A(_6281_), .B(_6282_), .Y(_6283_) );
OR2X2 OR2X2_604 ( .A(_5332__bF_buf1), .B(_6283_), .Y(_6284_) );
AND2X2 AND2X2_721 ( .A(_6284_), .B(_6280_), .Y(_6285_) );
OR2X2 OR2X2_605 ( .A(_5679_), .B(_6285_), .Y(_6286_) );
AND2X2 AND2X2_722 ( .A(_6045_), .B(_5681__bF_buf2), .Y(_6287_) );
AND2X2 AND2X2_723 ( .A(_6051_), .B(ULA_B_2_bF_buf4), .Y(_6288_) );
OR2X2 OR2X2_606 ( .A(_6287_), .B(_6288_), .Y(_6289_) );
OR2X2 OR2X2_607 ( .A(ULA_B_3_bF_buf1), .B(_6289_), .Y(_6290_) );
AND2X2 AND2X2_724 ( .A(_6290_), .B(_6280_), .Y(_6291_) );
OR2X2 OR2X2_608 ( .A(_5706_), .B(_6291_), .Y(_6292_) );
AND2X2 AND2X2_725 ( .A(_6025_), .B(ULA_B_2_bF_buf6), .Y(_6293_) );
AND2X2 AND2X2_726 ( .A(_6181_), .B(ULA_B_1_bF_buf1), .Y(_6294_) );
MUX2X1 MUX2X1_706 ( .A(ULA_A_6_), .B(ULA_A_7_), .S(ULA_B_0_bF_buf5), .Y(_6295_) );
AND2X2 AND2X2_727 ( .A(_6295_), .B(_5682__bF_buf6), .Y(_6296_) );
OR2X2 OR2X2_609 ( .A(_6294_), .B(_6296_), .Y(_6297_) );
AND2X2 AND2X2_728 ( .A(_6297_), .B(_5681__bF_buf1), .Y(_6298_) );
OR2X2 OR2X2_610 ( .A(_6293_), .B(_6298_), .Y(_6299_) );
OR2X2 OR2X2_611 ( .A(ULA_B_3_bF_buf3), .B(_6299_), .Y(_6300_) );
OR2X2 OR2X2_612 ( .A(_5945__bF_buf0), .B(_6300_), .Y(_6301_) );
OR2X2 OR2X2_613 ( .A(ULA_A_7_), .B(ULA_B_7_), .Y(_6302_) );
NAND2X1 NAND2X1_661 ( .A(ULA_A_7_), .B(ULA_B_7_), .Y(_6303_) );
AND2X2 AND2X2_729 ( .A(_5735__bF_buf3), .B(_6303_), .Y(_6304_) );
OAI21X1 OAI21X1_4 ( .A(_6304_), .B(_5734__bF_buf1), .C(_6302_), .Y(_6305_) );
NAND3X1 NAND3X1_36 ( .A(ULA_cin_bF_buf5), .B(ULA_A_7_), .C(ULA_B_7_), .Y(_6306_) );
NAND2X1 NAND2X1_662 ( .A(_5438__bF_buf2), .B(_6303_), .Y(_6307_) );
NAND3X1 NAND3X1_37 ( .A(_6307_), .B(_5740__bF_buf3), .C(_6306_), .Y(_6308_) );
AND2X2 AND2X2_730 ( .A(_6308_), .B(_6305_), .Y(_6309_) );
AND2X2 AND2X2_731 ( .A(_6309_), .B(_5739__bF_buf2), .Y(_6310_) );
AND2X2 AND2X2_732 ( .A(_6310_), .B(_6301_), .Y(_6311_) );
AND2X2 AND2X2_733 ( .A(_6311_), .B(_6292_), .Y(_6312_) );
MUX2X1 MUX2X1_707 ( .A(_6085_), .B(_6082_), .S(_5353__bF_buf2), .Y(_6313_) );
OR2X2 OR2X2_614 ( .A(_6144_), .B(_6313_), .Y(_6314_) );
AND2X2 AND2X2_734 ( .A(_6016_), .B(_5524__bF_buf1), .Y(_6315_) );
AND2X2 AND2X2_735 ( .A(_5417__bF_buf0), .B(_5822_), .Y(_6316_) );
AND2X2 AND2X2_736 ( .A(_5470__bF_buf2), .B(_5769_), .Y(_6317_) );
OR2X2 OR2X2_615 ( .A(_6316_), .B(_6317_), .Y(_6318_) );
AND2X2 AND2X2_737 ( .A(_6318_), .B(_5353__bF_buf2), .Y(_6319_) );
OR2X2 OR2X2_616 ( .A(_6315_), .B(_6319_), .Y(_6320_) );
OR2X2 OR2X2_617 ( .A(_6141_), .B(_6320_), .Y(_6321_) );
AND2X2 AND2X2_738 ( .A(_6314_), .B(_6321_), .Y(_6322_) );
AND2X2 AND2X2_739 ( .A(_6063_), .B(_5681__bF_buf4), .Y(_6323_) );
AND2X2 AND2X2_740 ( .A(_6069_), .B(ULA_B_2_bF_buf3), .Y(_6324_) );
OR2X2 OR2X2_618 ( .A(_6323_), .B(_6324_), .Y(_6325_) );
AND2X2 AND2X2_741 ( .A(_6325_), .B(_5289__bF_buf5), .Y(_6326_) );
AND2X2 AND2X2_742 ( .A(_6073_), .B(_5681__bF_buf2), .Y(_6327_) );
AND2X2 AND2X2_743 ( .A(_6041_), .B(ULA_B_2_bF_buf2), .Y(_6328_) );
OR2X2 OR2X2_619 ( .A(_6327_), .B(_6328_), .Y(_6329_) );
AND2X2 AND2X2_744 ( .A(_6329_), .B(ULA_B_3_bF_buf7), .Y(_6330_) );
OR2X2 OR2X2_620 ( .A(_6326_), .B(_6330_), .Y(_6331_) );
OR2X2 OR2X2_621 ( .A(_5730__bF_buf1), .B(_6331_), .Y(_6332_) );
AND2X2 AND2X2_745 ( .A(_6322_), .B(_6332_), .Y(_6333_) );
AND2X2 AND2X2_746 ( .A(_6333_), .B(_6312_), .Y(_6334_) );
AND2X2 AND2X2_747 ( .A(_6334_), .B(_6286_), .Y(_6335_) );
OR2X2 OR2X2_622 ( .A(_6278_), .B(_6335_), .Y(_6336_) );
INVX1 INVX1_25 ( .A(_6336_), .Y(ULA_ULA_OUT_7_) );
OR2X2 OR2X2_623 ( .A(_5672_), .B(_5332__bF_buf0), .Y(_6337_) );
OR2X2 OR2X2_624 ( .A(_6337_), .B(_5598_), .Y(_6338_) );
AND2X2 AND2X2_748 ( .A(_5666_), .B(_5332__bF_buf3), .Y(_6339_) );
AND2X2 AND2X2_749 ( .A(_5754_), .B(_5620__bF_buf3), .Y(_6340_) );
OR2X2 OR2X2_625 ( .A(_5760_), .B(_6340_), .Y(_6341_) );
OR2X2 OR2X2_626 ( .A(_6339_), .B(_6341_), .Y(_6342_) );
AND2X2 AND2X2_750 ( .A(_6342_), .B(_6338_), .Y(_6343_) );
OR2X2 OR2X2_627 ( .A(_5678_), .B(_6343_), .Y(_6344_) );
AND2X2 AND2X2_751 ( .A(_6107_), .B(ULA_B_2_bF_buf5), .Y(_6345_) );
AND2X2 AND2X2_752 ( .A(_6231_), .B(ULA_B_1_bF_buf3), .Y(_6346_) );
MUX2X1 MUX2X1_708 ( .A(ULA_A_7_), .B(ULA_A_8_), .S(ULA_B_0_bF_buf6), .Y(_6347_) );
AND2X2 AND2X2_753 ( .A(_6347_), .B(_5682__bF_buf3), .Y(_6348_) );
OR2X2 OR2X2_628 ( .A(_6346_), .B(_6348_), .Y(_6349_) );
AND2X2 AND2X2_754 ( .A(_6349_), .B(_5681__bF_buf6), .Y(_6350_) );
OR2X2 OR2X2_629 ( .A(_6345_), .B(_6350_), .Y(_6351_) );
OR2X2 OR2X2_630 ( .A(ULA_B_3_bF_buf4), .B(_6351_), .Y(_6352_) );
NAND3X1 NAND3X1_38 ( .A(_6279_), .B(ULA_A_0_), .C(ULA_B_3_bF_buf4), .Y(_6353_) );
AND2X2 AND2X2_755 ( .A(_6352_), .B(_6353_), .Y(_6354_) );
OR2X2 OR2X2_631 ( .A(_5945__bF_buf2), .B(_6354_), .Y(_6355_) );
INVX1 INVX1_26 ( .A(_5735__bF_buf4), .Y(_6356_) );
AND2X2 AND2X2_756 ( .A(ULA_A_8_), .B(ULA_B_8_), .Y(_6357_) );
OAI21X1 OAI21X1_5 ( .A(_6357_), .B(_6356_), .C(_5933_), .Y(_6358_) );
OAI21X1 OAI21X1_6 ( .A(ULA_A_8_), .B(ULA_B_8_), .C(_6358_), .Y(_6359_) );
NAND2X1 NAND2X1_663 ( .A(ULA_cin_bF_buf3), .B(_6357_), .Y(_6360_) );
OR2X2 OR2X2_632 ( .A(ULA_cin_bF_buf3), .B(_6357_), .Y(_6361_) );
NAND3X1 NAND3X1_39 ( .A(_5740__bF_buf2), .B(_6360_), .C(_6361_), .Y(_6362_) );
AND2X2 AND2X2_757 ( .A(_6362_), .B(_5739__bF_buf1), .Y(_6363_) );
AND2X2 AND2X2_758 ( .A(_6359_), .B(_6363_), .Y(_6364_) );
OR2X2 OR2X2_633 ( .A(ULA_B_3_bF_buf0), .B(_5720_), .Y(_6365_) );
OR2X2 OR2X2_634 ( .A(_5289__bF_buf3), .B(_5691_), .Y(_6366_) );
AND2X2 AND2X2_759 ( .A(_6366_), .B(_5669__bF_buf3), .Y(_6367_) );
AND2X2 AND2X2_760 ( .A(_6367_), .B(_6365_), .Y(_6368_) );
OR2X2 OR2X2_635 ( .A(ULA_B_3_bF_buf4), .B(_5701_), .Y(_6369_) );
AND2X2 AND2X2_761 ( .A(_6369_), .B(ULA_B_4_bF_buf1), .Y(_6370_) );
OR2X2 OR2X2_636 ( .A(_5799_), .B(_6370_), .Y(_6371_) );
OR2X2 OR2X2_637 ( .A(_6368_), .B(_6371_), .Y(_6372_) );
AND2X2 AND2X2_762 ( .A(_6364_), .B(_6372_), .Y(_6373_) );
AND2X2 AND2X2_763 ( .A(_6373_), .B(_6355_), .Y(_6374_) );
AND2X2 AND2X2_764 ( .A(_6344_), .B(_6374_), .Y(_6375_) );
NOR2X1 NOR2X1_36 ( .A(_5739__bF_buf5), .B(ULA_OUT_0__8_), .Y(_6376_) );
OR2X2 OR2X2_638 ( .A(_6376_), .B(_6375_), .Y(_6377_) );
INVX1 INVX1_27 ( .A(_6377_), .Y(ULA_ULA_OUT_8_) );
NOR2X1 NOR2X1_37 ( .A(_5739__bF_buf5), .B(ULA_OUT_0__9_), .Y(_6378_) );
OR2X2 OR2X2_639 ( .A(_6337_), .B(_5857_), .Y(_6379_) );
AND2X2 AND2X2_765 ( .A(_5861_), .B(_5332__bF_buf2), .Y(_6380_) );
AND2X2 AND2X2_766 ( .A(_5883_), .B(_5620__bF_buf1), .Y(_6381_) );
OR2X2 OR2X2_640 ( .A(_5760_), .B(_6381_), .Y(_6382_) );
OR2X2 OR2X2_641 ( .A(_6382_), .B(_6380_), .Y(_6383_) );
AND2X2 AND2X2_767 ( .A(_6383_), .B(_6379_), .Y(_6384_) );
OR2X2 OR2X2_642 ( .A(_5678_), .B(_6384_), .Y(_6385_) );
OR2X2 OR2X2_643 ( .A(ULA_B_3_bF_buf7), .B(_5826_), .Y(_6386_) );
OR2X2 OR2X2_644 ( .A(_5289__bF_buf1), .B(_5781_), .Y(_6387_) );
AND2X2 AND2X2_768 ( .A(_6387_), .B(_5669__bF_buf2), .Y(_6388_) );
AND2X2 AND2X2_769 ( .A(_6388_), .B(_6386_), .Y(_6389_) );
OR2X2 OR2X2_645 ( .A(ULA_B_3_bF_buf3), .B(_5795_), .Y(_6390_) );
AND2X2 AND2X2_770 ( .A(_6390_), .B(ULA_B_4_bF_buf0), .Y(_6391_) );
OR2X2 OR2X2_646 ( .A(_5799_), .B(_6391_), .Y(_6392_) );
OR2X2 OR2X2_647 ( .A(_6389_), .B(_6392_), .Y(_6393_) );
AND2X2 AND2X2_771 ( .A(_5843_), .B(ULA_B_3_bF_buf0), .Y(_6394_) );
AND2X2 AND2X2_772 ( .A(_6183_), .B(ULA_B_2_bF_buf6), .Y(_6395_) );
AND2X2 AND2X2_773 ( .A(_6295_), .B(ULA_B_1_bF_buf1), .Y(_6396_) );
MUX2X1 MUX2X1_709 ( .A(ULA_A_8_), .B(ULA_A_9_), .S(ULA_B_0_bF_buf5), .Y(_6397_) );
AND2X2 AND2X2_774 ( .A(_6397_), .B(_5682__bF_buf6), .Y(_6398_) );
OR2X2 OR2X2_648 ( .A(_6396_), .B(_6398_), .Y(_6399_) );
AND2X2 AND2X2_775 ( .A(_6399_), .B(_5681__bF_buf3), .Y(_6400_) );
OR2X2 OR2X2_649 ( .A(_6395_), .B(_6400_), .Y(_6401_) );
AND2X2 AND2X2_776 ( .A(_6401_), .B(_5289__bF_buf4), .Y(_6402_) );
OR2X2 OR2X2_650 ( .A(_6394_), .B(_6402_), .Y(_6403_) );
OR2X2 OR2X2_651 ( .A(_5945__bF_buf3), .B(_6403_), .Y(_6404_) );
OR2X2 OR2X2_652 ( .A(ULA_A_9_), .B(ULA_B_9_), .Y(_6405_) );
NAND2X1 NAND2X1_664 ( .A(ULA_A_9_), .B(ULA_B_9_), .Y(_6406_) );
AND2X2 AND2X2_777 ( .A(_5735__bF_buf2), .B(_6406_), .Y(_6407_) );
OAI21X1 OAI21X1_7 ( .A(_6407_), .B(_5734__bF_buf4), .C(_6405_), .Y(_6408_) );
NOR2X1 NOR2X1_38 ( .A(_6406_), .B(_5438__bF_buf3), .Y(_6409_) );
AOI21X1 AOI21X1_7 ( .A(ULA_A_9_), .B(ULA_B_9_), .C(ULA_cin_bF_buf5), .Y(_6410_) );
OR2X2 OR2X2_653 ( .A(_6410_), .B(_5940_), .Y(_6411_) );
OR2X2 OR2X2_654 ( .A(_6409_), .B(_6411_), .Y(_6412_) );
AND2X2 AND2X2_778 ( .A(_6412_), .B(_5739__bF_buf0), .Y(_6413_) );
AND2X2 AND2X2_779 ( .A(_6408_), .B(_6413_), .Y(_6414_) );
AND2X2 AND2X2_780 ( .A(_6404_), .B(_6414_), .Y(_6415_) );
AND2X2 AND2X2_781 ( .A(_6393_), .B(_6415_), .Y(_6416_) );
AND2X2 AND2X2_782 ( .A(_6385_), .B(_6416_), .Y(_6417_) );
OR2X2 OR2X2_655 ( .A(_6378_), .B(_6417_), .Y(_6418_) );
INVX1 INVX1_28 ( .A(_6418_), .Y(ULA_ULA_OUT_9_) );
OR2X2 OR2X2_656 ( .A(_5332__bF_buf3), .B(_5994_), .Y(_6419_) );
OR2X2 OR2X2_657 ( .A(_5620__bF_buf0), .B(_5972_), .Y(_6420_) );
AND2X2 AND2X2_783 ( .A(_6419_), .B(_6420_), .Y(_6421_) );
OR2X2 OR2X2_658 ( .A(_5761_), .B(_6421_), .Y(_6422_) );
OR2X2 OR2X2_659 ( .A(ULA_B_3_bF_buf5), .B(_5899_), .Y(_6423_) );
OR2X2 OR2X2_660 ( .A(_5289__bF_buf2), .B(_5921_), .Y(_6424_) );
AND2X2 AND2X2_784 ( .A(_6424_), .B(_5669__bF_buf3), .Y(_6425_) );
AND2X2 AND2X2_785 ( .A(_6425_), .B(_6423_), .Y(_6426_) );
OR2X2 OR2X2_661 ( .A(ULA_B_3_bF_buf4), .B(_5929_), .Y(_6427_) );
AND2X2 AND2X2_786 ( .A(_6427_), .B(ULA_B_4_bF_buf1), .Y(_6428_) );
OR2X2 OR2X2_662 ( .A(_5799_), .B(_6428_), .Y(_6429_) );
OR2X2 OR2X2_663 ( .A(_6426_), .B(_6429_), .Y(_6430_) );
OR2X2 OR2X2_664 ( .A(_5678_), .B(_6337_), .Y(_6431_) );
OR2X2 OR2X2_665 ( .A(_5962_), .B(_6431_), .Y(_6432_) );
AND2X2 AND2X2_787 ( .A(_5950_), .B(ULA_B_3_bF_buf6), .Y(_6433_) );
AND2X2 AND2X2_788 ( .A(_6233_), .B(ULA_B_2_bF_buf7), .Y(_6434_) );
AND2X2 AND2X2_789 ( .A(_6347_), .B(ULA_B_1_bF_buf3), .Y(_6435_) );
MUX2X1 MUX2X1_710 ( .A(ULA_A_9_), .B(ULA_A_10_), .S(ULA_B_0_bF_buf2), .Y(_6436_) );
AND2X2 AND2X2_790 ( .A(_6436_), .B(_5682__bF_buf3), .Y(_6437_) );
OR2X2 OR2X2_666 ( .A(_6435_), .B(_6437_), .Y(_6438_) );
AND2X2 AND2X2_791 ( .A(_6438_), .B(_5681__bF_buf6), .Y(_6439_) );
OR2X2 OR2X2_667 ( .A(_6434_), .B(_6439_), .Y(_6440_) );
AND2X2 AND2X2_792 ( .A(_6440_), .B(_5289__bF_buf6), .Y(_6441_) );
OR2X2 OR2X2_668 ( .A(_6433_), .B(_6441_), .Y(_6442_) );
OR2X2 OR2X2_669 ( .A(_5945__bF_buf2), .B(_6442_), .Y(_6443_) );
NOR2X1 NOR2X1_39 ( .A(ULA_A_10_), .B(ULA_B_10_), .Y(_6444_) );
NAND2X1 NAND2X1_665 ( .A(ULA_A_10_), .B(ULA_B_10_), .Y(_6445_) );
AOI21X1 AOI21X1_8 ( .A(_6445_), .B(_5735__bF_buf3), .C(_5734__bF_buf1), .Y(_6446_) );
OR2X2 OR2X2_670 ( .A(_6444_), .B(_6446_), .Y(_6447_) );
XOR2X1 XOR2X1_10 ( .A(ULA_cin_bF_buf0), .B(_6445_), .Y(_6448_) );
OR2X2 OR2X2_671 ( .A(_6448_), .B(_5940_), .Y(_6449_) );
AND2X2 AND2X2_793 ( .A(_6449_), .B(_5739__bF_buf0), .Y(_6450_) );
AND2X2 AND2X2_794 ( .A(_6447_), .B(_6450_), .Y(_6451_) );
AND2X2 AND2X2_795 ( .A(_6443_), .B(_6451_), .Y(_6452_) );
AND2X2 AND2X2_796 ( .A(_6452_), .B(_6432_), .Y(_6453_) );
AND2X2 AND2X2_797 ( .A(_6453_), .B(_6430_), .Y(_6454_) );
AND2X2 AND2X2_798 ( .A(_6454_), .B(_6422_), .Y(_6455_) );
NOR2X1 NOR2X1_40 ( .A(_5739__bF_buf5), .B(ULA_OUT_0__10_), .Y(_6456_) );
OR2X2 OR2X2_672 ( .A(_6456_), .B(_6455_), .Y(_6457_) );
INVX1 INVX1_29 ( .A(_6457_), .Y(ULA_ULA_OUT_10_) );
NOR2X1 NOR2X1_41 ( .A(_5739__bF_buf2), .B(ULA_OUT_0__11_), .Y(_6458_) );
OR2X2 OR2X2_673 ( .A(_6337_), .B(_6008_), .Y(_6459_) );
AND2X2 AND2X2_799 ( .A(_6018_), .B(_5332__bF_buf1), .Y(_6460_) );
AND2X2 AND2X2_800 ( .A(_6083_), .B(_5620__bF_buf2), .Y(_6461_) );
OR2X2 OR2X2_674 ( .A(_5760_), .B(_6461_), .Y(_6462_) );
OR2X2 OR2X2_675 ( .A(_6460_), .B(_6462_), .Y(_6463_) );
AND2X2 AND2X2_801 ( .A(_6463_), .B(_6459_), .Y(_6464_) );
OR2X2 OR2X2_676 ( .A(_5678_), .B(_6464_), .Y(_6465_) );
NOR3X1 NOR3X1_6 ( .A(_6070_), .B(ULA_B_3_bF_buf7), .C(_6074_), .Y(_6466_) );
NOR3X1 NOR3X1_7 ( .A(_6042_), .B(_5289__bF_buf0), .C(_6046_), .Y(_6467_) );
NOR3X1 NOR3X1_8 ( .A(_6466_), .B(ULA_B_4_bF_buf2), .C(_6467_), .Y(_6468_) );
AOI21X1 AOI21X1_9 ( .A(_6003_), .B(_6052_), .C(ULA_B_3_bF_buf1), .Y(_6469_) );
OAI21X1 OAI21X1_8 ( .A(_5669__bF_buf2), .B(_6469_), .C(_5705_), .Y(_6470_) );
OR2X2 OR2X2_677 ( .A(_6470_), .B(_6468_), .Y(_6471_) );
OR2X2 OR2X2_678 ( .A(ULA_B_2_bF_buf6), .B(_6025_), .Y(_6472_) );
AND2X2 AND2X2_802 ( .A(_6472_), .B(ULA_B_3_bF_buf3), .Y(_6473_) );
AND2X2 AND2X2_803 ( .A(_6297_), .B(ULA_B_2_bF_buf4), .Y(_6474_) );
AND2X2 AND2X2_804 ( .A(_6397_), .B(ULA_B_1_bF_buf1), .Y(_6475_) );
MUX2X1 MUX2X1_711 ( .A(ULA_A_10_), .B(ULA_A_11_), .S(ULA_B_0_bF_buf3), .Y(_6476_) );
AND2X2 AND2X2_805 ( .A(_6476_), .B(_5682__bF_buf5), .Y(_4959_) );
OR2X2 OR2X2_679 ( .A(_6475_), .B(_4959_), .Y(_4960_) );
AND2X2 AND2X2_806 ( .A(_4960_), .B(_5681__bF_buf2), .Y(_4961_) );
OR2X2 OR2X2_680 ( .A(_6474_), .B(_4961_), .Y(_4962_) );
AND2X2 AND2X2_807 ( .A(_4962_), .B(_5289__bF_buf1), .Y(_4963_) );
OR2X2 OR2X2_681 ( .A(_6473_), .B(_4963_), .Y(_4964_) );
OR2X2 OR2X2_682 ( .A(_5945__bF_buf0), .B(_4964_), .Y(_4965_) );
OR2X2 OR2X2_683 ( .A(ULA_A_11_), .B(ULA_B_11_), .Y(_4966_) );
NAND2X1 NAND2X1_666 ( .A(ULA_A_11_), .B(ULA_B_11_), .Y(_4967_) );
AND2X2 AND2X2_808 ( .A(_5735__bF_buf4), .B(_4967_), .Y(_4968_) );
OAI21X1 OAI21X1_9 ( .A(_4968_), .B(_5734__bF_buf2), .C(_4966_), .Y(_4969_) );
NAND3X1 NAND3X1_40 ( .A(ULA_cin_bF_buf6), .B(ULA_A_11_), .C(ULA_B_11_), .Y(_4970_) );
NAND2X1 NAND2X1_667 ( .A(_5438__bF_buf2), .B(_4967_), .Y(_4971_) );
NAND3X1 NAND3X1_41 ( .A(_4971_), .B(_5740__bF_buf3), .C(_4970_), .Y(_4972_) );
AND2X2 AND2X2_809 ( .A(_4972_), .B(_5739__bF_buf2), .Y(_4973_) );
AND2X2 AND2X2_810 ( .A(_4973_), .B(_4969_), .Y(_4974_) );
AND2X2 AND2X2_811 ( .A(_4965_), .B(_4974_), .Y(_4975_) );
AND2X2 AND2X2_812 ( .A(_6471_), .B(_4975_), .Y(_4976_) );
AND2X2 AND2X2_813 ( .A(_6465_), .B(_4976_), .Y(_4977_) );
OR2X2 OR2X2_684 ( .A(_6458_), .B(_4977_), .Y(_4978_) );
INVX1 INVX1_30 ( .A(_4978_), .Y(ULA_ULA_OUT_11_) );
OR2X2 OR2X2_685 ( .A(_6095_), .B(_6337_), .Y(_4979_) );
AND2X2 AND2X2_814 ( .A(_6099_), .B(_5332__bF_buf3), .Y(_4980_) );
AND2X2 AND2X2_815 ( .A(_6140_), .B(_5620__bF_buf3), .Y(_4981_) );
OR2X2 OR2X2_686 ( .A(_5760_), .B(_4981_), .Y(_4982_) );
OR2X2 OR2X2_687 ( .A(_4980_), .B(_4982_), .Y(_4983_) );
AND2X2 AND2X2_816 ( .A(_4983_), .B(_4979_), .Y(_4984_) );
OR2X2 OR2X2_688 ( .A(_5678_), .B(_4984_), .Y(_4985_) );
OR2X2 OR2X2_689 ( .A(ULA_B_3_bF_buf5), .B(_6130_), .Y(_4986_) );
OR2X2 OR2X2_690 ( .A(_5289__bF_buf3), .B(_6150_), .Y(_4987_) );
AND2X2 AND2X2_817 ( .A(_4987_), .B(_5669__bF_buf3), .Y(_4988_) );
AND2X2 AND2X2_818 ( .A(_4988_), .B(_4986_), .Y(_4989_) );
NOR3X1 NOR3X1_9 ( .A(_5693_), .B(ULA_B_2_bF_buf1), .C(_5694_), .Y(_4990_) );
AND2X2 AND2X2_819 ( .A(_4990_), .B(_5289__bF_buf3), .Y(_4991_) );
OAI21X1 OAI21X1_10 ( .A(_5669__bF_buf0), .B(_4991_), .C(_5705_), .Y(_4992_) );
OR2X2 OR2X2_691 ( .A(_4989_), .B(_4992_), .Y(_4993_) );
AND2X2 AND2X2_820 ( .A(_6109_), .B(ULA_B_3_bF_buf4), .Y(_4994_) );
AND2X2 AND2X2_821 ( .A(_6349_), .B(ULA_B_2_bF_buf5), .Y(_4995_) );
AND2X2 AND2X2_822 ( .A(_6436_), .B(ULA_B_1_bF_buf3), .Y(_4996_) );
MUX2X1 MUX2X1_712 ( .A(ULA_A_11_), .B(ULA_A_12_), .S(ULA_B_0_bF_buf2), .Y(_4997_) );
AND2X2 AND2X2_823 ( .A(_4997_), .B(_5682__bF_buf3), .Y(_4998_) );
OR2X2 OR2X2_692 ( .A(_4996_), .B(_4998_), .Y(_4999_) );
AND2X2 AND2X2_824 ( .A(_4999_), .B(_5681__bF_buf6), .Y(_5000_) );
OR2X2 OR2X2_693 ( .A(_4995_), .B(_5000_), .Y(_5001_) );
AND2X2 AND2X2_825 ( .A(_5001_), .B(_5289__bF_buf2), .Y(_5002_) );
OR2X2 OR2X2_694 ( .A(_4994_), .B(_5002_), .Y(_5003_) );
OR2X2 OR2X2_695 ( .A(_5945__bF_buf2), .B(_5003_), .Y(_5004_) );
OR2X2 OR2X2_696 ( .A(ULA_A_12_), .B(ULA_B_12_), .Y(_5005_) );
NAND2X1 NAND2X1_668 ( .A(ULA_A_12_), .B(ULA_B_12_), .Y(_5006_) );
AND2X2 AND2X2_826 ( .A(_5735__bF_buf3), .B(_5006_), .Y(_5007_) );
OAI21X1 OAI21X1_11 ( .A(_5007_), .B(_5734__bF_buf3), .C(_5005_), .Y(_5008_) );
NOR2X1 NOR2X1_42 ( .A(_5006_), .B(_5438__bF_buf1), .Y(_5009_) );
AOI21X1 AOI21X1_10 ( .A(ULA_A_12_), .B(ULA_B_12_), .C(ULA_cin_bF_buf4), .Y(_5010_) );
OR2X2 OR2X2_697 ( .A(_5010_), .B(_5940_), .Y(_5011_) );
OR2X2 OR2X2_698 ( .A(_5009_), .B(_5011_), .Y(_5012_) );
AND2X2 AND2X2_827 ( .A(_5012_), .B(_5739__bF_buf7), .Y(_5013_) );
AND2X2 AND2X2_828 ( .A(_5008_), .B(_5013_), .Y(_5014_) );
AND2X2 AND2X2_829 ( .A(_5004_), .B(_5014_), .Y(_5015_) );
AND2X2 AND2X2_830 ( .A(_4993_), .B(_5015_), .Y(_5016_) );
AND2X2 AND2X2_831 ( .A(_4985_), .B(_5016_), .Y(_5017_) );
NOR2X1 NOR2X1_43 ( .A(_5739__bF_buf0), .B(ULA_OUT_0__12_), .Y(_5018_) );
OR2X2 OR2X2_699 ( .A(_5018_), .B(_5017_), .Y(_5019_) );
INVX1 INVX1_31 ( .A(_5019_), .Y(ULA_ULA_OUT_12_) );
NOR2X1 NOR2X1_44 ( .A(_5739__bF_buf2), .B(ULA_OUT_0__13_), .Y(_5020_) );
NAND3X1 NAND3X1_42 ( .A(_6169_), .B(_5620__bF_buf1), .C(_5760_), .Y(_5021_) );
AND2X2 AND2X2_832 ( .A(_6172_), .B(_5332__bF_buf2), .Y(_5022_) );
AND2X2 AND2X2_833 ( .A(_6164_), .B(_5620__bF_buf2), .Y(_5023_) );
OR2X2 OR2X2_700 ( .A(_5760_), .B(_5023_), .Y(_5024_) );
OR2X2 OR2X2_701 ( .A(_5024_), .B(_5022_), .Y(_5025_) );
AND2X2 AND2X2_834 ( .A(_5025_), .B(_5021_), .Y(_5026_) );
OR2X2 OR2X2_702 ( .A(_5678_), .B(_5026_), .Y(_5027_) );
OR2X2 OR2X2_703 ( .A(ULA_B_3_bF_buf7), .B(_6210_), .Y(_5028_) );
OR2X2 OR2X2_704 ( .A(_5289__bF_buf1), .B(_6199_), .Y(_5029_) );
AND2X2 AND2X2_835 ( .A(_5029_), .B(_5669__bF_buf2), .Y(_5030_) );
AND2X2 AND2X2_836 ( .A(_5030_), .B(_5028_), .Y(_5031_) );
OR2X2 OR2X2_705 ( .A(ULA_B_3_bF_buf3), .B(_6201_), .Y(_5032_) );
AND2X2 AND2X2_837 ( .A(_5032_), .B(ULA_B_4_bF_buf0), .Y(_5033_) );
OR2X2 OR2X2_706 ( .A(_5799_), .B(_5033_), .Y(_5034_) );
OR2X2 OR2X2_707 ( .A(_5034_), .B(_5031_), .Y(_5035_) );
OR2X2 OR2X2_708 ( .A(_6179_), .B(_6184_), .Y(_5036_) );
AND2X2 AND2X2_838 ( .A(_5036_), .B(ULA_B_3_bF_buf1), .Y(_5037_) );
AND2X2 AND2X2_839 ( .A(_6399_), .B(ULA_B_2_bF_buf4), .Y(_5038_) );
AND2X2 AND2X2_840 ( .A(_6476_), .B(ULA_B_1_bF_buf5), .Y(_5039_) );
MUX2X1 MUX2X1_713 ( .A(ULA_A_12_), .B(ULA_A_13_), .S(ULA_B_0_bF_buf3), .Y(_5040_) );
AND2X2 AND2X2_841 ( .A(_5040_), .B(_5682__bF_buf5), .Y(_5041_) );
OR2X2 OR2X2_709 ( .A(_5039_), .B(_5041_), .Y(_5042_) );
AND2X2 AND2X2_842 ( .A(_5042_), .B(_5681__bF_buf1), .Y(_5043_) );
OR2X2 OR2X2_710 ( .A(_5038_), .B(_5043_), .Y(_5044_) );
AND2X2 AND2X2_843 ( .A(_5044_), .B(_5289__bF_buf4), .Y(_5045_) );
OR2X2 OR2X2_711 ( .A(_5037_), .B(_5045_), .Y(_5046_) );
OR2X2 OR2X2_712 ( .A(_5945__bF_buf0), .B(_5046_), .Y(_5047_) );
NOR2X1 NOR2X1_45 ( .A(ULA_A_13_), .B(ULA_B_13_), .Y(_5048_) );
NAND2X1 NAND2X1_669 ( .A(ULA_A_13_), .B(ULA_B_13_), .Y(_5049_) );
AOI21X1 AOI21X1_11 ( .A(_5049_), .B(_5735__bF_buf4), .C(_5734__bF_buf2), .Y(_5050_) );
OR2X2 OR2X2_713 ( .A(_5048_), .B(_5050_), .Y(_5051_) );
XOR2X1 XOR2X1_11 ( .A(_5438__bF_buf2), .B(_5049_), .Y(_5052_) );
NAND2X1 NAND2X1_670 ( .A(_5052_), .B(_5740__bF_buf3), .Y(_5053_) );
AND2X2 AND2X2_844 ( .A(_5053_), .B(_5739__bF_buf3), .Y(_5054_) );
AND2X2 AND2X2_845 ( .A(_5051_), .B(_5054_), .Y(_5055_) );
AND2X2 AND2X2_846 ( .A(_5055_), .B(_5047_), .Y(_5056_) );
AND2X2 AND2X2_847 ( .A(_5056_), .B(_5035_), .Y(_5057_) );
AND2X2 AND2X2_848 ( .A(_5027_), .B(_5057_), .Y(_5058_) );
OR2X2 OR2X2_714 ( .A(_5020_), .B(_5058_), .Y(_5059_) );
INVX1 INVX1_32 ( .A(_5059_), .Y(ULA_ULA_OUT_13_) );
NOR2X1 NOR2X1_46 ( .A(_5739__bF_buf0), .B(ULA_OUT_0__14_), .Y(_5060_) );
OR2X2 OR2X2_715 ( .A(ULA_B_3_bF_buf5), .B(_6258_), .Y(_5061_) );
OR2X2 OR2X2_716 ( .A(_5289__bF_buf2), .B(_6265_), .Y(_5062_) );
AND2X2 AND2X2_849 ( .A(_5062_), .B(_5669__bF_buf3), .Y(_5063_) );
AND2X2 AND2X2_850 ( .A(_5063_), .B(_5061_), .Y(_5064_) );
NOR3X1 NOR3X1_10 ( .A(_5534_), .B(ULA_B_1_bF_buf0), .C(ULA_B_2_bF_buf5), .Y(_5065_) );
AOI21X1 AOI21X1_12 ( .A(_5289__bF_buf3), .B(_5065_), .C(_5669__bF_buf3), .Y(_5066_) );
OR2X2 OR2X2_717 ( .A(_5799_), .B(_5066_), .Y(_5067_) );
OR2X2 OR2X2_718 ( .A(_5067_), .B(_5064_), .Y(_5068_) );
AND2X2 AND2X2_851 ( .A(_6235_), .B(ULA_B_3_bF_buf6), .Y(_5069_) );
AND2X2 AND2X2_852 ( .A(_6438_), .B(ULA_B_2_bF_buf7), .Y(_5070_) );
AND2X2 AND2X2_853 ( .A(_4997_), .B(ULA_B_1_bF_buf3), .Y(_5071_) );
MUX2X1 MUX2X1_714 ( .A(ULA_A_13_), .B(ULA_A_14_), .S(ULA_B_0_bF_buf2), .Y(_5072_) );
AND2X2 AND2X2_854 ( .A(_5072_), .B(_5682__bF_buf3), .Y(_5073_) );
OR2X2 OR2X2_719 ( .A(_5071_), .B(_5073_), .Y(_5074_) );
AND2X2 AND2X2_855 ( .A(_5074_), .B(_5681__bF_buf0), .Y(_5075_) );
OR2X2 OR2X2_720 ( .A(_5070_), .B(_5075_), .Y(_5076_) );
AND2X2 AND2X2_856 ( .A(_5076_), .B(_5289__bF_buf6), .Y(_5077_) );
OR2X2 OR2X2_721 ( .A(_5077_), .B(_5069_), .Y(_5078_) );
OR2X2 OR2X2_722 ( .A(_5945__bF_buf1), .B(_5078_), .Y(_5079_) );
NOR2X1 NOR2X1_47 ( .A(ULA_A_14_), .B(ULA_B_14_), .Y(_5080_) );
NAND2X1 NAND2X1_671 ( .A(ULA_A_14_), .B(ULA_B_14_), .Y(_5081_) );
AOI21X1 AOI21X1_13 ( .A(_5081_), .B(_5735__bF_buf2), .C(_5734__bF_buf4), .Y(_5082_) );
OR2X2 OR2X2_723 ( .A(_5080_), .B(_5082_), .Y(_5083_) );
NAND3X1 NAND3X1_43 ( .A(ULA_cin_bF_buf6), .B(ULA_A_14_), .C(ULA_B_14_), .Y(_5084_) );
NAND2X1 NAND2X1_672 ( .A(_5438__bF_buf2), .B(_5081_), .Y(_5085_) );
NAND3X1 NAND3X1_44 ( .A(_5085_), .B(_5740__bF_buf2), .C(_5084_), .Y(_5086_) );
AND2X2 AND2X2_857 ( .A(_5086_), .B(_5739__bF_buf0), .Y(_5087_) );
AND2X2 AND2X2_858 ( .A(_5083_), .B(_5087_), .Y(_5088_) );
AND2X2 AND2X2_859 ( .A(_5079_), .B(_5088_), .Y(_5089_) );
AND2X2 AND2X2_860 ( .A(_5089_), .B(_5068_), .Y(_5090_) );
OR2X2 OR2X2_724 ( .A(_6141_), .B(_6225_), .Y(_5091_) );
OR2X2 OR2X2_725 ( .A(_6221_), .B(_6431_), .Y(_5092_) );
OR2X2 OR2X2_726 ( .A(_6144_), .B(_6271_), .Y(_5093_) );
AND2X2 AND2X2_861 ( .A(_5093_), .B(_5092_), .Y(_5094_) );
AND2X2 AND2X2_862 ( .A(_5094_), .B(_5091_), .Y(_5095_) );
AND2X2 AND2X2_863 ( .A(_5090_), .B(_5095_), .Y(_5096_) );
OR2X2 OR2X2_727 ( .A(_5060_), .B(_5096_), .Y(_5097_) );
INVX1 INVX1_33 ( .A(_5097_), .Y(ULA_ULA_OUT_14_) );
NOR2X1 NOR2X1_48 ( .A(_5739__bF_buf2), .B(ULA_OUT_0__15_), .Y(_5098_) );
INVX1 INVX1_34 ( .A(ULA_A_31_), .Y(_5099_) );
NOR2X1 NOR2X1_49 ( .A(_5670_), .B(_5099_), .Y(_5100_) );
NAND2X1 NAND2X1_673 ( .A(ULA_B_4_bF_buf0), .B(_5100_), .Y(_5101_) );
AND2X2 AND2X2_864 ( .A(_6283_), .B(_5332__bF_buf1), .Y(_5102_) );
AND2X2 AND2X2_865 ( .A(_6320_), .B(_5620__bF_buf2), .Y(_5103_) );
OR2X2 OR2X2_728 ( .A(_5760_), .B(_5103_), .Y(_5104_) );
OR2X2 OR2X2_729 ( .A(_5102_), .B(_5104_), .Y(_5105_) );
AND2X2 AND2X2_866 ( .A(_5105_), .B(_5101_), .Y(_5106_) );
OR2X2 OR2X2_730 ( .A(_5678_), .B(_5106_), .Y(_5107_) );
AND2X2 AND2X2_867 ( .A(_6329_), .B(_5289__bF_buf0), .Y(_5108_) );
AND2X2 AND2X2_868 ( .A(_6289_), .B(ULA_B_3_bF_buf1), .Y(_5109_) );
OR2X2 OR2X2_731 ( .A(_5108_), .B(_5109_), .Y(_5110_) );
OR2X2 OR2X2_732 ( .A(_5730__bF_buf0), .B(_5110_), .Y(_5111_) );
AND2X2 AND2X2_869 ( .A(_6299_), .B(ULA_B_3_bF_buf3), .Y(_5112_) );
AND2X2 AND2X2_870 ( .A(_4960_), .B(ULA_B_2_bF_buf2), .Y(_5113_) );
AND2X2 AND2X2_871 ( .A(_5040_), .B(ULA_B_1_bF_buf5), .Y(_5114_) );
MUX2X1 MUX2X1_715 ( .A(ULA_A_14_), .B(ULA_A_15_), .S(ULA_B_0_bF_buf3), .Y(_5115_) );
AND2X2 AND2X2_872 ( .A(_5115_), .B(_5682__bF_buf5), .Y(_5116_) );
OR2X2 OR2X2_733 ( .A(_5114_), .B(_5116_), .Y(_5117_) );
AND2X2 AND2X2_873 ( .A(_5117_), .B(_5681__bF_buf2), .Y(_5118_) );
OR2X2 OR2X2_734 ( .A(_5113_), .B(_5118_), .Y(_5119_) );
AND2X2 AND2X2_874 ( .A(_5119_), .B(_5289__bF_buf1), .Y(_5120_) );
OR2X2 OR2X2_735 ( .A(_5112_), .B(_5120_), .Y(_5121_) );
OR2X2 OR2X2_736 ( .A(_5945__bF_buf0), .B(_5121_), .Y(_5122_) );
NOR2X1 NOR2X1_50 ( .A(ULA_A_15_), .B(ULA_B_15_), .Y(_5123_) );
NAND2X1 NAND2X1_674 ( .A(ULA_A_15_), .B(ULA_B_15_), .Y(_5124_) );
AOI21X1 AOI21X1_14 ( .A(_5124_), .B(_5735__bF_buf1), .C(_5734__bF_buf2), .Y(_5125_) );
OR2X2 OR2X2_737 ( .A(_5123_), .B(_5125_), .Y(_5126_) );
XOR2X1 XOR2X1_12 ( .A(_5438__bF_buf2), .B(_5124_), .Y(_5127_) );
NAND2X1 NAND2X1_675 ( .A(_5127_), .B(_5740__bF_buf3), .Y(_5128_) );
AND2X2 AND2X2_875 ( .A(_5128_), .B(_5739__bF_buf3), .Y(_5129_) );
AND2X2 AND2X2_876 ( .A(_5126_), .B(_5129_), .Y(_5130_) );
NAND3X1 NAND3X1_45 ( .A(_5100_), .B(ULA_B_4_bF_buf3), .C(_5705_), .Y(_5131_) );
AND2X2 AND2X2_877 ( .A(_5130_), .B(_5131_), .Y(_5132_) );
AND2X2 AND2X2_878 ( .A(_5132_), .B(_5122_), .Y(_5133_) );
AND2X2 AND2X2_879 ( .A(_5133_), .B(_5111_), .Y(_5134_) );
AND2X2 AND2X2_880 ( .A(_5107_), .B(_5134_), .Y(_5135_) );
OR2X2 OR2X2_738 ( .A(_5098_), .B(_5135_), .Y(_5136_) );
INVX1 INVX1_35 ( .A(_5136_), .Y(ULA_ULA_OUT_15_) );
NOR2X1 NOR2X1_51 ( .A(_5739__bF_buf3), .B(ULA_OUT_0__16_), .Y(_5137_) );
OR2X2 OR2X2_739 ( .A(_5761_), .B(_5668_), .Y(_5138_) );
AND2X2 AND2X2_881 ( .A(_6351_), .B(ULA_B_3_bF_buf4), .Y(_5139_) );
AND2X2 AND2X2_882 ( .A(_5072_), .B(ULA_B_1_bF_buf7), .Y(_5140_) );
MUX2X1 MUX2X1_716 ( .A(ULA_A_15_), .B(ULA_A_16_), .S(ULA_B_0_bF_buf2), .Y(_5141_) );
AND2X2 AND2X2_883 ( .A(_5141_), .B(_5682__bF_buf3), .Y(_5142_) );
OR2X2 OR2X2_740 ( .A(_5140_), .B(_5142_), .Y(_5143_) );
AND2X2 AND2X2_884 ( .A(_5143_), .B(_5681__bF_buf0), .Y(_5144_) );
AND2X2 AND2X2_885 ( .A(_4999_), .B(ULA_B_2_bF_buf7), .Y(_5145_) );
OR2X2 OR2X2_741 ( .A(_5144_), .B(_5145_), .Y(_5146_) );
AND2X2 AND2X2_886 ( .A(_5146_), .B(_5289__bF_buf6), .Y(_5147_) );
OR2X2 OR2X2_742 ( .A(_5945__bF_buf1), .B(_5147_), .Y(_5148_) );
OR2X2 OR2X2_743 ( .A(_5139_), .B(_5148_), .Y(_5149_) );
OR2X2 OR2X2_744 ( .A(_5730__bF_buf2), .B(_5703_), .Y(_5150_) );
NOR2X1 NOR2X1_52 ( .A(ULA_A_16_), .B(ULA_B_16_), .Y(_5151_) );
NAND2X1 NAND2X1_676 ( .A(ULA_A_16_), .B(ULA_B_16_), .Y(_5152_) );
AOI21X1 AOI21X1_15 ( .A(_5152_), .B(_5735__bF_buf1), .C(_5734__bF_buf3), .Y(_5153_) );
OR2X2 OR2X2_745 ( .A(_5151_), .B(_5153_), .Y(_5154_) );
XOR2X1 XOR2X1_13 ( .A(_5438__bF_buf0), .B(_5152_), .Y(_5155_) );
NAND2X1 NAND2X1_677 ( .A(_5155_), .B(_5740__bF_buf1), .Y(_5156_) );
AND2X2 AND2X2_887 ( .A(_5156_), .B(_5739__bF_buf3), .Y(_5157_) );
AND2X2 AND2X2_888 ( .A(_5154_), .B(_5157_), .Y(_5158_) );
NOR2X1 NOR2X1_53 ( .A(_5845_), .B(_5669__bF_buf0), .Y(_5159_) );
NAND3X1 NAND3X1_46 ( .A(_5159_), .B(ULA_A_0_), .C(_5745_), .Y(_5160_) );
AND2X2 AND2X2_889 ( .A(_5158_), .B(_5160_), .Y(_5161_) );
AND2X2 AND2X2_890 ( .A(_5161_), .B(_5150_), .Y(_5162_) );
AND2X2 AND2X2_891 ( .A(_5162_), .B(_5149_), .Y(_5163_) );
AND2X2 AND2X2_892 ( .A(_5163_), .B(_5138_), .Y(_5164_) );
OR2X2 OR2X2_746 ( .A(_5137_), .B(_5164_), .Y(_5165_) );
INVX1 INVX1_36 ( .A(_5165_), .Y(ULA_ULA_OUT_16_) );
NOR2X1 NOR2X1_54 ( .A(_5739__bF_buf3), .B(ULA_OUT_0__17_), .Y(_5166_) );
OR2X2 OR2X2_747 ( .A(_5761_), .B(_5863_), .Y(_5167_) );
MUX2X1 MUX2X1_717 ( .A(_6399_), .B(_6183_), .S(_5681__bF_buf3), .Y(_5168_) );
AND2X2 AND2X2_893 ( .A(_5115_), .B(ULA_B_1_bF_buf1), .Y(_5169_) );
MUX2X1 MUX2X1_718 ( .A(ULA_A_16_), .B(ULA_A_17_), .S(ULA_B_0_bF_buf3), .Y(_5170_) );
AND2X2 AND2X2_894 ( .A(_5170_), .B(_5682__bF_buf5), .Y(_5171_) );
OR2X2 OR2X2_748 ( .A(_5169_), .B(_5171_), .Y(_5172_) );
MUX2X1 MUX2X1_719 ( .A(_5172_), .B(_5042_), .S(_5681__bF_buf1), .Y(_5173_) );
MUX2X1 MUX2X1_720 ( .A(_5173_), .B(_5168_), .S(_5289__bF_buf4), .Y(_5174_) );
AND2X2 AND2X2_895 ( .A(_5174_), .B(_5669__bF_buf1), .Y(_5175_) );
OAI21X1 OAI21X1_12 ( .A(ULA_B_3_bF_buf0), .B(_5843_), .C(ULA_B_4_bF_buf2), .Y(_5176_) );
NAND2X1 NAND2X1_678 ( .A(_6178_), .B(_5176_), .Y(_5177_) );
OR2X2 OR2X2_749 ( .A(_5177_), .B(_5175_), .Y(_5178_) );
OR2X2 OR2X2_750 ( .A(_5730__bF_buf0), .B(_5797_), .Y(_5179_) );
NOR2X1 NOR2X1_55 ( .A(ULA_A_17_), .B(ULA_B_17_), .Y(_5180_) );
NAND2X1 NAND2X1_679 ( .A(ULA_A_17_), .B(ULA_B_17_), .Y(_5181_) );
AOI21X1 AOI21X1_16 ( .A(_5181_), .B(_5735__bF_buf1), .C(_5734__bF_buf3), .Y(_5182_) );
OR2X2 OR2X2_751 ( .A(_5180_), .B(_5182_), .Y(_5183_) );
NAND3X1 NAND3X1_47 ( .A(ULA_cin_bF_buf7), .B(ULA_A_17_), .C(ULA_B_17_), .Y(_5184_) );
NAND2X1 NAND2X1_680 ( .A(_5438__bF_buf0), .B(_5181_), .Y(_5185_) );
NAND3X1 NAND3X1_48 ( .A(_5185_), .B(_5740__bF_buf1), .C(_5184_), .Y(_5186_) );
AND2X2 AND2X2_896 ( .A(_5186_), .B(_5739__bF_buf4), .Y(_5187_) );
AND2X2 AND2X2_897 ( .A(_5183_), .B(_5187_), .Y(_5188_) );
AND2X2 AND2X2_898 ( .A(_5179_), .B(_5188_), .Y(_5189_) );
AND2X2 AND2X2_899 ( .A(_5178_), .B(_5189_), .Y(_5190_) );
AND2X2 AND2X2_900 ( .A(_5190_), .B(_5167_), .Y(_5191_) );
OR2X2 OR2X2_752 ( .A(_5166_), .B(_5191_), .Y(_5192_) );
INVX1 INVX1_37 ( .A(_5192_), .Y(ULA_ULA_OUT_17_) );
NOR2X1 NOR2X1_56 ( .A(_5739__bF_buf3), .B(ULA_OUT_0__18_), .Y(_5193_) );
OR2X2 OR2X2_753 ( .A(_5761_), .B(_5974_), .Y(_5194_) );
OR2X2 OR2X2_754 ( .A(_5730__bF_buf3), .B(_5931_), .Y(_5195_) );
AND2X2 AND2X2_901 ( .A(_6440_), .B(ULA_B_3_bF_buf2), .Y(_5196_) );
AND2X2 AND2X2_902 ( .A(_5141_), .B(ULA_B_1_bF_buf7), .Y(_5197_) );
MUX2X1 MUX2X1_721 ( .A(ULA_A_17_), .B(ULA_A_18_), .S(ULA_B_0_bF_buf4), .Y(_5198_) );
AND2X2 AND2X2_903 ( .A(_5198_), .B(_5682__bF_buf0), .Y(_5199_) );
OR2X2 OR2X2_755 ( .A(_5197_), .B(_5199_), .Y(_5200_) );
AND2X2 AND2X2_904 ( .A(_5200_), .B(_5681__bF_buf0), .Y(_5201_) );
AND2X2 AND2X2_905 ( .A(_5074_), .B(ULA_B_2_bF_buf7), .Y(_5202_) );
OR2X2 OR2X2_756 ( .A(_5201_), .B(_5202_), .Y(_5203_) );
AND2X2 AND2X2_906 ( .A(_5203_), .B(_5289__bF_buf6), .Y(_5204_) );
OR2X2 OR2X2_757 ( .A(_5945__bF_buf1), .B(_5204_), .Y(_5205_) );
OR2X2 OR2X2_758 ( .A(_5196_), .B(_5205_), .Y(_5206_) );
NOR2X1 NOR2X1_57 ( .A(ULA_A_18_), .B(ULA_B_18_), .Y(_5207_) );
OR2X2 OR2X2_759 ( .A(_5207_), .B(_5933_), .Y(_5208_) );
XOR2X1 XOR2X1_14 ( .A(ULA_A_18_), .B(ULA_B_18_), .Y(_5209_) );
NAND3X1 NAND3X1_49 ( .A(_5209_), .B(_5676_), .C(_5704_), .Y(_5210_) );
AND2X2 AND2X2_907 ( .A(_5208_), .B(_5210_), .Y(_5211_) );
NAND2X1 NAND2X1_681 ( .A(ULA_A_18_), .B(ULA_B_18_), .Y(_5212_) );
XOR2X1 XOR2X1_15 ( .A(ULA_cin_bF_buf1), .B(_5212_), .Y(_5213_) );
OR2X2 OR2X2_760 ( .A(_5213_), .B(_5940_), .Y(_5214_) );
AND2X2 AND2X2_908 ( .A(_5214_), .B(_5739__bF_buf0), .Y(_5215_) );
AND2X2 AND2X2_909 ( .A(_5211_), .B(_5215_), .Y(_5216_) );
INVX1 INVX1_38 ( .A(_5159_), .Y(_5217_) );
OR2X2 OR2X2_761 ( .A(_5217_), .B(_5951_), .Y(_5218_) );
AND2X2 AND2X2_910 ( .A(_5218_), .B(_5216_), .Y(_5219_) );
AND2X2 AND2X2_911 ( .A(_5206_), .B(_5219_), .Y(_5220_) );
AND2X2 AND2X2_912 ( .A(_5220_), .B(_5195_), .Y(_5221_) );
AND2X2 AND2X2_913 ( .A(_5221_), .B(_5194_), .Y(_5222_) );
OR2X2 OR2X2_762 ( .A(_5193_), .B(_5222_), .Y(_5223_) );
INVX1 INVX1_39 ( .A(_5223_), .Y(ULA_ULA_OUT_18_) );
NOR2X1 NOR2X1_58 ( .A(_5739__bF_buf3), .B(ULA_OUT_0__19_), .Y(_5224_) );
OR2X2 OR2X2_763 ( .A(_5761_), .B(_6020_), .Y(_5225_) );
AND2X2 AND2X2_914 ( .A(_4962_), .B(ULA_B_3_bF_buf7), .Y(_5226_) );
AND2X2 AND2X2_915 ( .A(_5117_), .B(ULA_B_2_bF_buf2), .Y(_5227_) );
AND2X2 AND2X2_916 ( .A(_5170_), .B(ULA_B_1_bF_buf5), .Y(_5228_) );
MUX2X1 MUX2X1_722 ( .A(ULA_A_18_), .B(ULA_A_19_), .S(ULA_B_0_bF_buf1), .Y(_5229_) );
AND2X2 AND2X2_917 ( .A(_5229_), .B(_5682__bF_buf5), .Y(_5230_) );
OR2X2 OR2X2_764 ( .A(_5228_), .B(_5230_), .Y(_5231_) );
AND2X2 AND2X2_918 ( .A(_5231_), .B(_5681__bF_buf2), .Y(_5232_) );
OR2X2 OR2X2_765 ( .A(_5227_), .B(_5232_), .Y(_5233_) );
AND2X2 AND2X2_919 ( .A(_5233_), .B(_5289__bF_buf0), .Y(_5234_) );
OR2X2 OR2X2_766 ( .A(_5226_), .B(_5234_), .Y(_5235_) );
AND2X2 AND2X2_920 ( .A(_5235_), .B(_5669__bF_buf2), .Y(_5236_) );
OAI21X1 OAI21X1_13 ( .A(_5669__bF_buf0), .B(_6026_), .C(_6178_), .Y(_5237_) );
OR2X2 OR2X2_767 ( .A(_5236_), .B(_5237_), .Y(_5238_) );
OR2X2 OR2X2_768 ( .A(_5730__bF_buf0), .B(_6055_), .Y(_5239_) );
NOR2X1 NOR2X1_59 ( .A(ULA_A_19_), .B(ULA_B_19_), .Y(_5240_) );
NAND2X1 NAND2X1_682 ( .A(ULA_A_19_), .B(ULA_B_19_), .Y(_5241_) );
AOI21X1 AOI21X1_17 ( .A(_5241_), .B(_5735__bF_buf0), .C(_5734__bF_buf0), .Y(_5242_) );
OR2X2 OR2X2_769 ( .A(_5240_), .B(_5242_), .Y(_5243_) );
XOR2X1 XOR2X1_16 ( .A(ULA_cin_bF_buf7), .B(_5241_), .Y(_5244_) );
OR2X2 OR2X2_770 ( .A(_5244_), .B(_5940_), .Y(_5245_) );
AND2X2 AND2X2_921 ( .A(_5245_), .B(_5739__bF_buf4), .Y(_5246_) );
AND2X2 AND2X2_922 ( .A(_5243_), .B(_5246_), .Y(_5247_) );
AND2X2 AND2X2_923 ( .A(_5239_), .B(_5247_), .Y(_5248_) );
AND2X2 AND2X2_924 ( .A(_5238_), .B(_5248_), .Y(_5249_) );
AND2X2 AND2X2_925 ( .A(_5249_), .B(_5225_), .Y(_5250_) );
OR2X2 OR2X2_771 ( .A(_5224_), .B(_5250_), .Y(_5251_) );
INVX1 INVX1_40 ( .A(_5251_), .Y(ULA_ULA_OUT_19_) );
NOR2X1 NOR2X1_60 ( .A(_5739__bF_buf7), .B(ULA_OUT_0__20_), .Y(_5252_) );
OR2X2 OR2X2_772 ( .A(_5761_), .B(_6101_), .Y(_5253_) );
AND2X2 AND2X2_926 ( .A(_5143_), .B(ULA_B_2_bF_buf7), .Y(_5254_) );
AND2X2 AND2X2_927 ( .A(_5198_), .B(ULA_B_1_bF_buf7), .Y(_5255_) );
MUX2X1 MUX2X1_723 ( .A(ULA_A_19_), .B(ULA_A_20_), .S(ULA_B_0_bF_buf4), .Y(_5256_) );
AND2X2 AND2X2_928 ( .A(_5256_), .B(_5682__bF_buf0), .Y(_5257_) );
OR2X2 OR2X2_773 ( .A(_5255_), .B(_5257_), .Y(_5258_) );
AND2X2 AND2X2_929 ( .A(_5258_), .B(_5681__bF_buf0), .Y(_5259_) );
OR2X2 OR2X2_774 ( .A(_5254_), .B(_5259_), .Y(_5260_) );
OR2X2 OR2X2_775 ( .A(ULA_B_3_bF_buf2), .B(_5260_), .Y(_5261_) );
OR2X2 OR2X2_776 ( .A(_5289__bF_buf2), .B(_5001_), .Y(_5262_) );
AND2X2 AND2X2_930 ( .A(_5261_), .B(_5262_), .Y(_5263_) );
OR2X2 OR2X2_777 ( .A(_5945__bF_buf2), .B(_5263_), .Y(_5264_) );
OR2X2 OR2X2_778 ( .A(_5730__bF_buf3), .B(_6152_), .Y(_5265_) );
NOR2X1 NOR2X1_61 ( .A(ULA_A_20_), .B(ULA_B_20_), .Y(_5266_) );
OR2X2 OR2X2_779 ( .A(_5266_), .B(_5933_), .Y(_5267_) );
XOR2X1 XOR2X1_17 ( .A(ULA_A_20_), .B(ULA_B_20_), .Y(_5268_) );
NAND3X1 NAND3X1_50 ( .A(_5268_), .B(_5676_), .C(_5704_), .Y(_5269_) );
AND2X2 AND2X2_931 ( .A(_5267_), .B(_5269_), .Y(_5270_) );
NAND2X1 NAND2X1_683 ( .A(ULA_A_20_), .B(ULA_B_20_), .Y(_5271_) );
XOR2X1 XOR2X1_18 ( .A(ULA_cin_bF_buf5), .B(_5271_), .Y(_5272_) );
OR2X2 OR2X2_780 ( .A(_5272_), .B(_5940_), .Y(_5273_) );
AND2X2 AND2X2_932 ( .A(_5273_), .B(_5739__bF_buf0), .Y(_5274_) );
AND2X2 AND2X2_933 ( .A(_5270_), .B(_5274_), .Y(_5275_) );
OR2X2 OR2X2_781 ( .A(_5217_), .B(_6110_), .Y(_5276_) );
AND2X2 AND2X2_934 ( .A(_5276_), .B(_5275_), .Y(_5277_) );
AND2X2 AND2X2_935 ( .A(_5265_), .B(_5277_), .Y(_5278_) );
AND2X2 AND2X2_936 ( .A(_5278_), .B(_5264_), .Y(_5279_) );
AND2X2 AND2X2_937 ( .A(_5279_), .B(_5253_), .Y(_5280_) );
OR2X2 OR2X2_782 ( .A(_5252_), .B(_5280_), .Y(_5281_) );
INVX1 INVX1_41 ( .A(_5281_), .Y(ULA_ULA_OUT_20_) );
NOR2X1 NOR2X1_62 ( .A(_5739__bF_buf0), .B(ULA_OUT_0__21_), .Y(_5282_) );
OR2X2 OR2X2_783 ( .A(_5761_), .B(_6174_), .Y(_5283_) );
MUX2X1 MUX2X1_724 ( .A(_5042_), .B(_6399_), .S(_5681__bF_buf1), .Y(_5284_) );
AND2X2 AND2X2_938 ( .A(_5229_), .B(ULA_B_1_bF_buf1), .Y(_5285_) );
MUX2X1 MUX2X1_725 ( .A(ULA_A_20_), .B(ULA_A_21_), .S(ULA_B_0_bF_buf7), .Y(_5286_) );
AND2X2 AND2X2_939 ( .A(_5286_), .B(_5682__bF_buf6), .Y(_5287_) );
OR2X2 OR2X2_784 ( .A(_5285_), .B(_5287_), .Y(_5288_) );
MUX2X1 MUX2X1_726 ( .A(_5288_), .B(_5172_), .S(_5681__bF_buf1), .Y(_5290_) );
MUX2X1 MUX2X1_727 ( .A(_5290_), .B(_5284_), .S(_5289__bF_buf5), .Y(_5291_) );
AND2X2 AND2X2_940 ( .A(_5291_), .B(_5669__bF_buf1), .Y(_5292_) );
OAI21X1 OAI21X1_14 ( .A(_5669__bF_buf1), .B(_6185_), .C(_6178_), .Y(_5293_) );
OR2X2 OR2X2_785 ( .A(_5293_), .B(_5292_), .Y(_5294_) );
OR2X2 OR2X2_786 ( .A(_5730__bF_buf1), .B(_6203_), .Y(_5295_) );
NOR2X1 NOR2X1_63 ( .A(ULA_A_21_), .B(ULA_B_21_), .Y(_5296_) );
NAND2X1 NAND2X1_684 ( .A(ULA_A_21_), .B(ULA_B_21_), .Y(_5297_) );
AOI21X1 AOI21X1_18 ( .A(_5297_), .B(_5735__bF_buf3), .C(_5734__bF_buf1), .Y(_5298_) );
OR2X2 OR2X2_787 ( .A(_5296_), .B(_5298_), .Y(_5299_) );
NAND3X1 NAND3X1_51 ( .A(ULA_cin_bF_buf0), .B(ULA_A_21_), .C(ULA_B_21_), .Y(_5301_) );
NAND2X1 NAND2X1_685 ( .A(_5438__bF_buf1), .B(_5297_), .Y(_5302_) );
NAND3X1 NAND3X1_52 ( .A(_5302_), .B(_5740__bF_buf0), .C(_5301_), .Y(_5303_) );
AND2X2 AND2X2_941 ( .A(_5303_), .B(_5739__bF_buf7), .Y(_5304_) );
AND2X2 AND2X2_942 ( .A(_5299_), .B(_5304_), .Y(_5305_) );
AND2X2 AND2X2_943 ( .A(_5305_), .B(_5295_), .Y(_5306_) );
AND2X2 AND2X2_944 ( .A(_5294_), .B(_5306_), .Y(_5307_) );
AND2X2 AND2X2_945 ( .A(_5307_), .B(_5283_), .Y(_5308_) );
OR2X2 OR2X2_788 ( .A(_5282_), .B(_5308_), .Y(_5309_) );
INVX1 INVX1_42 ( .A(_5309_), .Y(ULA_ULA_OUT_21_) );
NOR2X1 NOR2X1_64 ( .A(_5739__bF_buf6), .B(ULA_OUT_0__22_), .Y(_5311_) );
OR2X2 OR2X2_789 ( .A(_5761_), .B(_6227_), .Y(_5312_) );
AND2X2 AND2X2_946 ( .A(_5076_), .B(ULA_B_3_bF_buf2), .Y(_5313_) );
AND2X2 AND2X2_947 ( .A(_5200_), .B(ULA_B_2_bF_buf7), .Y(_5314_) );
AND2X2 AND2X2_948 ( .A(_5256_), .B(ULA_B_1_bF_buf7), .Y(_5315_) );
MUX2X1 MUX2X1_728 ( .A(ULA_A_21_), .B(ULA_A_22_), .S(ULA_B_0_bF_buf4), .Y(_5316_) );
AND2X2 AND2X2_949 ( .A(_5316_), .B(_5682__bF_buf0), .Y(_5317_) );
OR2X2 OR2X2_790 ( .A(_5315_), .B(_5317_), .Y(_5318_) );
AND2X2 AND2X2_950 ( .A(_5318_), .B(_5681__bF_buf0), .Y(_5319_) );
OR2X2 OR2X2_791 ( .A(_5314_), .B(_5319_), .Y(_5320_) );
AND2X2 AND2X2_951 ( .A(_5320_), .B(_5289__bF_buf6), .Y(_5322_) );
OR2X2 OR2X2_792 ( .A(_5945__bF_buf1), .B(_5322_), .Y(_5323_) );
OR2X2 OR2X2_793 ( .A(_5313_), .B(_5323_), .Y(_5324_) );
OR2X2 OR2X2_794 ( .A(_5730__bF_buf3), .B(_6267_), .Y(_5325_) );
NOR2X1 NOR2X1_65 ( .A(ULA_A_22_), .B(ULA_B_22_), .Y(_5326_) );
NAND2X1 NAND2X1_686 ( .A(ULA_A_22_), .B(ULA_B_22_), .Y(_5327_) );
AOI21X1 AOI21X1_19 ( .A(_5327_), .B(_5735__bF_buf3), .C(_5734__bF_buf1), .Y(_5328_) );
OR2X2 OR2X2_795 ( .A(_5326_), .B(_5328_), .Y(_5329_) );
XOR2X1 XOR2X1_19 ( .A(_5438__bF_buf1), .B(_5327_), .Y(_5330_) );
NAND2X1 NAND2X1_687 ( .A(_5330_), .B(_5740__bF_buf0), .Y(_5331_) );
AND2X2 AND2X2_952 ( .A(_5331_), .B(_5739__bF_buf6), .Y(_5333_) );
AND2X2 AND2X2_953 ( .A(_5329_), .B(_5333_), .Y(_5334_) );
OR2X2 OR2X2_796 ( .A(_5217_), .B(_6236_), .Y(_5335_) );
AND2X2 AND2X2_954 ( .A(_5334_), .B(_5335_), .Y(_5336_) );
AND2X2 AND2X2_955 ( .A(_5336_), .B(_5325_), .Y(_5337_) );
AND2X2 AND2X2_956 ( .A(_5337_), .B(_5324_), .Y(_5338_) );
AND2X2 AND2X2_957 ( .A(_5338_), .B(_5312_), .Y(_5339_) );
OR2X2 OR2X2_797 ( .A(_5311_), .B(_5339_), .Y(_5340_) );
INVX1 INVX1_43 ( .A(_5340_), .Y(ULA_ULA_OUT_22_) );
NOR2X1 NOR2X1_66 ( .A(_5739__bF_buf6), .B(ULA_OUT_0__23_), .Y(_5341_) );
OR2X2 OR2X2_798 ( .A(_5761_), .B(_6285_), .Y(_5343_) );
AND2X2 AND2X2_958 ( .A(_5119_), .B(ULA_B_3_bF_buf1), .Y(_5344_) );
AND2X2 AND2X2_959 ( .A(_5231_), .B(ULA_B_2_bF_buf2), .Y(_5345_) );
AND2X2 AND2X2_960 ( .A(_5286_), .B(ULA_B_1_bF_buf1), .Y(_5346_) );
MUX2X1 MUX2X1_729 ( .A(ULA_A_22_), .B(ULA_A_23_), .S(ULA_B_0_bF_buf6), .Y(_5347_) );
AND2X2 AND2X2_961 ( .A(_5347_), .B(_5682__bF_buf6), .Y(_5348_) );
OR2X2 OR2X2_799 ( .A(_5346_), .B(_5348_), .Y(_5349_) );
AND2X2 AND2X2_962 ( .A(_5349_), .B(_5681__bF_buf2), .Y(_5350_) );
OR2X2 OR2X2_800 ( .A(_5345_), .B(_5350_), .Y(_5351_) );
AND2X2 AND2X2_963 ( .A(_5351_), .B(_5289__bF_buf1), .Y(_5352_) );
OR2X2 OR2X2_801 ( .A(_5344_), .B(_5352_), .Y(_5354_) );
AND2X2 AND2X2_964 ( .A(_5354_), .B(_5669__bF_buf1), .Y(_5355_) );
AND2X2 AND2X2_965 ( .A(_6300_), .B(ULA_B_4_bF_buf0), .Y(_5356_) );
OR2X2 OR2X2_802 ( .A(_5845_), .B(_5356_), .Y(_5357_) );
OR2X2 OR2X2_803 ( .A(_5355_), .B(_5357_), .Y(_5358_) );
OR2X2 OR2X2_804 ( .A(_5730__bF_buf2), .B(_6291_), .Y(_5359_) );
NOR2X1 NOR2X1_67 ( .A(ULA_A_23_), .B(ULA_B_23_), .Y(_5360_) );
NAND2X1 NAND2X1_688 ( .A(ULA_A_23_), .B(ULA_B_23_), .Y(_5361_) );
AOI21X1 AOI21X1_20 ( .A(_5361_), .B(_5735__bF_buf1), .C(_5734__bF_buf3), .Y(_5362_) );
OR2X2 OR2X2_805 ( .A(_5360_), .B(_5362_), .Y(_5363_) );
INVX1 INVX1_44 ( .A(_5739__bF_buf4), .Y(_5365_) );
XOR2X1 XOR2X1_20 ( .A(_5438__bF_buf0), .B(_5361_), .Y(_5366_) );
AOI21X1 AOI21X1_21 ( .A(_5366_), .B(_5740__bF_buf1), .C(_5365_), .Y(_5367_) );
AND2X2 AND2X2_966 ( .A(_5367_), .B(_5363_), .Y(_5368_) );
AND2X2 AND2X2_967 ( .A(_5368_), .B(_5359_), .Y(_5369_) );
AND2X2 AND2X2_968 ( .A(_5369_), .B(_5358_), .Y(_5370_) );
AND2X2 AND2X2_969 ( .A(_5370_), .B(_5343_), .Y(_5371_) );
OR2X2 OR2X2_806 ( .A(_5341_), .B(_5371_), .Y(_5372_) );
INVX1 INVX1_45 ( .A(_5372_), .Y(ULA_ULA_OUT_23_) );
NOR2X1 NOR2X1_68 ( .A(_5739__bF_buf6), .B(ULA_OUT_0__24_), .Y(_5373_) );
OR2X2 OR2X2_807 ( .A(_5217_), .B(_6354_), .Y(_5375_) );
NAND2X1 NAND2X1_689 ( .A(ULA_B_3_bF_buf6), .B(_5146_), .Y(_5376_) );
AND2X2 AND2X2_970 ( .A(_5316_), .B(ULA_B_1_bF_buf7), .Y(_5377_) );
MUX2X1 MUX2X1_730 ( .A(ULA_A_23_), .B(ULA_A_24_), .S(ULA_B_0_bF_buf4), .Y(_5378_) );
AND2X2 AND2X2_971 ( .A(_5378_), .B(_5682__bF_buf0), .Y(_5379_) );
OR2X2 OR2X2_808 ( .A(_5377_), .B(_5379_), .Y(_5380_) );
MUX2X1 MUX2X1_731 ( .A(_5380_), .B(_5258_), .S(_5681__bF_buf0), .Y(_5381_) );
OR2X2 OR2X2_809 ( .A(ULA_B_3_bF_buf2), .B(_5381_), .Y(_5382_) );
NAND3X1 NAND3X1_53 ( .A(_5376_), .B(_5846_), .C(_5382_), .Y(_5383_) );
AND2X2 AND2X2_972 ( .A(_5383_), .B(_5375_), .Y(_5384_) );
OR2X2 OR2X2_810 ( .A(_6144_), .B(_5598_), .Y(_5386_) );
OR2X2 OR2X2_811 ( .A(_5730__bF_buf3), .B(_6369_), .Y(_5387_) );
NOR2X1 NOR2X1_69 ( .A(ULA_A_24_), .B(ULA_B_24_), .Y(_5388_) );
NAND2X1 NAND2X1_690 ( .A(ULA_A_24_), .B(ULA_B_24_), .Y(_5389_) );
AOI21X1 AOI21X1_22 ( .A(_5389_), .B(_5735__bF_buf3), .C(_5734__bF_buf1), .Y(_5390_) );
OR2X2 OR2X2_812 ( .A(_5388_), .B(_5390_), .Y(_5391_) );
XOR2X1 XOR2X1_21 ( .A(_5438__bF_buf1), .B(_5389_), .Y(_5392_) );
NAND2X1 NAND2X1_691 ( .A(_5392_), .B(_5740__bF_buf0), .Y(_5393_) );
AND2X2 AND2X2_973 ( .A(_5393_), .B(_5739__bF_buf6), .Y(_5394_) );
AND2X2 AND2X2_974 ( .A(_5391_), .B(_5394_), .Y(_5395_) );
AND2X2 AND2X2_975 ( .A(_5395_), .B(_5387_), .Y(_5397_) );
AND2X2 AND2X2_976 ( .A(_5397_), .B(_5386_), .Y(_5398_) );
AND2X2 AND2X2_977 ( .A(_5384_), .B(_5398_), .Y(_5399_) );
OR2X2 OR2X2_813 ( .A(_5373_), .B(_5399_), .Y(_5400_) );
INVX1 INVX1_46 ( .A(_5400_), .Y(ULA_ULA_OUT_24_) );
NOR2X1 NOR2X1_70 ( .A(_5739__bF_buf6), .B(ULA_OUT_0__25_), .Y(_5401_) );
OR2X2 OR2X2_814 ( .A(_5217_), .B(_6403_), .Y(_5402_) );
NAND2X1 NAND2X1_692 ( .A(ULA_B_2_bF_buf4), .B(_5042_), .Y(_5403_) );
NAND2X1 NAND2X1_693 ( .A(_5681__bF_buf1), .B(_5172_), .Y(_5404_) );
AOI21X1 AOI21X1_23 ( .A(_5403_), .B(_5404_), .C(_5289__bF_buf4), .Y(_5405_) );
AND2X2 AND2X2_978 ( .A(_5347_), .B(ULA_B_1_bF_buf4), .Y(_5407_) );
MUX2X1 MUX2X1_732 ( .A(ULA_A_24_), .B(ULA_A_25_), .S(ULA_B_0_bF_buf5), .Y(_5408_) );
AND2X2 AND2X2_979 ( .A(_5408_), .B(_5682__bF_buf6), .Y(_5409_) );
OR2X2 OR2X2_815 ( .A(_5407_), .B(_5409_), .Y(_5410_) );
AND2X2 AND2X2_980 ( .A(_5410_), .B(_5681__bF_buf3), .Y(_5411_) );
AND2X2 AND2X2_981 ( .A(_5288_), .B(ULA_B_2_bF_buf4), .Y(_5412_) );
OR2X2 OR2X2_816 ( .A(_5411_), .B(_5412_), .Y(_5413_) );
AND2X2 AND2X2_982 ( .A(_5413_), .B(_5289__bF_buf4), .Y(_5414_) );
OR2X2 OR2X2_817 ( .A(_5945__bF_buf3), .B(_5414_), .Y(_5415_) );
OR2X2 OR2X2_818 ( .A(_5415_), .B(_5405_), .Y(_5416_) );
AND2X2 AND2X2_983 ( .A(_5416_), .B(_5402_), .Y(_5418_) );
OR2X2 OR2X2_819 ( .A(_6144_), .B(_5857_), .Y(_5419_) );
OR2X2 OR2X2_820 ( .A(_5730__bF_buf2), .B(_6390_), .Y(_5420_) );
OR2X2 OR2X2_821 ( .A(ULA_A_25_), .B(ULA_B_25_), .Y(_5421_) );
NAND2X1 NAND2X1_694 ( .A(ULA_A_25_), .B(ULA_B_25_), .Y(_5422_) );
AND2X2 AND2X2_984 ( .A(_5735__bF_buf0), .B(_5422_), .Y(_5423_) );
OAI21X1 OAI21X1_15 ( .A(_5423_), .B(_5734__bF_buf0), .C(_5421_), .Y(_5424_) );
XOR2X1 XOR2X1_22 ( .A(ULA_cin_bF_buf4), .B(_5422_), .Y(_5425_) );
OR2X2 OR2X2_822 ( .A(_5425_), .B(_5940_), .Y(_5426_) );
AND2X2 AND2X2_985 ( .A(_5426_), .B(_5739__bF_buf7), .Y(_5427_) );
AND2X2 AND2X2_986 ( .A(_5424_), .B(_5427_), .Y(_5429_) );
AND2X2 AND2X2_987 ( .A(_5420_), .B(_5429_), .Y(_5430_) );
AND2X2 AND2X2_988 ( .A(_5430_), .B(_5419_), .Y(_5431_) );
AND2X2 AND2X2_989 ( .A(_5418_), .B(_5431_), .Y(_5432_) );
OR2X2 OR2X2_823 ( .A(_5401_), .B(_5432_), .Y(_5433_) );
INVX1 INVX1_47 ( .A(_5433_), .Y(ULA_ULA_OUT_25_) );
NOR2X1 NOR2X1_71 ( .A(_5739__bF_buf6), .B(ULA_OUT_0__26_), .Y(_5434_) );
OR2X2 OR2X2_824 ( .A(_5217_), .B(_6442_), .Y(_5435_) );
OR2X2 OR2X2_825 ( .A(_5730__bF_buf3), .B(_6427_), .Y(_5436_) );
OR2X2 OR2X2_826 ( .A(ULA_A_26_), .B(ULA_B_26_), .Y(_5437_) );
NAND2X1 NAND2X1_695 ( .A(ULA_A_26_), .B(ULA_B_26_), .Y(_5439_) );
AND2X2 AND2X2_990 ( .A(_5735__bF_buf0), .B(_5439_), .Y(_5440_) );
OAI21X1 OAI21X1_16 ( .A(_5440_), .B(_5734__bF_buf0), .C(_5437_), .Y(_5441_) );
XOR2X1 XOR2X1_23 ( .A(ULA_cin_bF_buf4), .B(_5439_), .Y(_5442_) );
OR2X2 OR2X2_827 ( .A(_5442_), .B(_5940_), .Y(_5443_) );
AND2X2 AND2X2_991 ( .A(_5443_), .B(_5739__bF_buf7), .Y(_5444_) );
AND2X2 AND2X2_992 ( .A(_5441_), .B(_5444_), .Y(_5445_) );
AND2X2 AND2X2_993 ( .A(_5436_), .B(_5445_), .Y(_5446_) );
AND2X2 AND2X2_994 ( .A(_5446_), .B(_5435_), .Y(_5447_) );
OR2X2 OR2X2_828 ( .A(_6144_), .B(_5962_), .Y(_5448_) );
AND2X2 AND2X2_995 ( .A(_5378_), .B(ULA_B_1_bF_buf7), .Y(_5450_) );
MUX2X1 MUX2X1_733 ( .A(ULA_A_25_), .B(ULA_A_26_), .S(ULA_B_0_bF_buf4), .Y(_5451_) );
AND2X2 AND2X2_996 ( .A(_5451_), .B(_5682__bF_buf0), .Y(_5452_) );
OR2X2 OR2X2_829 ( .A(_5450_), .B(_5452_), .Y(_5453_) );
AND2X2 AND2X2_997 ( .A(_5453_), .B(_5681__bF_buf0), .Y(_5454_) );
AND2X2 AND2X2_998 ( .A(_5318_), .B(ULA_B_2_bF_buf7), .Y(_5455_) );
OR2X2 OR2X2_830 ( .A(_5454_), .B(_5455_), .Y(_5456_) );
AND2X2 AND2X2_999 ( .A(_5456_), .B(_5289__bF_buf6), .Y(_5457_) );
AND2X2 AND2X2_1000 ( .A(_5203_), .B(ULA_B_3_bF_buf2), .Y(_5458_) );
OR2X2 OR2X2_831 ( .A(_5457_), .B(_5458_), .Y(_5459_) );
OR2X2 OR2X2_832 ( .A(_5945__bF_buf1), .B(_5459_), .Y(_5461_) );
AND2X2 AND2X2_1001 ( .A(_5461_), .B(_5448_), .Y(_5462_) );
AND2X2 AND2X2_1002 ( .A(_5447_), .B(_5462_), .Y(_5463_) );
OR2X2 OR2X2_833 ( .A(_5434_), .B(_5463_), .Y(_5464_) );
INVX1 INVX1_48 ( .A(_5464_), .Y(ULA_ULA_OUT_26_) );
NOR2X1 NOR2X1_72 ( .A(_5739__bF_buf6), .B(ULA_OUT_0__27_), .Y(_5465_) );
AND2X2 AND2X2_1003 ( .A(_5233_), .B(ULA_B_3_bF_buf7), .Y(_5466_) );
AND2X2 AND2X2_1004 ( .A(_5408_), .B(ULA_B_1_bF_buf4), .Y(_5467_) );
MUX2X1 MUX2X1_734 ( .A(ULA_A_26_), .B(ULA_A_27_), .S(ULA_B_0_bF_buf5), .Y(_5468_) );
AND2X2 AND2X2_1005 ( .A(_5468_), .B(_5682__bF_buf1), .Y(_5469_) );
OR2X2 OR2X2_834 ( .A(_5467_), .B(_5469_), .Y(_5471_) );
AND2X2 AND2X2_1006 ( .A(_5471_), .B(_5681__bF_buf1), .Y(_5472_) );
AND2X2 AND2X2_1007 ( .A(_5349_), .B(ULA_B_2_bF_buf2), .Y(_5473_) );
OR2X2 OR2X2_835 ( .A(_5472_), .B(_5473_), .Y(_5474_) );
AND2X2 AND2X2_1008 ( .A(_5474_), .B(_5289__bF_buf0), .Y(_5475_) );
OR2X2 OR2X2_836 ( .A(_5466_), .B(_5475_), .Y(_5476_) );
OR2X2 OR2X2_837 ( .A(_5945__bF_buf0), .B(_5476_), .Y(_5477_) );
OR2X2 OR2X2_838 ( .A(ULA_B_3_bF_buf3), .B(_6053_), .Y(_5478_) );
OR2X2 OR2X2_839 ( .A(_5730__bF_buf0), .B(_5478_), .Y(_5479_) );
NOR2X1 NOR2X1_73 ( .A(ULA_A_27_), .B(ULA_B_27_), .Y(_5480_) );
OR2X2 OR2X2_840 ( .A(_5480_), .B(_5933_), .Y(_5482_) );
XOR2X1 XOR2X1_24 ( .A(ULA_A_27_), .B(ULA_B_27_), .Y(_5483_) );
NAND3X1 NAND3X1_54 ( .A(_5483_), .B(_5676_), .C(_5704_), .Y(_5484_) );
AND2X2 AND2X2_1009 ( .A(_5482_), .B(_5484_), .Y(_5485_) );
NAND2X1 NAND2X1_696 ( .A(ULA_A_27_), .B(ULA_B_27_), .Y(_5486_) );
XOR2X1 XOR2X1_25 ( .A(ULA_cin_bF_buf1), .B(_5486_), .Y(_5487_) );
OR2X2 OR2X2_841 ( .A(_5487_), .B(_5940_), .Y(_5488_) );
AND2X2 AND2X2_1010 ( .A(_5488_), .B(_5739__bF_buf3), .Y(_5489_) );
AND2X2 AND2X2_1011 ( .A(_5485_), .B(_5489_), .Y(_5490_) );
AND2X2 AND2X2_1012 ( .A(_5479_), .B(_5490_), .Y(_5491_) );
AND2X2 AND2X2_1013 ( .A(_5477_), .B(_5491_), .Y(_5493_) );
OR2X2 OR2X2_842 ( .A(_5217_), .B(_4964_), .Y(_5494_) );
OR2X2 OR2X2_843 ( .A(_6144_), .B(_6008_), .Y(_5495_) );
AND2X2 AND2X2_1014 ( .A(_5494_), .B(_5495_), .Y(_5496_) );
AND2X2 AND2X2_1015 ( .A(_5493_), .B(_5496_), .Y(_5497_) );
OR2X2 OR2X2_844 ( .A(_5465_), .B(_5497_), .Y(_5498_) );
INVX1 INVX1_49 ( .A(_5498_), .Y(ULA_ULA_OUT_27_) );
NOR2X1 NOR2X1_74 ( .A(_5739__bF_buf7), .B(ULA_OUT_0__28_), .Y(_5499_) );
INVX1 INVX1_50 ( .A(_5380_), .Y(_5500_) );
MUX2X1 MUX2X1_735 ( .A(ULA_A_27_), .B(ULA_A_28_), .S(ULA_B_0_bF_buf4), .Y(_5501_) );
MUX2X1 MUX2X1_736 ( .A(_5501_), .B(_5451_), .S(_5682__bF_buf0), .Y(_5503_) );
MUX2X1 MUX2X1_737 ( .A(_5500_), .B(_5503_), .S(ULA_B_2_bF_buf7), .Y(_5504_) );
OR2X2 OR2X2_845 ( .A(ULA_B_3_bF_buf2), .B(_5504_), .Y(_5505_) );
OR2X2 OR2X2_846 ( .A(_5289__bF_buf6), .B(_5260_), .Y(_5506_) );
AND2X2 AND2X2_1016 ( .A(_5505_), .B(_5506_), .Y(_5507_) );
OR2X2 OR2X2_847 ( .A(_5945__bF_buf2), .B(_5507_), .Y(_5508_) );
NAND2X1 NAND2X1_697 ( .A(_6253_), .B(_4991_), .Y(_5509_) );
NOR2X1 NOR2X1_75 ( .A(ULA_A_28_), .B(ULA_B_28_), .Y(_5510_) );
NAND2X1 NAND2X1_698 ( .A(ULA_A_28_), .B(ULA_B_28_), .Y(_5511_) );
AOI21X1 AOI21X1_24 ( .A(_5511_), .B(_5735__bF_buf1), .C(_5734__bF_buf3), .Y(_5512_) );
OR2X2 OR2X2_848 ( .A(_5510_), .B(_5512_), .Y(_5514_) );
NAND3X1 NAND3X1_55 ( .A(ULA_cin_bF_buf7), .B(ULA_A_28_), .C(ULA_B_28_), .Y(_5515_) );
NAND2X1 NAND2X1_699 ( .A(_5438__bF_buf0), .B(_5511_), .Y(_5516_) );
NAND3X1 NAND3X1_56 ( .A(_5516_), .B(_5740__bF_buf1), .C(_5515_), .Y(_5517_) );
AND2X2 AND2X2_1017 ( .A(_5517_), .B(_5739__bF_buf4), .Y(_5518_) );
AND2X2 AND2X2_1018 ( .A(_5514_), .B(_5518_), .Y(_5519_) );
AND2X2 AND2X2_1019 ( .A(_5519_), .B(_5509_), .Y(_5520_) );
AND2X2 AND2X2_1020 ( .A(_5508_), .B(_5520_), .Y(_5521_) );
OR2X2 OR2X2_849 ( .A(_5217_), .B(_5003_), .Y(_5522_) );
OR2X2 OR2X2_850 ( .A(_6095_), .B(_6144_), .Y(_5523_) );
AND2X2 AND2X2_1021 ( .A(_5522_), .B(_5523_), .Y(_5525_) );
AND2X2 AND2X2_1022 ( .A(_5521_), .B(_5525_), .Y(_5526_) );
OR2X2 OR2X2_851 ( .A(_5499_), .B(_5526_), .Y(_5527_) );
INVX1 INVX1_51 ( .A(_5527_), .Y(ULA_ULA_OUT_28_) );
NOR2X1 NOR2X1_76 ( .A(_5739__bF_buf4), .B(ULA_OUT_0__29_), .Y(_5528_) );
NAND3X1 NAND3X1_57 ( .A(_6249_), .B(_5620__bF_buf1), .C(_6169_), .Y(_5529_) );
OR2X2 OR2X2_852 ( .A(_5730__bF_buf2), .B(_5032_), .Y(_5530_) );
NOR2X1 NOR2X1_77 ( .A(ULA_A_29_), .B(ULA_B_29_), .Y(_5531_) );
NAND2X1 NAND2X1_700 ( .A(ULA_A_29_), .B(ULA_B_29_), .Y(_5532_) );
AOI21X1 AOI21X1_25 ( .A(_5532_), .B(_5735__bF_buf0), .C(_5734__bF_buf0), .Y(_5533_) );
OR2X2 OR2X2_853 ( .A(_5531_), .B(_5533_), .Y(_5535_) );
XOR2X1 XOR2X1_26 ( .A(_5438__bF_buf0), .B(_5532_), .Y(_5536_) );
NAND2X1 NAND2X1_701 ( .A(_5536_), .B(_5740__bF_buf1), .Y(_5537_) );
AND2X2 AND2X2_1023 ( .A(_5537_), .B(_5739__bF_buf4), .Y(_5538_) );
AND2X2 AND2X2_1024 ( .A(_5535_), .B(_5538_), .Y(_5539_) );
AND2X2 AND2X2_1025 ( .A(_5539_), .B(_5530_), .Y(_5540_) );
AND2X2 AND2X2_1026 ( .A(_5529_), .B(_5540_), .Y(_5541_) );
OR2X2 OR2X2_854 ( .A(_5217_), .B(_5046_), .Y(_5542_) );
MUX2X1 MUX2X1_738 ( .A(_5170_), .B(_5115_), .S(_5682__bF_buf6), .Y(_5543_) );
MUX2X1 MUX2X1_739 ( .A(_5286_), .B(_5229_), .S(_5682__bF_buf6), .Y(_5544_) );
MUX2X1 MUX2X1_740 ( .A(_5544_), .B(_5543_), .S(_5681__bF_buf5), .Y(_5546_) );
AND2X2 AND2X2_1027 ( .A(_5546_), .B(ULA_B_3_bF_buf0), .Y(_5547_) );
MUX2X1 MUX2X1_741 ( .A(ULA_A_28_), .B(ULA_A_29_), .S(ULA_B_0_bF_buf5), .Y(_5548_) );
AND2X2 AND2X2_1028 ( .A(_5548_), .B(_5682__bF_buf1), .Y(_5549_) );
AND2X2 AND2X2_1029 ( .A(_5468_), .B(ULA_B_1_bF_buf0), .Y(_5550_) );
OR2X2 OR2X2_855 ( .A(_5549_), .B(_5550_), .Y(_5551_) );
AND2X2 AND2X2_1030 ( .A(_5551_), .B(_5681__bF_buf3), .Y(_5552_) );
AND2X2 AND2X2_1031 ( .A(_5410_), .B(ULA_B_2_bF_buf1), .Y(_5553_) );
OR2X2 OR2X2_856 ( .A(_5552_), .B(_5553_), .Y(_5554_) );
AND2X2 AND2X2_1032 ( .A(_5554_), .B(_5289__bF_buf4), .Y(_5555_) );
OR2X2 OR2X2_857 ( .A(_5945__bF_buf3), .B(_5555_), .Y(_5557_) );
OR2X2 OR2X2_858 ( .A(_5557_), .B(_5547_), .Y(_5558_) );
AND2X2 AND2X2_1033 ( .A(_5558_), .B(_5542_), .Y(_5559_) );
AND2X2 AND2X2_1034 ( .A(_5541_), .B(_5559_), .Y(_5560_) );
OR2X2 OR2X2_859 ( .A(_5528_), .B(_5560_), .Y(_5561_) );
INVX1 INVX1_52 ( .A(_5561_), .Y(ULA_ULA_OUT_29_) );
NOR2X1 NOR2X1_78 ( .A(_5739__bF_buf7), .B(ULA_OUT_0__30_), .Y(_5562_) );
MUX2X1 MUX2X1_742 ( .A(_5451_), .B(_5378_), .S(_5682__bF_buf0), .Y(_5563_) );
MUX2X1 MUX2X1_743 ( .A(ULA_A_29_), .B(ULA_A_30_), .S(ULA_B_0_bF_buf4), .Y(_5564_) );
MUX2X1 MUX2X1_744 ( .A(_5564_), .B(_5501_), .S(_5682__bF_buf0), .Y(_5565_) );
MUX2X1 MUX2X1_745 ( .A(_5565_), .B(_5563_), .S(_5681__bF_buf0), .Y(_5567_) );
AND2X2 AND2X2_1035 ( .A(_5567_), .B(_5289__bF_buf6), .Y(_5568_) );
AND2X2 AND2X2_1036 ( .A(_5320_), .B(ULA_B_3_bF_buf2), .Y(_5569_) );
OR2X2 OR2X2_860 ( .A(_5569_), .B(_5568_), .Y(_5570_) );
OR2X2 OR2X2_861 ( .A(_5945__bF_buf1), .B(_5570_), .Y(_5571_) );
NAND3X1 NAND3X1_58 ( .A(_6253_), .B(_5289__bF_buf2), .C(_5065_), .Y(_5572_) );
OR2X2 OR2X2_862 ( .A(ULA_A_30_), .B(ULA_B_30_), .Y(_5573_) );
NAND2X1 NAND2X1_702 ( .A(ULA_A_30_), .B(ULA_B_30_), .Y(_5574_) );
AND2X2 AND2X2_1037 ( .A(_5735__bF_buf1), .B(_5574_), .Y(_5575_) );
OAI21X1 OAI21X1_17 ( .A(_5575_), .B(_5734__bF_buf3), .C(_5573_), .Y(_5576_) );
NAND3X1 NAND3X1_59 ( .A(ULA_cin_bF_buf4), .B(ULA_A_30_), .C(ULA_B_30_), .Y(_5578_) );
NAND2X1 NAND2X1_703 ( .A(_5438__bF_buf1), .B(_5574_), .Y(_5579_) );
NAND3X1 NAND3X1_60 ( .A(_5579_), .B(_5740__bF_buf0), .C(_5578_), .Y(_5580_) );
AND2X2 AND2X2_1038 ( .A(_5580_), .B(_5739__bF_buf7), .Y(_5581_) );
AND2X2 AND2X2_1039 ( .A(_5581_), .B(_5576_), .Y(_5582_) );
AND2X2 AND2X2_1040 ( .A(_5572_), .B(_5582_), .Y(_5583_) );
AND2X2 AND2X2_1041 ( .A(_5571_), .B(_5583_), .Y(_5584_) );
OR2X2 OR2X2_863 ( .A(_5217_), .B(_5078_), .Y(_5585_) );
OR2X2 OR2X2_864 ( .A(_6221_), .B(_6144_), .Y(_5586_) );
AND2X2 AND2X2_1042 ( .A(_5585_), .B(_5586_), .Y(_5587_) );
AND2X2 AND2X2_1043 ( .A(_5584_), .B(_5587_), .Y(_5589_) );
OR2X2 OR2X2_865 ( .A(_5562_), .B(_5589_), .Y(_5590_) );
INVX1 INVX1_53 ( .A(_5590_), .Y(ULA_ULA_OUT_30_) );
NOR2X1 NOR2X1_79 ( .A(_5739__bF_buf4), .B(ULA_OUT_0__31_), .Y(_5591_) );
NOR2X1 NOR2X1_80 ( .A(ULA_A_31_), .B(ULA_B_31_), .Y(_5592_) );
NAND2X1 NAND2X1_704 ( .A(ULA_A_31_), .B(ULA_B_31_), .Y(_5593_) );
AOI21X1 AOI21X1_26 ( .A(_5593_), .B(_5735__bF_buf0), .C(_5734__bF_buf0), .Y(_5594_) );
OR2X2 OR2X2_866 ( .A(_5592_), .B(_5594_), .Y(_5595_) );
XOR2X1 XOR2X1_27 ( .A(ULA_cin_bF_buf7), .B(_5593_), .Y(_5596_) );
OR2X2 OR2X2_867 ( .A(_5596_), .B(_5940_), .Y(_5597_) );
AND2X2 AND2X2_1044 ( .A(_5597_), .B(_5739__bF_buf4), .Y(_5599_) );
AND2X2 AND2X2_1045 ( .A(_5595_), .B(_5599_), .Y(_5600_) );
INVX1 INVX1_54 ( .A(_5100_), .Y(_5601_) );
INVX1 INVX1_55 ( .A(_5675_), .Y(_5602_) );
AOI22X1 AOI22X1_1 ( .A(_5669__bF_buf0), .B(_5705_), .C(_5602_), .D(_5672_), .Y(_5603_) );
OR2X2 OR2X2_868 ( .A(_5601_), .B(_5603_), .Y(_5604_) );
AND2X2 AND2X2_1046 ( .A(_5604_), .B(_5600_), .Y(_5605_) );
OR2X2 OR2X2_869 ( .A(_5217_), .B(_5121_), .Y(_5606_) );
AND2X2 AND2X2_1047 ( .A(_5351_), .B(ULA_B_3_bF_buf1), .Y(_5607_) );
AOI21X1 AOI21X1_27 ( .A(ULA_B_0_bF_buf1), .B(ULA_A_30_), .C(ULA_B_1_bF_buf4), .Y(_5608_) );
AND2X2 AND2X2_1048 ( .A(_5548_), .B(ULA_B_1_bF_buf4), .Y(_5610_) );
OR2X2 OR2X2_870 ( .A(_5608_), .B(_5610_), .Y(_5611_) );
OR2X2 OR2X2_871 ( .A(_5300_), .B(_5099_), .Y(_5612_) );
AND2X2 AND2X2_1049 ( .A(_5612_), .B(_5681__bF_buf3), .Y(_5613_) );
AND2X2 AND2X2_1050 ( .A(_5611_), .B(_5613_), .Y(_5614_) );
AND2X2 AND2X2_1051 ( .A(_5471_), .B(ULA_B_2_bF_buf4), .Y(_5615_) );
OR2X2 OR2X2_872 ( .A(_5614_), .B(_5615_), .Y(_5616_) );
AND2X2 AND2X2_1052 ( .A(_5616_), .B(_5289__bF_buf4), .Y(_5617_) );
OR2X2 OR2X2_873 ( .A(_5945__bF_buf3), .B(_5617_), .Y(_5618_) );
OR2X2 OR2X2_874 ( .A(_5607_), .B(_5618_), .Y(_5619_) );
AND2X2 AND2X2_1053 ( .A(_5606_), .B(_5619_), .Y(_5621_) );
AND2X2 AND2X2_1054 ( .A(_5621_), .B(_5605_), .Y(_5622_) );
OR2X2 OR2X2_875 ( .A(_5591_), .B(_5622_), .Y(_5623_) );
INVX1 INVX1_56 ( .A(_5623_), .Y(ULA_ULA_OUT_31_) );
AND2X2 AND2X2_1055 ( .A(_6418_), .B(_6457_), .Y(_5624_) );
AND2X2 AND2X2_1056 ( .A(_4978_), .B(_5019_), .Y(_5625_) );
AND2X2 AND2X2_1057 ( .A(_5625_), .B(_5624_), .Y(_5626_) );
AND2X2 AND2X2_1058 ( .A(_5059_), .B(_5097_), .Y(_5627_) );
AND2X2 AND2X2_1059 ( .A(_5627_), .B(_5136_), .Y(_5628_) );
AND2X2 AND2X2_1060 ( .A(_5626_), .B(_5628_), .Y(_5629_) );
AND2X2 AND2X2_1061 ( .A(_5889_), .B(_6000_), .Y(_5631_) );
AND2X2 AND2X2_1062 ( .A(_6093_), .B(_6158_), .Y(_5632_) );
AND2X2 AND2X2_1063 ( .A(_5632_), .B(_5631_), .Y(_5633_) );
AND2X2 AND2X2_1064 ( .A(_6377_), .B(_6336_), .Y(_5634_) );
AND2X2 AND2X2_1065 ( .A(_6218_), .B(_6277_), .Y(_5635_) );
AND2X2 AND2X2_1066 ( .A(_5635_), .B(_5634_), .Y(_5636_) );
AND2X2 AND2X2_1067 ( .A(_5636_), .B(_5633_), .Y(_5637_) );
AND2X2 AND2X2_1068 ( .A(_5637_), .B(_5629_), .Y(_5638_) );
AND2X2 AND2X2_1069 ( .A(_5400_), .B(_5433_), .Y(_5639_) );
AND2X2 AND2X2_1070 ( .A(_5464_), .B(_5498_), .Y(_5640_) );
AND2X2 AND2X2_1071 ( .A(_5639_), .B(_5640_), .Y(_5642_) );
AND2X2 AND2X2_1072 ( .A(_5309_), .B(_5340_), .Y(_5643_) );
AND2X2 AND2X2_1073 ( .A(_5372_), .B(_5281_), .Y(_5644_) );
AND2X2 AND2X2_1074 ( .A(_5643_), .B(_5644_), .Y(_5645_) );
AND2X2 AND2X2_1075 ( .A(_5645_), .B(_5642_), .Y(_5646_) );
AND2X2 AND2X2_1076 ( .A(_5590_), .B(_5623_), .Y(_5647_) );
AND2X2 AND2X2_1077 ( .A(_5527_), .B(_5561_), .Y(_5648_) );
AND2X2 AND2X2_1078 ( .A(_5648_), .B(_5647_), .Y(_5649_) );
AND2X2 AND2X2_1079 ( .A(_5649_), .B(_5767_), .Y(_5650_) );
AND2X2 AND2X2_1080 ( .A(_5251_), .B(_5223_), .Y(_5651_) );
AND2X2 AND2X2_1081 ( .A(_5192_), .B(_5165_), .Y(_5653_) );
AND2X2 AND2X2_1082 ( .A(_5653_), .B(_5651_), .Y(_5654_) );
AND2X2 AND2X2_1083 ( .A(_5650_), .B(_5654_), .Y(_5655_) );
AND2X2 AND2X2_1084 ( .A(_5655_), .B(_5646_), .Y(_5656_) );
AND2X2 AND2X2_1085 ( .A(_5638_), .B(_5656_), .Y(ULA_zero) );
XOR2X1 XOR2X1_28 ( .A(ULA_B_0_bF_buf6), .B(ULA_A_0_), .Y(ULA_OUT_0__0_) );
MUX2X1 MUX2X1_746 ( .A(ULA_A_0_), .B(ULA_cin_bF_buf3), .S(ULA_B_0_bF_buf6), .Y(_6477_) );
XNOR2X1 XNOR2X1_3 ( .A(ULA_cin_bF_buf2), .B(ULA_B_1_bF_buf7), .Y(_6478_) );
XOR2X1 XOR2X1_29 ( .A(ULA_A_1_), .B(_6478_), .Y(_6479_) );
XOR2X1 XOR2X1_30 ( .A(_6477_), .B(_6479_), .Y(ULA_OUT_0__1_) );
INVX1 INVX1_57 ( .A(ULA_A_1_), .Y(_6480_) );
OR2X2 OR2X2_876 ( .A(_6480_), .B(_6478_), .Y(_6481_) );
OR2X2 OR2X2_877 ( .A(_6477_), .B(_6479_), .Y(_6482_) );
AND2X2 AND2X2_1086 ( .A(_6482_), .B(_6481_), .Y(_6483_) );
XNOR2X1 XNOR2X1_4 ( .A(ULA_cin_bF_buf2), .B(ULA_B_2_bF_buf7), .Y(_6484_) );
XOR2X1 XOR2X1_31 ( .A(ULA_A_2_), .B(_6484_), .Y(_6485_) );
XOR2X1 XOR2X1_32 ( .A(_6485_), .B(_6483_), .Y(ULA_OUT_0__2_) );
INVX1 INVX1_58 ( .A(ULA_A_2_), .Y(_6486_) );
OR2X2 OR2X2_878 ( .A(_6486_), .B(_6484_), .Y(_6487_) );
OR2X2 OR2X2_879 ( .A(_6485_), .B(_6483_), .Y(_6488_) );
AND2X2 AND2X2_1087 ( .A(_6488_), .B(_6487_), .Y(_6489_) );
INVX1 INVX1_59 ( .A(ULA_A_3_), .Y(_6490_) );
XNOR2X1 XNOR2X1_5 ( .A(ULA_cin_bF_buf6), .B(ULA_B_3_bF_buf6), .Y(_6491_) );
OR2X2 OR2X2_880 ( .A(_6490_), .B(_6491_), .Y(_6492_) );
NAND2X1 NAND2X1_705 ( .A(_6490_), .B(_6491_), .Y(_6493_) );
NAND2X1 NAND2X1_706 ( .A(_6492_), .B(_6493_), .Y(_6494_) );
XOR2X1 XOR2X1_33 ( .A(_6494_), .B(_6489_), .Y(ULA_OUT_0__3_) );
OR2X2 OR2X2_881 ( .A(_6494_), .B(_6489_), .Y(_6495_) );
AND2X2 AND2X2_1088 ( .A(_6495_), .B(_6492_), .Y(_6496_) );
INVX1 INVX1_60 ( .A(ULA_A_4_), .Y(_6497_) );
XNOR2X1 XNOR2X1_6 ( .A(ULA_cin_bF_buf6), .B(ULA_B_4_bF_buf3), .Y(_6498_) );
OR2X2 OR2X2_882 ( .A(_6497_), .B(_6498_), .Y(_6499_) );
NAND2X1 NAND2X1_707 ( .A(_6497_), .B(_6498_), .Y(_6500_) );
NAND2X1 NAND2X1_708 ( .A(_6499_), .B(_6500_), .Y(_6501_) );
XOR2X1 XOR2X1_34 ( .A(_6501_), .B(_6496_), .Y(ULA_OUT_0__4_) );
OR2X2 OR2X2_883 ( .A(_6501_), .B(_6496_), .Y(_6502_) );
AND2X2 AND2X2_1089 ( .A(_6502_), .B(_6499_), .Y(_6503_) );
INVX1 INVX1_61 ( .A(ULA_A_5_), .Y(_6504_) );
XNOR2X1 XNOR2X1_7 ( .A(ULA_cin_bF_buf3), .B(ULA_B_5_), .Y(_6505_) );
OR2X2 OR2X2_884 ( .A(_6504_), .B(_6505_), .Y(_6506_) );
NAND2X1 NAND2X1_709 ( .A(_6504_), .B(_6505_), .Y(_6507_) );
NAND2X1 NAND2X1_710 ( .A(_6506_), .B(_6507_), .Y(_6508_) );
XOR2X1 XOR2X1_35 ( .A(_6508_), .B(_6503_), .Y(ULA_OUT_0__5_) );
OR2X2 OR2X2_885 ( .A(_6508_), .B(_6503_), .Y(_6509_) );
AND2X2 AND2X2_1090 ( .A(_6509_), .B(_6506_), .Y(_6510_) );
INVX1 INVX1_62 ( .A(ULA_A_6_), .Y(_6511_) );
XNOR2X1 XNOR2X1_8 ( .A(ULA_cin_bF_buf5), .B(ULA_B_6_), .Y(_6512_) );
NOR2X1 NOR2X1_81 ( .A(_6512_), .B(_6511_), .Y(_6513_) );
INVX1 INVX1_63 ( .A(_6513_), .Y(_6514_) );
NAND2X1 NAND2X1_711 ( .A(_6511_), .B(_6512_), .Y(_6515_) );
NAND2X1 NAND2X1_712 ( .A(_6515_), .B(_6514_), .Y(_6516_) );
XOR2X1 XOR2X1_36 ( .A(_6516_), .B(_6510_), .Y(ULA_OUT_0__6_) );
OR2X2 OR2X2_886 ( .A(_6516_), .B(_6510_), .Y(_6517_) );
AND2X2 AND2X2_1091 ( .A(_6517_), .B(_6514_), .Y(_6518_) );
INVX1 INVX1_64 ( .A(ULA_A_7_), .Y(_6519_) );
XNOR2X1 XNOR2X1_9 ( .A(ULA_cin_bF_buf5), .B(ULA_B_7_), .Y(_6520_) );
NOR2X1 NOR2X1_82 ( .A(_6520_), .B(_6519_), .Y(_6521_) );
INVX1 INVX1_65 ( .A(_6521_), .Y(_6522_) );
NAND2X1 NAND2X1_713 ( .A(_6519_), .B(_6520_), .Y(_6523_) );
NAND2X1 NAND2X1_714 ( .A(_6523_), .B(_6522_), .Y(_6524_) );
XOR2X1 XOR2X1_37 ( .A(_6524_), .B(_6518_), .Y(ULA_OUT_0__7_) );
OR2X2 OR2X2_887 ( .A(_6524_), .B(_6518_), .Y(_6525_) );
AND2X2 AND2X2_1092 ( .A(_6525_), .B(_6522_), .Y(_6526_) );
XNOR2X1 XNOR2X1_10 ( .A(ULA_cin_bF_buf5), .B(ULA_B_8_), .Y(_6527_) );
XNOR2X1 XNOR2X1_11 ( .A(ULA_A_8_), .B(_6527_), .Y(_6528_) );
INVX1 INVX1_66 ( .A(_6528_), .Y(_6529_) );
XOR2X1 XOR2X1_38 ( .A(_6529_), .B(_6526_), .Y(ULA_OUT_0__8_) );
INVX1 INVX1_67 ( .A(ULA_A_8_), .Y(_6530_) );
NOR2X1 NOR2X1_83 ( .A(_6527_), .B(_6530_), .Y(_6531_) );
INVX1 INVX1_68 ( .A(_6531_), .Y(_6532_) );
OR2X2 OR2X2_888 ( .A(_6529_), .B(_6526_), .Y(_6533_) );
AND2X2 AND2X2_1093 ( .A(_6533_), .B(_6532_), .Y(_6534_) );
XNOR2X1 XNOR2X1_12 ( .A(ULA_cin_bF_buf5), .B(ULA_B_9_), .Y(_6535_) );
XNOR2X1 XNOR2X1_13 ( .A(ULA_A_9_), .B(_6535_), .Y(_6536_) );
INVX1 INVX1_69 ( .A(_6536_), .Y(_6537_) );
XOR2X1 XOR2X1_39 ( .A(_6537_), .B(_6534_), .Y(ULA_OUT_0__9_) );
INVX1 INVX1_70 ( .A(ULA_A_9_), .Y(_6538_) );
NOR2X1 NOR2X1_84 ( .A(_6535_), .B(_6538_), .Y(_6539_) );
INVX1 INVX1_71 ( .A(_6539_), .Y(_6540_) );
OR2X2 OR2X2_889 ( .A(_6537_), .B(_6534_), .Y(_6541_) );
AND2X2 AND2X2_1094 ( .A(_6541_), .B(_6540_), .Y(_6542_) );
XNOR2X1 XNOR2X1_14 ( .A(ULA_cin_bF_buf5), .B(ULA_B_10_), .Y(_6543_) );
XNOR2X1 XNOR2X1_15 ( .A(ULA_A_10_), .B(_6543_), .Y(_6544_) );
INVX1 INVX1_72 ( .A(_6544_), .Y(_6545_) );
XOR2X1 XOR2X1_40 ( .A(_6545_), .B(_6542_), .Y(ULA_OUT_0__10_) );
INVX1 INVX1_73 ( .A(ULA_A_10_), .Y(_6546_) );
NOR2X1 NOR2X1_85 ( .A(_6543_), .B(_6546_), .Y(_6547_) );
INVX1 INVX1_74 ( .A(_6547_), .Y(_6548_) );
OR2X2 OR2X2_890 ( .A(_6545_), .B(_6542_), .Y(_6549_) );
AND2X2 AND2X2_1095 ( .A(_6549_), .B(_6548_), .Y(_6550_) );
XNOR2X1 XNOR2X1_16 ( .A(ULA_cin_bF_buf6), .B(ULA_B_11_), .Y(_6551_) );
XNOR2X1 XNOR2X1_17 ( .A(ULA_A_11_), .B(_6551_), .Y(_6552_) );
INVX1 INVX1_75 ( .A(_6552_), .Y(_6553_) );
XOR2X1 XOR2X1_41 ( .A(_6553_), .B(_6550_), .Y(ULA_OUT_0__11_) );
INVX1 INVX1_76 ( .A(ULA_A_11_), .Y(_6554_) );
NOR2X1 NOR2X1_86 ( .A(_6551_), .B(_6554_), .Y(_6555_) );
INVX1 INVX1_77 ( .A(_6555_), .Y(_6556_) );
OR2X2 OR2X2_891 ( .A(_6553_), .B(_6550_), .Y(_6557_) );
AND2X2 AND2X2_1096 ( .A(_6557_), .B(_6556_), .Y(_6558_) );
XNOR2X1 XNOR2X1_18 ( .A(ULA_cin_bF_buf1), .B(ULA_B_12_), .Y(_6559_) );
XNOR2X1 XNOR2X1_19 ( .A(ULA_A_12_), .B(_6559_), .Y(_6560_) );
INVX1 INVX1_78 ( .A(_6560_), .Y(_6561_) );
XOR2X1 XOR2X1_42 ( .A(_6561_), .B(_6558_), .Y(ULA_OUT_0__12_) );
INVX1 INVX1_79 ( .A(ULA_A_12_), .Y(_6562_) );
NOR2X1 NOR2X1_87 ( .A(_6559_), .B(_6562_), .Y(_6563_) );
INVX1 INVX1_80 ( .A(_6563_), .Y(_6564_) );
OR2X2 OR2X2_892 ( .A(_6561_), .B(_6558_), .Y(_6565_) );
AND2X2 AND2X2_1097 ( .A(_6565_), .B(_6564_), .Y(_6566_) );
XNOR2X1 XNOR2X1_20 ( .A(ULA_cin_bF_buf1), .B(ULA_B_13_), .Y(_6567_) );
XNOR2X1 XNOR2X1_21 ( .A(ULA_A_13_), .B(_6567_), .Y(_6568_) );
INVX1 INVX1_81 ( .A(_6568_), .Y(_6569_) );
XOR2X1 XOR2X1_43 ( .A(_6569_), .B(_6566_), .Y(ULA_OUT_0__13_) );
INVX1 INVX1_82 ( .A(ULA_A_13_), .Y(_6570_) );
NOR2X1 NOR2X1_88 ( .A(_6567_), .B(_6570_), .Y(_6571_) );
INVX1 INVX1_83 ( .A(_6571_), .Y(_6572_) );
OR2X2 OR2X2_893 ( .A(_6569_), .B(_6566_), .Y(_6573_) );
AND2X2 AND2X2_1098 ( .A(_6573_), .B(_6572_), .Y(_6574_) );
XNOR2X1 XNOR2X1_22 ( .A(ULA_cin_bF_buf6), .B(ULA_B_14_), .Y(_6575_) );
XNOR2X1 XNOR2X1_23 ( .A(ULA_A_14_), .B(_6575_), .Y(_6576_) );
INVX1 INVX1_84 ( .A(_6576_), .Y(_6577_) );
XOR2X1 XOR2X1_44 ( .A(_6577_), .B(_6574_), .Y(ULA_OUT_0__14_) );
INVX1 INVX1_85 ( .A(ULA_A_14_), .Y(_6578_) );
NOR2X1 NOR2X1_89 ( .A(_6575_), .B(_6578_), .Y(_6579_) );
INVX1 INVX1_86 ( .A(_6579_), .Y(_6580_) );
OR2X2 OR2X2_894 ( .A(_6577_), .B(_6574_), .Y(_6581_) );
AND2X2 AND2X2_1099 ( .A(_6581_), .B(_6580_), .Y(_6582_) );
XNOR2X1 XNOR2X1_24 ( .A(ULA_cin_bF_buf1), .B(ULA_B_15_), .Y(_6583_) );
XNOR2X1 XNOR2X1_25 ( .A(ULA_A_15_), .B(_6583_), .Y(_6584_) );
INVX1 INVX1_87 ( .A(_6584_), .Y(_6585_) );
XOR2X1 XOR2X1_45 ( .A(_6585_), .B(_6582_), .Y(ULA_OUT_0__15_) );
INVX1 INVX1_88 ( .A(ULA_A_15_), .Y(_6586_) );
NOR2X1 NOR2X1_90 ( .A(_6583_), .B(_6586_), .Y(_6587_) );
INVX1 INVX1_89 ( .A(_6587_), .Y(_6588_) );
OR2X2 OR2X2_895 ( .A(_6585_), .B(_6582_), .Y(_6589_) );
AND2X2 AND2X2_1100 ( .A(_6589_), .B(_6588_), .Y(_6590_) );
XNOR2X1 XNOR2X1_26 ( .A(ULA_cin_bF_buf1), .B(ULA_B_16_), .Y(_6591_) );
XNOR2X1 XNOR2X1_27 ( .A(ULA_A_16_), .B(_6591_), .Y(_6592_) );
INVX1 INVX1_90 ( .A(_6592_), .Y(_6593_) );
XOR2X1 XOR2X1_46 ( .A(_6593_), .B(_6590_), .Y(ULA_OUT_0__16_) );
INVX1 INVX1_91 ( .A(ULA_A_16_), .Y(_6594_) );
NOR2X1 NOR2X1_91 ( .A(_6591_), .B(_6594_), .Y(_6595_) );
INVX1 INVX1_92 ( .A(_6595_), .Y(_6596_) );
OR2X2 OR2X2_896 ( .A(_6593_), .B(_6590_), .Y(_6597_) );
AND2X2 AND2X2_1101 ( .A(_6597_), .B(_6596_), .Y(_6598_) );
XNOR2X1 XNOR2X1_28 ( .A(ULA_cin_bF_buf7), .B(ULA_B_17_), .Y(_6599_) );
XNOR2X1 XNOR2X1_29 ( .A(ULA_A_17_), .B(_6599_), .Y(_6600_) );
INVX1 INVX1_93 ( .A(_6600_), .Y(_6601_) );
XOR2X1 XOR2X1_47 ( .A(_6601_), .B(_6598_), .Y(ULA_OUT_0__17_) );
INVX1 INVX1_94 ( .A(ULA_A_17_), .Y(_6602_) );
NOR2X1 NOR2X1_92 ( .A(_6599_), .B(_6602_), .Y(_6603_) );
INVX1 INVX1_95 ( .A(_6603_), .Y(_6604_) );
OR2X2 OR2X2_897 ( .A(_6601_), .B(_6598_), .Y(_6605_) );
AND2X2 AND2X2_1102 ( .A(_6605_), .B(_6604_), .Y(_6606_) );
XNOR2X1 XNOR2X1_30 ( .A(ULA_cin_bF_buf7), .B(ULA_B_18_), .Y(_6607_) );
XNOR2X1 XNOR2X1_31 ( .A(ULA_A_18_), .B(_6607_), .Y(_6608_) );
INVX1 INVX1_96 ( .A(_6608_), .Y(_6609_) );
XOR2X1 XOR2X1_48 ( .A(_6609_), .B(_6606_), .Y(ULA_OUT_0__18_) );
INVX1 INVX1_97 ( .A(ULA_A_18_), .Y(_6610_) );
NOR2X1 NOR2X1_93 ( .A(_6607_), .B(_6610_), .Y(_6611_) );
INVX1 INVX1_98 ( .A(_6611_), .Y(_6612_) );
OR2X2 OR2X2_898 ( .A(_6609_), .B(_6606_), .Y(_6613_) );
AND2X2 AND2X2_1103 ( .A(_6613_), .B(_6612_), .Y(_6614_) );
XNOR2X1 XNOR2X1_32 ( .A(ULA_cin_bF_buf7), .B(ULA_B_19_), .Y(_6615_) );
XNOR2X1 XNOR2X1_33 ( .A(ULA_A_19_), .B(_6615_), .Y(_6616_) );
INVX1 INVX1_99 ( .A(_6616_), .Y(_6617_) );
XOR2X1 XOR2X1_49 ( .A(_6617_), .B(_6614_), .Y(ULA_OUT_0__19_) );
INVX1 INVX1_100 ( .A(ULA_A_19_), .Y(_6618_) );
NOR2X1 NOR2X1_94 ( .A(_6615_), .B(_6618_), .Y(_6619_) );
INVX1 INVX1_101 ( .A(_6619_), .Y(_6620_) );
OR2X2 OR2X2_899 ( .A(_6617_), .B(_6614_), .Y(_6621_) );
AND2X2 AND2X2_1104 ( .A(_6621_), .B(_6620_), .Y(_6622_) );
XNOR2X1 XNOR2X1_34 ( .A(ULA_cin_bF_buf1), .B(ULA_B_20_), .Y(_6623_) );
XNOR2X1 XNOR2X1_35 ( .A(ULA_A_20_), .B(_6623_), .Y(_6624_) );
INVX1 INVX1_102 ( .A(_6624_), .Y(_6625_) );
XOR2X1 XOR2X1_50 ( .A(_6625_), .B(_6622_), .Y(ULA_OUT_0__20_) );
INVX1 INVX1_103 ( .A(ULA_A_20_), .Y(_6626_) );
NOR2X1 NOR2X1_95 ( .A(_6623_), .B(_6626_), .Y(_6627_) );
INVX1 INVX1_104 ( .A(_6627_), .Y(_6628_) );
OR2X2 OR2X2_900 ( .A(_6625_), .B(_6622_), .Y(_6629_) );
AND2X2 AND2X2_1105 ( .A(_6629_), .B(_6628_), .Y(_6630_) );
XNOR2X1 XNOR2X1_36 ( .A(ULA_cin_bF_buf0), .B(ULA_B_21_), .Y(_6631_) );
XNOR2X1 XNOR2X1_37 ( .A(ULA_A_21_), .B(_6631_), .Y(_6632_) );
INVX1 INVX1_105 ( .A(_6632_), .Y(_6633_) );
XOR2X1 XOR2X1_51 ( .A(_6633_), .B(_6630_), .Y(ULA_OUT_0__21_) );
INVX1 INVX1_106 ( .A(ULA_A_21_), .Y(_6634_) );
NOR2X1 NOR2X1_96 ( .A(_6631_), .B(_6634_), .Y(_6635_) );
INVX1 INVX1_107 ( .A(_6635_), .Y(_6636_) );
OR2X2 OR2X2_901 ( .A(_6633_), .B(_6630_), .Y(_6637_) );
AND2X2 AND2X2_1106 ( .A(_6637_), .B(_6636_), .Y(_6638_) );
XNOR2X1 XNOR2X1_38 ( .A(ULA_cin_bF_buf0), .B(ULA_B_22_), .Y(_6639_) );
XNOR2X1 XNOR2X1_39 ( .A(ULA_A_22_), .B(_6639_), .Y(_6640_) );
INVX1 INVX1_108 ( .A(_6640_), .Y(_6641_) );
XOR2X1 XOR2X1_52 ( .A(_6641_), .B(_6638_), .Y(ULA_OUT_0__22_) );
INVX1 INVX1_109 ( .A(ULA_A_22_), .Y(_6642_) );
NOR2X1 NOR2X1_97 ( .A(_6639_), .B(_6642_), .Y(_6643_) );
INVX1 INVX1_110 ( .A(_6643_), .Y(_6644_) );
OR2X2 OR2X2_902 ( .A(_6641_), .B(_6638_), .Y(_6645_) );
AND2X2 AND2X2_1107 ( .A(_6645_), .B(_6644_), .Y(_6646_) );
XNOR2X1 XNOR2X1_40 ( .A(ULA_cin_bF_buf4), .B(ULA_B_23_), .Y(_6647_) );
XNOR2X1 XNOR2X1_41 ( .A(ULA_A_23_), .B(_6647_), .Y(_6648_) );
INVX1 INVX1_111 ( .A(_6648_), .Y(_6649_) );
XOR2X1 XOR2X1_53 ( .A(_6649_), .B(_6646_), .Y(ULA_OUT_0__23_) );
INVX1 INVX1_112 ( .A(ULA_A_23_), .Y(_6650_) );
NOR2X1 NOR2X1_98 ( .A(_6647_), .B(_6650_), .Y(_6651_) );
INVX1 INVX1_113 ( .A(_6651_), .Y(_6652_) );
OR2X2 OR2X2_903 ( .A(_6649_), .B(_6646_), .Y(_6653_) );
AND2X2 AND2X2_1108 ( .A(_6653_), .B(_6652_), .Y(_6654_) );
XNOR2X1 XNOR2X1_42 ( .A(ULA_cin_bF_buf0), .B(ULA_B_24_), .Y(_6655_) );
XNOR2X1 XNOR2X1_43 ( .A(ULA_A_24_), .B(_6655_), .Y(_6656_) );
INVX1 INVX1_114 ( .A(_6656_), .Y(_6657_) );
XOR2X1 XOR2X1_54 ( .A(_6657_), .B(_6654_), .Y(ULA_OUT_0__24_) );
INVX1 INVX1_115 ( .A(ULA_A_24_), .Y(_6658_) );
NOR2X1 NOR2X1_99 ( .A(_6655_), .B(_6658_), .Y(_6659_) );
INVX1 INVX1_116 ( .A(_6659_), .Y(_6660_) );
OR2X2 OR2X2_904 ( .A(_6657_), .B(_6654_), .Y(_6661_) );
AND2X2 AND2X2_1109 ( .A(_6661_), .B(_6660_), .Y(_6662_) );
XNOR2X1 XNOR2X1_44 ( .A(ULA_cin_bF_buf0), .B(ULA_B_25_), .Y(_6663_) );
XNOR2X1 XNOR2X1_45 ( .A(ULA_A_25_), .B(_6663_), .Y(_6664_) );
INVX1 INVX1_117 ( .A(_6664_), .Y(_6665_) );
XOR2X1 XOR2X1_55 ( .A(_6665_), .B(_6662_), .Y(ULA_OUT_0__25_) );
INVX1 INVX1_118 ( .A(ULA_A_25_), .Y(_6666_) );
NOR2X1 NOR2X1_100 ( .A(_6663_), .B(_6666_), .Y(_6667_) );
INVX1 INVX1_119 ( .A(_6667_), .Y(_6668_) );
OR2X2 OR2X2_905 ( .A(_6665_), .B(_6662_), .Y(_6669_) );
AND2X2 AND2X2_1110 ( .A(_6669_), .B(_6668_), .Y(_6670_) );
XNOR2X1 XNOR2X1_46 ( .A(ULA_cin_bF_buf0), .B(ULA_B_26_), .Y(_6671_) );
XNOR2X1 XNOR2X1_47 ( .A(ULA_A_26_), .B(_6671_), .Y(_6672_) );
INVX1 INVX1_120 ( .A(_6672_), .Y(_6673_) );
XOR2X1 XOR2X1_56 ( .A(_6673_), .B(_6670_), .Y(ULA_OUT_0__26_) );
INVX1 INVX1_121 ( .A(ULA_A_26_), .Y(_6674_) );
NOR2X1 NOR2X1_101 ( .A(_6671_), .B(_6674_), .Y(_6675_) );
INVX1 INVX1_122 ( .A(_6675_), .Y(_6676_) );
OR2X2 OR2X2_906 ( .A(_6673_), .B(_6670_), .Y(_6677_) );
AND2X2 AND2X2_1111 ( .A(_6677_), .B(_6676_), .Y(_6678_) );
XNOR2X1 XNOR2X1_48 ( .A(ULA_cin_bF_buf4), .B(ULA_B_27_), .Y(_6679_) );
XNOR2X1 XNOR2X1_49 ( .A(ULA_A_27_), .B(_6679_), .Y(_6680_) );
INVX1 INVX1_123 ( .A(_6680_), .Y(_6681_) );
XOR2X1 XOR2X1_57 ( .A(_6681_), .B(_6678_), .Y(ULA_OUT_0__27_) );
INVX1 INVX1_124 ( .A(ULA_A_27_), .Y(_6682_) );
NOR2X1 NOR2X1_102 ( .A(_6679_), .B(_6682_), .Y(_6683_) );
INVX1 INVX1_125 ( .A(_6683_), .Y(_6684_) );
OR2X2 OR2X2_907 ( .A(_6681_), .B(_6678_), .Y(_6685_) );
AND2X2 AND2X2_1112 ( .A(_6685_), .B(_6684_), .Y(_6686_) );
XNOR2X1 XNOR2X1_50 ( .A(ULA_cin_bF_buf4), .B(ULA_B_28_), .Y(_6687_) );
XNOR2X1 XNOR2X1_51 ( .A(ULA_A_28_), .B(_6687_), .Y(_6688_) );
INVX1 INVX1_126 ( .A(_6688_), .Y(_6689_) );
XOR2X1 XOR2X1_58 ( .A(_6689_), .B(_6686_), .Y(ULA_OUT_0__28_) );
INVX1 INVX1_127 ( .A(ULA_A_28_), .Y(_6690_) );
NOR2X1 NOR2X1_103 ( .A(_6687_), .B(_6690_), .Y(_6691_) );
INVX1 INVX1_128 ( .A(_6691_), .Y(_6692_) );
OR2X2 OR2X2_908 ( .A(_6689_), .B(_6686_), .Y(_6693_) );
AND2X2 AND2X2_1113 ( .A(_6693_), .B(_6692_), .Y(_6694_) );
XNOR2X1 XNOR2X1_52 ( .A(ULA_cin_bF_buf4), .B(ULA_B_29_), .Y(_6695_) );
XNOR2X1 XNOR2X1_53 ( .A(ULA_A_29_), .B(_6695_), .Y(_6696_) );
INVX1 INVX1_129 ( .A(_6696_), .Y(_6697_) );
XOR2X1 XOR2X1_59 ( .A(_6697_), .B(_6694_), .Y(ULA_OUT_0__29_) );
INVX1 INVX1_130 ( .A(ULA_A_29_), .Y(_6698_) );
NOR2X1 NOR2X1_104 ( .A(_6695_), .B(_6698_), .Y(_6699_) );
INVX1 INVX1_131 ( .A(_6699_), .Y(_6700_) );
OR2X2 OR2X2_909 ( .A(_6697_), .B(_6694_), .Y(_6701_) );
AND2X2 AND2X2_1114 ( .A(_6701_), .B(_6700_), .Y(_6702_) );
XNOR2X1 XNOR2X1_54 ( .A(ULA_cin_bF_buf0), .B(ULA_B_30_), .Y(_6703_) );
XNOR2X1 XNOR2X1_55 ( .A(ULA_A_30_), .B(_6703_), .Y(_6704_) );
INVX1 INVX1_132 ( .A(_6704_), .Y(_6705_) );
XOR2X1 XOR2X1_60 ( .A(_6705_), .B(_6702_), .Y(ULA_OUT_0__30_) );
INVX1 INVX1_133 ( .A(ULA_A_30_), .Y(_6706_) );
NOR2X1 NOR2X1_105 ( .A(_6703_), .B(_6706_), .Y(_6707_) );
INVX1 INVX1_134 ( .A(_6707_), .Y(_6708_) );
OR2X2 OR2X2_910 ( .A(_6705_), .B(_6702_), .Y(_6709_) );
AND2X2 AND2X2_1115 ( .A(_6709_), .B(_6708_), .Y(_6710_) );
XNOR2X1 XNOR2X1_56 ( .A(ULA_cin_bF_buf7), .B(ULA_A_31_), .Y(_6711_) );
XOR2X1 XOR2X1_61 ( .A(ULA_B_31_), .B(_6711_), .Y(_6712_) );
XOR2X1 XOR2X1_62 ( .A(_6712_), .B(_6710_), .Y(ULA_OUT_0__31_) );
INVX1 INVX1_135 ( .A(PC_ULA_OUT_0_), .Y(_0_) );
NAND2X1 NAND2X1_715 ( .A(DDATA_CORE_out[0]), .B(CORE_DATA_REGMux_exec_pipe_bF_buf4), .Y(_1_) );
OAI21X1 OAI21X1_18 ( .A(_0_), .B(CORE_DATA_REGMux_exec_pipe_bF_buf2), .C(_1_), .Y(REG_RD_wb_pipe_0_) );
INVX1 INVX1_136 ( .A(PC_ULA_OUT_1_), .Y(_2_) );
NAND2X1 NAND2X1_716 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(DDATA_CORE_out[1]), .Y(_3_) );
OAI21X1 OAI21X1_19 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_2_), .C(_3_), .Y(REG_RD_wb_pipe_1_) );
INVX1 INVX1_137 ( .A(PC_ULA_OUT_2_), .Y(_4_) );
NAND2X1 NAND2X1_717 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[2]), .Y(_5_) );
OAI21X1 OAI21X1_20 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_4_), .C(_5_), .Y(REG_RD_wb_pipe_2_) );
INVX1 INVX1_138 ( .A(PC_ULA_OUT_3_), .Y(_6_) );
NAND2X1 NAND2X1_718 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(DDATA_CORE_out[3]), .Y(_7_) );
OAI21X1 OAI21X1_21 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_6_), .C(_7_), .Y(REG_RD_wb_pipe_3_) );
INVX1 INVX1_139 ( .A(PC_ULA_OUT_4_), .Y(_8_) );
NAND2X1 NAND2X1_719 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[4]), .Y(_9_) );
OAI21X1 OAI21X1_22 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(_8_), .C(_9_), .Y(REG_RD_wb_pipe_4_) );
INVX1 INVX1_140 ( .A(PC_ULA_OUT_5_), .Y(_10_) );
NAND2X1 NAND2X1_720 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(DDATA_CORE_out[5]), .Y(_11_) );
OAI21X1 OAI21X1_23 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_10_), .C(_11_), .Y(REG_RD_wb_pipe_5_) );
INVX1 INVX1_141 ( .A(PC_ULA_OUT_6_), .Y(_12_) );
NAND2X1 NAND2X1_721 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[6]), .Y(_13_) );
OAI21X1 OAI21X1_24 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(_12_), .C(_13_), .Y(REG_RD_wb_pipe_6_) );
INVX1 INVX1_142 ( .A(PC_ULA_OUT_7_), .Y(_14_) );
NAND2X1 NAND2X1_722 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[7]), .Y(_15_) );
OAI21X1 OAI21X1_25 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(_14_), .C(_15_), .Y(REG_RD_wb_pipe_7_) );
INVX1 INVX1_143 ( .A(ULA_out_exec_pipe_8_), .Y(_16_) );
NAND2X1 NAND2X1_723 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(DDATA_CORE_out[8]), .Y(_17_) );
OAI21X1 OAI21X1_26 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(_16_), .C(_17_), .Y(REG_RD_wb_pipe_8_) );
INVX1 INVX1_144 ( .A(ULA_out_exec_pipe_9_), .Y(_18_) );
NAND2X1 NAND2X1_724 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(DDATA_CORE_out[9]), .Y(_19_) );
OAI21X1 OAI21X1_27 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(_18_), .C(_19_), .Y(REG_RD_wb_pipe_9_) );
INVX1 INVX1_145 ( .A(ULA_out_exec_pipe_10_), .Y(_20_) );
NAND2X1 NAND2X1_725 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(DDATA_CORE_out[10]), .Y(_21_) );
OAI21X1 OAI21X1_28 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(_20_), .C(_21_), .Y(REG_RD_wb_pipe_10_) );
INVX1 INVX1_146 ( .A(ULA_out_exec_pipe_11_), .Y(_22_) );
NAND2X1 NAND2X1_726 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(DDATA_CORE_out[11]), .Y(_23_) );
OAI21X1 OAI21X1_29 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(_22_), .C(_23_), .Y(REG_RD_wb_pipe_11_) );
INVX1 INVX1_147 ( .A(ULA_out_exec_pipe_12_), .Y(_24_) );
NAND2X1 NAND2X1_727 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[12]), .Y(_25_) );
OAI21X1 OAI21X1_30 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(_24_), .C(_25_), .Y(REG_RD_wb_pipe_12_) );
INVX1 INVX1_148 ( .A(ULA_out_exec_pipe_13_), .Y(_26_) );
NAND2X1 NAND2X1_728 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(DDATA_CORE_out[13]), .Y(_27_) );
OAI21X1 OAI21X1_31 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(_26_), .C(_27_), .Y(REG_RD_wb_pipe_13_) );
INVX1 INVX1_149 ( .A(ULA_out_exec_pipe_14_), .Y(_28_) );
NAND2X1 NAND2X1_729 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(DDATA_CORE_out[14]), .Y(_29_) );
OAI21X1 OAI21X1_32 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(_28_), .C(_29_), .Y(REG_RD_wb_pipe_14_) );
INVX1 INVX1_150 ( .A(ULA_out_exec_pipe_15_), .Y(_30_) );
NAND2X1 NAND2X1_730 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(DDATA_CORE_out[15]), .Y(_31_) );
OAI21X1 OAI21X1_33 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(_30_), .C(_31_), .Y(REG_RD_wb_pipe_15_) );
INVX1 INVX1_151 ( .A(ULA_out_exec_pipe_16_), .Y(_32_) );
NAND2X1 NAND2X1_731 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(DDATA_CORE_out[16]), .Y(_33_) );
OAI21X1 OAI21X1_34 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(_32_), .C(_33_), .Y(REG_RD_wb_pipe_16_) );
INVX1 INVX1_152 ( .A(ULA_out_exec_pipe_17_), .Y(_34_) );
NAND2X1 NAND2X1_732 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[17]), .Y(_35_) );
OAI21X1 OAI21X1_35 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(_34_), .C(_35_), .Y(REG_RD_wb_pipe_17_) );
INVX1 INVX1_153 ( .A(ULA_out_exec_pipe_18_), .Y(_36_) );
NAND2X1 NAND2X1_733 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(DDATA_CORE_out[18]), .Y(_37_) );
OAI21X1 OAI21X1_36 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(_36_), .C(_37_), .Y(REG_RD_wb_pipe_18_) );
INVX1 INVX1_154 ( .A(ULA_out_exec_pipe_19_), .Y(_38_) );
NAND2X1 NAND2X1_734 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(DDATA_CORE_out[19]), .Y(_39_) );
OAI21X1 OAI21X1_37 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(_38_), .C(_39_), .Y(REG_RD_wb_pipe_19_) );
INVX1 INVX1_155 ( .A(ULA_out_exec_pipe_20_), .Y(_40_) );
NAND2X1 NAND2X1_735 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(DDATA_CORE_out[20]), .Y(_41_) );
OAI21X1 OAI21X1_38 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(_40_), .C(_41_), .Y(REG_RD_wb_pipe_20_) );
INVX1 INVX1_156 ( .A(ULA_out_exec_pipe_21_), .Y(_42_) );
NAND2X1 NAND2X1_736 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(DDATA_CORE_out[21]), .Y(_43_) );
OAI21X1 OAI21X1_39 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(_42_), .C(_43_), .Y(REG_RD_wb_pipe_21_) );
INVX1 INVX1_157 ( .A(ULA_out_exec_pipe_22_), .Y(_44_) );
NAND2X1 NAND2X1_737 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[22]), .Y(_45_) );
OAI21X1 OAI21X1_40 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(_44_), .C(_45_), .Y(REG_RD_wb_pipe_22_) );
INVX1 INVX1_158 ( .A(ULA_out_exec_pipe_23_), .Y(_46_) );
NAND2X1 NAND2X1_738 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(DDATA_CORE_out[23]), .Y(_47_) );
OAI21X1 OAI21X1_41 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(_46_), .C(_47_), .Y(REG_RD_wb_pipe_23_) );
INVX1 INVX1_159 ( .A(ULA_out_exec_pipe_24_), .Y(_48_) );
NAND2X1 NAND2X1_739 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf3), .B(DDATA_CORE_out[24]), .Y(_49_) );
OAI21X1 OAI21X1_42 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf2), .B(_48_), .C(_49_), .Y(REG_RD_wb_pipe_24_) );
INVX1 INVX1_160 ( .A(ULA_out_exec_pipe_25_), .Y(_50_) );
NAND2X1 NAND2X1_740 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(DDATA_CORE_out[25]), .Y(_51_) );
OAI21X1 OAI21X1_43 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(_50_), .C(_51_), .Y(REG_RD_wb_pipe_25_) );
INVX1 INVX1_161 ( .A(ULA_out_exec_pipe_26_), .Y(_52_) );
NAND2X1 NAND2X1_741 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf0), .B(DDATA_CORE_out[26]), .Y(_53_) );
OAI21X1 OAI21X1_44 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(_52_), .C(_53_), .Y(REG_RD_wb_pipe_26_) );
INVX1 INVX1_162 ( .A(ULA_out_exec_pipe_27_), .Y(_54_) );
NAND2X1 NAND2X1_742 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(DDATA_CORE_out[27]), .Y(_55_) );
OAI21X1 OAI21X1_45 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf4), .B(_54_), .C(_55_), .Y(REG_RD_wb_pipe_27_) );
INVX1 INVX1_163 ( .A(ULA_out_exec_pipe_28_), .Y(_56_) );
NAND2X1 NAND2X1_743 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(DDATA_CORE_out[28]), .Y(_57_) );
OAI21X1 OAI21X1_46 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf1), .B(_56_), .C(_57_), .Y(REG_RD_wb_pipe_28_) );
INVX1 INVX1_164 ( .A(ULA_out_exec_pipe_29_), .Y(_58_) );
NAND2X1 NAND2X1_744 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(DDATA_CORE_out[29]), .Y(_59_) );
OAI21X1 OAI21X1_47 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_58_), .C(_59_), .Y(REG_RD_wb_pipe_29_) );
INVX1 INVX1_165 ( .A(ULA_out_exec_pipe_30_), .Y(_60_) );
NAND2X1 NAND2X1_745 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf7), .B(DDATA_CORE_out[30]), .Y(_61_) );
OAI21X1 OAI21X1_48 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_60_), .C(_61_), .Y(REG_RD_wb_pipe_30_) );
INVX1 INVX1_166 ( .A(ULA_out_exec_pipe_31_), .Y(_62_) );
NAND2X1 NAND2X1_746 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf6), .B(DDATA_CORE_out[31]), .Y(_63_) );
OAI21X1 OAI21X1_49 ( .A(CORE_DATA_REGMux_exec_pipe_bF_buf5), .B(_62_), .C(_63_), .Y(REG_RD_wb_pipe_31_) );
MUX2X1 MUX2X1_747 ( .A(PC_ULA_OUT_0_), .B(REG_B_0_), .S(CORE_ULA_REGB_Stall_bF_buf4), .Y(_64_) );
INVX1 INVX1_167 ( .A(_64_), .Y(_143__0_) );
MUX2X1 MUX2X1_748 ( .A(PC_ULA_OUT_1_), .B(REG_B_1_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_65_) );
INVX1 INVX1_168 ( .A(_65_), .Y(_143__1_) );
MUX2X1 MUX2X1_749 ( .A(PC_ULA_OUT_2_), .B(REG_B_2_), .S(CORE_ULA_REGB_Stall_bF_buf1), .Y(_66_) );
INVX1 INVX1_169 ( .A(_66_), .Y(_143__2_) );
MUX2X1 MUX2X1_750 ( .A(PC_ULA_OUT_3_), .B(REG_B_3_), .S(CORE_ULA_REGB_Stall_bF_buf1), .Y(_67_) );
INVX1 INVX1_170 ( .A(_67_), .Y(_143__3_) );
MUX2X1 MUX2X1_751 ( .A(PC_ULA_OUT_4_), .B(REG_B_4_), .S(CORE_ULA_REGB_Stall_bF_buf1), .Y(_68_) );
INVX1 INVX1_171 ( .A(_68_), .Y(_143__4_) );
MUX2X1 MUX2X1_752 ( .A(PC_ULA_OUT_5_), .B(REG_B_5_), .S(CORE_ULA_REGB_Stall_bF_buf1), .Y(_69_) );
INVX1 INVX1_172 ( .A(_69_), .Y(_143__5_) );
MUX2X1 MUX2X1_753 ( .A(PC_ULA_OUT_6_), .B(REG_B_6_), .S(CORE_ULA_REGB_Stall_bF_buf1), .Y(_70_) );
INVX1 INVX1_173 ( .A(_70_), .Y(_143__6_) );
MUX2X1 MUX2X1_754 ( .A(PC_ULA_OUT_7_), .B(REG_B_7_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_71_) );
INVX1 INVX1_174 ( .A(_71_), .Y(_143__7_) );
MUX2X1 MUX2X1_755 ( .A(ULA_out_exec_pipe_8_), .B(REG_B_8_), .S(CORE_ULA_REGB_Stall_bF_buf4), .Y(_72_) );
INVX1 INVX1_175 ( .A(_72_), .Y(_143__8_) );
MUX2X1 MUX2X1_756 ( .A(ULA_out_exec_pipe_9_), .B(REG_B_9_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_73_) );
INVX1 INVX1_176 ( .A(_73_), .Y(_143__9_) );
MUX2X1 MUX2X1_757 ( .A(ULA_out_exec_pipe_10_), .B(REG_B_10_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_74_) );
INVX1 INVX1_177 ( .A(_74_), .Y(_143__10_) );
MUX2X1 MUX2X1_758 ( .A(ULA_out_exec_pipe_11_), .B(REG_B_11_), .S(CORE_ULA_REGB_Stall_bF_buf4), .Y(_75_) );
INVX1 INVX1_178 ( .A(_75_), .Y(_143__11_) );
MUX2X1 MUX2X1_759 ( .A(ULA_out_exec_pipe_12_), .B(REG_B_12_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_76_) );
INVX1 INVX1_179 ( .A(_76_), .Y(_143__12_) );
MUX2X1 MUX2X1_760 ( .A(ULA_out_exec_pipe_13_), .B(REG_B_13_), .S(CORE_ULA_REGB_Stall_bF_buf0), .Y(_77_) );
INVX1 INVX1_180 ( .A(_77_), .Y(_143__13_) );
MUX2X1 MUX2X1_761 ( .A(ULA_out_exec_pipe_14_), .B(REG_B_14_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_78_) );
INVX1 INVX1_181 ( .A(_78_), .Y(_143__14_) );
MUX2X1 MUX2X1_762 ( .A(ULA_out_exec_pipe_15_), .B(REG_B_15_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_79_) );
INVX1 INVX1_182 ( .A(_79_), .Y(_143__15_) );
MUX2X1 MUX2X1_763 ( .A(ULA_out_exec_pipe_16_), .B(REG_B_16_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_80_) );
INVX1 INVX1_183 ( .A(_80_), .Y(_143__16_) );
MUX2X1 MUX2X1_764 ( .A(ULA_out_exec_pipe_17_), .B(REG_B_17_), .S(CORE_ULA_REGB_Stall_bF_buf0), .Y(_81_) );
INVX1 INVX1_184 ( .A(_81_), .Y(_143__17_) );
MUX2X1 MUX2X1_765 ( .A(ULA_out_exec_pipe_18_), .B(REG_B_18_), .S(CORE_ULA_REGB_Stall_bF_buf4), .Y(_82_) );
INVX1 INVX1_185 ( .A(_82_), .Y(_143__18_) );
MUX2X1 MUX2X1_766 ( .A(ULA_out_exec_pipe_19_), .B(REG_B_19_), .S(CORE_ULA_REGB_Stall_bF_buf4), .Y(_83_) );
INVX1 INVX1_186 ( .A(_83_), .Y(_143__19_) );
MUX2X1 MUX2X1_767 ( .A(ULA_out_exec_pipe_20_), .B(REG_B_20_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_84_) );
INVX1 INVX1_187 ( .A(_84_), .Y(_143__20_) );
MUX2X1 MUX2X1_768 ( .A(ULA_out_exec_pipe_21_), .B(REG_B_21_), .S(CORE_ULA_REGB_Stall_bF_buf0), .Y(_85_) );
INVX1 INVX1_188 ( .A(_85_), .Y(_143__21_) );
MUX2X1 MUX2X1_769 ( .A(ULA_out_exec_pipe_22_), .B(REG_B_22_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_86_) );
INVX1 INVX1_189 ( .A(_86_), .Y(_143__22_) );
MUX2X1 MUX2X1_770 ( .A(ULA_out_exec_pipe_23_), .B(REG_B_23_), .S(CORE_ULA_REGB_Stall_bF_buf4), .Y(_87_) );
INVX1 INVX1_190 ( .A(_87_), .Y(_143__23_) );
MUX2X1 MUX2X1_771 ( .A(ULA_out_exec_pipe_24_), .B(REG_B_24_), .S(CORE_ULA_REGB_Stall_bF_buf0), .Y(_88_) );
INVX1 INVX1_191 ( .A(_88_), .Y(_143__24_) );
MUX2X1 MUX2X1_772 ( .A(ULA_out_exec_pipe_25_), .B(REG_B_25_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_89_) );
INVX1 INVX1_192 ( .A(_89_), .Y(_143__25_) );
MUX2X1 MUX2X1_773 ( .A(ULA_out_exec_pipe_26_), .B(REG_B_26_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_90_) );
INVX1 INVX1_193 ( .A(_90_), .Y(_143__26_) );
MUX2X1 MUX2X1_774 ( .A(ULA_out_exec_pipe_27_), .B(REG_B_27_), .S(CORE_ULA_REGB_Stall_bF_buf3), .Y(_91_) );
INVX1 INVX1_194 ( .A(_91_), .Y(_143__27_) );
MUX2X1 MUX2X1_775 ( .A(ULA_out_exec_pipe_28_), .B(REG_B_28_), .S(CORE_ULA_REGB_Stall_bF_buf2), .Y(_92_) );
INVX1 INVX1_195 ( .A(_92_), .Y(_143__28_) );
MUX2X1 MUX2X1_776 ( .A(ULA_out_exec_pipe_29_), .B(REG_B_29_), .S(CORE_ULA_REGB_Stall_bF_buf0), .Y(_93_) );
INVX1 INVX1_196 ( .A(_93_), .Y(_143__29_) );
MUX2X1 MUX2X1_777 ( .A(ULA_out_exec_pipe_30_), .B(REG_B_30_), .S(CORE_ULA_REGB_Stall_bF_buf0), .Y(_94_) );
INVX1 INVX1_197 ( .A(_94_), .Y(_143__30_) );
OR2X2 OR2X2_911 ( .A(CORE_ULA_REGB_Stall_bF_buf1), .B(REG_B_31_), .Y(_95_) );
INVX1 INVX1_198 ( .A(CORE_ULA_REGB_Stall_bF_buf4), .Y(_96_) );
OR2X2 OR2X2_912 ( .A(ULA_out_exec_pipe_31_), .B(_96_), .Y(_97_) );
AND2X2 AND2X2_1116 ( .A(_97_), .B(_95_), .Y(_143__31_) );
OR2X2 OR2X2_913 ( .A(CORE_InstructionToULAMux_0_), .B(CORE_InstructionToULAMux_1_), .Y(_98_) );
OAI21X1 OAI21X1_50 ( .A(CORE_InstructionToULAMux_0_), .B(CORE_InstructionToULAMux_1_), .C(InstructionIN_0_), .Y(_99_) );
OAI21X1 OAI21X1_51 ( .A(_98__bF_buf3), .B(_64_), .C(_99_), .Y(ULA_B_0_) );
OAI21X1 OAI21X1_52 ( .A(CORE_InstructionToULAMux_0_), .B(CORE_InstructionToULAMux_1_), .C(InstructionIN_1_), .Y(_100_) );
OAI21X1 OAI21X1_53 ( .A(_98__bF_buf3), .B(_65_), .C(_100_), .Y(ULA_B_1_) );
OAI21X1 OAI21X1_54 ( .A(CORE_InstructionToULAMux_0_), .B(CORE_InstructionToULAMux_1_), .C(InstructionIN_2_), .Y(_101_) );
OAI21X1 OAI21X1_55 ( .A(_98__bF_buf3), .B(_66_), .C(_101_), .Y(ULA_B_2_) );
OAI21X1 OAI21X1_56 ( .A(CORE_InstructionToULAMux_0_), .B(CORE_InstructionToULAMux_1_), .C(InstructionIN_3_), .Y(_102_) );
OAI21X1 OAI21X1_57 ( .A(_98__bF_buf3), .B(_67_), .C(_102_), .Y(ULA_B_3_) );
NAND2X1 NAND2X1_747 ( .A(CORE_InstructionToULAMux_1_), .B(InstructionIN_4_), .Y(_103_) );
OAI21X1 OAI21X1_58 ( .A(_98__bF_buf3), .B(_68_), .C(_103_), .Y(ULA_B_4_) );
NAND2X1 NAND2X1_748 ( .A(CORE_InstructionToULAMux_1_), .B(InstructionIN_5_), .Y(_104_) );
OAI21X1 OAI21X1_59 ( .A(_98__bF_buf3), .B(_69_), .C(_104_), .Y(ULA_B_5_) );
NAND2X1 NAND2X1_749 ( .A(CORE_InstructionToULAMux_1_), .B(InstructionIN_6_), .Y(_105_) );
OAI21X1 OAI21X1_60 ( .A(_98__bF_buf3), .B(_70_), .C(_105_), .Y(ULA_B_6_) );
NAND2X1 NAND2X1_750 ( .A(CORE_InstructionToULAMux_1_), .B(InstructionIN_7_), .Y(_106_) );
OAI21X1 OAI21X1_61 ( .A(_98__bF_buf2), .B(_71_), .C(_106_), .Y(ULA_B_7_) );
NAND3X1 NAND3X1_61 ( .A(CORE_InstructionToULAMux_0_), .B(CORE_InstructionToULAMux_1_), .C(InstructionIN_7_), .Y(_107_) );
OAI21X1 OAI21X1_62 ( .A(_98__bF_buf0), .B(_72_), .C(_107__bF_buf1), .Y(ULA_B_8_) );
OAI21X1 OAI21X1_63 ( .A(_98__bF_buf0), .B(_73_), .C(_107__bF_buf1), .Y(ULA_B_9_) );
OAI21X1 OAI21X1_64 ( .A(_98__bF_buf2), .B(_74_), .C(_107__bF_buf3), .Y(ULA_B_10_) );
OAI21X1 OAI21X1_65 ( .A(_98__bF_buf0), .B(_75_), .C(_107__bF_buf1), .Y(ULA_B_11_) );
OAI21X1 OAI21X1_66 ( .A(_98__bF_buf4), .B(_76_), .C(_107__bF_buf0), .Y(ULA_B_12_) );
OAI21X1 OAI21X1_67 ( .A(_98__bF_buf0), .B(_77_), .C(_107__bF_buf1), .Y(ULA_B_13_) );
OAI21X1 OAI21X1_68 ( .A(_98__bF_buf0), .B(_78_), .C(_107__bF_buf1), .Y(ULA_B_14_) );
OAI21X1 OAI21X1_69 ( .A(_98__bF_buf0), .B(_79_), .C(_107__bF_buf1), .Y(ULA_B_15_) );
OAI21X1 OAI21X1_70 ( .A(_98__bF_buf2), .B(_80_), .C(_107__bF_buf3), .Y(ULA_B_16_) );
OAI21X1 OAI21X1_71 ( .A(_98__bF_buf4), .B(_81_), .C(_107__bF_buf3), .Y(ULA_B_17_) );
OAI21X1 OAI21X1_72 ( .A(_98__bF_buf2), .B(_82_), .C(_107__bF_buf3), .Y(ULA_B_18_) );
OAI21X1 OAI21X1_73 ( .A(_98__bF_buf1), .B(_83_), .C(_107__bF_buf2), .Y(ULA_B_19_) );
OAI21X1 OAI21X1_74 ( .A(_98__bF_buf2), .B(_84_), .C(_107__bF_buf3), .Y(ULA_B_20_) );
OAI21X1 OAI21X1_75 ( .A(_98__bF_buf2), .B(_85_), .C(_107__bF_buf3), .Y(ULA_B_21_) );
OAI21X1 OAI21X1_76 ( .A(_98__bF_buf1), .B(_86_), .C(_107__bF_buf2), .Y(ULA_B_22_) );
OAI21X1 OAI21X1_77 ( .A(_98__bF_buf4), .B(_87_), .C(_107__bF_buf0), .Y(ULA_B_23_) );
OAI21X1 OAI21X1_78 ( .A(_98__bF_buf1), .B(_88_), .C(_107__bF_buf2), .Y(ULA_B_24_) );
OAI21X1 OAI21X1_79 ( .A(_98__bF_buf4), .B(_89_), .C(_107__bF_buf0), .Y(ULA_B_25_) );
OAI21X1 OAI21X1_80 ( .A(_98__bF_buf1), .B(_90_), .C(_107__bF_buf2), .Y(ULA_B_26_) );
OAI21X1 OAI21X1_81 ( .A(_98__bF_buf4), .B(_91_), .C(_107__bF_buf0), .Y(ULA_B_27_) );
OAI21X1 OAI21X1_82 ( .A(_98__bF_buf1), .B(_92_), .C(_107__bF_buf2), .Y(ULA_B_28_) );
OAI21X1 OAI21X1_83 ( .A(_98__bF_buf4), .B(_93_), .C(_107__bF_buf0), .Y(ULA_B_29_) );
OAI21X1 OAI21X1_84 ( .A(_98__bF_buf1), .B(_94_), .C(_107__bF_buf2), .Y(ULA_B_30_) );
INVX1 INVX1_199 ( .A(_98__bF_buf4), .Y(_108_) );
AND2X2 AND2X2_1117 ( .A(_143__31_), .B(_108_), .Y(ULA_B_31_) );
INVX1 INVX1_200 ( .A(REG_A_0_), .Y(_109_) );
INVX2 INVX2_5 ( .A(CORE_ULA_REGA_Stall), .Y(_110_) );
MUX2X1 MUX2X1_778 ( .A(_109_), .B(_0_), .S(_110__bF_buf2), .Y(ULA_A_0_) );
INVX1 INVX1_201 ( .A(REG_A_1_), .Y(_111_) );
MUX2X1 MUX2X1_779 ( .A(_111_), .B(_2_), .S(_110__bF_buf4), .Y(ULA_A_1_) );
INVX1 INVX1_202 ( .A(REG_A_2_), .Y(_112_) );
MUX2X1 MUX2X1_780 ( .A(_112_), .B(_4_), .S(_110__bF_buf2), .Y(ULA_A_2_) );
INVX1 INVX1_203 ( .A(REG_A_3_), .Y(_113_) );
MUX2X1 MUX2X1_781 ( .A(_113_), .B(_6_), .S(_110__bF_buf0), .Y(ULA_A_3_) );
INVX1 INVX1_204 ( .A(REG_A_4_), .Y(_114_) );
MUX2X1 MUX2X1_782 ( .A(_114_), .B(_8_), .S(_110__bF_buf0), .Y(ULA_A_4_) );
INVX1 INVX1_205 ( .A(REG_A_5_), .Y(_115_) );
MUX2X1 MUX2X1_783 ( .A(_115_), .B(_10_), .S(_110__bF_buf4), .Y(ULA_A_5_) );
INVX1 INVX1_206 ( .A(REG_A_6_), .Y(_116_) );
MUX2X1 MUX2X1_784 ( .A(_116_), .B(_12_), .S(_110__bF_buf0), .Y(ULA_A_6_) );
INVX1 INVX1_207 ( .A(REG_A_7_), .Y(_117_) );
MUX2X1 MUX2X1_785 ( .A(_117_), .B(_14_), .S(_110__bF_buf0), .Y(ULA_A_7_) );
INVX1 INVX1_208 ( .A(REG_A_8_), .Y(_118_) );
MUX2X1 MUX2X1_786 ( .A(_118_), .B(_16_), .S(_110__bF_buf4), .Y(ULA_A_8_) );
INVX1 INVX1_209 ( .A(REG_A_9_), .Y(_119_) );
MUX2X1 MUX2X1_787 ( .A(_119_), .B(_18_), .S(_110__bF_buf1), .Y(ULA_A_9_) );
INVX1 INVX1_210 ( .A(REG_A_10_), .Y(_120_) );
MUX2X1 MUX2X1_788 ( .A(_120_), .B(_20_), .S(_110__bF_buf1), .Y(ULA_A_10_) );
INVX1 INVX1_211 ( .A(REG_A_11_), .Y(_121_) );
MUX2X1 MUX2X1_789 ( .A(_121_), .B(_22_), .S(_110__bF_buf4), .Y(ULA_A_11_) );
INVX1 INVX1_212 ( .A(REG_A_12_), .Y(_122_) );
MUX2X1 MUX2X1_790 ( .A(_122_), .B(_24_), .S(_110__bF_buf3), .Y(ULA_A_12_) );
INVX1 INVX1_213 ( .A(REG_A_13_), .Y(_123_) );
MUX2X1 MUX2X1_791 ( .A(_123_), .B(_26_), .S(_110__bF_buf3), .Y(ULA_A_13_) );
INVX1 INVX1_214 ( .A(REG_A_14_), .Y(_124_) );
MUX2X1 MUX2X1_792 ( .A(_124_), .B(_28_), .S(_110__bF_buf1), .Y(ULA_A_14_) );
INVX1 INVX1_215 ( .A(REG_A_15_), .Y(_125_) );
MUX2X1 MUX2X1_793 ( .A(_125_), .B(_30_), .S(_110__bF_buf1), .Y(ULA_A_15_) );
INVX1 INVX1_216 ( .A(REG_A_16_), .Y(_126_) );
MUX2X1 MUX2X1_794 ( .A(_126_), .B(_32_), .S(_110__bF_buf1), .Y(ULA_A_16_) );
INVX1 INVX1_217 ( .A(REG_A_17_), .Y(_127_) );
MUX2X1 MUX2X1_795 ( .A(_127_), .B(_34_), .S(_110__bF_buf3), .Y(ULA_A_17_) );
INVX1 INVX1_218 ( .A(REG_A_18_), .Y(_128_) );
MUX2X1 MUX2X1_796 ( .A(_128_), .B(_36_), .S(_110__bF_buf4), .Y(ULA_A_18_) );
INVX1 INVX1_219 ( .A(REG_A_19_), .Y(_129_) );
MUX2X1 MUX2X1_797 ( .A(_129_), .B(_38_), .S(_110__bF_buf2), .Y(ULA_A_19_) );
INVX1 INVX1_220 ( .A(REG_A_20_), .Y(_130_) );
MUX2X1 MUX2X1_798 ( .A(_130_), .B(_40_), .S(_110__bF_buf0), .Y(ULA_A_20_) );
INVX1 INVX1_221 ( .A(REG_A_21_), .Y(_131_) );
MUX2X1 MUX2X1_799 ( .A(_131_), .B(_42_), .S(_110__bF_buf4), .Y(ULA_A_21_) );
INVX1 INVX1_222 ( .A(REG_A_22_), .Y(_132_) );
MUX2X1 MUX2X1_800 ( .A(_132_), .B(_44_), .S(_110__bF_buf3), .Y(ULA_A_22_) );
INVX1 INVX1_223 ( .A(REG_A_23_), .Y(_133_) );
MUX2X1 MUX2X1_801 ( .A(_133_), .B(_46_), .S(_110__bF_buf1), .Y(ULA_A_23_) );
INVX1 INVX1_224 ( .A(REG_A_24_), .Y(_134_) );
MUX2X1 MUX2X1_802 ( .A(_134_), .B(_48_), .S(_110__bF_buf2), .Y(ULA_A_24_) );
INVX1 INVX1_225 ( .A(REG_A_25_), .Y(_135_) );
MUX2X1 MUX2X1_803 ( .A(_135_), .B(_50_), .S(_110__bF_buf3), .Y(ULA_A_25_) );
INVX1 INVX1_226 ( .A(REG_A_26_), .Y(_136_) );
MUX2X1 MUX2X1_804 ( .A(_136_), .B(_52_), .S(_110__bF_buf3), .Y(ULA_A_26_) );
INVX1 INVX1_227 ( .A(REG_A_27_), .Y(_137_) );
MUX2X1 MUX2X1_805 ( .A(_137_), .B(_54_), .S(_110__bF_buf0), .Y(ULA_A_27_) );
INVX1 INVX1_228 ( .A(REG_A_28_), .Y(_138_) );
MUX2X1 MUX2X1_806 ( .A(_138_), .B(_56_), .S(_110__bF_buf4), .Y(ULA_A_28_) );
INVX1 INVX1_229 ( .A(REG_A_29_), .Y(_139_) );
MUX2X1 MUX2X1_807 ( .A(_139_), .B(_58_), .S(_110__bF_buf2), .Y(ULA_A_29_) );
INVX1 INVX1_230 ( .A(REG_A_30_), .Y(_140_) );
MUX2X1 MUX2X1_808 ( .A(_140_), .B(_60_), .S(_110__bF_buf3), .Y(ULA_A_30_) );
INVX1 INVX1_231 ( .A(REG_A_31_), .Y(_141_) );
MUX2X1 MUX2X1_809 ( .A(_141_), .B(_62_), .S(_110__bF_buf2), .Y(ULA_A_31_) );
BUFX2 BUFX2_862 ( .A(_undef), .Y(DDATA_CORE_addr[0]) );
BUFX2 BUFX2_863 ( .A(_undef), .Y(DDATA_CORE_addr[1]) );
BUFX2 BUFX2_864 ( .A(_undef), .Y(DDATA_CORE_addr[2]) );
BUFX2 BUFX2_865 ( .A(_undef), .Y(DDATA_CORE_addr[3]) );
BUFX2 BUFX2_866 ( .A(_undef), .Y(DDATA_CORE_addr[4]) );
BUFX2 BUFX2_867 ( .A(_undef), .Y(DDATA_CORE_addr[5]) );
BUFX2 BUFX2_868 ( .A(_undef), .Y(DDATA_CORE_addr[6]) );
BUFX2 BUFX2_869 ( .A(_undef), .Y(DDATA_CORE_addr[7]) );
BUFX2 BUFX2_870 ( .A(_142__0_), .Y(DDATA_CORE_ctrl[0]) );
BUFX2 BUFX2_871 ( .A(_142__1_), .Y(DDATA_CORE_ctrl[1]) );
BUFX2 BUFX2_872 ( .A(_142__2_), .Y(DDATA_CORE_ctrl[2]) );
BUFX2 BUFX2_873 ( .A(_143__0_), .Y(DDATA_CORE_in[0]) );
BUFX2 BUFX2_874 ( .A(_143__1_), .Y(DDATA_CORE_in[1]) );
BUFX2 BUFX2_875 ( .A(_143__2_), .Y(DDATA_CORE_in[2]) );
BUFX2 BUFX2_876 ( .A(_143__3_), .Y(DDATA_CORE_in[3]) );
BUFX2 BUFX2_877 ( .A(_143__4_), .Y(DDATA_CORE_in[4]) );
BUFX2 BUFX2_878 ( .A(_143__5_), .Y(DDATA_CORE_in[5]) );
BUFX2 BUFX2_879 ( .A(_143__6_), .Y(DDATA_CORE_in[6]) );
BUFX2 BUFX2_880 ( .A(_143__7_), .Y(DDATA_CORE_in[7]) );
BUFX2 BUFX2_881 ( .A(_143__8_), .Y(DDATA_CORE_in[8]) );
BUFX2 BUFX2_882 ( .A(_143__9_), .Y(DDATA_CORE_in[9]) );
BUFX2 BUFX2_883 ( .A(_143__10_), .Y(DDATA_CORE_in[10]) );
BUFX2 BUFX2_884 ( .A(_143__11_), .Y(DDATA_CORE_in[11]) );
BUFX2 BUFX2_885 ( .A(_143__12_), .Y(DDATA_CORE_in[12]) );
BUFX2 BUFX2_886 ( .A(_143__13_), .Y(DDATA_CORE_in[13]) );
BUFX2 BUFX2_887 ( .A(_143__14_), .Y(DDATA_CORE_in[14]) );
BUFX2 BUFX2_888 ( .A(_143__15_), .Y(DDATA_CORE_in[15]) );
BUFX2 BUFX2_889 ( .A(_143__16_), .Y(DDATA_CORE_in[16]) );
BUFX2 BUFX2_890 ( .A(_143__17_), .Y(DDATA_CORE_in[17]) );
BUFX2 BUFX2_891 ( .A(_143__18_), .Y(DDATA_CORE_in[18]) );
BUFX2 BUFX2_892 ( .A(_143__19_), .Y(DDATA_CORE_in[19]) );
BUFX2 BUFX2_893 ( .A(_143__20_), .Y(DDATA_CORE_in[20]) );
BUFX2 BUFX2_894 ( .A(_143__21_), .Y(DDATA_CORE_in[21]) );
BUFX2 BUFX2_895 ( .A(_143__22_), .Y(DDATA_CORE_in[22]) );
BUFX2 BUFX2_896 ( .A(_143__23_), .Y(DDATA_CORE_in[23]) );
BUFX2 BUFX2_897 ( .A(_143__24_), .Y(DDATA_CORE_in[24]) );
BUFX2 BUFX2_898 ( .A(_143__25_), .Y(DDATA_CORE_in[25]) );
BUFX2 BUFX2_899 ( .A(_143__26_), .Y(DDATA_CORE_in[26]) );
BUFX2 BUFX2_900 ( .A(_143__27_), .Y(DDATA_CORE_in[27]) );
BUFX2 BUFX2_901 ( .A(_143__28_), .Y(DDATA_CORE_in[28]) );
BUFX2 BUFX2_902 ( .A(_143__29_), .Y(DDATA_CORE_in[29]) );
BUFX2 BUFX2_903 ( .A(_143__30_), .Y(DDATA_CORE_in[30]) );
BUFX2 BUFX2_904 ( .A(_143__31_), .Y(DDATA_CORE_in[31]) );
BUFX2 BUFX2_905 ( .A(_144_), .Y(DDATA_CORE_load) );
BUFX2 BUFX2_906 ( .A(_145_), .Y(DDATA_CORE_write) );
BUFX2 BUFX2_907 ( .A(_146__0_), .Y(IDATA_CORE_addr[0]) );
BUFX2 BUFX2_908 ( .A(_146__1_), .Y(IDATA_CORE_addr[1]) );
BUFX2 BUFX2_909 ( .A(_146__2_), .Y(IDATA_CORE_addr[2]) );
BUFX2 BUFX2_910 ( .A(_146__3_), .Y(IDATA_CORE_addr[3]) );
BUFX2 BUFX2_911 ( .A(_146__4_), .Y(IDATA_CORE_addr[4]) );
BUFX2 BUFX2_912 ( .A(_146__5_), .Y(IDATA_CORE_addr[5]) );
BUFX2 BUFX2_913 ( .A(_146__6_), .Y(IDATA_CORE_addr[6]) );
BUFX2 BUFX2_914 ( .A(_146__7_), .Y(IDATA_CORE_addr[7]) );
BUFX2 BUFX2_915 ( .A(_147_), .Y(IDATA_CORE_clk) );
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf87), .D(CORE_InstructionIN_0_), .Q(InstructionIN_0_) );
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf53), .D(CORE_InstructionIN_1_), .Q(InstructionIN_1_) );
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf81), .D(CORE_InstructionIN_2_), .Q(InstructionIN_2_) );
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf69), .D(CORE_InstructionIN_3_), .Q(InstructionIN_3_) );
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf65), .D(CORE_InstructionIN_4_), .Q(InstructionIN_4_) );
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf65), .D(CORE_InstructionIN_5_), .Q(InstructionIN_5_) );
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf87), .D(CORE_InstructionIN_6_), .Q(InstructionIN_6_) );
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf27), .D(CORE_InstructionIN_7_), .Q(InstructionIN_7_) );
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf19), .D(CORE_REG_RFD_0_), .Q(REG_RFD_exec_pipe_0_) );
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf53), .D(CORE_REG_RFD_1_), .Q(REG_RFD_exec_pipe_1_) );
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf6), .D(CORE_REG_RFD_2_), .Q(REG_RFD_exec_pipe_2_) );
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf6), .D(CORE_REG_RFD_3_), .Q(REG_RFD_exec_pipe_3_) );
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf77), .D(CORE_REG_write), .Q(REG_Write_exec_pipe) );
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf19), .D(CORE_DATA_REGMux), .Q(CORE_DATA_REGMux_exec_pipe) );
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf5), .D(ULA_ULA_OUT_0_), .Q(PC_ULA_OUT_0_) );
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_1_), .Q(PC_ULA_OUT_1_) );
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf7), .D(ULA_ULA_OUT_2_), .Q(PC_ULA_OUT_2_) );
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf5), .D(ULA_ULA_OUT_3_), .Q(PC_ULA_OUT_3_) );
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf56), .D(ULA_ULA_OUT_4_), .Q(PC_ULA_OUT_4_) );
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf5), .D(ULA_ULA_OUT_5_), .Q(PC_ULA_OUT_5_) );
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf13), .D(ULA_ULA_OUT_6_), .Q(PC_ULA_OUT_6_) );
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_7_), .Q(PC_ULA_OUT_7_) );
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_8_), .Q(ULA_out_exec_pipe_8_) );
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_9_), .Q(ULA_out_exec_pipe_9_) );
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_10_), .Q(ULA_out_exec_pipe_10_) );
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_11_), .Q(ULA_out_exec_pipe_11_) );
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_12_), .Q(ULA_out_exec_pipe_12_) );
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf31), .D(ULA_ULA_OUT_13_), .Q(ULA_out_exec_pipe_13_) );
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_14_), .Q(ULA_out_exec_pipe_14_) );
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_15_), .Q(ULA_out_exec_pipe_15_) );
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_16_), .Q(ULA_out_exec_pipe_16_) );
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_17_), .Q(ULA_out_exec_pipe_17_) );
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf31), .D(ULA_ULA_OUT_18_), .Q(ULA_out_exec_pipe_18_) );
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf5), .D(ULA_ULA_OUT_19_), .Q(ULA_out_exec_pipe_19_) );
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_20_), .Q(ULA_out_exec_pipe_20_) );
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_21_), .Q(ULA_out_exec_pipe_21_) );
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_22_), .Q(ULA_out_exec_pipe_22_) );
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf5), .D(ULA_ULA_OUT_23_), .Q(ULA_out_exec_pipe_23_) );
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf31), .D(ULA_ULA_OUT_24_), .Q(ULA_out_exec_pipe_24_) );
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_25_), .Q(ULA_out_exec_pipe_25_) );
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_26_), .Q(ULA_out_exec_pipe_26_) );
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_27_), .Q(ULA_out_exec_pipe_27_) );
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf40), .D(ULA_ULA_OUT_28_), .Q(ULA_out_exec_pipe_28_) );
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf31), .D(ULA_ULA_OUT_29_), .Q(ULA_out_exec_pipe_29_) );
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf72), .D(ULA_ULA_OUT_30_), .Q(ULA_out_exec_pipe_30_) );
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf31), .D(ULA_ULA_OUT_31_), .Q(ULA_out_exec_pipe_31_) );
DFFNEGX1 DFFNEGX1_1 ( .CLK(clk_bF_buf19), .D(REG_Write_exec_pipe), .Q(REG_Write_wb_pipe) );
INVX1 INVX1_232 ( .A(rst_bF_buf4), .Y(_164_) );
AND2X2 AND2X2_1118 ( .A(_164_), .B(ID_old_rd1_0_), .Y(_163__0_) );
AND2X2 AND2X2_1119 ( .A(_164_), .B(ID_old_rd1_1_), .Y(_163__1_) );
AND2X2 AND2X2_1120 ( .A(_164_), .B(ID_old_rd1_2_), .Y(_163__2_) );
AND2X2 AND2X2_1121 ( .A(_164_), .B(ID_old_rd1_3_), .Y(_163__3_) );
INVX1 INVX1_233 ( .A(CORE_InstructionIN_5_), .Y(_165_) );
INVX1 INVX1_234 ( .A(CORE_InstructionIN_4_), .Y(_166_) );
AOI21X1 AOI21X1_28 ( .A(CORE_InstructionIN_8_), .B(CORE_InstructionIN_9_), .C(CORE_InstructionIN_10_), .Y(_167_) );
INVX1 INVX1_235 ( .A(CORE_InstructionIN_1_), .Y(_168_) );
NOR2X1 NOR2X1_106 ( .A(CORE_InstructionIN_2_), .B(CORE_InstructionIN_3_), .Y(_169_) );
NAND3X1 NAND3X1_62 ( .A(_169_), .B(_168_), .C(CORE_InstructionIN_0_), .Y(_170_) );
OR2X2 OR2X2_914 ( .A(CORE_InstructionIN_13_), .B(CORE_InstructionIN_12_), .Y(_171_) );
OR2X2 OR2X2_915 ( .A(CORE_InstructionIN_14_), .B(_171_), .Y(_172_) );
INVX1 INVX1_236 ( .A(CORE_InstructionIN_0_), .Y(_173_) );
NAND3X1 NAND3X1_63 ( .A(_169_), .B(_168_), .C(_173_), .Y(_174_) );
INVX1 INVX1_237 ( .A(_174_), .Y(_175_) );
INVX1 INVX1_238 ( .A(CORE_InstructionIN_8_), .Y(_176_) );
INVX1 INVX1_239 ( .A(CORE_InstructionIN_9_), .Y(_177_) );
INVX1 INVX1_240 ( .A(CORE_InstructionIN_10_), .Y(_178_) );
NAND2X1 NAND2X1_751 ( .A(CORE_InstructionIN_0_), .B(_169_), .Y(_179_) );
NOR3X1 NOR3X1_11 ( .A(CORE_InstructionIN_14_), .B(CORE_InstructionIN_13_), .C(CORE_InstructionIN_12_), .Y(_180_) );
NAND2X1 NAND2X1_752 ( .A(CORE_InstructionIN_11_), .B(_180_), .Y(_181_) );
INVX1 INVX1_241 ( .A(CORE_InstructionIN_15_), .Y(_182_) );
AND2X2 AND2X2_1122 ( .A(CORE_InstructionIN_8_), .B(CORE_InstructionIN_9_), .Y(_183_) );
AND2X2 AND2X2_1123 ( .A(_171_), .B(CORE_InstructionIN_14_), .Y(_184_) );
INVX1 INVX1_242 ( .A(_184_), .Y(_185_) );
OAI21X1 OAI21X1_85 ( .A(CORE_InstructionIN_14_), .B(CORE_InstructionIN_13_), .C(_185_), .Y(_186_) );
NAND2X1 NAND2X1_753 ( .A(_182_), .B(_186_), .Y(_187_) );
MUX2X1 MUX2X1_810 ( .A(CORE_InstructionIN_8_), .B(CORE_REG_RFD_0_), .S(_187_), .Y(_188_) );
INVX1 INVX1_243 ( .A(CORE_InstructionIN_14_), .Y(_189_) );
INVX1 INVX1_244 ( .A(CORE_InstructionIN_12_), .Y(_190_) );
NAND3X1 NAND3X1_64 ( .A(_189_), .B(CORE_InstructionIN_13_), .C(_190_), .Y(_191_) );
OAI21X1 OAI21X1_86 ( .A(_191_), .B(_174_), .C(_182_), .Y(_192_) );
NAND2X1 NAND2X1_754 ( .A(_164_), .B(_192_), .Y(_193_) );
NOR2X1 NOR2X1_107 ( .A(_188_), .B(_193_), .Y(_162__0_) );
MUX2X1 MUX2X1_811 ( .A(CORE_InstructionIN_9_), .B(CORE_REG_RFD_1_), .S(_187_), .Y(_194_) );
NOR2X1 NOR2X1_108 ( .A(_194_), .B(_193_), .Y(_162__1_) );
MUX2X1 MUX2X1_812 ( .A(CORE_InstructionIN_10_), .B(CORE_REG_RFD_2_), .S(_187_), .Y(_195_) );
NOR2X1 NOR2X1_109 ( .A(_195_), .B(_193_), .Y(_162__2_) );
MUX2X1 MUX2X1_813 ( .A(CORE_REG_RFD_3_), .B(CORE_InstructionIN_11_), .S(_186_), .Y(_196_) );
AOI21X1 AOI21X1_29 ( .A(_182_), .B(_196_), .C(rst_bF_buf3), .Y(_154__3_) );
AND2X2 AND2X2_1124 ( .A(_154__3_), .B(_192_), .Y(_162__3_) );
NOR2X1 NOR2X1_110 ( .A(rst_bF_buf2), .B(CORE_InstructionIN_15_), .Y(_197_) );
NOR2X1 NOR2X1_111 ( .A(_177_), .B(CORE_InstructionIN_10_), .Y(_198_) );
OR2X2 OR2X2_916 ( .A(CORE_InstructionIN_10_), .B(_183_), .Y(_199_) );
INVX1 INVX1_245 ( .A(_197_), .Y(_200_) );
INVX1 INVX1_246 ( .A(CORE_InstructionIN_11_), .Y(_201_) );
NAND3X1 NAND3X1_65 ( .A(_177_), .B(CORE_InstructionIN_8_), .C(ULA_zero), .Y(_202_) );
NAND2X1 NAND2X1_755 ( .A(gnd), .B(_183_), .Y(_203_) );
OAI21X1 OAI21X1_87 ( .A(gnd), .B(_177_), .C(_176_), .Y(_204_) );
NAND3X1 NAND3X1_66 ( .A(_204_), .B(_203_), .C(_202_), .Y(_205_) );
INVX1 INVX1_247 ( .A(CORE_InstructionIN_13_), .Y(_206_) );
AND2X2 AND2X2_1125 ( .A(_189_), .B(CORE_InstructionIN_12_), .Y(_207_) );
AND2X2 AND2X2_1126 ( .A(_207_), .B(_206_), .Y(_208_) );
NAND3X1 NAND3X1_67 ( .A(_205_), .B(_201_), .C(_208_), .Y(_209_) );
NOR2X1 NOR2X1_112 ( .A(_177_), .B(_178_), .Y(_210_) );
NOR2X1 NOR2X1_113 ( .A(_167_), .B(CORE_PC_ctrl_0_), .Y(_211_) );
NOR3X1 NOR3X1_12 ( .A(_181_), .B(_210_), .C(_211_), .Y(_212_) );
NAND2X1 NAND2X1_756 ( .A(CORE_InstructionIN_11_), .B(_208_), .Y(_213_) );
NAND2X1 NAND2X1_757 ( .A(_185_), .B(_213_), .Y(_214_) );
AOI21X1 AOI21X1_30 ( .A(CORE_PC_ctrl_0_), .B(_214_), .C(_212_), .Y(_215_) );
AOI21X1 AOI21X1_31 ( .A(_209_), .B(_215_), .C(_200_), .Y(_153__0_) );
NOR2X1 NOR2X1_114 ( .A(_181_), .B(_167_), .Y(_216_) );
AOI21X1 AOI21X1_32 ( .A(CORE_PC_ctrl_1_), .B(_214_), .C(_216_), .Y(_217_) );
OAI21X1 OAI21X1_88 ( .A(CORE_PC_ctrl_1_), .B(_210_), .C(_197_), .Y(_218_) );
NOR2X1 NOR2X1_115 ( .A(_217_), .B(_218_), .Y(_153__1_) );
NOR2X1 NOR2X1_116 ( .A(_172_), .B(_201_), .Y(_219_) );
INVX1 INVX1_248 ( .A(CORE_STACK_ctrl_0_), .Y(_220_) );
OAI21X1 OAI21X1_89 ( .A(_220_), .B(_210_), .C(_199_), .Y(_221_) );
AOI22X1 AOI22X1_2 ( .A(CORE_STACK_ctrl_0_), .B(_184_), .C(_221_), .D(_219_), .Y(_222_) );
NOR2X1 NOR2X1_117 ( .A(_222_), .B(_200_), .Y(_158__0_) );
AOI21X1 AOI21X1_33 ( .A(_210_), .B(_219_), .C(CORE_STACK_ctrl_1_), .Y(_223_) );
OAI21X1 OAI21X1_90 ( .A(_184_), .B(_216_), .C(_197_), .Y(_224_) );
NOR2X1 NOR2X1_118 ( .A(_224_), .B(_223_), .Y(_158__1_) );
OAI21X1 OAI21X1_91 ( .A(_191_), .B(_175_), .C(_185_), .Y(_225_) );
AND2X2 AND2X2_1127 ( .A(_225_), .B(CORE_DATA_REGMux), .Y(_226_) );
NAND2X1 NAND2X1_758 ( .A(_168_), .B(_173_), .Y(_227_) );
AND2X2 AND2X2_1128 ( .A(_227_), .B(_169_), .Y(_228_) );
INVX1 INVX1_249 ( .A(_228_), .Y(_229_) );
INVX1 INVX1_250 ( .A(CORE_InstructionIN_3_), .Y(_230_) );
NAND3X1 NAND3X1_68 ( .A(_168_), .B(CORE_InstructionIN_2_), .C(_230_), .Y(_231_) );
AOI21X1 AOI21X1_34 ( .A(_231_), .B(_229_), .C(_191_), .Y(_232_) );
OR2X2 OR2X2_917 ( .A(_232_), .B(_226_), .Y(_233_) );
AND2X2 AND2X2_1129 ( .A(_233_), .B(_197_), .Y(_148_) );
INVX1 INVX1_251 ( .A(_142__0_), .Y(_234_) );
NOR3X1 NOR3X1_13 ( .A(_206_), .B(CORE_InstructionIN_14_), .C(CORE_InstructionIN_12_), .Y(_235_) );
NAND3X1 NAND3X1_69 ( .A(_170_), .B(_231_), .C(_235_), .Y(_236_) );
AOI21X1 AOI21X1_35 ( .A(_234_), .B(_229_), .C(_236_), .Y(_237_) );
NAND2X1 NAND2X1_759 ( .A(CORE_InstructionIN_13_), .B(_207_), .Y(_238_) );
NOR3X1 NOR3X1_14 ( .A(_178_), .B(_142__0_), .C(_201_), .Y(_239_) );
NOR2X1 NOR2X1_119 ( .A(CORE_InstructionIN_8_), .B(CORE_InstructionIN_11_), .Y(_240_) );
NOR3X1 NOR3X1_15 ( .A(_238_), .B(_239_), .C(_240_), .Y(_241_) );
OR2X2 OR2X2_918 ( .A(_241_), .B(_237_), .Y(_242_) );
AND2X2 AND2X2_1130 ( .A(_242_), .B(_197_), .Y(_243_) );
NOR2X1 NOR2X1_120 ( .A(_186_), .B(CORE_InstructionIN_15_), .Y(_244_) );
NOR3X1 NOR3X1_16 ( .A(_244_), .B(rst_bF_buf2), .C(_234_), .Y(_245_) );
OR2X2 OR2X2_919 ( .A(_245_), .B(_243_), .Y(_149__0_) );
INVX1 INVX1_252 ( .A(_238_), .Y(_246_) );
OAI21X1 OAI21X1_92 ( .A(CORE_InstructionIN_10_), .B(_177_), .C(_201_), .Y(_247_) );
INVX1 INVX1_253 ( .A(_142__1_), .Y(_248_) );
NAND3X1 NAND3X1_70 ( .A(_248_), .B(CORE_InstructionIN_10_), .C(CORE_InstructionIN_11_), .Y(_249_) );
NAND3X1 NAND3X1_71 ( .A(_246_), .B(_249_), .C(_247_), .Y(_250_) );
NAND2X1 NAND2X1_760 ( .A(_248_), .B(_231_), .Y(_251_) );
NAND3X1 NAND3X1_72 ( .A(_229_), .B(_235_), .C(_251_), .Y(_252_) );
AOI21X1 AOI21X1_36 ( .A(_250_), .B(_252_), .C(_200_), .Y(_253_) );
NOR3X1 NOR3X1_17 ( .A(_244_), .B(rst_bF_buf2), .C(_248_), .Y(_254_) );
OR2X2 OR2X2_920 ( .A(_254_), .B(_253_), .Y(_149__1_) );
NOR3X1 NOR3X1_18 ( .A(_178_), .B(_142__2_), .C(_201_), .Y(_255_) );
OR2X2 OR2X2_921 ( .A(CORE_InstructionIN_10_), .B(CORE_InstructionIN_11_), .Y(_256_) );
INVX1 INVX1_254 ( .A(_256_), .Y(_257_) );
NOR3X1 NOR3X1_19 ( .A(_238_), .B(_255_), .C(_257_), .Y(_258_) );
NOR2X1 NOR2X1_121 ( .A(_231_), .B(_173_), .Y(_259_) );
INVX1 INVX1_255 ( .A(CORE_InstructionIN_2_), .Y(_260_) );
NOR3X1 NOR3X1_20 ( .A(_260_), .B(CORE_InstructionIN_1_), .C(CORE_InstructionIN_3_), .Y(_261_) );
NOR3X1 NOR3X1_21 ( .A(_228_), .B(_142__2_), .C(_261_), .Y(_262_) );
NAND2X1 NAND2X1_761 ( .A(_235_), .B(_179_), .Y(_263_) );
NOR3X1 NOR3X1_22 ( .A(_262_), .B(_259_), .C(_263_), .Y(_264_) );
OR2X2 OR2X2_922 ( .A(_258_), .B(_264_), .Y(_265_) );
AND2X2 AND2X2_1131 ( .A(_265_), .B(_197_), .Y(_266_) );
INVX1 INVX1_256 ( .A(_142__2_), .Y(_267_) );
NOR3X1 NOR3X1_23 ( .A(_244_), .B(rst_bF_buf2), .C(_267_), .Y(_268_) );
OR2X2 OR2X2_923 ( .A(_268_), .B(_266_), .Y(_149__2_) );
AND2X2 AND2X2_1132 ( .A(_225_), .B(_144_), .Y(_269_) );
OR2X2 OR2X2_924 ( .A(_232_), .B(_269_), .Y(_270_) );
AND2X2 AND2X2_1133 ( .A(_270_), .B(_197_), .Y(_150_) );
NAND2X1 NAND2X1_762 ( .A(_145_), .B(_184_), .Y(_271_) );
AOI21X1 AOI21X1_37 ( .A(_271_), .B(_238_), .C(_200_), .Y(_151_) );
OAI21X1 OAI21X1_93 ( .A(_184_), .B(_216_), .C(CORE_REG_write), .Y(_272_) );
NOR2X1 NOR2X1_122 ( .A(_189_), .B(_171_), .Y(_273_) );
NOR3X1 NOR3X1_24 ( .A(_235_), .B(CORE_InstructionIN_15_), .C(_273_), .Y(_274_) );
AOI21X1 AOI21X1_38 ( .A(_274_), .B(_272_), .C(rst_bF_buf2), .Y(_157_) );
NOR3X1 NOR3X1_25 ( .A(_199_), .B(_201_), .C(_172_), .Y(_275_) );
OR2X2 OR2X2_925 ( .A(CORE_InstructionIN_15_), .B(_207_), .Y(_276_) );
OR2X2 OR2X2_926 ( .A(_276_), .B(_275_), .Y(_277_) );
OR2X2 OR2X2_927 ( .A(_201_), .B(_199_), .Y(_278_) );
AND2X2 AND2X2_1134 ( .A(_278_), .B(_180_), .Y(_279_) );
OR2X2 OR2X2_928 ( .A(CORE_InstructionIN_14_), .B(_279_), .Y(_280_) );
AND2X2 AND2X2_1135 ( .A(_182_), .B(CORE_REG_RF2_0_), .Y(_281_) );
AOI22X1 AOI22X1_3 ( .A(_280_), .B(_281_), .C(_277_), .D(CORE_InstructionIN_0_), .Y(_282_) );
NOR2X1 NOR2X1_123 ( .A(_282_), .B(rst_bF_buf4), .Y(_156__0_) );
AND2X2 AND2X2_1136 ( .A(_277_), .B(CORE_InstructionIN_1_), .Y(_283_) );
AND2X2 AND2X2_1137 ( .A(_182_), .B(CORE_REG_RF2_1_), .Y(_284_) );
AND2X2 AND2X2_1138 ( .A(_280_), .B(_284_), .Y(_285_) );
OR2X2 OR2X2_929 ( .A(_285_), .B(_283_), .Y(_286_) );
AND2X2 AND2X2_1139 ( .A(_286_), .B(_164_), .Y(_156__1_) );
AND2X2 AND2X2_1140 ( .A(_182_), .B(CORE_REG_RF2_2_), .Y(_287_) );
AOI22X1 AOI22X1_4 ( .A(_280_), .B(_287_), .C(_277_), .D(CORE_InstructionIN_2_), .Y(_288_) );
NOR2X1 NOR2X1_124 ( .A(_288_), .B(rst_bF_buf3), .Y(_156__2_) );
AND2X2 AND2X2_1141 ( .A(_277_), .B(CORE_InstructionIN_3_), .Y(_289_) );
AND2X2 AND2X2_1142 ( .A(_182_), .B(CORE_REG_RF2_3_), .Y(_290_) );
AND2X2 AND2X2_1143 ( .A(_280_), .B(_290_), .Y(_291_) );
OR2X2 OR2X2_930 ( .A(_291_), .B(_289_), .Y(_292_) );
AND2X2 AND2X2_1144 ( .A(_292_), .B(_164_), .Y(_156__3_) );
NAND2X1 NAND2X1_763 ( .A(CORE_InstructionIN_15_), .B(_166_), .Y(_293_) );
NOR3X1 NOR3X1_26 ( .A(_166_), .B(CORE_InstructionIN_14_), .C(_206_), .Y(_294_) );
OR2X2 OR2X2_931 ( .A(CORE_InstructionIN_4_), .B(_256_), .Y(_295_) );
OR2X2 OR2X2_932 ( .A(CORE_REG_RF1_0_), .B(_201_), .Y(_296_) );
AND2X2 AND2X2_1145 ( .A(_208_), .B(_296_), .Y(_297_) );
AND2X2 AND2X2_1146 ( .A(_297_), .B(_295_), .Y(_298_) );
OR2X2 OR2X2_933 ( .A(_294_), .B(_298_), .Y(_299_) );
NAND2X1 NAND2X1_764 ( .A(CORE_InstructionIN_8_), .B(_166_), .Y(_300_) );
AND2X2 AND2X2_1147 ( .A(_275_), .B(_300_), .Y(_301_) );
OR2X2 OR2X2_934 ( .A(_301_), .B(_299_), .Y(_302_) );
OR2X2 OR2X2_935 ( .A(_184_), .B(_279_), .Y(_303_) );
AND2X2 AND2X2_1148 ( .A(_303_), .B(CORE_REG_RF1_0_), .Y(_304_) );
OR2X2 OR2X2_936 ( .A(CORE_InstructionIN_15_), .B(_304_), .Y(_305_) );
OR2X2 OR2X2_937 ( .A(_305_), .B(_302_), .Y(_306_) );
AND2X2 AND2X2_1149 ( .A(_306_), .B(_293_), .Y(_307_) );
AND2X2 AND2X2_1150 ( .A(_307_), .B(_164_), .Y(_155__0_) );
AND2X2 AND2X2_1151 ( .A(_257_), .B(CORE_InstructionIN_5_), .Y(_308_) );
AND2X2 AND2X2_1152 ( .A(CORE_InstructionIN_11_), .B(CORE_REG_RF1_1_), .Y(_309_) );
OR2X2 OR2X2_938 ( .A(_309_), .B(_308_), .Y(_310_) );
AND2X2 AND2X2_1153 ( .A(_310_), .B(_208_), .Y(_311_) );
NOR3X1 NOR3X1_27 ( .A(_165_), .B(CORE_InstructionIN_14_), .C(_206_), .Y(_312_) );
OR2X2 OR2X2_939 ( .A(_312_), .B(_311_), .Y(_313_) );
AND2X2 AND2X2_1154 ( .A(_167_), .B(CORE_InstructionIN_8_), .Y(_314_) );
AND2X2 AND2X2_1155 ( .A(_219_), .B(_314_), .Y(_315_) );
AND2X2 AND2X2_1156 ( .A(_315_), .B(CORE_InstructionIN_5_), .Y(_316_) );
OR2X2 OR2X2_940 ( .A(_316_), .B(_313_), .Y(_317_) );
AND2X2 AND2X2_1157 ( .A(_303_), .B(CORE_REG_RF1_1_), .Y(_318_) );
OR2X2 OR2X2_941 ( .A(CORE_InstructionIN_15_), .B(_318_), .Y(_319_) );
OR2X2 OR2X2_942 ( .A(_319_), .B(_317_), .Y(_320_) );
NAND2X1 NAND2X1_765 ( .A(CORE_InstructionIN_15_), .B(_165_), .Y(_321_) );
AND2X2 AND2X2_1158 ( .A(_320_), .B(_321_), .Y(_322_) );
AND2X2 AND2X2_1159 ( .A(_322_), .B(_164_), .Y(_155__1_) );
AND2X2 AND2X2_1160 ( .A(_208_), .B(CORE_InstructionIN_11_), .Y(_323_) );
AND2X2 AND2X2_1161 ( .A(_182_), .B(CORE_REG_RF1_2_), .Y(_324_) );
OAI21X1 OAI21X1_94 ( .A(_323_), .B(_303_), .C(_324_), .Y(_325_) );
INVX1 INVX1_257 ( .A(CORE_InstructionIN_6_), .Y(_326_) );
NAND2X1 NAND2X1_766 ( .A(CORE_InstructionIN_13_), .B(_189_), .Y(_327_) );
NAND3X1 NAND3X1_73 ( .A(_314_), .B(CORE_InstructionIN_11_), .C(_180_), .Y(_328_) );
AND2X2 AND2X2_1162 ( .A(_328_), .B(_327_), .Y(_329_) );
AOI21X1 AOI21X1_39 ( .A(_257_), .B(_208_), .C(CORE_InstructionIN_15_), .Y(_330_) );
AND2X2 AND2X2_1163 ( .A(_329_), .B(_330_), .Y(_331_) );
OR2X2 OR2X2_943 ( .A(_326_), .B(_331_), .Y(_332_) );
AND2X2 AND2X2_1164 ( .A(_332_), .B(_325_), .Y(_333_) );
NOR2X1 NOR2X1_125 ( .A(_333_), .B(rst_bF_buf3), .Y(_155__2_) );
OR2X2 OR2X2_944 ( .A(_323_), .B(_303_), .Y(_334_) );
AND2X2 AND2X2_1165 ( .A(_182_), .B(CORE_REG_RF1_3_), .Y(_335_) );
AND2X2 AND2X2_1166 ( .A(_334_), .B(_335_), .Y(_336_) );
NOR2X1 NOR2X1_126 ( .A(_206_), .B(CORE_InstructionIN_14_), .Y(_337_) );
OR2X2 OR2X2_945 ( .A(_337_), .B(_315_), .Y(_338_) );
AND2X2 AND2X2_1167 ( .A(_208_), .B(_257_), .Y(_339_) );
OR2X2 OR2X2_946 ( .A(CORE_InstructionIN_15_), .B(_339_), .Y(_340_) );
OR2X2 OR2X2_947 ( .A(_340_), .B(_338_), .Y(_341_) );
AND2X2 AND2X2_1168 ( .A(_341_), .B(CORE_InstructionIN_7_), .Y(_342_) );
OR2X2 OR2X2_948 ( .A(_336_), .B(_342_), .Y(_343_) );
AND2X2 AND2X2_1169 ( .A(_343_), .B(_164_), .Y(_155__3_) );
NOR2X1 NOR2X1_127 ( .A(_188_), .B(rst_bF_buf4), .Y(_154__0_) );
NOR2X1 NOR2X1_128 ( .A(_194_), .B(rst_bF_buf3), .Y(_154__1_) );
NOR2X1 NOR2X1_129 ( .A(_195_), .B(rst_bF_buf4), .Y(_154__2_) );
XOR2X1 XOR2X1_63 ( .A(ID_old_rd_0_), .B(_282_), .Y(_344_) );
INVX1 INVX1_258 ( .A(ID_old_rd_0_), .Y(_345_) );
NOR3X1 NOR3X1_28 ( .A(ID_old_rd_3_), .B(ID_old_rd_2_), .C(ID_old_rd_1_), .Y(_346_) );
AOI21X1 AOI21X1_40 ( .A(_345_), .B(_346_), .C(rst_bF_buf4), .Y(_347_) );
INVX1 INVX1_259 ( .A(ID_old_rd_1_), .Y(_348_) );
XOR2X1 XOR2X1_64 ( .A(_348_), .B(_286_), .Y(_349_) );
AND2X2 AND2X2_1170 ( .A(_349_), .B(_347_), .Y(_350_) );
INVX1 INVX1_260 ( .A(ID_old_rd_3_), .Y(_351_) );
XOR2X1 XOR2X1_65 ( .A(_351_), .B(_292_), .Y(_352_) );
AND2X2 AND2X2_1171 ( .A(_350_), .B(_352_), .Y(_353_) );
XOR2X1 XOR2X1_66 ( .A(ID_old_rd_2_), .B(_288_), .Y(_354_) );
AND2X2 AND2X2_1172 ( .A(_353_), .B(_354_), .Y(_355_) );
AND2X2 AND2X2_1173 ( .A(_355_), .B(_344_), .Y(_160_) );
OR2X2 OR2X2_949 ( .A(ID_old_rd_2_), .B(_333_), .Y(_356_) );
AND2X2 AND2X2_1174 ( .A(_356_), .B(_347_), .Y(_357_) );
INVX1 INVX1_261 ( .A(ID_old_rd_2_), .Y(_358_) );
AND2X2 AND2X2_1175 ( .A(_334_), .B(_324_), .Y(_359_) );
AND2X2 AND2X2_1176 ( .A(_341_), .B(CORE_InstructionIN_6_), .Y(_360_) );
OR2X2 OR2X2_950 ( .A(_359_), .B(_360_), .Y(_361_) );
OR2X2 OR2X2_951 ( .A(_358_), .B(_361_), .Y(_362_) );
XOR2X1 XOR2X1_67 ( .A(_351_), .B(_343_), .Y(_363_) );
AND2X2 AND2X2_1177 ( .A(_363_), .B(_362_), .Y(_364_) );
AND2X2 AND2X2_1178 ( .A(_364_), .B(_357_), .Y(_365_) );
XOR2X1 XOR2X1_68 ( .A(_345_), .B(_307_), .Y(_366_) );
XOR2X1 XOR2X1_69 ( .A(_348_), .B(_322_), .Y(_367_) );
AND2X2 AND2X2_1179 ( .A(_367_), .B(_366_), .Y(_368_) );
AND2X2 AND2X2_1180 ( .A(_365_), .B(_368_), .Y(_159_) );
NAND2X1 NAND2X1_767 ( .A(CORE_InstructionIN_13_), .B(CORE_InstructionIN_12_), .Y(_369_) );
INVX1 INVX1_262 ( .A(_279_), .Y(_370_) );
NAND3X1 NAND3X1_74 ( .A(_370_), .B(_185_), .C(_369_), .Y(_371_) );
NAND3X1 NAND3X1_75 ( .A(_371_), .B(_182_), .C(ULA_cin_bF_buf2), .Y(_372_) );
NOR2X1 NOR2X1_130 ( .A(_191_), .B(_201_), .Y(_373_) );
OAI21X1 OAI21X1_95 ( .A(_208_), .B(_373_), .C(CORE_InstructionIN_15_), .Y(_374_) );
AOI21X1 AOI21X1_41 ( .A(_374_), .B(_372_), .C(rst_bF_buf4), .Y(_161__0_) );
NAND2X1 NAND2X1_768 ( .A(CORE_InstructionIN_14_), .B(CORE_InstructionIN_12_), .Y(_375_) );
AOI22X1 AOI22X1_5 ( .A(_201_), .B(_207_), .C(_327_), .D(_375_), .Y(_376_) );
NAND2X1 NAND2X1_769 ( .A(CORE_InstructionIN_15_), .B(_376_), .Y(_377_) );
NAND3X1 NAND3X1_76 ( .A(_371_), .B(_182_), .C(CORE_ULA_ctrl_1_), .Y(_378_) );
AOI21X1 AOI21X1_42 ( .A(_377_), .B(_378_), .C(rst_bF_buf3), .Y(_161__1_) );
NAND3X1 NAND3X1_77 ( .A(_371_), .B(_182_), .C(CORE_ULA_ctrl_2_), .Y(_379_) );
NAND2X1 NAND2X1_770 ( .A(_189_), .B(_190_), .Y(_380_) );
NAND3X1 NAND3X1_78 ( .A(_380_), .B(CORE_InstructionIN_13_), .C(CORE_InstructionIN_15_), .Y(_381_) );
AOI21X1 AOI21X1_43 ( .A(_381_), .B(_379_), .C(rst_bF_buf3), .Y(_161__2_) );
NAND2X1 NAND2X1_771 ( .A(CORE_InstructionIN_14_), .B(CORE_InstructionIN_15_), .Y(_382_) );
NAND3X1 NAND3X1_79 ( .A(_371_), .B(_182_), .C(CORE_ULA_ctrl_3_), .Y(_383_) );
AOI21X1 AOI21X1_44 ( .A(_382_), .B(_383_), .C(rst_bF_buf3), .Y(_161__3_) );
INVX1 INVX1_263 ( .A(CORE_InstructionToULAMux_0_), .Y(_384_) );
AOI21X1 AOI21X1_45 ( .A(CORE_InstructionIN_13_), .B(CORE_InstructionIN_12_), .C(_303_), .Y(_385_) );
AOI21X1 AOI21X1_46 ( .A(_213_), .B(_385_), .C(_384_), .Y(_386_) );
AOI21X1 AOI21X1_47 ( .A(_176_), .B(_198_), .C(CORE_InstructionIN_14_), .Y(_387_) );
NOR3X1 NOR3X1_29 ( .A(_387_), .B(_201_), .C(_171_), .Y(_388_) );
OR2X2 OR2X2_952 ( .A(_388_), .B(_386_), .Y(_389_) );
AND2X2 AND2X2_1181 ( .A(_389_), .B(_197_), .Y(_390_) );
NAND3X1 NAND3X1_80 ( .A(_164_), .B(CORE_InstructionIN_11_), .C(CORE_InstructionIN_15_), .Y(_391_) );
NOR2X1 NOR2X1_131 ( .A(_337_), .B(_391_), .Y(_392_) );
OR2X2 OR2X2_953 ( .A(_392_), .B(_390_), .Y(_152__0_) );
NAND2X1 NAND2X1_772 ( .A(_172_), .B(_369_), .Y(_393_) );
OAI21X1 OAI21X1_96 ( .A(_393_), .B(_214_), .C(CORE_InstructionToULAMux_1_), .Y(_394_) );
NOR2X1 NOR2X1_132 ( .A(_275_), .B(_273_), .Y(_395_) );
AOI21X1 AOI21X1_48 ( .A(_395_), .B(_394_), .C(_200_), .Y(_152__1_) );
DFFNEGX1 DFFNEGX1_2 ( .CLK(clk_bF_buf28), .D(_163__0_), .Q(ID_old_rd_0_) );
DFFNEGX1 DFFNEGX1_3 ( .CLK(clk_bF_buf6), .D(_163__1_), .Q(ID_old_rd_1_) );
DFFNEGX1 DFFNEGX1_4 ( .CLK(clk_bF_buf28), .D(_163__2_), .Q(ID_old_rd_2_) );
DFFNEGX1 DFFNEGX1_5 ( .CLK(clk_bF_buf28), .D(_163__3_), .Q(ID_old_rd_3_) );
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf65), .D(_152__0_), .Q(CORE_InstructionToULAMux_0_) );
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf65), .D(_152__1_), .Q(CORE_InstructionToULAMux_1_) );
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf77), .D(_157_), .Q(CORE_REG_write) );
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf28), .D(_155__0_), .Q(CORE_REG_RF1_0_) );
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf28), .D(_155__1_), .Q(CORE_REG_RF1_1_) );
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf19), .D(_155__2_), .Q(CORE_REG_RF1_2_) );
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf53), .D(_155__3_), .Q(CORE_REG_RF1_3_) );
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf53), .D(_156__0_), .Q(CORE_REG_RF2_0_) );
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf69), .D(_156__1_), .Q(CORE_REG_RF2_1_) );
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf19), .D(_156__2_), .Q(CORE_REG_RF2_2_) );
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf53), .D(_156__3_), .Q(CORE_REG_RF2_3_) );
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf87), .D(_161__0_), .Q(ULA_cin) );
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf19), .D(_161__1_), .Q(CORE_ULA_ctrl_1_) );
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf53), .D(_161__2_), .Q(CORE_ULA_ctrl_2_) );
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf19), .D(_161__3_), .Q(CORE_ULA_ctrl_3_) );
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf0), .D(_159_), .Q(CORE_ULA_REGA_Stall) );
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf85), .D(_160_), .Q(CORE_ULA_REGB_Stall) );
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf77), .D(_158__0_), .Q(CORE_STACK_ctrl_0_) );
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf77), .D(_158__1_), .Q(CORE_STACK_ctrl_1_) );
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf65), .D(_153__0_), .Q(CORE_PC_ctrl_0_) );
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf77), .D(_153__1_), .Q(CORE_PC_ctrl_1_) );
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf65), .D(_148_), .Q(CORE_DATA_REGMux) );
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf28), .D(_154__0_), .Q(CORE_REG_RFD_0_) );
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf53), .D(_154__1_), .Q(CORE_REG_RFD_1_) );
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf28), .D(_154__2_), .Q(CORE_REG_RFD_2_) );
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf53), .D(_154__3_), .Q(CORE_REG_RFD_3_) );
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf77), .D(_151_), .Q(_145_) );
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf65), .D(_150_), .Q(_144_) );
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf65), .D(_149__0_), .Q(_142__0_) );
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf65), .D(_149__1_), .Q(_142__1_) );
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf65), .D(_149__2_), .Q(_142__2_) );
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf28), .D(_162__0_), .Q(ID_old_rd1_0_) );
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf6), .D(_162__1_), .Q(ID_old_rd1_1_) );
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf28), .D(_162__2_), .Q(ID_old_rd1_2_) );
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf53), .D(_162__3_), .Q(ID_old_rd1_3_) );
INVX1 INVX1_264 ( .A(PC_delay_0_), .Y(_404_) );
NOR2X1 NOR2X1_133 ( .A(_404_), .B(rst_bF_buf2), .Y(_403__1_) );
INVX1 INVX1_265 ( .A(CORE_PC_ctrl_1_), .Y(_405_) );
INVX1 INVX1_266 ( .A(CORE_PC_ctrl_0_), .Y(_406_) );
NAND2X1 NAND2X1_773 ( .A(_405_), .B(_406_), .Y(_407_) );
INVX1 INVX1_267 ( .A(_407_), .Y(_408_) );
NOR2X1 NOR2X1_134 ( .A(_408_), .B(rst_bF_buf2), .Y(_403__0_) );
INVX2 INVX2_6 ( .A(rst_bF_buf1), .Y(_409_) );
AND2X2 AND2X2_1182 ( .A(_409__bF_buf4), .B(PC_ADDR_stack_0__0_), .Y(_397__0_) );
AND2X2 AND2X2_1183 ( .A(_409__bF_buf4), .B(PC_ADDR_stack_0__1_), .Y(_397__1_) );
AND2X2 AND2X2_1184 ( .A(_409__bF_buf4), .B(PC_ADDR_stack_0__2_), .Y(_397__2_) );
AND2X2 AND2X2_1185 ( .A(_409__bF_buf1), .B(PC_ADDR_stack_0__3_), .Y(_397__3_) );
AND2X2 AND2X2_1186 ( .A(_409__bF_buf2), .B(PC_ADDR_stack_0__4_), .Y(_397__4_) );
AND2X2 AND2X2_1187 ( .A(_409__bF_buf4), .B(PC_ADDR_stack_0__5_), .Y(_397__5_) );
AND2X2 AND2X2_1188 ( .A(_409__bF_buf3), .B(PC_ADDR_stack_0__6_), .Y(_397__6_) );
AND2X2 AND2X2_1189 ( .A(_409__bF_buf3), .B(PC_ADDR_stack_0__7_), .Y(_397__7_) );
INVX1 INVX1_268 ( .A(PC_PC_pointer_0_), .Y(_410_) );
NOR2X1 NOR2X1_135 ( .A(_410_), .B(PC_PC_pointer_1_), .Y(_411_) );
INVX1 INVX1_269 ( .A(PC_PC_pointer_1_), .Y(_412_) );
NOR2X1 NOR2X1_136 ( .A(_410_), .B(_412_), .Y(_413_) );
AOI22X1 AOI22X1_6 ( .A(PC_PC_STACK_1__0_), .B(_411_), .C(PC_PC_STACK_3__0_), .D(_413_), .Y(_414_) );
NOR2X1 NOR2X1_137 ( .A(PC_PC_pointer_0_), .B(PC_PC_pointer_1_), .Y(_415_) );
NAND2X1 NAND2X1_774 ( .A(PC_PC_STACK_0__0_), .B(_415_), .Y(_416_) );
NOR2X1 NOR2X1_138 ( .A(_412_), .B(PC_PC_pointer_0_), .Y(_417_) );
NAND2X1 NAND2X1_775 ( .A(PC_PC_STACK_2__0_), .B(_417_), .Y(_418_) );
NAND3X1 NAND3X1_81 ( .A(_414_), .B(_416_), .C(_418_), .Y(_146__0_) );
AND2X2 AND2X2_1190 ( .A(_146__0_), .B(_409__bF_buf4), .Y(_396__0_) );
AOI22X1 AOI22X1_7 ( .A(PC_PC_STACK_1__1_), .B(_411_), .C(PC_PC_STACK_2__1_), .D(_417_), .Y(_419_) );
AOI22X1 AOI22X1_8 ( .A(PC_PC_STACK_0__1_), .B(_415_), .C(_413_), .D(PC_PC_STACK_3__1_), .Y(_420_) );
NAND2X1 NAND2X1_776 ( .A(_420_), .B(_419_), .Y(_146__1_) );
AOI21X1 AOI21X1_49 ( .A(_420_), .B(_419_), .C(rst_bF_buf0), .Y(_396__1_) );
AOI22X1 AOI22X1_9 ( .A(PC_PC_STACK_1__2_), .B(_411_), .C(PC_PC_STACK_2__2_), .D(_417_), .Y(_421_) );
AOI22X1 AOI22X1_10 ( .A(PC_PC_STACK_0__2_), .B(_415_), .C(_413_), .D(PC_PC_STACK_3__2_), .Y(_422_) );
NAND2X1 NAND2X1_777 ( .A(_422_), .B(_421_), .Y(_146__2_) );
AOI21X1 AOI21X1_50 ( .A(_422_), .B(_421_), .C(rst_bF_buf0), .Y(_396__2_) );
NAND2X1 NAND2X1_778 ( .A(PC_PC_STACK_0__3_), .B(_415_), .Y(_423_) );
NAND2X1 NAND2X1_779 ( .A(PC_PC_STACK_3__3_), .B(_413_), .Y(_424_) );
AOI22X1 AOI22X1_11 ( .A(PC_PC_STACK_1__3_), .B(_411_), .C(PC_PC_STACK_2__3_), .D(_417_), .Y(_425_) );
NAND3X1 NAND3X1_82 ( .A(_425_), .B(_423_), .C(_424_), .Y(_146__3_) );
AND2X2 AND2X2_1191 ( .A(_146__3_), .B(_409__bF_buf1), .Y(_396__3_) );
AOI22X1 AOI22X1_12 ( .A(PC_PC_STACK_1__4_), .B(_411_), .C(PC_PC_STACK_2__4_), .D(_417_), .Y(_426_) );
AOI22X1 AOI22X1_13 ( .A(PC_PC_STACK_0__4_), .B(_415_), .C(_413_), .D(PC_PC_STACK_3__4_), .Y(_427_) );
NAND2X1 NAND2X1_780 ( .A(_427_), .B(_426_), .Y(_146__4_) );
AOI21X1 AOI21X1_51 ( .A(_427_), .B(_426_), .C(rst_bF_buf0), .Y(_396__4_) );
NAND2X1 NAND2X1_781 ( .A(PC_PC_STACK_0__5_), .B(_415_), .Y(_428_) );
NAND2X1 NAND2X1_782 ( .A(PC_PC_STACK_2__5_), .B(_417_), .Y(_429_) );
AOI22X1 AOI22X1_14 ( .A(PC_PC_STACK_1__5_), .B(_411_), .C(PC_PC_STACK_3__5_), .D(_413_), .Y(_430_) );
NAND3X1 NAND3X1_83 ( .A(_430_), .B(_428_), .C(_429_), .Y(_146__5_) );
AND2X2 AND2X2_1192 ( .A(_146__5_), .B(_409__bF_buf4), .Y(_396__5_) );
NAND2X1 NAND2X1_783 ( .A(PC_PC_STACK_0__6_), .B(_415_), .Y(_431_) );
NAND2X1 NAND2X1_784 ( .A(PC_PC_STACK_3__6_), .B(_413_), .Y(_432_) );
AOI22X1 AOI22X1_15 ( .A(PC_PC_STACK_1__6_), .B(_411_), .C(PC_PC_STACK_2__6_), .D(_417_), .Y(_433_) );
NAND3X1 NAND3X1_84 ( .A(_433_), .B(_431_), .C(_432_), .Y(_146__6_) );
AND2X2 AND2X2_1193 ( .A(_146__6_), .B(_409__bF_buf3), .Y(_396__6_) );
NAND2X1 NAND2X1_785 ( .A(PC_PC_STACK_0__7_), .B(_415_), .Y(_434_) );
NAND2X1 NAND2X1_786 ( .A(PC_PC_STACK_3__7_), .B(_413_), .Y(_435_) );
AOI22X1 AOI22X1_16 ( .A(PC_PC_STACK_1__7_), .B(_411_), .C(PC_PC_STACK_2__7_), .D(_417_), .Y(_436_) );
NAND3X1 NAND3X1_85 ( .A(_436_), .B(_434_), .C(_435_), .Y(_146__7_) );
AND2X2 AND2X2_1194 ( .A(_146__7_), .B(_409__bF_buf3), .Y(_396__7_) );
XNOR2X1 XNOR2X1_57 ( .A(CORE_STACK_ctrl_0_), .B(INTERRUPT_flag_bF_buf14_bF_buf3), .Y(_437_) );
OR2X2 OR2X2_954 ( .A(CORE_STACK_ctrl_1_), .B(_437_), .Y(_438_) );
INVX1 INVX1_270 ( .A(CORE_STACK_ctrl_1_), .Y(_439_) );
OR2X2 OR2X2_955 ( .A(CORE_STACK_ctrl_0_), .B(INTERRUPT_flag_bF_buf13_bF_buf0), .Y(_440_) );
OR2X2 OR2X2_956 ( .A(_440_), .B(_439_), .Y(_441_) );
AND2X2 AND2X2_1195 ( .A(_438_), .B(_441_), .Y(_442_) );
XOR2X1 XOR2X1_70 ( .A(PC_PC_pointer_0_), .B(_442_), .Y(_443_) );
NOR2X1 NOR2X1_139 ( .A(_443_), .B(rst_bF_buf1), .Y(_402__0_) );
NAND3X1 NAND3X1_86 ( .A(_438_), .B(PC_PC_pointer_1_), .C(_441_), .Y(_444_) );
XNOR2X1 XNOR2X1_58 ( .A(PC_PC_pointer_0_), .B(PC_PC_pointer_1_), .Y(_445_) );
AND2X2 AND2X2_1196 ( .A(_441_), .B(_445_), .Y(_446_) );
XOR2X1 XOR2X1_71 ( .A(PC_PC_pointer_0_), .B(PC_PC_pointer_1_), .Y(_447_) );
AND2X2 AND2X2_1197 ( .A(_438_), .B(_447_), .Y(_448_) );
OR2X2 OR2X2_957 ( .A(_446_), .B(_448_), .Y(_449_) );
AND2X2 AND2X2_1198 ( .A(_444_), .B(_449_), .Y(_450_) );
NOR2X1 NOR2X1_140 ( .A(_450_), .B(rst_bF_buf1), .Y(_402__1_) );
AND2X2 AND2X2_1199 ( .A(_450_), .B(_443_), .Y(_451_) );
AND2X2 AND2X2_1200 ( .A(_451__bF_buf3), .B(PC_PC_STACK_0__0_), .Y(_452_) );
INVX1 INVX1_271 ( .A(_452_), .Y(_453_) );
INVX1 INVX1_272 ( .A(INTERRUPT_flag_bF_buf12_bF_buf2), .Y(_454_) );
NAND2X1 NAND2X1_787 ( .A(_406_), .B(_454_), .Y(_455_) );
INVX1 INVX1_273 ( .A(_455_), .Y(_456_) );
OR2X2 OR2X2_958 ( .A(PC_PC_STACK_0__0_), .B(_451__bF_buf3), .Y(_457_) );
NAND3X1 NAND3X1_87 ( .A(_453_), .B(_456__bF_buf3), .C(_457_), .Y(_458_) );
NAND2X1 NAND2X1_788 ( .A(CORE_PC_ctrl_0_), .B(INTERRUPT_flag_bF_buf11_bF_buf1), .Y(_459_) );
INVX1 INVX1_274 ( .A(_459_), .Y(_460_) );
NAND2X1 NAND2X1_789 ( .A(PC_PC_STACK_0__0_), .B(_460_), .Y(_461_) );
INVX1 INVX1_275 ( .A(INTERRUPT_ch[0]), .Y(_462_) );
NAND2X1 NAND2X1_790 ( .A(INTERRUPT_flag_bF_buf10_bF_buf3), .B(_406_), .Y(_463_) );
AOI21X1 AOI21X1_52 ( .A(_462_), .B(_451__bF_buf3), .C(_463_), .Y(_464_) );
INVX1 INVX1_276 ( .A(PC_ULA_OUT_0_), .Y(_465_) );
NAND2X1 NAND2X1_791 ( .A(CORE_PC_ctrl_0_), .B(_454_), .Y(_466_) );
AOI21X1 AOI21X1_53 ( .A(_465_), .B(_451__bF_buf3), .C(_466__bF_buf2), .Y(_467_) );
OAI21X1 OAI21X1_97 ( .A(_464_), .B(_467_), .C(_457_), .Y(_468_) );
NAND3X1 NAND3X1_88 ( .A(_468_), .B(_461_), .C(_458_), .Y(_469_) );
AND2X2 AND2X2_1201 ( .A(_469_), .B(_409__bF_buf1), .Y(_398__0_) );
INVX1 INVX1_277 ( .A(_451__bF_buf2), .Y(_470_) );
NAND2X1 NAND2X1_792 ( .A(PC_PC_STACK_0__1_), .B(_470__bF_buf3), .Y(_471_) );
XOR2X1 XOR2X1_72 ( .A(_410_), .B(_442_), .Y(_472_) );
AND2X2 AND2X2_1202 ( .A(_450_), .B(_472_), .Y(_473_) );
AND2X2 AND2X2_1203 ( .A(_473__bF_buf0), .B(PC_PC_STACK_1__0_), .Y(_474_) );
AND2X2 AND2X2_1204 ( .A(_442_), .B(PC_PC_pointer_1_), .Y(_475_) );
AOI21X1 AOI21X1_54 ( .A(CORE_STACK_ctrl_0_), .B(INTERRUPT_flag_bF_buf9_bF_buf0), .C(CORE_STACK_ctrl_1_), .Y(_476_) );
AND2X2 AND2X2_1205 ( .A(_476_), .B(_440_), .Y(_477_) );
AND2X2 AND2X2_1206 ( .A(_477_), .B(_447_), .Y(_478_) );
INVX1 INVX1_278 ( .A(_440_), .Y(_479_) );
AND2X2 AND2X2_1207 ( .A(_479_), .B(CORE_STACK_ctrl_1_), .Y(_480_) );
AND2X2 AND2X2_1208 ( .A(_480_), .B(_445_), .Y(_481_) );
OR2X2 OR2X2_959 ( .A(_478_), .B(_481_), .Y(_482_) );
OR2X2 OR2X2_960 ( .A(_475_), .B(_482_), .Y(_483_) );
AND2X2 AND2X2_1209 ( .A(_483_), .B(_443_), .Y(_484_) );
AND2X2 AND2X2_1210 ( .A(_484__bF_buf2), .B(PC_PC_STACK_2__0_), .Y(_485_) );
OR2X2 OR2X2_961 ( .A(_474_), .B(_485_), .Y(_486_) );
AND2X2 AND2X2_1211 ( .A(_483_), .B(_472_), .Y(_487_) );
AND2X2 AND2X2_1212 ( .A(_487__bF_buf0), .B(PC_PC_STACK_3__0_), .Y(_488_) );
OR2X2 OR2X2_962 ( .A(_452_), .B(_488_), .Y(_489_) );
OR2X2 OR2X2_963 ( .A(_486_), .B(_489_), .Y(_490_) );
AND2X2 AND2X2_1213 ( .A(_484__bF_buf3), .B(PC_PC_STACK_2__1_), .Y(_491_) );
AND2X2 AND2X2_1214 ( .A(_487__bF_buf3), .B(PC_PC_STACK_3__1_), .Y(_492_) );
OR2X2 OR2X2_964 ( .A(_491_), .B(_492_), .Y(_493_) );
AND2X2 AND2X2_1215 ( .A(_451__bF_buf0), .B(PC_PC_STACK_0__1_), .Y(_494_) );
AND2X2 AND2X2_1216 ( .A(_473__bF_buf2), .B(PC_PC_STACK_1__1_), .Y(_495_) );
OR2X2 OR2X2_965 ( .A(_494_), .B(_495_), .Y(_496_) );
OR2X2 OR2X2_966 ( .A(_493_), .B(_496_), .Y(_497_) );
XOR2X1 XOR2X1_73 ( .A(_490_), .B(_497_), .Y(_498_) );
NAND2X1 NAND2X1_793 ( .A(_451__bF_buf0), .B(_498_), .Y(_499_) );
NAND2X1 NAND2X1_794 ( .A(_471_), .B(_499_), .Y(_500_) );
NAND2X1 NAND2X1_795 ( .A(_456__bF_buf3), .B(_500_), .Y(_501_) );
NAND2X1 NAND2X1_796 ( .A(_463_), .B(_466__bF_buf1), .Y(_502_) );
NAND3X1 NAND3X1_89 ( .A(_470__bF_buf3), .B(PC_PC_STACK_0__1_), .C(_502_), .Y(_503_) );
INVX1 INVX1_279 ( .A(PC_ULA_OUT_1_), .Y(_504_) );
INVX1 INVX1_280 ( .A(_463_), .Y(_505_) );
NAND2X1 NAND2X1_797 ( .A(INTERRUPT_ch[1]), .B(_505__bF_buf3), .Y(_506_) );
OAI21X1 OAI21X1_98 ( .A(_504_), .B(_466__bF_buf2), .C(_506_), .Y(_507_) );
AOI22X1 AOI22X1_17 ( .A(PC_PC_STACK_0__1_), .B(_460_), .C(_507_), .D(_451__bF_buf0), .Y(_508_) );
AND2X2 AND2X2_1217 ( .A(_508_), .B(_503_), .Y(_509_) );
AOI21X1 AOI21X1_55 ( .A(_509_), .B(_501_), .C(rst_bF_buf1), .Y(_398__1_) );
NAND2X1 NAND2X1_798 ( .A(PC_PC_STACK_0__2_), .B(_470__bF_buf3), .Y(_510_) );
AND2X2 AND2X2_1218 ( .A(_490_), .B(_497_), .Y(_511_) );
AND2X2 AND2X2_1219 ( .A(_473__bF_buf2), .B(PC_PC_STACK_1__2_), .Y(_512_) );
AND2X2 AND2X2_1220 ( .A(_487__bF_buf0), .B(PC_PC_STACK_3__2_), .Y(_513_) );
OR2X2 OR2X2_967 ( .A(_512_), .B(_513_), .Y(_514_) );
AND2X2 AND2X2_1221 ( .A(_451__bF_buf3), .B(PC_PC_STACK_0__2_), .Y(_515_) );
AND2X2 AND2X2_1222 ( .A(_484__bF_buf3), .B(PC_PC_STACK_2__2_), .Y(_516_) );
OR2X2 OR2X2_968 ( .A(_515_), .B(_516_), .Y(_517_) );
OR2X2 OR2X2_969 ( .A(_514_), .B(_517_), .Y(_518_) );
XNOR2X1 XNOR2X1_59 ( .A(_518_), .B(_511_), .Y(_519_) );
OAI21X1 OAI21X1_99 ( .A(_470__bF_buf3), .B(_519_), .C(_510_), .Y(_520_) );
NAND2X1 NAND2X1_799 ( .A(_456__bF_buf3), .B(_520_), .Y(_521_) );
NAND2X1 NAND2X1_800 ( .A(PC_PC_STACK_0__2_), .B(_460_), .Y(_522_) );
INVX1 INVX1_281 ( .A(_466__bF_buf0), .Y(_523_) );
NAND2X1 NAND2X1_801 ( .A(PC_ULA_OUT_2_), .B(_451__bF_buf3), .Y(_524_) );
NAND2X1 NAND2X1_802 ( .A(_524_), .B(_510_), .Y(_525_) );
INVX1 INVX1_282 ( .A(INTERRUPT_ch[2]), .Y(_526_) );
OAI21X1 OAI21X1_100 ( .A(_526_), .B(_470__bF_buf1), .C(_510_), .Y(_527_) );
AOI22X1 AOI22X1_18 ( .A(_523_), .B(_525_), .C(_505__bF_buf3), .D(_527_), .Y(_528_) );
NAND3X1 NAND3X1_90 ( .A(_521_), .B(_522_), .C(_528_), .Y(_529_) );
AND2X2 AND2X2_1223 ( .A(_529_), .B(_409__bF_buf1), .Y(_398__2_) );
NAND2X1 NAND2X1_803 ( .A(PC_PC_STACK_0__3_), .B(_470__bF_buf2), .Y(_530_) );
AND2X2 AND2X2_1224 ( .A(_511_), .B(_518_), .Y(_531_) );
AND2X2 AND2X2_1225 ( .A(_451__bF_buf2), .B(PC_PC_STACK_0__3_), .Y(_532_) );
AND2X2 AND2X2_1226 ( .A(_484__bF_buf2), .B(PC_PC_STACK_2__3_), .Y(_533_) );
OR2X2 OR2X2_970 ( .A(_532_), .B(_533_), .Y(_534_) );
AND2X2 AND2X2_1227 ( .A(_473__bF_buf1), .B(PC_PC_STACK_1__3_), .Y(_535_) );
AND2X2 AND2X2_1228 ( .A(_487__bF_buf1), .B(PC_PC_STACK_3__3_), .Y(_536_) );
OR2X2 OR2X2_971 ( .A(_535_), .B(_536_), .Y(_537_) );
OR2X2 OR2X2_972 ( .A(_534_), .B(_537_), .Y(_538_) );
XOR2X1 XOR2X1_74 ( .A(_538_), .B(_531_), .Y(_539_) );
NAND2X1 NAND2X1_804 ( .A(_451__bF_buf2), .B(_539_), .Y(_540_) );
AOI21X1 AOI21X1_56 ( .A(_530_), .B(_540_), .C(_455_), .Y(_541_) );
NAND2X1 NAND2X1_805 ( .A(PC_PC_STACK_0__3_), .B(_460_), .Y(_542_) );
INVX1 INVX1_283 ( .A(PC_ULA_OUT_3_), .Y(_543_) );
OAI21X1 OAI21X1_101 ( .A(_543_), .B(_470__bF_buf2), .C(_530_), .Y(_544_) );
INVX1 INVX1_284 ( .A(INTERRUPT_ch[3]), .Y(_545_) );
OAI21X1 OAI21X1_102 ( .A(_545_), .B(_470__bF_buf2), .C(_530_), .Y(_546_) );
AOI22X1 AOI22X1_19 ( .A(_505__bF_buf0), .B(_546_), .C(_523_), .D(_544_), .Y(_547_) );
NAND2X1 NAND2X1_806 ( .A(_542_), .B(_547_), .Y(_548_) );
OR2X2 OR2X2_973 ( .A(_541_), .B(_548_), .Y(_549_) );
AND2X2 AND2X2_1229 ( .A(_549_), .B(_409__bF_buf5), .Y(_398__3_) );
NAND2X1 NAND2X1_807 ( .A(PC_PC_STACK_0__4_), .B(_470__bF_buf0), .Y(_550_) );
AND2X2 AND2X2_1230 ( .A(_531_), .B(_538_), .Y(_551_) );
AOI22X1 AOI22X1_20 ( .A(PC_PC_STACK_3__4_), .B(_487__bF_buf1), .C(PC_PC_STACK_2__4_), .D(_484__bF_buf0), .Y(_552_) );
NAND2X1 NAND2X1_808 ( .A(PC_PC_STACK_0__4_), .B(_451__bF_buf1), .Y(_553_) );
NAND2X1 NAND2X1_809 ( .A(PC_PC_STACK_1__4_), .B(_473__bF_buf1), .Y(_554_) );
NAND3X1 NAND3X1_91 ( .A(_552_), .B(_553_), .C(_554_), .Y(_555_) );
XNOR2X1 XNOR2X1_60 ( .A(_555_), .B(_551_), .Y(_556_) );
OAI21X1 OAI21X1_103 ( .A(_470__bF_buf0), .B(_556_), .C(_550_), .Y(_557_) );
NAND2X1 NAND2X1_810 ( .A(_456__bF_buf3), .B(_557_), .Y(_558_) );
NAND2X1 NAND2X1_811 ( .A(PC_PC_STACK_0__4_), .B(_460_), .Y(_559_) );
INVX1 INVX1_285 ( .A(INTERRUPT_ch[4]), .Y(_560_) );
OAI21X1 OAI21X1_104 ( .A(_560_), .B(_470__bF_buf0), .C(_550_), .Y(_561_) );
NAND2X1 NAND2X1_812 ( .A(PC_ULA_OUT_4_), .B(_451__bF_buf2), .Y(_562_) );
NAND2X1 NAND2X1_813 ( .A(_562_), .B(_550_), .Y(_563_) );
AOI22X1 AOI22X1_21 ( .A(_523_), .B(_563_), .C(_505__bF_buf2), .D(_561_), .Y(_564_) );
AND2X2 AND2X2_1231 ( .A(_564_), .B(_559_), .Y(_565_) );
AOI21X1 AOI21X1_57 ( .A(_565_), .B(_558_), .C(rst_bF_buf0), .Y(_398__4_) );
AND2X2 AND2X2_1232 ( .A(_551_), .B(_555_), .Y(_566_) );
AOI22X1 AOI22X1_22 ( .A(PC_PC_STACK_1__5_), .B(_473__bF_buf1), .C(PC_PC_STACK_2__5_), .D(_484__bF_buf2), .Y(_567_) );
AOI22X1 AOI22X1_23 ( .A(PC_PC_STACK_3__5_), .B(_487__bF_buf3), .C(PC_PC_STACK_0__5_), .D(_451__bF_buf2), .Y(_568_) );
NAND2X1 NAND2X1_814 ( .A(_567_), .B(_568_), .Y(_569_) );
XOR2X1 XOR2X1_75 ( .A(_569_), .B(_566_), .Y(_570_) );
MUX2X1 MUX2X1_814 ( .A(_570_), .B(PC_PC_STACK_0__5_), .S(_451__bF_buf2), .Y(_571_) );
OR2X2 OR2X2_974 ( .A(_455_), .B(_571_), .Y(_572_) );
NAND2X1 NAND2X1_815 ( .A(PC_PC_STACK_0__5_), .B(_460_), .Y(_573_) );
INVX1 INVX1_286 ( .A(PC_ULA_OUT_5_), .Y(_574_) );
NAND2X1 NAND2X1_816 ( .A(PC_PC_STACK_0__5_), .B(_470__bF_buf1), .Y(_575_) );
OAI21X1 OAI21X1_105 ( .A(_574_), .B(_470__bF_buf1), .C(_575_), .Y(_576_) );
INVX1 INVX1_287 ( .A(INTERRUPT_ch[5]), .Y(_577_) );
OAI21X1 OAI21X1_106 ( .A(_577_), .B(_470__bF_buf1), .C(_575_), .Y(_578_) );
AOI22X1 AOI22X1_24 ( .A(_505__bF_buf2), .B(_578_), .C(_523_), .D(_576_), .Y(_579_) );
NAND3X1 NAND3X1_92 ( .A(_572_), .B(_573_), .C(_579_), .Y(_580_) );
AND2X2 AND2X2_1233 ( .A(_580_), .B(_409__bF_buf5), .Y(_398__5_) );
NAND2X1 NAND2X1_817 ( .A(PC_PC_STACK_0__6_), .B(_470__bF_buf2), .Y(_581_) );
AND2X2 AND2X2_1234 ( .A(_566_), .B(_569_), .Y(_582_) );
AOI22X1 AOI22X1_25 ( .A(PC_PC_STACK_3__6_), .B(_487__bF_buf2), .C(PC_PC_STACK_2__6_), .D(_484__bF_buf0), .Y(_583_) );
NAND2X1 NAND2X1_818 ( .A(PC_PC_STACK_0__6_), .B(_451__bF_buf1), .Y(_584_) );
NAND2X1 NAND2X1_819 ( .A(PC_PC_STACK_1__6_), .B(_473__bF_buf1), .Y(_585_) );
NAND3X1 NAND3X1_93 ( .A(_583_), .B(_584_), .C(_585_), .Y(_586_) );
XNOR2X1 XNOR2X1_61 ( .A(_586_), .B(_582_), .Y(_587_) );
OAI21X1 OAI21X1_107 ( .A(_470__bF_buf2), .B(_587_), .C(_581_), .Y(_588_) );
AND2X2 AND2X2_1235 ( .A(_588_), .B(_456__bF_buf2), .Y(_589_) );
MUX2X1 MUX2X1_815 ( .A(INTERRUPT_ch[6]), .B(PC_PC_STACK_0__6_), .S(_451__bF_buf1), .Y(_590_) );
NAND2X1 NAND2X1_820 ( .A(PC_ULA_OUT_6_), .B(_451__bF_buf1), .Y(_591_) );
NAND2X1 NAND2X1_821 ( .A(_591_), .B(_581_), .Y(_592_) );
AOI22X1 AOI22X1_26 ( .A(PC_PC_STACK_0__6_), .B(_460_), .C(_592_), .D(_523_), .Y(_593_) );
OAI21X1 OAI21X1_108 ( .A(_463_), .B(_590_), .C(_593_), .Y(_594_) );
OR2X2 OR2X2_975 ( .A(_594_), .B(_589_), .Y(_595_) );
AND2X2 AND2X2_1236 ( .A(_595_), .B(_409__bF_buf0), .Y(_398__6_) );
NAND2X1 NAND2X1_822 ( .A(PC_PC_STACK_0__7_), .B(_470__bF_buf0), .Y(_596_) );
INVX1 INVX1_288 ( .A(_596_), .Y(_597_) );
AND2X2 AND2X2_1237 ( .A(_582_), .B(_586_), .Y(_598_) );
INVX1 INVX1_289 ( .A(PC_PC_STACK_0__7_), .Y(_599_) );
NAND2X1 NAND2X1_823 ( .A(PC_PC_STACK_1__7_), .B(_473__bF_buf3), .Y(_600_) );
INVX1 INVX1_290 ( .A(_484__bF_buf0), .Y(_601_) );
INVX1 INVX1_291 ( .A(PC_PC_STACK_3__7_), .Y(_602_) );
OAI21X1 OAI21X1_109 ( .A(_602_), .B(_450_), .C(_472_), .Y(_603_) );
OAI21X1 OAI21X1_110 ( .A(PC_PC_STACK_2__7_), .B(_601__bF_buf3), .C(_603_), .Y(_604_) );
AOI22X1 AOI22X1_27 ( .A(_599_), .B(_451__bF_buf0), .C(_604_), .D(_600_), .Y(_605_) );
XOR2X1 XOR2X1_76 ( .A(_605_), .B(_598_), .Y(_606_) );
AND2X2 AND2X2_1238 ( .A(_606_), .B(_451__bF_buf0), .Y(_607_) );
OR2X2 OR2X2_976 ( .A(_597_), .B(_607_), .Y(_608_) );
AND2X2 AND2X2_1239 ( .A(_608_), .B(_456__bF_buf3), .Y(_609_) );
NAND2X1 NAND2X1_824 ( .A(INTERRUPT_ch[7]), .B(_451__bF_buf1), .Y(_610_) );
NAND2X1 NAND2X1_825 ( .A(_610_), .B(_596_), .Y(_611_) );
INVX1 INVX1_292 ( .A(PC_ULA_OUT_7_), .Y(_612_) );
OAI21X1 OAI21X1_111 ( .A(_612_), .B(_470__bF_buf3), .C(_596_), .Y(_613_) );
AOI22X1 AOI22X1_28 ( .A(_505__bF_buf3), .B(_611_), .C(_523_), .D(_613_), .Y(_614_) );
OAI21X1 OAI21X1_112 ( .A(_599_), .B(_459_), .C(_614_), .Y(_615_) );
OR2X2 OR2X2_977 ( .A(_615_), .B(_609_), .Y(_616_) );
AND2X2 AND2X2_1240 ( .A(_616_), .B(_409__bF_buf2), .Y(_398__7_) );
NAND2X1 NAND2X1_826 ( .A(_409__bF_buf2), .B(_459_), .Y(_617_) );
NAND2X1 NAND2X1_827 ( .A(PC_PC_STACK_3__0_), .B(_617__bF_buf1), .Y(_618_) );
NOR2X1 NOR2X1_141 ( .A(_488_), .B(_455_), .Y(_619_) );
NAND2X1 NAND2X1_828 ( .A(_462_), .B(_466__bF_buf2), .Y(_620_) );
OAI21X1 OAI21X1_113 ( .A(PC_ULA_OUT_0_), .B(_505__bF_buf3), .C(_620_), .Y(_621_) );
NAND2X1 NAND2X1_829 ( .A(_487__bF_buf0), .B(_621_), .Y(_622_) );
AOI21X1 AOI21X1_58 ( .A(_502_), .B(_622_), .C(_619_), .Y(_623_) );
OAI21X1 OAI21X1_114 ( .A(PC_PC_STACK_3__0_), .B(_487__bF_buf0), .C(_409__bF_buf5), .Y(_624_) );
OAI21X1 OAI21X1_115 ( .A(_624_), .B(_623_), .C(_618_), .Y(_401__0_) );
NAND2X1 NAND2X1_830 ( .A(PC_PC_STACK_3__1_), .B(_617__bF_buf0), .Y(_625_) );
INVX1 INVX1_293 ( .A(_487__bF_buf1), .Y(_626_) );
AOI22X1 AOI22X1_29 ( .A(INTERRUPT_ch[1]), .B(_505__bF_buf3), .C(_498_), .D(_456__bF_buf3), .Y(_627_) );
OR2X2 OR2X2_978 ( .A(_626__bF_buf3), .B(_627_), .Y(_628_) );
NAND2X1 NAND2X1_831 ( .A(PC_PC_STACK_3__1_), .B(_626__bF_buf3), .Y(_629_) );
OAI21X1 OAI21X1_116 ( .A(_504_), .B(_626__bF_buf3), .C(_629_), .Y(_630_) );
AND2X2 AND2X2_1241 ( .A(_406_), .B(PC_PC_STACK_3__1_), .Y(_631_) );
AOI22X1 AOI22X1_30 ( .A(_626__bF_buf3), .B(_631_), .C(_630_), .D(_523_), .Y(_632_) );
AND2X2 AND2X2_1242 ( .A(_632_), .B(_628_), .Y(_633_) );
OAI21X1 OAI21X1_117 ( .A(rst_bF_buf1), .B(_633_), .C(_625_), .Y(_401__1_) );
NAND2X1 NAND2X1_832 ( .A(PC_PC_STACK_3__2_), .B(_617__bF_buf0), .Y(_634_) );
NOR3X1 NOR3X1_30 ( .A(_519_), .B(_455_), .C(_626__bF_buf3), .Y(_635_) );
AND2X2 AND2X2_1243 ( .A(_626__bF_buf1), .B(PC_PC_STACK_3__2_), .Y(_636_) );
AOI21X1 AOI21X1_59 ( .A(PC_ULA_OUT_2_), .B(_487__bF_buf3), .C(_636_), .Y(_637_) );
NOR2X1 NOR2X1_142 ( .A(_463_), .B(_526_), .Y(_638_) );
AOI22X1 AOI22X1_31 ( .A(_487__bF_buf3), .B(_638_), .C(_636_), .D(_406_), .Y(_639_) );
OAI21X1 OAI21X1_118 ( .A(_466__bF_buf2), .B(_637_), .C(_639_), .Y(_640_) );
OAI21X1 OAI21X1_119 ( .A(_640_), .B(_635_), .C(_409__bF_buf1), .Y(_641_) );
NAND2X1 NAND2X1_833 ( .A(_634_), .B(_641_), .Y(_401__2_) );
INVX1 INVX1_294 ( .A(PC_PC_STACK_3__3_), .Y(_642_) );
INVX1 INVX1_295 ( .A(_617__bF_buf3), .Y(_643_) );
NOR2X1 NOR2X1_143 ( .A(_643_), .B(_642_), .Y(_644_) );
OR2X2 OR2X2_979 ( .A(_626__bF_buf0), .B(_539_), .Y(_645_) );
NAND2X1 NAND2X1_834 ( .A(_642_), .B(_626__bF_buf0), .Y(_646_) );
NAND3X1 NAND3X1_94 ( .A(_645_), .B(_456__bF_buf1), .C(_646_), .Y(_647_) );
NAND2X1 NAND2X1_835 ( .A(PC_PC_STACK_3__3_), .B(_626__bF_buf0), .Y(_648_) );
OAI21X1 OAI21X1_120 ( .A(_545_), .B(_626__bF_buf0), .C(_648_), .Y(_649_) );
NAND2X1 NAND2X1_836 ( .A(_505__bF_buf0), .B(_649_), .Y(_650_) );
OAI21X1 OAI21X1_121 ( .A(_543_), .B(_626__bF_buf0), .C(_648_), .Y(_651_) );
NAND2X1 NAND2X1_837 ( .A(_523_), .B(_651_), .Y(_652_) );
NAND3X1 NAND3X1_95 ( .A(_647_), .B(_650_), .C(_652_), .Y(_653_) );
AND2X2 AND2X2_1244 ( .A(_653_), .B(_409__bF_buf0), .Y(_654_) );
OR2X2 OR2X2_980 ( .A(_644_), .B(_654_), .Y(_401__3_) );
AND2X2 AND2X2_1245 ( .A(_617__bF_buf3), .B(PC_PC_STACK_3__4_), .Y(_655_) );
NAND2X1 NAND2X1_838 ( .A(PC_PC_STACK_3__4_), .B(_626__bF_buf2), .Y(_656_) );
OAI21X1 OAI21X1_122 ( .A(_626__bF_buf2), .B(_556_), .C(_656_), .Y(_657_) );
AND2X2 AND2X2_1246 ( .A(_657_), .B(_456__bF_buf0), .Y(_658_) );
OAI21X1 OAI21X1_123 ( .A(_560_), .B(_626__bF_buf2), .C(_656_), .Y(_659_) );
NAND2X1 NAND2X1_839 ( .A(_505__bF_buf0), .B(_659_), .Y(_660_) );
MUX2X1 MUX2X1_816 ( .A(PC_ULA_OUT_4_), .B(PC_PC_STACK_3__4_), .S(_487__bF_buf1), .Y(_661_) );
OAI21X1 OAI21X1_124 ( .A(_466__bF_buf0), .B(_661_), .C(_660_), .Y(_662_) );
OR2X2 OR2X2_981 ( .A(_658_), .B(_662_), .Y(_663_) );
AND2X2 AND2X2_1247 ( .A(_663_), .B(_409__bF_buf0), .Y(_664_) );
OR2X2 OR2X2_982 ( .A(_655_), .B(_664_), .Y(_401__4_) );
NAND2X1 NAND2X1_840 ( .A(PC_PC_STACK_3__5_), .B(_617__bF_buf3), .Y(_665_) );
OR2X2 OR2X2_983 ( .A(PC_PC_STACK_3__5_), .B(_487__bF_buf3), .Y(_666_) );
OAI21X1 OAI21X1_125 ( .A(_626__bF_buf1), .B(_570_), .C(_666_), .Y(_667_) );
OR2X2 OR2X2_984 ( .A(_455_), .B(_667_), .Y(_668_) );
NAND2X1 NAND2X1_841 ( .A(PC_PC_STACK_3__5_), .B(_626__bF_buf1), .Y(_669_) );
OAI21X1 OAI21X1_126 ( .A(_577_), .B(_626__bF_buf1), .C(_669_), .Y(_670_) );
OAI21X1 OAI21X1_127 ( .A(_574_), .B(_626__bF_buf1), .C(_669_), .Y(_671_) );
AOI22X1 AOI22X1_32 ( .A(_505__bF_buf2), .B(_670_), .C(_523_), .D(_671_), .Y(_672_) );
AND2X2 AND2X2_1248 ( .A(_668_), .B(_672_), .Y(_673_) );
OAI21X1 OAI21X1_128 ( .A(rst_bF_buf0), .B(_673_), .C(_665_), .Y(_401__5_) );
AND2X2 AND2X2_1249 ( .A(_617__bF_buf2), .B(PC_PC_STACK_3__6_), .Y(_674_) );
NAND2X1 NAND2X1_842 ( .A(PC_PC_STACK_3__6_), .B(_626__bF_buf2), .Y(_675_) );
OAI21X1 OAI21X1_129 ( .A(_626__bF_buf2), .B(_587_), .C(_675_), .Y(_676_) );
AND2X2 AND2X2_1250 ( .A(_676_), .B(_456__bF_buf0), .Y(_677_) );
INVX1 INVX1_296 ( .A(INTERRUPT_ch[6]), .Y(_678_) );
OAI21X1 OAI21X1_130 ( .A(_678_), .B(_626__bF_buf2), .C(_675_), .Y(_679_) );
NAND2X1 NAND2X1_843 ( .A(_505__bF_buf1), .B(_679_), .Y(_680_) );
MUX2X1 MUX2X1_817 ( .A(PC_ULA_OUT_6_), .B(PC_PC_STACK_3__6_), .S(_487__bF_buf2), .Y(_681_) );
OAI21X1 OAI21X1_131 ( .A(_466__bF_buf3), .B(_681_), .C(_680_), .Y(_682_) );
OR2X2 OR2X2_985 ( .A(_682_), .B(_677_), .Y(_683_) );
AND2X2 AND2X2_1251 ( .A(_683_), .B(_409__bF_buf3), .Y(_684_) );
OR2X2 OR2X2_986 ( .A(_674_), .B(_684_), .Y(_401__6_) );
NOR2X1 NOR2X1_144 ( .A(_643_), .B(_602_), .Y(_685_) );
NOR2X1 NOR2X1_145 ( .A(_487__bF_buf2), .B(_602_), .Y(_686_) );
AND2X2 AND2X2_1252 ( .A(_606_), .B(_487__bF_buf2), .Y(_687_) );
OR2X2 OR2X2_987 ( .A(_686_), .B(_687_), .Y(_688_) );
AND2X2 AND2X2_1253 ( .A(_688_), .B(_456__bF_buf2), .Y(_689_) );
NOR2X1 NOR2X1_146 ( .A(_626__bF_buf3), .B(_612_), .Y(_690_) );
OAI21X1 OAI21X1_132 ( .A(_686_), .B(_690_), .C(_523_), .Y(_691_) );
AOI21X1 AOI21X1_60 ( .A(INTERRUPT_ch[7]), .B(_487__bF_buf2), .C(_686_), .Y(_692_) );
OAI21X1 OAI21X1_133 ( .A(_463_), .B(_692_), .C(_691_), .Y(_693_) );
OR2X2 OR2X2_988 ( .A(_693_), .B(_689_), .Y(_694_) );
AND2X2 AND2X2_1254 ( .A(_694_), .B(_409__bF_buf2), .Y(_695_) );
OR2X2 OR2X2_989 ( .A(_685_), .B(_695_), .Y(_401__7_) );
NAND2X1 NAND2X1_844 ( .A(PC_PC_STACK_2__0_), .B(_617__bF_buf1), .Y(_696_) );
NOR2X1 NOR2X1_147 ( .A(_485_), .B(_455_), .Y(_697_) );
NAND2X1 NAND2X1_845 ( .A(_484__bF_buf3), .B(_621_), .Y(_698_) );
AOI21X1 AOI21X1_61 ( .A(_502_), .B(_698_), .C(_697_), .Y(_699_) );
OAI21X1 OAI21X1_134 ( .A(PC_PC_STACK_2__0_), .B(_484__bF_buf2), .C(_409__bF_buf5), .Y(_700_) );
OAI21X1 OAI21X1_135 ( .A(_700_), .B(_699_), .C(_696_), .Y(_400__0_) );
NAND2X1 NAND2X1_846 ( .A(PC_PC_STACK_2__1_), .B(_617__bF_buf0), .Y(_701_) );
OR2X2 OR2X2_990 ( .A(_601__bF_buf3), .B(_627_), .Y(_702_) );
NAND2X1 NAND2X1_847 ( .A(PC_PC_STACK_2__1_), .B(_601__bF_buf3), .Y(_703_) );
OAI21X1 OAI21X1_136 ( .A(_504_), .B(_601__bF_buf3), .C(_703_), .Y(_704_) );
OAI21X1 OAI21X1_137 ( .A(CORE_PC_ctrl_0_), .B(_703_), .C(_466__bF_buf2), .Y(_705_) );
NAND2X1 NAND2X1_848 ( .A(_704_), .B(_705_), .Y(_706_) );
AND2X2 AND2X2_1255 ( .A(_706_), .B(_702_), .Y(_707_) );
OAI21X1 OAI21X1_138 ( .A(rst_bF_buf1), .B(_707_), .C(_701_), .Y(_400__1_) );
NAND2X1 NAND2X1_849 ( .A(PC_PC_STACK_2__2_), .B(_617__bF_buf1), .Y(_708_) );
NOR3X1 NOR3X1_31 ( .A(_519_), .B(_455_), .C(_601__bF_buf3), .Y(_709_) );
AND2X2 AND2X2_1256 ( .A(_601__bF_buf3), .B(PC_PC_STACK_2__2_), .Y(_710_) );
AOI21X1 AOI21X1_62 ( .A(PC_ULA_OUT_2_), .B(_484__bF_buf3), .C(_710_), .Y(_711_) );
AOI22X1 AOI22X1_33 ( .A(_484__bF_buf3), .B(_638_), .C(_710_), .D(_406_), .Y(_712_) );
OAI21X1 OAI21X1_139 ( .A(_466__bF_buf1), .B(_711_), .C(_712_), .Y(_713_) );
OAI21X1 OAI21X1_140 ( .A(_713_), .B(_709_), .C(_409__bF_buf1), .Y(_714_) );
NAND2X1 NAND2X1_850 ( .A(_708_), .B(_714_), .Y(_400__2_) );
INVX1 INVX1_297 ( .A(PC_PC_STACK_2__3_), .Y(_715_) );
NOR2X1 NOR2X1_148 ( .A(_643_), .B(_715_), .Y(_716_) );
NAND2X1 NAND2X1_851 ( .A(_715_), .B(_601__bF_buf1), .Y(_717_) );
OR2X2 OR2X2_991 ( .A(_601__bF_buf1), .B(_539_), .Y(_718_) );
NAND3X1 NAND3X1_96 ( .A(_718_), .B(_456__bF_buf1), .C(_717_), .Y(_719_) );
NAND2X1 NAND2X1_852 ( .A(PC_PC_STACK_2__3_), .B(_601__bF_buf1), .Y(_720_) );
OAI21X1 OAI21X1_141 ( .A(_545_), .B(_601__bF_buf1), .C(_720_), .Y(_721_) );
NAND2X1 NAND2X1_853 ( .A(_505__bF_buf0), .B(_721_), .Y(_722_) );
OAI21X1 OAI21X1_142 ( .A(_543_), .B(_601__bF_buf1), .C(_720_), .Y(_723_) );
NAND2X1 NAND2X1_854 ( .A(_523_), .B(_723_), .Y(_724_) );
NAND3X1 NAND3X1_97 ( .A(_719_), .B(_722_), .C(_724_), .Y(_725_) );
AND2X2 AND2X2_1257 ( .A(_725_), .B(_409__bF_buf0), .Y(_726_) );
OR2X2 OR2X2_992 ( .A(_716_), .B(_726_), .Y(_400__3_) );
AND2X2 AND2X2_1258 ( .A(_617__bF_buf2), .B(PC_PC_STACK_2__4_), .Y(_727_) );
NAND2X1 NAND2X1_855 ( .A(PC_PC_STACK_2__4_), .B(_601__bF_buf2), .Y(_728_) );
OAI21X1 OAI21X1_143 ( .A(_601__bF_buf0), .B(_556_), .C(_728_), .Y(_729_) );
AND2X2 AND2X2_1259 ( .A(_729_), .B(_456__bF_buf2), .Y(_730_) );
OAI21X1 OAI21X1_144 ( .A(_560_), .B(_601__bF_buf2), .C(_728_), .Y(_731_) );
NAND2X1 NAND2X1_856 ( .A(_505__bF_buf1), .B(_731_), .Y(_732_) );
MUX2X1 MUX2X1_818 ( .A(PC_ULA_OUT_4_), .B(PC_PC_STACK_2__4_), .S(_484__bF_buf1), .Y(_733_) );
OAI21X1 OAI21X1_145 ( .A(_466__bF_buf3), .B(_733_), .C(_732_), .Y(_734_) );
OR2X2 OR2X2_993 ( .A(_730_), .B(_734_), .Y(_735_) );
AND2X2 AND2X2_1260 ( .A(_735_), .B(_409__bF_buf2), .Y(_736_) );
OR2X2 OR2X2_994 ( .A(_727_), .B(_736_), .Y(_400__4_) );
AND2X2 AND2X2_1261 ( .A(_617__bF_buf3), .B(PC_PC_STACK_2__5_), .Y(_737_) );
XNOR2X1 XNOR2X1_62 ( .A(_569_), .B(_566_), .Y(_738_) );
NAND2X1 NAND2X1_857 ( .A(PC_PC_STACK_2__5_), .B(_601__bF_buf2), .Y(_739_) );
OAI21X1 OAI21X1_146 ( .A(_601__bF_buf2), .B(_738_), .C(_739_), .Y(_740_) );
AND2X2 AND2X2_1262 ( .A(_740_), .B(_456__bF_buf1), .Y(_741_) );
OAI21X1 OAI21X1_147 ( .A(_577_), .B(_601__bF_buf2), .C(_739_), .Y(_742_) );
NAND2X1 NAND2X1_858 ( .A(_505__bF_buf2), .B(_742_), .Y(_743_) );
MUX2X1 MUX2X1_819 ( .A(PC_ULA_OUT_5_), .B(PC_PC_STACK_2__5_), .S(_484__bF_buf2), .Y(_744_) );
OAI21X1 OAI21X1_148 ( .A(_466__bF_buf0), .B(_744_), .C(_743_), .Y(_745_) );
OR2X2 OR2X2_995 ( .A(_741_), .B(_745_), .Y(_746_) );
AND2X2 AND2X2_1263 ( .A(_746_), .B(_409__bF_buf5), .Y(_747_) );
OR2X2 OR2X2_996 ( .A(_737_), .B(_747_), .Y(_400__5_) );
AND2X2 AND2X2_1264 ( .A(_617__bF_buf2), .B(PC_PC_STACK_2__6_), .Y(_748_) );
NAND2X1 NAND2X1_859 ( .A(PC_PC_STACK_2__6_), .B(_601__bF_buf0), .Y(_749_) );
OAI21X1 OAI21X1_149 ( .A(_601__bF_buf0), .B(_587_), .C(_749_), .Y(_750_) );
AND2X2 AND2X2_1265 ( .A(_750_), .B(_456__bF_buf0), .Y(_751_) );
OAI21X1 OAI21X1_150 ( .A(_678_), .B(_601__bF_buf0), .C(_749_), .Y(_752_) );
NAND2X1 NAND2X1_860 ( .A(_505__bF_buf1), .B(_752_), .Y(_753_) );
MUX2X1 MUX2X1_820 ( .A(PC_ULA_OUT_6_), .B(PC_PC_STACK_2__6_), .S(_484__bF_buf0), .Y(_754_) );
OAI21X1 OAI21X1_151 ( .A(_466__bF_buf3), .B(_754_), .C(_753_), .Y(_755_) );
OR2X2 OR2X2_997 ( .A(_755_), .B(_751_), .Y(_756_) );
AND2X2 AND2X2_1266 ( .A(_756_), .B(_409__bF_buf3), .Y(_757_) );
OR2X2 OR2X2_998 ( .A(_748_), .B(_757_), .Y(_400__6_) );
INVX1 INVX1_298 ( .A(PC_PC_STACK_2__7_), .Y(_758_) );
NOR2X1 NOR2X1_149 ( .A(_643_), .B(_758_), .Y(_759_) );
NOR2X1 NOR2X1_150 ( .A(_484__bF_buf1), .B(_758_), .Y(_760_) );
AND2X2 AND2X2_1267 ( .A(_606_), .B(_484__bF_buf1), .Y(_761_) );
OR2X2 OR2X2_999 ( .A(_760_), .B(_761_), .Y(_762_) );
AND2X2 AND2X2_1268 ( .A(_762_), .B(_456__bF_buf2), .Y(_763_) );
NOR2X1 NOR2X1_151 ( .A(_601__bF_buf0), .B(_612_), .Y(_764_) );
OAI21X1 OAI21X1_152 ( .A(_760_), .B(_764_), .C(_523_), .Y(_765_) );
AOI21X1 AOI21X1_63 ( .A(INTERRUPT_ch[7]), .B(_484__bF_buf1), .C(_760_), .Y(_766_) );
OAI21X1 OAI21X1_153 ( .A(_463_), .B(_766_), .C(_765_), .Y(_767_) );
OR2X2 OR2X2_1000 ( .A(_767_), .B(_763_), .Y(_768_) );
AND2X2 AND2X2_1269 ( .A(_768_), .B(_409__bF_buf2), .Y(_769_) );
OR2X2 OR2X2_1001 ( .A(_759_), .B(_769_), .Y(_400__7_) );
NAND2X1 NAND2X1_861 ( .A(PC_PC_STACK_1__0_), .B(_617__bF_buf1), .Y(_770_) );
NOR2X1 NOR2X1_152 ( .A(_474_), .B(_455_), .Y(_771_) );
NAND2X1 NAND2X1_862 ( .A(_473__bF_buf0), .B(_621_), .Y(_772_) );
AOI21X1 AOI21X1_64 ( .A(_502_), .B(_772_), .C(_771_), .Y(_773_) );
OAI21X1 OAI21X1_154 ( .A(PC_PC_STACK_1__0_), .B(_473__bF_buf0), .C(_409__bF_buf5), .Y(_774_) );
OAI21X1 OAI21X1_155 ( .A(_774_), .B(_773_), .C(_770_), .Y(_399__0_) );
NAND2X1 NAND2X1_863 ( .A(PC_PC_STACK_1__1_), .B(_617__bF_buf0), .Y(_775_) );
INVX1 INVX1_299 ( .A(_473__bF_buf2), .Y(_776_) );
OR2X2 OR2X2_1002 ( .A(_776__bF_buf2), .B(_627_), .Y(_777_) );
NAND2X1 NAND2X1_864 ( .A(PC_PC_STACK_1__1_), .B(_776__bF_buf2), .Y(_778_) );
OAI21X1 OAI21X1_156 ( .A(_504_), .B(_776__bF_buf2), .C(_778_), .Y(_779_) );
OAI21X1 OAI21X1_157 ( .A(CORE_PC_ctrl_0_), .B(_778_), .C(_466__bF_buf1), .Y(_780_) );
NAND2X1 NAND2X1_865 ( .A(_779_), .B(_780_), .Y(_781_) );
AND2X2 AND2X2_1270 ( .A(_781_), .B(_777_), .Y(_782_) );
OAI21X1 OAI21X1_158 ( .A(rst_bF_buf0), .B(_782_), .C(_775_), .Y(_399__1_) );
NAND2X1 NAND2X1_866 ( .A(PC_PC_STACK_1__2_), .B(_617__bF_buf1), .Y(_783_) );
NOR3X1 NOR3X1_32 ( .A(_519_), .B(_455_), .C(_776__bF_buf2), .Y(_784_) );
AND2X2 AND2X2_1271 ( .A(_776__bF_buf2), .B(PC_PC_STACK_1__2_), .Y(_785_) );
AOI21X1 AOI21X1_65 ( .A(PC_ULA_OUT_2_), .B(_473__bF_buf2), .C(_785_), .Y(_786_) );
AOI22X1 AOI22X1_34 ( .A(_473__bF_buf2), .B(_638_), .C(_785_), .D(_406_), .Y(_787_) );
OAI21X1 OAI21X1_159 ( .A(_466__bF_buf1), .B(_786_), .C(_787_), .Y(_788_) );
OAI21X1 OAI21X1_160 ( .A(_788_), .B(_784_), .C(_409__bF_buf4), .Y(_789_) );
NAND2X1 NAND2X1_867 ( .A(_783_), .B(_789_), .Y(_399__2_) );
INVX1 INVX1_300 ( .A(PC_PC_STACK_1__3_), .Y(_790_) );
NOR2X1 NOR2X1_153 ( .A(_643_), .B(_790_), .Y(_791_) );
NAND2X1 NAND2X1_868 ( .A(_790_), .B(_776__bF_buf0), .Y(_792_) );
OR2X2 OR2X2_1003 ( .A(_776__bF_buf0), .B(_539_), .Y(_793_) );
NAND3X1 NAND3X1_98 ( .A(_793_), .B(_456__bF_buf1), .C(_792_), .Y(_794_) );
NAND2X1 NAND2X1_869 ( .A(PC_PC_STACK_1__3_), .B(_776__bF_buf0), .Y(_795_) );
OAI21X1 OAI21X1_161 ( .A(_545_), .B(_776__bF_buf0), .C(_795_), .Y(_796_) );
NAND2X1 NAND2X1_870 ( .A(_505__bF_buf0), .B(_796_), .Y(_797_) );
OAI21X1 OAI21X1_162 ( .A(_543_), .B(_776__bF_buf0), .C(_795_), .Y(_798_) );
NAND2X1 NAND2X1_871 ( .A(_523_), .B(_798_), .Y(_799_) );
NAND3X1 NAND3X1_99 ( .A(_794_), .B(_797_), .C(_799_), .Y(_800_) );
AND2X2 AND2X2_1272 ( .A(_800_), .B(_409__bF_buf0), .Y(_801_) );
OR2X2 OR2X2_1004 ( .A(_791_), .B(_801_), .Y(_399__3_) );
AND2X2 AND2X2_1273 ( .A(_617__bF_buf2), .B(PC_PC_STACK_1__4_), .Y(_802_) );
NAND2X1 NAND2X1_872 ( .A(PC_PC_STACK_1__4_), .B(_776__bF_buf1), .Y(_803_) );
OAI21X1 OAI21X1_163 ( .A(_776__bF_buf3), .B(_556_), .C(_803_), .Y(_804_) );
AND2X2 AND2X2_1274 ( .A(_804_), .B(_456__bF_buf0), .Y(_805_) );
OAI21X1 OAI21X1_164 ( .A(_560_), .B(_776__bF_buf1), .C(_803_), .Y(_806_) );
NAND2X1 NAND2X1_873 ( .A(_505__bF_buf1), .B(_806_), .Y(_807_) );
MUX2X1 MUX2X1_821 ( .A(PC_ULA_OUT_4_), .B(PC_PC_STACK_1__4_), .S(_473__bF_buf1), .Y(_808_) );
OAI21X1 OAI21X1_165 ( .A(_466__bF_buf3), .B(_808_), .C(_807_), .Y(_809_) );
OR2X2 OR2X2_1005 ( .A(_805_), .B(_809_), .Y(_810_) );
AND2X2 AND2X2_1275 ( .A(_810_), .B(_409__bF_buf0), .Y(_811_) );
OR2X2 OR2X2_1006 ( .A(_802_), .B(_811_), .Y(_399__4_) );
AND2X2 AND2X2_1276 ( .A(_617__bF_buf3), .B(PC_PC_STACK_1__5_), .Y(_812_) );
NAND2X1 NAND2X1_874 ( .A(PC_PC_STACK_1__5_), .B(_776__bF_buf3), .Y(_813_) );
OAI21X1 OAI21X1_166 ( .A(_776__bF_buf3), .B(_738_), .C(_813_), .Y(_814_) );
AND2X2 AND2X2_1277 ( .A(_814_), .B(_456__bF_buf1), .Y(_815_) );
OAI21X1 OAI21X1_167 ( .A(_577_), .B(_776__bF_buf3), .C(_813_), .Y(_816_) );
NAND2X1 NAND2X1_875 ( .A(_505__bF_buf2), .B(_816_), .Y(_817_) );
MUX2X1 MUX2X1_822 ( .A(PC_ULA_OUT_5_), .B(PC_PC_STACK_1__5_), .S(_473__bF_buf0), .Y(_818_) );
OAI21X1 OAI21X1_168 ( .A(_466__bF_buf0), .B(_818_), .C(_817_), .Y(_819_) );
OR2X2 OR2X2_1007 ( .A(_815_), .B(_819_), .Y(_820_) );
AND2X2 AND2X2_1278 ( .A(_820_), .B(_409__bF_buf5), .Y(_821_) );
OR2X2 OR2X2_1008 ( .A(_812_), .B(_821_), .Y(_399__5_) );
AND2X2 AND2X2_1279 ( .A(_617__bF_buf2), .B(PC_PC_STACK_1__6_), .Y(_822_) );
NAND2X1 NAND2X1_876 ( .A(PC_PC_STACK_1__6_), .B(_776__bF_buf1), .Y(_823_) );
OAI21X1 OAI21X1_169 ( .A(_776__bF_buf1), .B(_587_), .C(_823_), .Y(_824_) );
AND2X2 AND2X2_1280 ( .A(_824_), .B(_456__bF_buf0), .Y(_825_) );
OAI21X1 OAI21X1_170 ( .A(_678_), .B(_776__bF_buf1), .C(_823_), .Y(_826_) );
NAND2X1 NAND2X1_877 ( .A(_505__bF_buf1), .B(_826_), .Y(_827_) );
MUX2X1 MUX2X1_823 ( .A(PC_ULA_OUT_6_), .B(PC_PC_STACK_1__6_), .S(_473__bF_buf3), .Y(_828_) );
OAI21X1 OAI21X1_171 ( .A(_466__bF_buf3), .B(_828_), .C(_827_), .Y(_829_) );
OR2X2 OR2X2_1009 ( .A(_829_), .B(_825_), .Y(_830_) );
AND2X2 AND2X2_1281 ( .A(_830_), .B(_409__bF_buf3), .Y(_831_) );
OR2X2 OR2X2_1010 ( .A(_822_), .B(_831_), .Y(_399__6_) );
INVX1 INVX1_301 ( .A(PC_PC_STACK_1__7_), .Y(_832_) );
NOR2X1 NOR2X1_154 ( .A(_643_), .B(_832_), .Y(_833_) );
NOR2X1 NOR2X1_155 ( .A(_473__bF_buf3), .B(_832_), .Y(_834_) );
AND2X2 AND2X2_1282 ( .A(_606_), .B(_473__bF_buf3), .Y(_835_) );
OR2X2 OR2X2_1011 ( .A(_834_), .B(_835_), .Y(_836_) );
AND2X2 AND2X2_1283 ( .A(_836_), .B(_456__bF_buf2), .Y(_837_) );
NOR2X1 NOR2X1_156 ( .A(_776__bF_buf3), .B(_612_), .Y(_838_) );
OAI21X1 OAI21X1_172 ( .A(_834_), .B(_838_), .C(_523_), .Y(_839_) );
AOI21X1 AOI21X1_66 ( .A(INTERRUPT_ch[7]), .B(_473__bF_buf3), .C(_834_), .Y(_840_) );
OAI21X1 OAI21X1_173 ( .A(_463_), .B(_840_), .C(_839_), .Y(_841_) );
OR2X2 OR2X2_1012 ( .A(_841_), .B(_837_), .Y(_842_) );
AND2X2 AND2X2_1284 ( .A(_842_), .B(_409__bF_buf2), .Y(_843_) );
OR2X2 OR2X2_1013 ( .A(_833_), .B(_843_), .Y(_399__7_) );
INVX1 INVX1_302 ( .A(IDATA_CORE_out[0]), .Y(_844_) );
INVX1 INVX1_303 ( .A(PC_delay_1_), .Y(_845_) );
NAND3X1 NAND3X1_100 ( .A(_408_), .B(_404_), .C(_845_), .Y(_846_) );
NOR2X1 NOR2X1_157 ( .A(_846_), .B(_844_), .Y(CORE_InstructionIN_0_) );
INVX1 INVX1_304 ( .A(IDATA_CORE_out[1]), .Y(_847_) );
NOR2X1 NOR2X1_158 ( .A(_846_), .B(_847_), .Y(CORE_InstructionIN_1_) );
INVX1 INVX1_305 ( .A(IDATA_CORE_out[2]), .Y(_848_) );
NOR2X1 NOR2X1_159 ( .A(_846_), .B(_848_), .Y(CORE_InstructionIN_2_) );
INVX1 INVX1_306 ( .A(IDATA_CORE_out[3]), .Y(_849_) );
NOR2X1 NOR2X1_160 ( .A(_846_), .B(_849_), .Y(CORE_InstructionIN_3_) );
INVX1 INVX1_307 ( .A(IDATA_CORE_out[4]), .Y(_850_) );
NOR2X1 NOR2X1_161 ( .A(_846_), .B(_850_), .Y(CORE_InstructionIN_4_) );
INVX1 INVX1_308 ( .A(IDATA_CORE_out[5]), .Y(_851_) );
NOR2X1 NOR2X1_162 ( .A(_846_), .B(_851_), .Y(CORE_InstructionIN_5_) );
INVX1 INVX1_309 ( .A(IDATA_CORE_out[6]), .Y(_852_) );
NOR2X1 NOR2X1_163 ( .A(_846_), .B(_852_), .Y(CORE_InstructionIN_6_) );
INVX1 INVX1_310 ( .A(IDATA_CORE_out[7]), .Y(_853_) );
NOR2X1 NOR2X1_164 ( .A(_846_), .B(_853_), .Y(CORE_InstructionIN_7_) );
INVX1 INVX1_311 ( .A(IDATA_CORE_out[8]), .Y(_854_) );
NOR2X1 NOR2X1_165 ( .A(_846_), .B(_854_), .Y(CORE_InstructionIN_8_) );
INVX1 INVX1_312 ( .A(IDATA_CORE_out[9]), .Y(_855_) );
NOR2X1 NOR2X1_166 ( .A(_846_), .B(_855_), .Y(CORE_InstructionIN_9_) );
INVX1 INVX1_313 ( .A(IDATA_CORE_out[10]), .Y(_856_) );
NOR2X1 NOR2X1_167 ( .A(_846_), .B(_856_), .Y(CORE_InstructionIN_10_) );
INVX1 INVX1_314 ( .A(IDATA_CORE_out[11]), .Y(_857_) );
NOR2X1 NOR2X1_168 ( .A(_846_), .B(_857_), .Y(CORE_InstructionIN_11_) );
INVX1 INVX1_315 ( .A(IDATA_CORE_out[12]), .Y(_858_) );
NOR2X1 NOR2X1_169 ( .A(_846_), .B(_858_), .Y(CORE_InstructionIN_12_) );
INVX1 INVX1_316 ( .A(IDATA_CORE_out[13]), .Y(_859_) );
NOR2X1 NOR2X1_170 ( .A(_846_), .B(_859_), .Y(CORE_InstructionIN_13_) );
INVX1 INVX1_317 ( .A(IDATA_CORE_out[14]), .Y(_860_) );
NOR2X1 NOR2X1_171 ( .A(_846_), .B(_860_), .Y(CORE_InstructionIN_14_) );
INVX1 INVX1_318 ( .A(IDATA_CORE_out[15]), .Y(_861_) );
NOR2X1 NOR2X1_172 ( .A(_846_), .B(_861_), .Y(CORE_InstructionIN_15_) );
NAND2X1 NAND2X1_878 ( .A(clk_bF_buf51), .B(_404_), .Y(_862_) );
NOR2X1 NOR2X1_173 ( .A(_407_), .B(_862_), .Y(_147_) );
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf51), .D(_403__0_), .Q(PC_delay_0_) );
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf51), .D(_403__1_), .Q(PC_delay_1_) );
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf48), .D(_402__0_), .Q(PC_PC_pointer_0_) );
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf21), .D(_402__1_), .Q(PC_PC_pointer_1_) );
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf8), .D(_396__0_), .Q(PC_ADDR_stack_0__0_) );
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf61), .D(_396__1_), .Q(PC_ADDR_stack_0__1_) );
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf61), .D(_396__2_), .Q(PC_ADDR_stack_0__2_) );
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf21), .D(_396__3_), .Q(PC_ADDR_stack_0__3_) );
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf57), .D(_396__4_), .Q(PC_ADDR_stack_0__4_) );
DFFPOSX1 DFFPOSX1_795 ( .CLK(clk_bF_buf61), .D(_396__5_), .Q(PC_ADDR_stack_0__5_) );
DFFPOSX1 DFFPOSX1_796 ( .CLK(clk_bF_buf36), .D(_396__6_), .Q(PC_ADDR_stack_0__6_) );
DFFPOSX1 DFFPOSX1_797 ( .CLK(clk_bF_buf36), .D(_396__7_), .Q(PC_ADDR_stack_0__7_) );
DFFPOSX1 DFFPOSX1_798 ( .CLK(clk_bF_buf61), .D(_397__0_), .Q(PC_ADDR_stack_1__0_) );
DFFPOSX1 DFFPOSX1_799 ( .CLK(clk_bF_buf60), .D(_397__1_), .Q(PC_ADDR_stack_1__1_) );
DFFPOSX1 DFFPOSX1_800 ( .CLK(clk_bF_buf61), .D(_397__2_), .Q(PC_ADDR_stack_1__2_) );
DFFPOSX1 DFFPOSX1_801 ( .CLK(clk_bF_buf61), .D(_397__3_), .Q(PC_ADDR_stack_1__3_) );
DFFPOSX1 DFFPOSX1_802 ( .CLK(clk_bF_buf57), .D(_397__4_), .Q(PC_ADDR_stack_1__4_) );
DFFPOSX1 DFFPOSX1_803 ( .CLK(clk_bF_buf60), .D(_397__5_), .Q(PC_ADDR_stack_1__5_) );
DFFPOSX1 DFFPOSX1_804 ( .CLK(clk_bF_buf36), .D(_397__6_), .Q(PC_ADDR_stack_1__6_) );
DFFPOSX1 DFFPOSX1_805 ( .CLK(clk_bF_buf57), .D(_397__7_), .Q(PC_ADDR_stack_1__7_) );
DFFPOSX1 DFFPOSX1_806 ( .CLK(clk_bF_buf21), .D(_398__0_), .Q(PC_PC_STACK_0__0_) );
DFFPOSX1 DFFPOSX1_807 ( .CLK(clk_bF_buf21), .D(_398__1_), .Q(PC_PC_STACK_0__1_) );
DFFPOSX1 DFFPOSX1_808 ( .CLK(clk_bF_buf21), .D(_398__2_), .Q(PC_PC_STACK_0__2_) );
DFFPOSX1 DFFPOSX1_809 ( .CLK(clk_bF_buf17), .D(_398__3_), .Q(PC_PC_STACK_0__3_) );
DFFPOSX1 DFFPOSX1_810 ( .CLK(clk_bF_buf21), .D(_398__4_), .Q(PC_PC_STACK_0__4_) );
DFFPOSX1 DFFPOSX1_811 ( .CLK(clk_bF_buf8), .D(_398__5_), .Q(PC_PC_STACK_0__5_) );
DFFPOSX1 DFFPOSX1_812 ( .CLK(clk_bF_buf17), .D(_398__6_), .Q(PC_PC_STACK_0__6_) );
DFFPOSX1 DFFPOSX1_813 ( .CLK(clk_bF_buf21), .D(_398__7_), .Q(PC_PC_STACK_0__7_) );
DFFPOSX1 DFFPOSX1_814 ( .CLK(clk_bF_buf8), .D(_399__0_), .Q(PC_PC_STACK_1__0_) );
DFFPOSX1 DFFPOSX1_815 ( .CLK(clk_bF_buf61), .D(_399__1_), .Q(PC_PC_STACK_1__1_) );
DFFPOSX1 DFFPOSX1_816 ( .CLK(clk_bF_buf8), .D(_399__2_), .Q(PC_PC_STACK_1__2_) );
DFFPOSX1 DFFPOSX1_817 ( .CLK(clk_bF_buf17), .D(_399__3_), .Q(PC_PC_STACK_1__3_) );
DFFPOSX1 DFFPOSX1_818 ( .CLK(clk_bF_buf17), .D(_399__4_), .Q(PC_PC_STACK_1__4_) );
DFFPOSX1 DFFPOSX1_819 ( .CLK(clk_bF_buf8), .D(_399__5_), .Q(PC_PC_STACK_1__5_) );
DFFPOSX1 DFFPOSX1_820 ( .CLK(clk_bF_buf36), .D(_399__6_), .Q(PC_PC_STACK_1__6_) );
DFFPOSX1 DFFPOSX1_821 ( .CLK(clk_bF_buf36), .D(_399__7_), .Q(PC_PC_STACK_1__7_) );
DFFPOSX1 DFFPOSX1_822 ( .CLK(clk_bF_buf8), .D(_400__0_), .Q(PC_PC_STACK_2__0_) );
DFFPOSX1 DFFPOSX1_823 ( .CLK(clk_bF_buf43), .D(_400__1_), .Q(PC_PC_STACK_2__1_) );
DFFPOSX1 DFFPOSX1_824 ( .CLK(clk_bF_buf8), .D(_400__2_), .Q(PC_PC_STACK_2__2_) );
DFFPOSX1 DFFPOSX1_825 ( .CLK(clk_bF_buf17), .D(_400__3_), .Q(PC_PC_STACK_2__3_) );
DFFPOSX1 DFFPOSX1_826 ( .CLK(clk_bF_buf36), .D(_400__4_), .Q(PC_PC_STACK_2__4_) );
DFFPOSX1 DFFPOSX1_827 ( .CLK(clk_bF_buf17), .D(_400__5_), .Q(PC_PC_STACK_2__5_) );
DFFPOSX1 DFFPOSX1_828 ( .CLK(clk_bF_buf36), .D(_400__6_), .Q(PC_PC_STACK_2__6_) );
DFFPOSX1 DFFPOSX1_829 ( .CLK(clk_bF_buf57), .D(_400__7_), .Q(PC_PC_STACK_2__7_) );
DFFPOSX1 DFFPOSX1_830 ( .CLK(clk_bF_buf8), .D(_401__0_), .Q(PC_PC_STACK_3__0_) );
DFFPOSX1 DFFPOSX1_831 ( .CLK(clk_bF_buf21), .D(_401__1_), .Q(PC_PC_STACK_3__1_) );
DFFPOSX1 DFFPOSX1_832 ( .CLK(clk_bF_buf8), .D(_401__2_), .Q(PC_PC_STACK_3__2_) );
DFFPOSX1 DFFPOSX1_833 ( .CLK(clk_bF_buf17), .D(_401__3_), .Q(PC_PC_STACK_3__3_) );
DFFPOSX1 DFFPOSX1_834 ( .CLK(clk_bF_buf17), .D(_401__4_), .Q(PC_PC_STACK_3__4_) );
DFFPOSX1 DFFPOSX1_835 ( .CLK(clk_bF_buf17), .D(_401__5_), .Q(PC_PC_STACK_3__5_) );
DFFPOSX1 DFFPOSX1_836 ( .CLK(clk_bF_buf36), .D(_401__6_), .Q(PC_PC_STACK_3__6_) );
DFFPOSX1 DFFPOSX1_837 ( .CLK(clk_bF_buf21), .D(_401__7_), .Q(PC_PC_STACK_3__7_) );
INVX2 INVX2_7 ( .A(REG_RD_wb_pipe_0_), .Y(_1567_) );
INVX8 INVX8_1 ( .A(INTERRUPT_flag_bF_buf8_bF_buf2), .Y(_1568_) );
NAND3X1 NAND3X1_101 ( .A(_1568__bF_buf15_bF_buf1), .B(REG_RFD_exec_pipe_3_), .C(REG_Write_wb_pipe), .Y(_1569_) );
INVX1 INVX1_319 ( .A(REG_RFD_exec_pipe_0_), .Y(_1570_) );
NAND3X1 NAND3X1_102 ( .A(_1570_), .B(REG_RFD_exec_pipe_1_), .C(REG_RFD_exec_pipe_2_), .Y(_1571_) );
NOR2X1 NOR2X1_174 ( .A(_1569_), .B(_1571_), .Y(_1572_) );
INVX8 INVX8_2 ( .A(rst_bF_buf4), .Y(_1573_) );
NAND2X1 NAND2X1_879 ( .A(REGs_USR_REGS_6__0_), .B(_1573__bF_buf39), .Y(_1574_) );
MUX2X1 MUX2X1_824 ( .A(_1567__bF_buf0), .B(_1574_), .S(_1572__bF_buf0), .Y(_863_) );
INVX2 INVX2_8 ( .A(REG_RD_wb_pipe_1_), .Y(_1575_) );
NAND2X1 NAND2X1_880 ( .A(REGs_USR_REGS_6__1_), .B(_1573__bF_buf53), .Y(_1576_) );
MUX2X1 MUX2X1_825 ( .A(_1575__bF_buf0), .B(_1576_), .S(_1572__bF_buf0), .Y(_864_) );
INVX2 INVX2_9 ( .A(REG_RD_wb_pipe_2_), .Y(_1577_) );
NAND2X1 NAND2X1_881 ( .A(REGs_USR_REGS_6__2_), .B(_1573__bF_buf61), .Y(_1578_) );
MUX2X1 MUX2X1_826 ( .A(_1577__bF_buf2), .B(_1578_), .S(_1572__bF_buf4), .Y(_865_) );
INVX2 INVX2_10 ( .A(REG_RD_wb_pipe_3_), .Y(_1579_) );
NAND2X1 NAND2X1_882 ( .A(REGs_USR_REGS_6__3_), .B(_1573__bF_buf56), .Y(_1580_) );
MUX2X1 MUX2X1_827 ( .A(_1579__bF_buf3), .B(_1580_), .S(_1572__bF_buf4), .Y(_866_) );
INVX2 INVX2_11 ( .A(REG_RD_wb_pipe_4_), .Y(_1581_) );
NAND2X1 NAND2X1_883 ( .A(REGs_USR_REGS_6__4_), .B(_1573__bF_buf27), .Y(_1582_) );
MUX2X1 MUX2X1_828 ( .A(_1581__bF_buf2), .B(_1582_), .S(_1572__bF_buf4), .Y(_867_) );
INVX2 INVX2_12 ( .A(REG_RD_wb_pipe_5_), .Y(_1583_) );
NAND2X1 NAND2X1_884 ( .A(REGs_USR_REGS_6__5_), .B(_1573__bF_buf78), .Y(_1584_) );
MUX2X1 MUX2X1_829 ( .A(_1583__bF_buf1), .B(_1584_), .S(_1572__bF_buf2), .Y(_868_) );
INVX2 INVX2_13 ( .A(REG_RD_wb_pipe_6_), .Y(_1585_) );
NAND2X1 NAND2X1_885 ( .A(REGs_USR_REGS_6__6_), .B(_1573__bF_buf57), .Y(_1586_) );
MUX2X1 MUX2X1_830 ( .A(_1585__bF_buf2), .B(_1586_), .S(_1572__bF_buf3), .Y(_869_) );
INVX2 INVX2_14 ( .A(REG_RD_wb_pipe_7_), .Y(_1587_) );
NAND2X1 NAND2X1_886 ( .A(REGs_USR_REGS_6__7_), .B(_1573__bF_buf48), .Y(_1588_) );
MUX2X1 MUX2X1_831 ( .A(_1587__bF_buf2), .B(_1588_), .S(_1572__bF_buf4), .Y(_870_) );
INVX2 INVX2_15 ( .A(REG_RD_wb_pipe_8_), .Y(_1589_) );
NAND2X1 NAND2X1_887 ( .A(REGs_USR_REGS_6__8_), .B(_1573__bF_buf31), .Y(_1590_) );
MUX2X1 MUX2X1_832 ( .A(_1589__bF_buf0), .B(_1590_), .S(_1572__bF_buf0), .Y(_871_) );
INVX2 INVX2_16 ( .A(REG_RD_wb_pipe_9_), .Y(_1591_) );
NAND2X1 NAND2X1_888 ( .A(REGs_USR_REGS_6__9_), .B(_1573__bF_buf78), .Y(_1592_) );
MUX2X1 MUX2X1_833 ( .A(_1591__bF_buf1), .B(_1592_), .S(_1572__bF_buf2), .Y(_872_) );
INVX2 INVX2_17 ( .A(REG_RD_wb_pipe_10_), .Y(_1593_) );
NAND2X1 NAND2X1_889 ( .A(REGs_USR_REGS_6__10_), .B(_1573__bF_buf21), .Y(_1594_) );
MUX2X1 MUX2X1_834 ( .A(_1593__bF_buf3), .B(_1594_), .S(_1572__bF_buf1), .Y(_873_) );
INVX2 INVX2_18 ( .A(REG_RD_wb_pipe_11_), .Y(_1595_) );
NAND2X1 NAND2X1_890 ( .A(REGs_USR_REGS_6__11_), .B(_1573__bF_buf78), .Y(_1596_) );
MUX2X1 MUX2X1_835 ( .A(_1595__bF_buf3), .B(_1596_), .S(_1572__bF_buf2), .Y(_874_) );
INVX2 INVX2_19 ( .A(REG_RD_wb_pipe_12_), .Y(_1597_) );
NAND2X1 NAND2X1_891 ( .A(REGs_USR_REGS_6__12_), .B(_1573__bF_buf57), .Y(_1598_) );
MUX2X1 MUX2X1_836 ( .A(_1597__bF_buf3), .B(_1598_), .S(_1572__bF_buf3), .Y(_875_) );
INVX2 INVX2_20 ( .A(REG_RD_wb_pipe_13_), .Y(_1599_) );
NAND2X1 NAND2X1_892 ( .A(REGs_USR_REGS_6__13_), .B(_1573__bF_buf6), .Y(_1600_) );
MUX2X1 MUX2X1_837 ( .A(_1599__bF_buf0), .B(_1600_), .S(_1572__bF_buf3), .Y(_876_) );
INVX2 INVX2_21 ( .A(REG_RD_wb_pipe_14_), .Y(_1601_) );
NAND2X1 NAND2X1_893 ( .A(REGs_USR_REGS_6__14_), .B(_1573__bF_buf9), .Y(_1602_) );
MUX2X1 MUX2X1_838 ( .A(_1601__bF_buf3), .B(_1602_), .S(_1572__bF_buf1), .Y(_877_) );
INVX2 INVX2_22 ( .A(REG_RD_wb_pipe_15_), .Y(_1603_) );
NAND2X1 NAND2X1_894 ( .A(REGs_USR_REGS_6__15_), .B(_1573__bF_buf78), .Y(_1604_) );
MUX2X1 MUX2X1_839 ( .A(_1603__bF_buf3), .B(_1604_), .S(_1572__bF_buf2), .Y(_878_) );
INVX2 INVX2_23 ( .A(REG_RD_wb_pipe_16_), .Y(_1605_) );
NAND2X1 NAND2X1_895 ( .A(REGs_USR_REGS_6__16_), .B(_1573__bF_buf45), .Y(_1606_) );
MUX2X1 MUX2X1_840 ( .A(_1605__bF_buf0), .B(_1606_), .S(_1572__bF_buf1), .Y(_879_) );
INVX2 INVX2_24 ( .A(REG_RD_wb_pipe_17_), .Y(_1607_) );
NAND2X1 NAND2X1_896 ( .A(REGs_USR_REGS_6__17_), .B(_1573__bF_buf6), .Y(_1608_) );
MUX2X1 MUX2X1_841 ( .A(_1607__bF_buf1), .B(_1608_), .S(_1572__bF_buf3), .Y(_880_) );
INVX2 INVX2_25 ( .A(REG_RD_wb_pipe_18_), .Y(_1609_) );
NAND2X1 NAND2X1_897 ( .A(REGs_USR_REGS_6__18_), .B(_1573__bF_buf70), .Y(_1610_) );
MUX2X1 MUX2X1_842 ( .A(_1609__bF_buf3), .B(_1610_), .S(_1572__bF_buf2), .Y(_881_) );
INVX2 INVX2_26 ( .A(REG_RD_wb_pipe_19_), .Y(_1611_) );
NAND2X1 NAND2X1_898 ( .A(REGs_USR_REGS_6__19_), .B(_1573__bF_buf16), .Y(_1612_) );
MUX2X1 MUX2X1_843 ( .A(_1611__bF_buf1), .B(_1612_), .S(_1572__bF_buf0), .Y(_882_) );
INVX2 INVX2_27 ( .A(REG_RD_wb_pipe_20_), .Y(_1613_) );
NAND2X1 NAND2X1_899 ( .A(REGs_USR_REGS_6__20_), .B(_1573__bF_buf7), .Y(_1614_) );
MUX2X1 MUX2X1_844 ( .A(_1613__bF_buf0), .B(_1614_), .S(_1572__bF_buf3), .Y(_883_) );
INVX2 INVX2_28 ( .A(REG_RD_wb_pipe_21_), .Y(_1615_) );
NAND2X1 NAND2X1_900 ( .A(REGs_USR_REGS_6__21_), .B(_1573__bF_buf21), .Y(_1616_) );
MUX2X1 MUX2X1_845 ( .A(_1615__bF_buf0), .B(_1616_), .S(_1572__bF_buf1), .Y(_884_) );
INVX2 INVX2_29 ( .A(REG_RD_wb_pipe_22_), .Y(_1617_) );
NAND2X1 NAND2X1_901 ( .A(REGs_USR_REGS_6__22_), .B(_1573__bF_buf27), .Y(_1618_) );
MUX2X1 MUX2X1_846 ( .A(_1617__bF_buf3), .B(_1618_), .S(_1572__bF_buf4), .Y(_885_) );
INVX2 INVX2_30 ( .A(REG_RD_wb_pipe_23_), .Y(_1619_) );
NAND2X1 NAND2X1_902 ( .A(REGs_USR_REGS_6__23_), .B(_1573__bF_buf21), .Y(_1620_) );
MUX2X1 MUX2X1_847 ( .A(_1619__bF_buf2), .B(_1620_), .S(_1572__bF_buf1), .Y(_886_) );
INVX2 INVX2_31 ( .A(REG_RD_wb_pipe_24_), .Y(_1621_) );
NAND2X1 NAND2X1_903 ( .A(REGs_USR_REGS_6__24_), .B(_1573__bF_buf30), .Y(_1622_) );
MUX2X1 MUX2X1_848 ( .A(_1621__bF_buf3), .B(_1622_), .S(_1572__bF_buf0), .Y(_887_) );
INVX2 INVX2_32 ( .A(REG_RD_wb_pipe_25_), .Y(_1623_) );
NAND2X1 NAND2X1_904 ( .A(REGs_USR_REGS_6__25_), .B(_1573__bF_buf6), .Y(_1624_) );
MUX2X1 MUX2X1_849 ( .A(_1623__bF_buf0), .B(_1624_), .S(_1572__bF_buf3), .Y(_888_) );
INVX2 INVX2_33 ( .A(REG_RD_wb_pipe_26_), .Y(_1625_) );
NAND2X1 NAND2X1_905 ( .A(REGs_USR_REGS_6__26_), .B(_1573__bF_buf55), .Y(_1626_) );
MUX2X1 MUX2X1_850 ( .A(_1625__bF_buf2), .B(_1626_), .S(_1572__bF_buf4), .Y(_889_) );
INVX2 INVX2_34 ( .A(REG_RD_wb_pipe_27_), .Y(_1627_) );
NAND2X1 NAND2X1_906 ( .A(REGs_USR_REGS_6__27_), .B(_1573__bF_buf55), .Y(_1628_) );
MUX2X1 MUX2X1_851 ( .A(_1627__bF_buf2), .B(_1628_), .S(_1572__bF_buf4), .Y(_890_) );
INVX2 INVX2_35 ( .A(REG_RD_wb_pipe_28_), .Y(_1629_) );
NAND2X1 NAND2X1_907 ( .A(REGs_USR_REGS_6__28_), .B(_1573__bF_buf21), .Y(_1630_) );
MUX2X1 MUX2X1_852 ( .A(_1629__bF_buf0), .B(_1630_), .S(_1572__bF_buf1), .Y(_891_) );
INVX2 INVX2_36 ( .A(REG_RD_wb_pipe_29_), .Y(_1631_) );
NAND2X1 NAND2X1_908 ( .A(REGs_USR_REGS_6__29_), .B(_1573__bF_buf18), .Y(_1632_) );
MUX2X1 MUX2X1_853 ( .A(_1631__bF_buf0), .B(_1632_), .S(_1572__bF_buf0), .Y(_892_) );
INVX2 INVX2_37 ( .A(REG_RD_wb_pipe_30_), .Y(_1633_) );
NAND2X1 NAND2X1_909 ( .A(REGs_USR_REGS_6__30_), .B(_1573__bF_buf55), .Y(_1634_) );
MUX2X1 MUX2X1_854 ( .A(_1633__bF_buf0), .B(_1634_), .S(_1572__bF_buf3), .Y(_893_) );
INVX2 INVX2_38 ( .A(REG_RD_wb_pipe_31_), .Y(_1635_) );
NAND2X1 NAND2X1_910 ( .A(REGs_USR_REGS_6__31_), .B(_1573__bF_buf70), .Y(_1636_) );
MUX2X1 MUX2X1_855 ( .A(_1635__bF_buf2), .B(_1636_), .S(_1572__bF_buf2), .Y(_894_) );
INVX1 INVX1_320 ( .A(REG_RFD_exec_pipe_3_), .Y(_1637_) );
INVX1 INVX1_321 ( .A(REG_Write_wb_pipe), .Y(_1638_) );
NOR3X1 NOR3X1_33 ( .A(_1637_), .B(INTERRUPT_flag_bF_buf7_bF_buf1), .C(_1638_), .Y(_1639_) );
OR2X2 OR2X2_1014 ( .A(REG_RFD_exec_pipe_1_), .B(REG_RFD_exec_pipe_2_), .Y(_1640_) );
INVX1 INVX1_322 ( .A(_1640_), .Y(_1641_) );
NAND3X1 NAND3X1_103 ( .A(_1639_), .B(_1570_), .C(_1641_), .Y(_1642_) );
NAND2X1 NAND2X1_911 ( .A(REGs_USR_REGS_0__0_), .B(_1573__bF_buf6), .Y(_1643_) );
MUX2X1 MUX2X1_856 ( .A(_1643_), .B(_1567__bF_buf2), .S(_1642__bF_buf3), .Y(_895_) );
NAND2X1 NAND2X1_912 ( .A(REGs_USR_REGS_0__1_), .B(_1573__bF_buf24), .Y(_1644_) );
MUX2X1 MUX2X1_857 ( .A(_1644_), .B(_1575__bF_buf2), .S(_1642__bF_buf0), .Y(_896_) );
NAND2X1 NAND2X1_913 ( .A(REGs_USR_REGS_0__2_), .B(_1573__bF_buf7), .Y(_1645_) );
MUX2X1 MUX2X1_858 ( .A(_1645_), .B(_1577__bF_buf3), .S(_1642__bF_buf3), .Y(_897_) );
NAND2X1 NAND2X1_914 ( .A(REGs_USR_REGS_0__3_), .B(_1573__bF_buf56), .Y(_1646_) );
MUX2X1 MUX2X1_859 ( .A(_1646_), .B(_1579__bF_buf3), .S(_1642__bF_buf4), .Y(_898_) );
NAND2X1 NAND2X1_915 ( .A(REGs_USR_REGS_0__4_), .B(_1573__bF_buf3), .Y(_1647_) );
MUX2X1 MUX2X1_860 ( .A(_1647_), .B(_1581__bF_buf1), .S(_1642__bF_buf4), .Y(_899_) );
NAND2X1 NAND2X1_916 ( .A(REGs_USR_REGS_0__5_), .B(_1573__bF_buf25), .Y(_1648_) );
MUX2X1 MUX2X1_861 ( .A(_1648_), .B(_1583__bF_buf0), .S(_1642__bF_buf0), .Y(_900_) );
NAND2X1 NAND2X1_917 ( .A(REGs_USR_REGS_0__6_), .B(_1573__bF_buf3), .Y(_1649_) );
MUX2X1 MUX2X1_862 ( .A(_1649_), .B(_1585__bF_buf0), .S(_1642__bF_buf4), .Y(_901_) );
NAND2X1 NAND2X1_918 ( .A(REGs_USR_REGS_0__7_), .B(_1573__bF_buf17), .Y(_1650_) );
MUX2X1 MUX2X1_863 ( .A(_1650_), .B(_1587__bF_buf1), .S(_1642__bF_buf3), .Y(_902_) );
NAND2X1 NAND2X1_919 ( .A(REGs_USR_REGS_0__8_), .B(_1573__bF_buf18), .Y(_1651_) );
MUX2X1 MUX2X1_864 ( .A(_1651_), .B(_1589__bF_buf2), .S(_1642__bF_buf2), .Y(_903_) );
NAND2X1 NAND2X1_920 ( .A(REGs_USR_REGS_0__9_), .B(_1573__bF_buf31), .Y(_1652_) );
MUX2X1 MUX2X1_865 ( .A(_1652_), .B(_1591__bF_buf3), .S(_1642__bF_buf1), .Y(_904_) );
NAND2X1 NAND2X1_921 ( .A(REGs_USR_REGS_0__10_), .B(_1573__bF_buf31), .Y(_1653_) );
MUX2X1 MUX2X1_866 ( .A(_1653_), .B(_1593__bF_buf1), .S(_1642__bF_buf1), .Y(_905_) );
NAND2X1 NAND2X1_922 ( .A(REGs_USR_REGS_0__11_), .B(_1573__bF_buf40), .Y(_1654_) );
MUX2X1 MUX2X1_867 ( .A(_1654_), .B(_1595__bF_buf1), .S(_1642__bF_buf2), .Y(_906_) );
NAND2X1 NAND2X1_923 ( .A(REGs_USR_REGS_0__12_), .B(_1573__bF_buf3), .Y(_1655_) );
MUX2X1 MUX2X1_868 ( .A(_1655_), .B(_1597__bF_buf2), .S(_1642__bF_buf4), .Y(_907_) );
NAND2X1 NAND2X1_924 ( .A(REGs_USR_REGS_0__13_), .B(_1573__bF_buf32), .Y(_1656_) );
MUX2X1 MUX2X1_869 ( .A(_1656_), .B(_1599__bF_buf0), .S(_1642__bF_buf2), .Y(_908_) );
NAND2X1 NAND2X1_925 ( .A(REGs_USR_REGS_0__14_), .B(_1573__bF_buf77), .Y(_1657_) );
MUX2X1 MUX2X1_870 ( .A(_1657_), .B(_1601__bF_buf0), .S(_1642__bF_buf0), .Y(_909_) );
NAND2X1 NAND2X1_926 ( .A(REGs_USR_REGS_0__15_), .B(_1573__bF_buf74), .Y(_1658_) );
MUX2X1 MUX2X1_871 ( .A(_1658_), .B(_1603__bF_buf0), .S(_1642__bF_buf1), .Y(_910_) );
NAND2X1 NAND2X1_927 ( .A(REGs_USR_REGS_0__16_), .B(_1573__bF_buf31), .Y(_1659_) );
MUX2X1 MUX2X1_872 ( .A(_1659_), .B(_1605__bF_buf1), .S(_1642__bF_buf1), .Y(_911_) );
NAND2X1 NAND2X1_928 ( .A(REGs_USR_REGS_0__17_), .B(_1573__bF_buf57), .Y(_1660_) );
MUX2X1 MUX2X1_873 ( .A(_1660_), .B(_1607__bF_buf2), .S(_1642__bF_buf3), .Y(_912_) );
NAND2X1 NAND2X1_929 ( .A(REGs_USR_REGS_0__18_), .B(_1573__bF_buf64), .Y(_1661_) );
MUX2X1 MUX2X1_874 ( .A(_1661_), .B(_1609__bF_buf0), .S(_1642__bF_buf0), .Y(_913_) );
NAND2X1 NAND2X1_930 ( .A(REGs_USR_REGS_0__19_), .B(_1573__bF_buf43), .Y(_1662_) );
MUX2X1 MUX2X1_875 ( .A(_1662_), .B(_1611__bF_buf2), .S(_1642__bF_buf2), .Y(_914_) );
NAND2X1 NAND2X1_931 ( .A(REGs_USR_REGS_0__20_), .B(_1573__bF_buf48), .Y(_1663_) );
MUX2X1 MUX2X1_876 ( .A(_1663_), .B(_1613__bF_buf2), .S(_1642__bF_buf4), .Y(_915_) );
NAND2X1 NAND2X1_932 ( .A(REGs_USR_REGS_0__21_), .B(_1573__bF_buf8), .Y(_1664_) );
MUX2X1 MUX2X1_877 ( .A(_1664_), .B(_1615__bF_buf3), .S(_1642__bF_buf1), .Y(_916_) );
NAND2X1 NAND2X1_933 ( .A(REGs_USR_REGS_0__22_), .B(_1573__bF_buf11), .Y(_1665_) );
MUX2X1 MUX2X1_878 ( .A(_1665_), .B(_1617__bF_buf3), .S(_1642__bF_buf4), .Y(_917_) );
NAND2X1 NAND2X1_934 ( .A(REGs_USR_REGS_0__23_), .B(_1573__bF_buf25), .Y(_1666_) );
MUX2X1 MUX2X1_879 ( .A(_1666_), .B(_1619__bF_buf0), .S(_1642__bF_buf0), .Y(_918_) );
NAND2X1 NAND2X1_935 ( .A(REGs_USR_REGS_0__24_), .B(_1573__bF_buf30), .Y(_1667_) );
MUX2X1 MUX2X1_880 ( .A(_1667_), .B(_1621__bF_buf3), .S(_1642__bF_buf2), .Y(_919_) );
NAND2X1 NAND2X1_936 ( .A(REGs_USR_REGS_0__25_), .B(_1573__bF_buf76), .Y(_1668_) );
MUX2X1 MUX2X1_881 ( .A(_1668_), .B(_1623__bF_buf3), .S(_1642__bF_buf3), .Y(_920_) );
NAND2X1 NAND2X1_937 ( .A(REGs_USR_REGS_0__26_), .B(_1573__bF_buf69), .Y(_1669_) );
MUX2X1 MUX2X1_882 ( .A(_1669_), .B(_1625__bF_buf3), .S(_1642__bF_buf3), .Y(_921_) );
NAND2X1 NAND2X1_938 ( .A(REGs_USR_REGS_0__27_), .B(_1573__bF_buf57), .Y(_1670_) );
MUX2X1 MUX2X1_883 ( .A(_1670_), .B(_1627__bF_buf2), .S(_1642__bF_buf3), .Y(_922_) );
NAND2X1 NAND2X1_939 ( .A(REGs_USR_REGS_0__28_), .B(_1573__bF_buf26), .Y(_1671_) );
MUX2X1 MUX2X1_884 ( .A(_1671_), .B(_1629__bF_buf1), .S(_1642__bF_buf1), .Y(_923_) );
NAND2X1 NAND2X1_940 ( .A(REGs_USR_REGS_0__29_), .B(_1573__bF_buf58), .Y(_1672_) );
MUX2X1 MUX2X1_885 ( .A(_1672_), .B(_1631__bF_buf3), .S(_1642__bF_buf0), .Y(_924_) );
NAND2X1 NAND2X1_941 ( .A(REGs_USR_REGS_0__30_), .B(_1573__bF_buf56), .Y(_1673_) );
MUX2X1 MUX2X1_886 ( .A(_1673_), .B(_1633__bF_buf3), .S(_1642__bF_buf4), .Y(_925_) );
NAND2X1 NAND2X1_942 ( .A(REGs_USR_REGS_0__31_), .B(_1573__bF_buf32), .Y(_1674_) );
MUX2X1 MUX2X1_887 ( .A(_1674_), .B(_1635__bF_buf3), .S(_1642__bF_buf2), .Y(_926_) );
INVX1 INVX1_323 ( .A(CORE_REG_RF2_3_), .Y(_1675_) );
AND2X2 AND2X2_1285 ( .A(_1675_), .B(CORE_REG_RF2_2_), .Y(_1676_) );
NOR2X1 NOR2X1_175 ( .A(CORE_REG_RF2_1_), .B(CORE_REG_RF2_0_), .Y(_1677_) );
AND2X2 AND2X2_1286 ( .A(_1676_), .B(_1677_), .Y(_1678_) );
AND2X2 AND2X2_1287 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__0_), .Y(_1679_) );
INVX1 INVX1_324 ( .A(CORE_REG_RF2_1_), .Y(_1680_) );
AND2X2 AND2X2_1288 ( .A(_1680_), .B(CORE_REG_RF2_0_), .Y(_1681_) );
AND2X2 AND2X2_1289 ( .A(_1676_), .B(_1681_), .Y(_1682_) );
AND2X2 AND2X2_1290 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__0_), .Y(_1683_) );
OR2X2 OR2X2_1015 ( .A(_1679_), .B(_1683_), .Y(_1684_) );
INVX1 INVX1_325 ( .A(CORE_REG_RF2_0_), .Y(_1685_) );
AND2X2 AND2X2_1291 ( .A(_1685_), .B(CORE_REG_RF2_1_), .Y(_1686_) );
AND2X2 AND2X2_1292 ( .A(_1676_), .B(_1686_), .Y(_1687_) );
AND2X2 AND2X2_1293 ( .A(_1687__bF_buf0), .B(REGs_REGS_6__0_), .Y(_1688_) );
AND2X2 AND2X2_1294 ( .A(CORE_REG_RF2_1_), .B(CORE_REG_RF2_0_), .Y(_1689_) );
AND2X2 AND2X2_1295 ( .A(_1676_), .B(_1689_), .Y(_1690_) );
AND2X2 AND2X2_1296 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__0_), .Y(_1691_) );
OR2X2 OR2X2_1016 ( .A(_1691_), .B(_1688_), .Y(_1692_) );
OR2X2 OR2X2_1017 ( .A(_1684_), .B(_1692_), .Y(_1693_) );
NOR2X1 NOR2X1_176 ( .A(CORE_REG_RF2_3_), .B(CORE_REG_RF2_2_), .Y(_1694_) );
AND2X2 AND2X2_1297 ( .A(_1681_), .B(_1694_), .Y(_1695_) );
AND2X2 AND2X2_1298 ( .A(_1695__bF_buf4), .B(PC_ADDR_stack_1__0_), .Y(_1696_) );
AND2X2 AND2X2_1299 ( .A(_1694_), .B(_1689_), .Y(_1697_) );
AND2X2 AND2X2_1300 ( .A(_1697__bF_buf0), .B(REGs_REGS_3__0_), .Y(_1698_) );
AND2X2 AND2X2_1301 ( .A(_1686_), .B(_1694_), .Y(_1699_) );
AND2X2 AND2X2_1302 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__0_), .Y(_1700_) );
OR2X2 OR2X2_1018 ( .A(_1698_), .B(_1700_), .Y(_1701_) );
OR2X2 OR2X2_1019 ( .A(_1696_), .B(_1701_), .Y(_1702_) );
OR2X2 OR2X2_1020 ( .A(_1702_), .B(_1693_), .Y(_1703_) );
AND2X2 AND2X2_1303 ( .A(CORE_REG_RF2_3_), .B(CORE_REG_RF2_2_), .Y(_1704_) );
AND2X2 AND2X2_1304 ( .A(_1681_), .B(_1704_), .Y(_1705_) );
OR2X2 OR2X2_1021 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_5__0_), .Y(_1706_) );
OR2X2 OR2X2_1022 ( .A(REGs_FIRQ_REGS_5__0_), .B(_1568__bF_buf13), .Y(_1707_) );
AND2X2 AND2X2_1305 ( .A(_1707_), .B(_1706_), .Y(_1708_) );
AND2X2 AND2X2_1306 ( .A(_1708_), .B(_1705__bF_buf0), .Y(_1709_) );
AND2X2 AND2X2_1307 ( .A(_1677_), .B(_1704_), .Y(_1710_) );
OR2X2 OR2X2_1023 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_4__0_), .Y(_1711_) );
OR2X2 OR2X2_1024 ( .A(REGs_FIRQ_REGS_4__0_), .B(_1568__bF_buf6), .Y(_1712_) );
AND2X2 AND2X2_1308 ( .A(_1712_), .B(_1711_), .Y(_1713_) );
AND2X2 AND2X2_1309 ( .A(_1713_), .B(_1710__bF_buf2), .Y(_1714_) );
OR2X2 OR2X2_1025 ( .A(_1714_), .B(_1709_), .Y(_1715_) );
AND2X2 AND2X2_1310 ( .A(_1686_), .B(_1704_), .Y(_1716_) );
OR2X2 OR2X2_1026 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_6__0_), .Y(_1717_) );
OR2X2 OR2X2_1027 ( .A(REGs_FIRQ_REGS_6__0_), .B(_1568__bF_buf6), .Y(_1718_) );
AND2X2 AND2X2_1311 ( .A(_1718_), .B(_1717_), .Y(_1719_) );
AND2X2 AND2X2_1312 ( .A(_1719_), .B(_1716__bF_buf0), .Y(_1720_) );
AND2X2 AND2X2_1313 ( .A(_1689_), .B(_1704_), .Y(_1721_) );
OR2X2 OR2X2_1028 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_7__0_), .Y(_1722_) );
OR2X2 OR2X2_1029 ( .A(REGs_FIRQ_REGS_7__0_), .B(_1568__bF_buf13), .Y(_1723_) );
AND2X2 AND2X2_1314 ( .A(_1723_), .B(_1722_), .Y(_1724_) );
AND2X2 AND2X2_1315 ( .A(_1724_), .B(_1721__bF_buf2), .Y(_1725_) );
OR2X2 OR2X2_1030 ( .A(_1725_), .B(_1720_), .Y(_1726_) );
OR2X2 OR2X2_1031 ( .A(_1715_), .B(_1726_), .Y(_1727_) );
INVX1 INVX1_326 ( .A(CORE_REG_RF2_2_), .Y(_1728_) );
AND2X2 AND2X2_1316 ( .A(_1728_), .B(CORE_REG_RF2_3_), .Y(_1729_) );
AND2X2 AND2X2_1317 ( .A(_1729_), .B(_1677_), .Y(_1730_) );
OR2X2 OR2X2_1032 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_0__0_), .Y(_1731_) );
OR2X2 OR2X2_1033 ( .A(REGs_FIRQ_REGS_0__0_), .B(_1568__bF_buf4), .Y(_1732_) );
AND2X2 AND2X2_1318 ( .A(_1732_), .B(_1731_), .Y(_1733_) );
AND2X2 AND2X2_1319 ( .A(_1730__bF_buf2), .B(_1733_), .Y(_1734_) );
AND2X2 AND2X2_1320 ( .A(_1681_), .B(_1729_), .Y(_1735_) );
OR2X2 OR2X2_1034 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_1__0_), .Y(_1736_) );
OR2X2 OR2X2_1035 ( .A(REGs_FIRQ_REGS_1__0_), .B(_1568__bF_buf9), .Y(_1737_) );
AND2X2 AND2X2_1321 ( .A(_1737_), .B(_1736_), .Y(_1738_) );
AND2X2 AND2X2_1322 ( .A(_1735__bF_buf0), .B(_1738_), .Y(_1739_) );
OR2X2 OR2X2_1036 ( .A(_1734_), .B(_1739_), .Y(_1740_) );
AND2X2 AND2X2_1323 ( .A(_1729_), .B(_1689_), .Y(_1741_) );
OR2X2 OR2X2_1037 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_3__0_), .Y(_1742_) );
OR2X2 OR2X2_1038 ( .A(REGs_FIRQ_REGS_3__0_), .B(_1568__bF_buf9), .Y(_1743_) );
AND2X2 AND2X2_1324 ( .A(_1743_), .B(_1742_), .Y(_1744_) );
AND2X2 AND2X2_1325 ( .A(_1744_), .B(_1741__bF_buf1), .Y(_1745_) );
AND2X2 AND2X2_1326 ( .A(_1729_), .B(_1686_), .Y(_1746_) );
OR2X2 OR2X2_1039 ( .A(INTERRUPT_flag_bF_buf15_bF_buf3), .B(REGs_USR_REGS_2__0_), .Y(_1747_) );
OR2X2 OR2X2_1040 ( .A(REGs_FIRQ_REGS_2__0_), .B(_1568__bF_buf6), .Y(_1748_) );
AND2X2 AND2X2_1327 ( .A(_1748_), .B(_1747_), .Y(_1749_) );
AND2X2 AND2X2_1328 ( .A(_1746__bF_buf0), .B(_1749_), .Y(_1750_) );
OR2X2 OR2X2_1041 ( .A(_1745_), .B(_1750_), .Y(_1751_) );
OR2X2 OR2X2_1042 ( .A(_1751_), .B(_1740_), .Y(_1752_) );
OR2X2 OR2X2_1043 ( .A(_1727_), .B(_1752_), .Y(_1753_) );
OR2X2 OR2X2_1044 ( .A(_1703_), .B(_1753_), .Y(REG_B_0_) );
AND2X2 AND2X2_1329 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__1_), .Y(_1754_) );
AND2X2 AND2X2_1330 ( .A(_1682__bF_buf2), .B(REGs_REGS_5__1_), .Y(_1755_) );
OR2X2 OR2X2_1045 ( .A(_1754_), .B(_1755_), .Y(_1756_) );
AND2X2 AND2X2_1331 ( .A(_1687__bF_buf0), .B(REGs_REGS_6__1_), .Y(_1757_) );
AND2X2 AND2X2_1332 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__1_), .Y(_1758_) );
OR2X2 OR2X2_1046 ( .A(_1758_), .B(_1757_), .Y(_1759_) );
OR2X2 OR2X2_1047 ( .A(_1756_), .B(_1759_), .Y(_1760_) );
AND2X2 AND2X2_1333 ( .A(_1695__bF_buf4), .B(PC_ADDR_stack_1__1_), .Y(_1761_) );
AND2X2 AND2X2_1334 ( .A(_1697__bF_buf0), .B(REGs_REGS_3__1_), .Y(_1762_) );
AND2X2 AND2X2_1335 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__1_), .Y(_1763_) );
OR2X2 OR2X2_1048 ( .A(_1762_), .B(_1763_), .Y(_1764_) );
OR2X2 OR2X2_1049 ( .A(_1761_), .B(_1764_), .Y(_1765_) );
OR2X2 OR2X2_1050 ( .A(_1765_), .B(_1760_), .Y(_1766_) );
OR2X2 OR2X2_1051 ( .A(INTERRUPT_flag_bF_buf14_bF_buf1), .B(REGs_USR_REGS_5__1_), .Y(_1767_) );
OR2X2 OR2X2_1052 ( .A(REGs_FIRQ_REGS_5__1_), .B(_1568__bF_buf5), .Y(_1768_) );
AND2X2 AND2X2_1336 ( .A(_1768_), .B(_1767_), .Y(_1769_) );
AND2X2 AND2X2_1337 ( .A(_1769_), .B(_1705__bF_buf2), .Y(_1770_) );
OR2X2 OR2X2_1053 ( .A(INTERRUPT_flag_bF_buf13_bF_buf1), .B(REGs_USR_REGS_4__1_), .Y(_1771_) );
OR2X2 OR2X2_1054 ( .A(REGs_FIRQ_REGS_4__1_), .B(_1568__bF_buf5), .Y(_1772_) );
AND2X2 AND2X2_1338 ( .A(_1772_), .B(_1771_), .Y(_1773_) );
AND2X2 AND2X2_1339 ( .A(_1773_), .B(_1710__bF_buf1), .Y(_1774_) );
OR2X2 OR2X2_1055 ( .A(_1774_), .B(_1770_), .Y(_1775_) );
OR2X2 OR2X2_1056 ( .A(INTERRUPT_flag_bF_buf12_bF_buf3), .B(REGs_USR_REGS_6__1_), .Y(_1776_) );
OR2X2 OR2X2_1057 ( .A(REGs_FIRQ_REGS_6__1_), .B(_1568__bF_buf12), .Y(_1777_) );
AND2X2 AND2X2_1340 ( .A(_1777_), .B(_1776_), .Y(_1778_) );
AND2X2 AND2X2_1341 ( .A(_1778_), .B(_1716__bF_buf1), .Y(_1779_) );
OR2X2 OR2X2_1058 ( .A(INTERRUPT_flag_bF_buf11_bF_buf2), .B(REGs_USR_REGS_7__1_), .Y(_1780_) );
OR2X2 OR2X2_1059 ( .A(REGs_FIRQ_REGS_7__1_), .B(_1568__bF_buf5), .Y(_1781_) );
AND2X2 AND2X2_1342 ( .A(_1781_), .B(_1780_), .Y(_1782_) );
AND2X2 AND2X2_1343 ( .A(_1782_), .B(_1721__bF_buf1), .Y(_1783_) );
OR2X2 OR2X2_1060 ( .A(_1783_), .B(_1779_), .Y(_1784_) );
OR2X2 OR2X2_1061 ( .A(_1775_), .B(_1784_), .Y(_1785_) );
OR2X2 OR2X2_1062 ( .A(INTERRUPT_flag_bF_buf10_bF_buf3), .B(REGs_USR_REGS_0__1_), .Y(_1786_) );
OR2X2 OR2X2_1063 ( .A(REGs_FIRQ_REGS_0__1_), .B(_1568__bF_buf3), .Y(_1787_) );
AND2X2 AND2X2_1344 ( .A(_1787_), .B(_1786_), .Y(_1788_) );
AND2X2 AND2X2_1345 ( .A(_1730__bF_buf0), .B(_1788_), .Y(_1789_) );
OR2X2 OR2X2_1064 ( .A(INTERRUPT_flag_bF_buf9_bF_buf3), .B(REGs_USR_REGS_1__1_), .Y(_1790_) );
OR2X2 OR2X2_1065 ( .A(REGs_FIRQ_REGS_1__1_), .B(_1568__bF_buf7), .Y(_1791_) );
AND2X2 AND2X2_1346 ( .A(_1791_), .B(_1790_), .Y(_1792_) );
AND2X2 AND2X2_1347 ( .A(_1735__bF_buf2), .B(_1792_), .Y(_1793_) );
OR2X2 OR2X2_1066 ( .A(_1789_), .B(_1793_), .Y(_1794_) );
OR2X2 OR2X2_1067 ( .A(INTERRUPT_flag_bF_buf8_bF_buf2), .B(REGs_USR_REGS_3__1_), .Y(_1795_) );
OR2X2 OR2X2_1068 ( .A(REGs_FIRQ_REGS_3__1_), .B(_1568__bF_buf6), .Y(_1796_) );
AND2X2 AND2X2_1348 ( .A(_1796_), .B(_1795_), .Y(_1797_) );
AND2X2 AND2X2_1349 ( .A(_1797_), .B(_1741__bF_buf4), .Y(_1798_) );
OR2X2 OR2X2_1069 ( .A(INTERRUPT_flag_bF_buf7_bF_buf0), .B(REGs_USR_REGS_2__1_), .Y(_1799_) );
OR2X2 OR2X2_1070 ( .A(REGs_FIRQ_REGS_2__1_), .B(_1568__bF_buf15_bF_buf1), .Y(_1800_) );
AND2X2 AND2X2_1350 ( .A(_1800_), .B(_1799_), .Y(_1801_) );
AND2X2 AND2X2_1351 ( .A(_1746__bF_buf4), .B(_1801_), .Y(_1802_) );
OR2X2 OR2X2_1071 ( .A(_1798_), .B(_1802_), .Y(_1803_) );
OR2X2 OR2X2_1072 ( .A(_1803_), .B(_1794_), .Y(_1804_) );
OR2X2 OR2X2_1073 ( .A(_1785_), .B(_1804_), .Y(_1805_) );
OR2X2 OR2X2_1074 ( .A(_1766_), .B(_1805_), .Y(REG_B_1_) );
AND2X2 AND2X2_1352 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__2_), .Y(_1806_) );
AND2X2 AND2X2_1353 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__2_), .Y(_1807_) );
OR2X2 OR2X2_1075 ( .A(_1806_), .B(_1807_), .Y(_1808_) );
AND2X2 AND2X2_1354 ( .A(_1687__bF_buf1), .B(REGs_REGS_6__2_), .Y(_1809_) );
AND2X2 AND2X2_1355 ( .A(_1690__bF_buf2), .B(REGs_REGS_7__2_), .Y(_1810_) );
OR2X2 OR2X2_1076 ( .A(_1810_), .B(_1809_), .Y(_1811_) );
OR2X2 OR2X2_1077 ( .A(_1808_), .B(_1811_), .Y(_1812_) );
AND2X2 AND2X2_1356 ( .A(_1695__bF_buf0), .B(PC_ADDR_stack_1__2_), .Y(_1813_) );
AND2X2 AND2X2_1357 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__2_), .Y(_1814_) );
AND2X2 AND2X2_1358 ( .A(_1699__bF_buf0), .B(REGs_REGS_2__2_), .Y(_1815_) );
OR2X2 OR2X2_1078 ( .A(_1814_), .B(_1815_), .Y(_1816_) );
OR2X2 OR2X2_1079 ( .A(_1813_), .B(_1816_), .Y(_1817_) );
OR2X2 OR2X2_1080 ( .A(_1817_), .B(_1812_), .Y(_1818_) );
OR2X2 OR2X2_1081 ( .A(INTERRUPT_flag_bF_buf15), .B(REGs_USR_REGS_5__2_), .Y(_1819_) );
OR2X2 OR2X2_1082 ( .A(REGs_FIRQ_REGS_5__2_), .B(_1568__bF_buf0), .Y(_1820_) );
AND2X2 AND2X2_1359 ( .A(_1820_), .B(_1819_), .Y(_1821_) );
AND2X2 AND2X2_1360 ( .A(_1821_), .B(_1705__bF_buf4), .Y(_1822_) );
OR2X2 OR2X2_1083 ( .A(INTERRUPT_flag_bF_buf15), .B(REGs_USR_REGS_4__2_), .Y(_1823_) );
OR2X2 OR2X2_1084 ( .A(REGs_FIRQ_REGS_4__2_), .B(_1568__bF_buf13), .Y(_1824_) );
AND2X2 AND2X2_1361 ( .A(_1824_), .B(_1823_), .Y(_1825_) );
AND2X2 AND2X2_1362 ( .A(_1825_), .B(_1710__bF_buf3), .Y(_1826_) );
OR2X2 OR2X2_1085 ( .A(_1826_), .B(_1822_), .Y(_1827_) );
OR2X2 OR2X2_1086 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_6__2_), .Y(_1828_) );
OR2X2 OR2X2_1087 ( .A(REGs_FIRQ_REGS_6__2_), .B(_1568__bF_buf1), .Y(_1829_) );
AND2X2 AND2X2_1363 ( .A(_1829_), .B(_1828_), .Y(_1830_) );
AND2X2 AND2X2_1364 ( .A(_1830_), .B(_1716__bF_buf4), .Y(_1831_) );
OR2X2 OR2X2_1088 ( .A(INTERRUPT_flag_bF_buf15), .B(REGs_USR_REGS_7__2_), .Y(_1832_) );
OR2X2 OR2X2_1089 ( .A(REGs_FIRQ_REGS_7__2_), .B(_1568__bF_buf6), .Y(_1833_) );
AND2X2 AND2X2_1365 ( .A(_1833_), .B(_1832_), .Y(_1834_) );
AND2X2 AND2X2_1366 ( .A(_1834_), .B(_1721__bF_buf0), .Y(_1835_) );
OR2X2 OR2X2_1090 ( .A(_1835_), .B(_1831_), .Y(_1836_) );
OR2X2 OR2X2_1091 ( .A(_1827_), .B(_1836_), .Y(_1837_) );
OR2X2 OR2X2_1092 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_0__2_), .Y(_1838_) );
OR2X2 OR2X2_1093 ( .A(REGs_FIRQ_REGS_0__2_), .B(_1568__bF_buf1), .Y(_1839_) );
AND2X2 AND2X2_1367 ( .A(_1839_), .B(_1838_), .Y(_1840_) );
AND2X2 AND2X2_1368 ( .A(_1730__bF_buf3), .B(_1840_), .Y(_1841_) );
OR2X2 OR2X2_1094 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_1__2_), .Y(_1842_) );
OR2X2 OR2X2_1095 ( .A(REGs_FIRQ_REGS_1__2_), .B(_1568__bF_buf1), .Y(_1843_) );
AND2X2 AND2X2_1369 ( .A(_1843_), .B(_1842_), .Y(_1844_) );
AND2X2 AND2X2_1370 ( .A(_1735__bF_buf1), .B(_1844_), .Y(_1845_) );
OR2X2 OR2X2_1096 ( .A(_1841_), .B(_1845_), .Y(_1846_) );
OR2X2 OR2X2_1097 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_3__2_), .Y(_1847_) );
OR2X2 OR2X2_1098 ( .A(REGs_FIRQ_REGS_3__2_), .B(_1568__bF_buf1), .Y(_1848_) );
AND2X2 AND2X2_1371 ( .A(_1848_), .B(_1847_), .Y(_1849_) );
AND2X2 AND2X2_1372 ( .A(_1849_), .B(_1741__bF_buf3), .Y(_1850_) );
OR2X2 OR2X2_1099 ( .A(INTERRUPT_flag_bF_buf15_bF_buf1), .B(REGs_USR_REGS_2__2_), .Y(_1851_) );
OR2X2 OR2X2_1100 ( .A(REGs_FIRQ_REGS_2__2_), .B(_1568__bF_buf1), .Y(_1852_) );
AND2X2 AND2X2_1373 ( .A(_1852_), .B(_1851_), .Y(_1853_) );
AND2X2 AND2X2_1374 ( .A(_1746__bF_buf0), .B(_1853_), .Y(_1854_) );
OR2X2 OR2X2_1101 ( .A(_1850_), .B(_1854_), .Y(_1855_) );
OR2X2 OR2X2_1102 ( .A(_1855_), .B(_1846_), .Y(_1856_) );
OR2X2 OR2X2_1103 ( .A(_1837_), .B(_1856_), .Y(_1857_) );
OR2X2 OR2X2_1104 ( .A(_1818_), .B(_1857_), .Y(REG_B_2_) );
AND2X2 AND2X2_1375 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__3_), .Y(_1858_) );
AND2X2 AND2X2_1376 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__3_), .Y(_1859_) );
OR2X2 OR2X2_1105 ( .A(_1858_), .B(_1859_), .Y(_1860_) );
AND2X2 AND2X2_1377 ( .A(_1687__bF_buf1), .B(REGs_REGS_6__3_), .Y(_1861_) );
AND2X2 AND2X2_1378 ( .A(_1690__bF_buf2), .B(REGs_REGS_7__3_), .Y(_1862_) );
OR2X2 OR2X2_1106 ( .A(_1862_), .B(_1861_), .Y(_1863_) );
OR2X2 OR2X2_1107 ( .A(_1860_), .B(_1863_), .Y(_1864_) );
AND2X2 AND2X2_1379 ( .A(_1695__bF_buf0), .B(PC_ADDR_stack_1__3_), .Y(_1865_) );
AND2X2 AND2X2_1380 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__3_), .Y(_1866_) );
AND2X2 AND2X2_1381 ( .A(_1699__bF_buf0), .B(REGs_REGS_2__3_), .Y(_1867_) );
OR2X2 OR2X2_1108 ( .A(_1866_), .B(_1867_), .Y(_1868_) );
OR2X2 OR2X2_1109 ( .A(_1865_), .B(_1868_), .Y(_1869_) );
OR2X2 OR2X2_1110 ( .A(_1869_), .B(_1864_), .Y(_1870_) );
OR2X2 OR2X2_1111 ( .A(INTERRUPT_flag_bF_buf14_bF_buf3), .B(REGs_USR_REGS_5__3_), .Y(_1871_) );
OR2X2 OR2X2_1112 ( .A(REGs_FIRQ_REGS_5__3_), .B(_1568__bF_buf15), .Y(_1872_) );
AND2X2 AND2X2_1382 ( .A(_1872_), .B(_1871_), .Y(_1873_) );
AND2X2 AND2X2_1383 ( .A(_1873_), .B(_1705__bF_buf4), .Y(_1874_) );
OR2X2 OR2X2_1113 ( .A(INTERRUPT_flag_bF_buf13_bF_buf0), .B(REGs_USR_REGS_4__3_), .Y(_1875_) );
OR2X2 OR2X2_1114 ( .A(REGs_FIRQ_REGS_4__3_), .B(_1568__bF_buf0), .Y(_1876_) );
AND2X2 AND2X2_1384 ( .A(_1876_), .B(_1875_), .Y(_1877_) );
AND2X2 AND2X2_1385 ( .A(_1877_), .B(_1710__bF_buf3), .Y(_1878_) );
OR2X2 OR2X2_1115 ( .A(_1878_), .B(_1874_), .Y(_1879_) );
OR2X2 OR2X2_1116 ( .A(INTERRUPT_flag_bF_buf12_bF_buf2), .B(REGs_USR_REGS_6__3_), .Y(_1880_) );
OR2X2 OR2X2_1117 ( .A(REGs_FIRQ_REGS_6__3_), .B(_1568__bF_buf0), .Y(_1881_) );
AND2X2 AND2X2_1386 ( .A(_1881_), .B(_1880_), .Y(_1882_) );
AND2X2 AND2X2_1387 ( .A(_1882_), .B(_1716__bF_buf4), .Y(_1883_) );
OR2X2 OR2X2_1118 ( .A(INTERRUPT_flag_bF_buf11_bF_buf1), .B(REGs_USR_REGS_7__3_), .Y(_1884_) );
OR2X2 OR2X2_1119 ( .A(REGs_FIRQ_REGS_7__3_), .B(_1568__bF_buf0), .Y(_1885_) );
AND2X2 AND2X2_1388 ( .A(_1885_), .B(_1884_), .Y(_1886_) );
AND2X2 AND2X2_1389 ( .A(_1886_), .B(_1721__bF_buf0), .Y(_1887_) );
OR2X2 OR2X2_1120 ( .A(_1887_), .B(_1883_), .Y(_1888_) );
OR2X2 OR2X2_1121 ( .A(_1879_), .B(_1888_), .Y(_1889_) );
OR2X2 OR2X2_1122 ( .A(INTERRUPT_flag_bF_buf10_bF_buf3), .B(REGs_USR_REGS_0__3_), .Y(_1890_) );
OR2X2 OR2X2_1123 ( .A(REGs_FIRQ_REGS_0__3_), .B(_1568__bF_buf0), .Y(_1891_) );
AND2X2 AND2X2_1390 ( .A(_1891_), .B(_1890_), .Y(_1892_) );
AND2X2 AND2X2_1391 ( .A(_1730__bF_buf3), .B(_1892_), .Y(_1893_) );
OR2X2 OR2X2_1124 ( .A(INTERRUPT_flag_bF_buf9_bF_buf0), .B(REGs_USR_REGS_1__3_), .Y(_1894_) );
OR2X2 OR2X2_1125 ( .A(REGs_FIRQ_REGS_1__3_), .B(_1568__bF_buf0), .Y(_1895_) );
AND2X2 AND2X2_1392 ( .A(_1895_), .B(_1894_), .Y(_1896_) );
AND2X2 AND2X2_1393 ( .A(_1735__bF_buf1), .B(_1896_), .Y(_1897_) );
OR2X2 OR2X2_1126 ( .A(_1893_), .B(_1897_), .Y(_1898_) );
OR2X2 OR2X2_1127 ( .A(INTERRUPT_flag_bF_buf8_bF_buf0), .B(REGs_USR_REGS_3__3_), .Y(_1899_) );
OR2X2 OR2X2_1128 ( .A(REGs_FIRQ_REGS_3__3_), .B(_1568__bF_buf15), .Y(_1900_) );
AND2X2 AND2X2_1394 ( .A(_1900_), .B(_1899_), .Y(_1901_) );
AND2X2 AND2X2_1395 ( .A(_1901_), .B(_1741__bF_buf3), .Y(_1902_) );
OR2X2 OR2X2_1129 ( .A(INTERRUPT_flag_bF_buf7_bF_buf2), .B(REGs_USR_REGS_2__3_), .Y(_1903_) );
OR2X2 OR2X2_1130 ( .A(REGs_FIRQ_REGS_2__3_), .B(_1568__bF_buf15_bF_buf2), .Y(_1904_) );
AND2X2 AND2X2_1396 ( .A(_1904_), .B(_1903_), .Y(_1905_) );
AND2X2 AND2X2_1397 ( .A(_1746__bF_buf1), .B(_1905_), .Y(_1906_) );
OR2X2 OR2X2_1131 ( .A(_1902_), .B(_1906_), .Y(_1907_) );
OR2X2 OR2X2_1132 ( .A(_1907_), .B(_1898_), .Y(_1908_) );
OR2X2 OR2X2_1133 ( .A(_1889_), .B(_1908_), .Y(_1909_) );
OR2X2 OR2X2_1134 ( .A(_1870_), .B(_1909_), .Y(REG_B_3_) );
AND2X2 AND2X2_1398 ( .A(_1678__bF_buf0), .B(REGs_REGS_4__4_), .Y(_1910_) );
AND2X2 AND2X2_1399 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__4_), .Y(_1911_) );
OR2X2 OR2X2_1135 ( .A(_1910_), .B(_1911_), .Y(_1912_) );
AND2X2 AND2X2_1400 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__4_), .Y(_1913_) );
AND2X2 AND2X2_1401 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__4_), .Y(_1914_) );
OR2X2 OR2X2_1136 ( .A(_1914_), .B(_1913_), .Y(_1915_) );
OR2X2 OR2X2_1137 ( .A(_1912_), .B(_1915_), .Y(_1916_) );
AND2X2 AND2X2_1402 ( .A(_1695__bF_buf2), .B(PC_ADDR_stack_1__4_), .Y(_1917_) );
AND2X2 AND2X2_1403 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__4_), .Y(_1918_) );
AND2X2 AND2X2_1404 ( .A(_1699__bF_buf2), .B(REGs_REGS_2__4_), .Y(_1919_) );
OR2X2 OR2X2_1138 ( .A(_1918_), .B(_1919_), .Y(_1920_) );
OR2X2 OR2X2_1139 ( .A(_1917_), .B(_1920_), .Y(_1921_) );
OR2X2 OR2X2_1140 ( .A(_1921_), .B(_1916_), .Y(_1922_) );
OR2X2 OR2X2_1141 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_5__4_), .Y(_1923_) );
OR2X2 OR2X2_1142 ( .A(REGs_FIRQ_REGS_5__4_), .B(_1568__bF_buf14), .Y(_1924_) );
AND2X2 AND2X2_1405 ( .A(_1924_), .B(_1923_), .Y(_1925_) );
AND2X2 AND2X2_1406 ( .A(_1925_), .B(_1705__bF_buf4), .Y(_1926_) );
OR2X2 OR2X2_1143 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_4__4_), .Y(_1927_) );
OR2X2 OR2X2_1144 ( .A(REGs_FIRQ_REGS_4__4_), .B(_1568__bF_buf14), .Y(_1928_) );
AND2X2 AND2X2_1407 ( .A(_1928_), .B(_1927_), .Y(_1929_) );
AND2X2 AND2X2_1408 ( .A(_1929_), .B(_1710__bF_buf3), .Y(_1930_) );
OR2X2 OR2X2_1145 ( .A(_1930_), .B(_1926_), .Y(_1931_) );
OR2X2 OR2X2_1146 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_6__4_), .Y(_1932_) );
OR2X2 OR2X2_1147 ( .A(REGs_FIRQ_REGS_6__4_), .B(_1568__bF_buf14), .Y(_1933_) );
AND2X2 AND2X2_1409 ( .A(_1933_), .B(_1932_), .Y(_1934_) );
AND2X2 AND2X2_1410 ( .A(_1934_), .B(_1716__bF_buf4), .Y(_1935_) );
OR2X2 OR2X2_1148 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_7__4_), .Y(_1936_) );
OR2X2 OR2X2_1149 ( .A(REGs_FIRQ_REGS_7__4_), .B(_1568__bF_buf14), .Y(_1937_) );
AND2X2 AND2X2_1411 ( .A(_1937_), .B(_1936_), .Y(_1938_) );
AND2X2 AND2X2_1412 ( .A(_1938_), .B(_1721__bF_buf0), .Y(_1939_) );
OR2X2 OR2X2_1150 ( .A(_1939_), .B(_1935_), .Y(_1940_) );
OR2X2 OR2X2_1151 ( .A(_1931_), .B(_1940_), .Y(_1941_) );
OR2X2 OR2X2_1152 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_0__4_), .Y(_1942_) );
OR2X2 OR2X2_1153 ( .A(REGs_FIRQ_REGS_0__4_), .B(_1568__bF_buf14), .Y(_1943_) );
AND2X2 AND2X2_1413 ( .A(_1943_), .B(_1942_), .Y(_1944_) );
AND2X2 AND2X2_1414 ( .A(_1730__bF_buf3), .B(_1944_), .Y(_1945_) );
OR2X2 OR2X2_1154 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_1__4_), .Y(_1946_) );
OR2X2 OR2X2_1155 ( .A(REGs_FIRQ_REGS_1__4_), .B(_1568__bF_buf14), .Y(_1947_) );
AND2X2 AND2X2_1415 ( .A(_1947_), .B(_1946_), .Y(_1948_) );
AND2X2 AND2X2_1416 ( .A(_1735__bF_buf1), .B(_1948_), .Y(_1949_) );
OR2X2 OR2X2_1156 ( .A(_1945_), .B(_1949_), .Y(_1950_) );
OR2X2 OR2X2_1157 ( .A(INTERRUPT_flag_bF_buf13), .B(REGs_USR_REGS_3__4_), .Y(_1951_) );
OR2X2 OR2X2_1158 ( .A(REGs_FIRQ_REGS_3__4_), .B(_1568__bF_buf11), .Y(_1952_) );
AND2X2 AND2X2_1417 ( .A(_1952_), .B(_1951_), .Y(_1953_) );
AND2X2 AND2X2_1418 ( .A(_1953_), .B(_1741__bF_buf3), .Y(_1954_) );
OR2X2 OR2X2_1159 ( .A(INTERRUPT_flag_bF_buf15_bF_buf2), .B(REGs_USR_REGS_2__4_), .Y(_1955_) );
OR2X2 OR2X2_1160 ( .A(REGs_FIRQ_REGS_2__4_), .B(_1568__bF_buf11), .Y(_1956_) );
AND2X2 AND2X2_1419 ( .A(_1956_), .B(_1955_), .Y(_1957_) );
AND2X2 AND2X2_1420 ( .A(_1746__bF_buf1), .B(_1957_), .Y(_1958_) );
OR2X2 OR2X2_1161 ( .A(_1954_), .B(_1958_), .Y(_1959_) );
OR2X2 OR2X2_1162 ( .A(_1959_), .B(_1950_), .Y(_1960_) );
OR2X2 OR2X2_1163 ( .A(_1941_), .B(_1960_), .Y(_1961_) );
OR2X2 OR2X2_1164 ( .A(_1922_), .B(_1961_), .Y(REG_B_4_) );
AND2X2 AND2X2_1421 ( .A(_1678__bF_buf1), .B(REGs_REGS_4__5_), .Y(_1962_) );
AND2X2 AND2X2_1422 ( .A(_1682__bF_buf0), .B(REGs_REGS_5__5_), .Y(_1963_) );
OR2X2 OR2X2_1165 ( .A(_1962_), .B(_1963_), .Y(_1964_) );
AND2X2 AND2X2_1423 ( .A(_1687__bF_buf0), .B(REGs_REGS_6__5_), .Y(_1965_) );
AND2X2 AND2X2_1424 ( .A(_1690__bF_buf1), .B(REGs_REGS_7__5_), .Y(_1966_) );
OR2X2 OR2X2_1166 ( .A(_1966_), .B(_1965_), .Y(_1967_) );
OR2X2 OR2X2_1167 ( .A(_1964_), .B(_1967_), .Y(_1968_) );
AND2X2 AND2X2_1425 ( .A(_1695__bF_buf1), .B(PC_ADDR_stack_1__5_), .Y(_1969_) );
AND2X2 AND2X2_1426 ( .A(_1697__bF_buf2), .B(REGs_REGS_3__5_), .Y(_1970_) );
AND2X2 AND2X2_1427 ( .A(_1699__bF_buf1), .B(REGs_REGS_2__5_), .Y(_1971_) );
OR2X2 OR2X2_1168 ( .A(_1970_), .B(_1971_), .Y(_1972_) );
OR2X2 OR2X2_1169 ( .A(_1969_), .B(_1972_), .Y(_1973_) );
OR2X2 OR2X2_1170 ( .A(_1973_), .B(_1968_), .Y(_1974_) );
OR2X2 OR2X2_1171 ( .A(INTERRUPT_flag_bF_buf14_bF_buf1), .B(REGs_USR_REGS_5__5_), .Y(_1975_) );
OR2X2 OR2X2_1172 ( .A(REGs_FIRQ_REGS_5__5_), .B(_1568__bF_buf12), .Y(_1976_) );
AND2X2 AND2X2_1428 ( .A(_1976_), .B(_1975_), .Y(_1977_) );
AND2X2 AND2X2_1429 ( .A(_1977_), .B(_1705__bF_buf1), .Y(_1978_) );
OR2X2 OR2X2_1173 ( .A(INTERRUPT_flag_bF_buf13_bF_buf1), .B(REGs_USR_REGS_4__5_), .Y(_1979_) );
OR2X2 OR2X2_1174 ( .A(REGs_FIRQ_REGS_4__5_), .B(_1568__bF_buf5), .Y(_1980_) );
AND2X2 AND2X2_1430 ( .A(_1980_), .B(_1979_), .Y(_1981_) );
AND2X2 AND2X2_1431 ( .A(_1981_), .B(_1710__bF_buf0), .Y(_1982_) );
OR2X2 OR2X2_1175 ( .A(_1982_), .B(_1978_), .Y(_1983_) );
OR2X2 OR2X2_1176 ( .A(INTERRUPT_flag_bF_buf12_bF_buf1), .B(REGs_USR_REGS_6__5_), .Y(_1984_) );
OR2X2 OR2X2_1177 ( .A(REGs_FIRQ_REGS_6__5_), .B(_1568__bF_buf8), .Y(_1985_) );
AND2X2 AND2X2_1432 ( .A(_1985_), .B(_1984_), .Y(_1986_) );
AND2X2 AND2X2_1433 ( .A(_1986_), .B(_1716__bF_buf2), .Y(_1987_) );
OR2X2 OR2X2_1178 ( .A(INTERRUPT_flag_bF_buf11_bF_buf0), .B(REGs_USR_REGS_7__5_), .Y(_1988_) );
OR2X2 OR2X2_1179 ( .A(REGs_FIRQ_REGS_7__5_), .B(_1568__bF_buf12), .Y(_1989_) );
AND2X2 AND2X2_1434 ( .A(_1989_), .B(_1988_), .Y(_1990_) );
AND2X2 AND2X2_1435 ( .A(_1990_), .B(_1721__bF_buf4), .Y(_1991_) );
OR2X2 OR2X2_1180 ( .A(_1991_), .B(_1987_), .Y(_1992_) );
OR2X2 OR2X2_1181 ( .A(_1983_), .B(_1992_), .Y(_1993_) );
OR2X2 OR2X2_1182 ( .A(INTERRUPT_flag_bF_buf10_bF_buf3), .B(REGs_USR_REGS_0__5_), .Y(_1994_) );
OR2X2 OR2X2_1183 ( .A(REGs_FIRQ_REGS_0__5_), .B(_1568__bF_buf3), .Y(_1995_) );
AND2X2 AND2X2_1436 ( .A(_1995_), .B(_1994_), .Y(_1996_) );
AND2X2 AND2X2_1437 ( .A(_1730__bF_buf0), .B(_1996_), .Y(_1997_) );
OR2X2 OR2X2_1184 ( .A(INTERRUPT_flag_bF_buf9_bF_buf3), .B(REGs_USR_REGS_1__5_), .Y(_1998_) );
OR2X2 OR2X2_1185 ( .A(REGs_FIRQ_REGS_1__5_), .B(_1568__bF_buf3), .Y(_1999_) );
AND2X2 AND2X2_1438 ( .A(_1999_), .B(_1998_), .Y(_2000_) );
AND2X2 AND2X2_1439 ( .A(_1735__bF_buf2), .B(_2000_), .Y(_2001_) );
OR2X2 OR2X2_1186 ( .A(_1997_), .B(_2001_), .Y(_2002_) );
OR2X2 OR2X2_1187 ( .A(INTERRUPT_flag_bF_buf8_bF_buf1), .B(REGs_USR_REGS_3__5_), .Y(_2003_) );
OR2X2 OR2X2_1188 ( .A(REGs_FIRQ_REGS_3__5_), .B(_1568__bF_buf7), .Y(_2004_) );
AND2X2 AND2X2_1440 ( .A(_2004_), .B(_2003_), .Y(_2005_) );
AND2X2 AND2X2_1441 ( .A(_2005_), .B(_1741__bF_buf4), .Y(_2006_) );
OR2X2 OR2X2_1189 ( .A(INTERRUPT_flag_bF_buf7_bF_buf1), .B(REGs_USR_REGS_2__5_), .Y(_2007_) );
OR2X2 OR2X2_1190 ( .A(REGs_FIRQ_REGS_2__5_), .B(_1568__bF_buf15_bF_buf1), .Y(_2008_) );
AND2X2 AND2X2_1442 ( .A(_2008_), .B(_2007_), .Y(_2009_) );
AND2X2 AND2X2_1443 ( .A(_1746__bF_buf4), .B(_2009_), .Y(_2010_) );
OR2X2 OR2X2_1191 ( .A(_2006_), .B(_2010_), .Y(_2011_) );
OR2X2 OR2X2_1192 ( .A(_2011_), .B(_2002_), .Y(_2012_) );
OR2X2 OR2X2_1193 ( .A(_1993_), .B(_2012_), .Y(_2013_) );
OR2X2 OR2X2_1194 ( .A(_1974_), .B(_2013_), .Y(REG_B_5_) );
AND2X2 AND2X2_1444 ( .A(_1678__bF_buf0), .B(REGs_REGS_4__6_), .Y(_2014_) );
AND2X2 AND2X2_1445 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__6_), .Y(_2015_) );
OR2X2 OR2X2_1195 ( .A(_2014_), .B(_2015_), .Y(_2016_) );
AND2X2 AND2X2_1446 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__6_), .Y(_2017_) );
AND2X2 AND2X2_1447 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__6_), .Y(_2018_) );
OR2X2 OR2X2_1196 ( .A(_2018_), .B(_2017_), .Y(_2019_) );
OR2X2 OR2X2_1197 ( .A(_2016_), .B(_2019_), .Y(_2020_) );
AND2X2 AND2X2_1448 ( .A(_1695__bF_buf2), .B(PC_ADDR_stack_1__6_), .Y(_2021_) );
AND2X2 AND2X2_1449 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__6_), .Y(_2022_) );
AND2X2 AND2X2_1450 ( .A(_1699__bF_buf2), .B(REGs_REGS_2__6_), .Y(_2023_) );
OR2X2 OR2X2_1198 ( .A(_2022_), .B(_2023_), .Y(_2024_) );
OR2X2 OR2X2_1199 ( .A(_2021_), .B(_2024_), .Y(_2025_) );
OR2X2 OR2X2_1200 ( .A(_2025_), .B(_2020_), .Y(_2026_) );
OR2X2 OR2X2_1201 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_5__6_), .Y(_2027_) );
OR2X2 OR2X2_1202 ( .A(REGs_FIRQ_REGS_5__6_), .B(_1568__bF_buf14), .Y(_2028_) );
AND2X2 AND2X2_1451 ( .A(_2028_), .B(_2027_), .Y(_2029_) );
AND2X2 AND2X2_1452 ( .A(_2029_), .B(_1705__bF_buf4), .Y(_2030_) );
OR2X2 OR2X2_1203 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_4__6_), .Y(_2031_) );
OR2X2 OR2X2_1204 ( .A(REGs_FIRQ_REGS_4__6_), .B(_1568__bF_buf14), .Y(_2032_) );
AND2X2 AND2X2_1453 ( .A(_2032_), .B(_2031_), .Y(_2033_) );
AND2X2 AND2X2_1454 ( .A(_2033_), .B(_1710__bF_buf3), .Y(_2034_) );
OR2X2 OR2X2_1205 ( .A(_2034_), .B(_2030_), .Y(_2035_) );
OR2X2 OR2X2_1206 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_6__6_), .Y(_2036_) );
OR2X2 OR2X2_1207 ( .A(REGs_FIRQ_REGS_6__6_), .B(_1568__bF_buf11), .Y(_2037_) );
AND2X2 AND2X2_1455 ( .A(_2037_), .B(_2036_), .Y(_2038_) );
AND2X2 AND2X2_1456 ( .A(_2038_), .B(_1716__bF_buf4), .Y(_2039_) );
OR2X2 OR2X2_1208 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_7__6_), .Y(_2040_) );
OR2X2 OR2X2_1209 ( .A(REGs_FIRQ_REGS_7__6_), .B(_1568__bF_buf14), .Y(_2041_) );
AND2X2 AND2X2_1457 ( .A(_2041_), .B(_2040_), .Y(_2042_) );
AND2X2 AND2X2_1458 ( .A(_2042_), .B(_1721__bF_buf0), .Y(_2043_) );
OR2X2 OR2X2_1210 ( .A(_2043_), .B(_2039_), .Y(_2044_) );
OR2X2 OR2X2_1211 ( .A(_2035_), .B(_2044_), .Y(_2045_) );
OR2X2 OR2X2_1212 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_0__6_), .Y(_2046_) );
OR2X2 OR2X2_1213 ( .A(REGs_FIRQ_REGS_0__6_), .B(_1568__bF_buf14), .Y(_2047_) );
AND2X2 AND2X2_1459 ( .A(_2047_), .B(_2046_), .Y(_2048_) );
AND2X2 AND2X2_1460 ( .A(_1730__bF_buf3), .B(_2048_), .Y(_2049_) );
OR2X2 OR2X2_1214 ( .A(INTERRUPT_flag_bF_buf13), .B(REGs_USR_REGS_1__6_), .Y(_2050_) );
OR2X2 OR2X2_1215 ( .A(REGs_FIRQ_REGS_1__6_), .B(_1568__bF_buf11), .Y(_2051_) );
AND2X2 AND2X2_1461 ( .A(_2051_), .B(_2050_), .Y(_2052_) );
AND2X2 AND2X2_1462 ( .A(_1735__bF_buf1), .B(_2052_), .Y(_2053_) );
OR2X2 OR2X2_1216 ( .A(_2049_), .B(_2053_), .Y(_2054_) );
OR2X2 OR2X2_1217 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_3__6_), .Y(_2055_) );
OR2X2 OR2X2_1218 ( .A(REGs_FIRQ_REGS_3__6_), .B(_1568__bF_buf11), .Y(_2056_) );
AND2X2 AND2X2_1463 ( .A(_2056_), .B(_2055_), .Y(_2057_) );
AND2X2 AND2X2_1464 ( .A(_2057_), .B(_1741__bF_buf3), .Y(_2058_) );
OR2X2 OR2X2_1219 ( .A(INTERRUPT_flag_bF_buf15_bF_buf2), .B(REGs_USR_REGS_2__6_), .Y(_2059_) );
OR2X2 OR2X2_1220 ( .A(REGs_FIRQ_REGS_2__6_), .B(_1568__bF_buf9), .Y(_2060_) );
AND2X2 AND2X2_1465 ( .A(_2060_), .B(_2059_), .Y(_2061_) );
AND2X2 AND2X2_1466 ( .A(_1746__bF_buf1), .B(_2061_), .Y(_2062_) );
OR2X2 OR2X2_1221 ( .A(_2058_), .B(_2062_), .Y(_2063_) );
OR2X2 OR2X2_1222 ( .A(_2063_), .B(_2054_), .Y(_2064_) );
OR2X2 OR2X2_1223 ( .A(_2045_), .B(_2064_), .Y(_2065_) );
OR2X2 OR2X2_1224 ( .A(_2026_), .B(_2065_), .Y(REG_B_6_) );
AND2X2 AND2X2_1467 ( .A(_1678__bF_buf0), .B(REGs_REGS_4__7_), .Y(_2066_) );
AND2X2 AND2X2_1468 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__7_), .Y(_2067_) );
OR2X2 OR2X2_1225 ( .A(_2066_), .B(_2067_), .Y(_2068_) );
AND2X2 AND2X2_1469 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__7_), .Y(_2069_) );
AND2X2 AND2X2_1470 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__7_), .Y(_2070_) );
OR2X2 OR2X2_1226 ( .A(_2070_), .B(_2069_), .Y(_2071_) );
OR2X2 OR2X2_1227 ( .A(_2068_), .B(_2071_), .Y(_2072_) );
AND2X2 AND2X2_1471 ( .A(_1695__bF_buf2), .B(PC_ADDR_stack_1__7_), .Y(_2073_) );
AND2X2 AND2X2_1472 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__7_), .Y(_2074_) );
AND2X2 AND2X2_1473 ( .A(_1699__bF_buf2), .B(REGs_REGS_2__7_), .Y(_2075_) );
OR2X2 OR2X2_1228 ( .A(_2074_), .B(_2075_), .Y(_2076_) );
OR2X2 OR2X2_1229 ( .A(_2073_), .B(_2076_), .Y(_2077_) );
OR2X2 OR2X2_1230 ( .A(_2077_), .B(_2072_), .Y(_2078_) );
OR2X2 OR2X2_1231 ( .A(INTERRUPT_flag_bF_buf14_bF_buf3), .B(REGs_USR_REGS_5__7_), .Y(_2079_) );
OR2X2 OR2X2_1232 ( .A(REGs_FIRQ_REGS_5__7_), .B(_1568__bF_buf0), .Y(_2080_) );
AND2X2 AND2X2_1474 ( .A(_2080_), .B(_2079_), .Y(_2081_) );
AND2X2 AND2X2_1475 ( .A(_2081_), .B(_1705__bF_buf3), .Y(_2082_) );
OR2X2 OR2X2_1233 ( .A(INTERRUPT_flag_bF_buf13_bF_buf3), .B(REGs_USR_REGS_4__7_), .Y(_2083_) );
OR2X2 OR2X2_1234 ( .A(REGs_FIRQ_REGS_4__7_), .B(_1568__bF_buf2), .Y(_2084_) );
AND2X2 AND2X2_1476 ( .A(_2084_), .B(_2083_), .Y(_2085_) );
AND2X2 AND2X2_1477 ( .A(_2085_), .B(_1710__bF_buf4), .Y(_2086_) );
OR2X2 OR2X2_1235 ( .A(_2086_), .B(_2082_), .Y(_2087_) );
OR2X2 OR2X2_1236 ( .A(INTERRUPT_flag_bF_buf12_bF_buf2), .B(REGs_USR_REGS_6__7_), .Y(_2088_) );
OR2X2 OR2X2_1237 ( .A(REGs_FIRQ_REGS_6__7_), .B(_1568__bF_buf1), .Y(_2089_) );
AND2X2 AND2X2_1478 ( .A(_2089_), .B(_2088_), .Y(_2090_) );
AND2X2 AND2X2_1479 ( .A(_2090_), .B(_1716__bF_buf3), .Y(_2091_) );
OR2X2 OR2X2_1238 ( .A(INTERRUPT_flag_bF_buf11_bF_buf3), .B(REGs_USR_REGS_7__7_), .Y(_2092_) );
OR2X2 OR2X2_1239 ( .A(REGs_FIRQ_REGS_7__7_), .B(_1568__bF_buf2), .Y(_2093_) );
AND2X2 AND2X2_1480 ( .A(_2093_), .B(_2092_), .Y(_2094_) );
AND2X2 AND2X2_1481 ( .A(_2094_), .B(_1721__bF_buf3), .Y(_2095_) );
OR2X2 OR2X2_1240 ( .A(_2095_), .B(_2091_), .Y(_2096_) );
OR2X2 OR2X2_1241 ( .A(_2087_), .B(_2096_), .Y(_2097_) );
OR2X2 OR2X2_1242 ( .A(INTERRUPT_flag_bF_buf10_bF_buf2), .B(REGs_USR_REGS_0__7_), .Y(_2098_) );
OR2X2 OR2X2_1243 ( .A(REGs_FIRQ_REGS_0__7_), .B(_1568__bF_buf9), .Y(_2099_) );
AND2X2 AND2X2_1482 ( .A(_2099_), .B(_2098_), .Y(_2100_) );
AND2X2 AND2X2_1483 ( .A(_1730__bF_buf4), .B(_2100_), .Y(_2101_) );
OR2X2 OR2X2_1244 ( .A(INTERRUPT_flag_bF_buf9_bF_buf1), .B(REGs_USR_REGS_1__7_), .Y(_2102_) );
OR2X2 OR2X2_1245 ( .A(REGs_FIRQ_REGS_1__7_), .B(_1568__bF_buf2), .Y(_2103_) );
AND2X2 AND2X2_1484 ( .A(_2103_), .B(_2102_), .Y(_2104_) );
AND2X2 AND2X2_1485 ( .A(_1735__bF_buf4), .B(_2104_), .Y(_2105_) );
OR2X2 OR2X2_1246 ( .A(_2101_), .B(_2105_), .Y(_2106_) );
OR2X2 OR2X2_1247 ( .A(INTERRUPT_flag_bF_buf8_bF_buf3), .B(REGs_USR_REGS_3__7_), .Y(_2107_) );
OR2X2 OR2X2_1248 ( .A(REGs_FIRQ_REGS_3__7_), .B(_1568__bF_buf2), .Y(_2108_) );
AND2X2 AND2X2_1486 ( .A(_2108_), .B(_2107_), .Y(_2109_) );
AND2X2 AND2X2_1487 ( .A(_2109_), .B(_1741__bF_buf0), .Y(_2110_) );
OR2X2 OR2X2_1249 ( .A(INTERRUPT_flag_bF_buf7_bF_buf3), .B(REGs_USR_REGS_2__7_), .Y(_2111_) );
OR2X2 OR2X2_1250 ( .A(REGs_FIRQ_REGS_2__7_), .B(_1568__bF_buf15_bF_buf3), .Y(_2112_) );
AND2X2 AND2X2_1488 ( .A(_2112_), .B(_2111_), .Y(_2113_) );
AND2X2 AND2X2_1489 ( .A(_1746__bF_buf3), .B(_2113_), .Y(_2114_) );
OR2X2 OR2X2_1251 ( .A(_2110_), .B(_2114_), .Y(_2115_) );
OR2X2 OR2X2_1252 ( .A(_2115_), .B(_2106_), .Y(_2116_) );
OR2X2 OR2X2_1253 ( .A(_2097_), .B(_2116_), .Y(_2117_) );
OR2X2 OR2X2_1254 ( .A(_2078_), .B(_2117_), .Y(REG_B_7_) );
AND2X2 AND2X2_1490 ( .A(_1678__bF_buf1), .B(REGs_REGS_4__8_), .Y(_2118_) );
AND2X2 AND2X2_1491 ( .A(_1682__bF_buf0), .B(REGs_REGS_5__8_), .Y(_2119_) );
OR2X2 OR2X2_1255 ( .A(_2118_), .B(_2119_), .Y(_2120_) );
AND2X2 AND2X2_1492 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__8_), .Y(_2121_) );
AND2X2 AND2X2_1493 ( .A(_1690__bF_buf1), .B(REGs_REGS_7__8_), .Y(_2122_) );
OR2X2 OR2X2_1256 ( .A(_2122_), .B(_2121_), .Y(_2123_) );
OR2X2 OR2X2_1257 ( .A(_2120_), .B(_2123_), .Y(_2124_) );
AND2X2 AND2X2_1494 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2125_) );
AND2X2 AND2X2_1495 ( .A(_1697__bF_buf2), .B(REGs_REGS_3__8_), .Y(_2126_) );
AND2X2 AND2X2_1496 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__8_), .Y(_2127_) );
OR2X2 OR2X2_1258 ( .A(_2126_), .B(_2127_), .Y(_2128_) );
OR2X2 OR2X2_1259 ( .A(_2125_), .B(_2128_), .Y(_2129_) );
OR2X2 OR2X2_1260 ( .A(_2129_), .B(_2124_), .Y(_2130_) );
OR2X2 OR2X2_1261 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_5__8_), .Y(_2131_) );
OR2X2 OR2X2_1262 ( .A(REGs_FIRQ_REGS_5__8_), .B(_1568__bF_buf7), .Y(_2132_) );
AND2X2 AND2X2_1497 ( .A(_2132_), .B(_2131_), .Y(_2133_) );
AND2X2 AND2X2_1498 ( .A(_2133_), .B(_1705__bF_buf0), .Y(_2134_) );
OR2X2 OR2X2_1263 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_4__8_), .Y(_2135_) );
OR2X2 OR2X2_1264 ( .A(REGs_FIRQ_REGS_4__8_), .B(_1568__bF_buf10), .Y(_2136_) );
AND2X2 AND2X2_1499 ( .A(_2136_), .B(_2135_), .Y(_2137_) );
AND2X2 AND2X2_1500 ( .A(_2137_), .B(_1710__bF_buf2), .Y(_2138_) );
OR2X2 OR2X2_1265 ( .A(_2138_), .B(_2134_), .Y(_2139_) );
OR2X2 OR2X2_1266 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_6__8_), .Y(_2140_) );
OR2X2 OR2X2_1267 ( .A(REGs_FIRQ_REGS_6__8_), .B(_1568__bF_buf10), .Y(_2141_) );
AND2X2 AND2X2_1501 ( .A(_2141_), .B(_2140_), .Y(_2142_) );
AND2X2 AND2X2_1502 ( .A(_2142_), .B(_1716__bF_buf0), .Y(_2143_) );
OR2X2 OR2X2_1268 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_7__8_), .Y(_2144_) );
OR2X2 OR2X2_1269 ( .A(REGs_FIRQ_REGS_7__8_), .B(_1568__bF_buf3), .Y(_2145_) );
AND2X2 AND2X2_1503 ( .A(_2145_), .B(_2144_), .Y(_2146_) );
AND2X2 AND2X2_1504 ( .A(_2146_), .B(_1721__bF_buf2), .Y(_2147_) );
OR2X2 OR2X2_1270 ( .A(_2147_), .B(_2143_), .Y(_2148_) );
OR2X2 OR2X2_1271 ( .A(_2139_), .B(_2148_), .Y(_2149_) );
OR2X2 OR2X2_1272 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_0__8_), .Y(_2150_) );
OR2X2 OR2X2_1273 ( .A(REGs_FIRQ_REGS_0__8_), .B(_1568__bF_buf4), .Y(_2151_) );
AND2X2 AND2X2_1505 ( .A(_2151_), .B(_2150_), .Y(_2152_) );
AND2X2 AND2X2_1506 ( .A(_1730__bF_buf2), .B(_2152_), .Y(_2153_) );
OR2X2 OR2X2_1274 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_1__8_), .Y(_2154_) );
OR2X2 OR2X2_1275 ( .A(REGs_FIRQ_REGS_1__8_), .B(_1568__bF_buf13), .Y(_2155_) );
AND2X2 AND2X2_1507 ( .A(_2155_), .B(_2154_), .Y(_2156_) );
AND2X2 AND2X2_1508 ( .A(_1735__bF_buf2), .B(_2156_), .Y(_2157_) );
OR2X2 OR2X2_1276 ( .A(_2153_), .B(_2157_), .Y(_2158_) );
OR2X2 OR2X2_1277 ( .A(INTERRUPT_flag_bF_buf12), .B(REGs_USR_REGS_3__8_), .Y(_2159_) );
OR2X2 OR2X2_1278 ( .A(REGs_FIRQ_REGS_3__8_), .B(_1568__bF_buf7), .Y(_2160_) );
AND2X2 AND2X2_1509 ( .A(_2160_), .B(_2159_), .Y(_2161_) );
AND2X2 AND2X2_1510 ( .A(_2161_), .B(_1741__bF_buf4), .Y(_2162_) );
OR2X2 OR2X2_1279 ( .A(INTERRUPT_flag_bF_buf15_bF_buf3), .B(REGs_USR_REGS_2__8_), .Y(_2163_) );
OR2X2 OR2X2_1280 ( .A(REGs_FIRQ_REGS_2__8_), .B(_1568__bF_buf6), .Y(_2164_) );
AND2X2 AND2X2_1511 ( .A(_2164_), .B(_2163_), .Y(_2165_) );
AND2X2 AND2X2_1512 ( .A(_1746__bF_buf4), .B(_2165_), .Y(_2166_) );
OR2X2 OR2X2_1281 ( .A(_2162_), .B(_2166_), .Y(_2167_) );
OR2X2 OR2X2_1282 ( .A(_2167_), .B(_2158_), .Y(_2168_) );
OR2X2 OR2X2_1283 ( .A(_2149_), .B(_2168_), .Y(_2169_) );
OR2X2 OR2X2_1284 ( .A(_2130_), .B(_2169_), .Y(REG_B_8_) );
AND2X2 AND2X2_1513 ( .A(_1678__bF_buf2), .B(REGs_REGS_4__9_), .Y(_2170_) );
AND2X2 AND2X2_1514 ( .A(_1682__bF_buf1), .B(REGs_REGS_5__9_), .Y(_2171_) );
OR2X2 OR2X2_1285 ( .A(_2170_), .B(_2171_), .Y(_2172_) );
AND2X2 AND2X2_1515 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__9_), .Y(_2173_) );
AND2X2 AND2X2_1516 ( .A(_1690__bF_buf0), .B(REGs_REGS_7__9_), .Y(_2174_) );
OR2X2 OR2X2_1286 ( .A(_2174_), .B(_2173_), .Y(_2175_) );
OR2X2 OR2X2_1287 ( .A(_2172_), .B(_2175_), .Y(_2176_) );
AND2X2 AND2X2_1517 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2177_) );
AND2X2 AND2X2_1518 ( .A(_1697__bF_buf1), .B(REGs_REGS_3__9_), .Y(_2178_) );
AND2X2 AND2X2_1519 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__9_), .Y(_2179_) );
OR2X2 OR2X2_1288 ( .A(_2178_), .B(_2179_), .Y(_2180_) );
OR2X2 OR2X2_1289 ( .A(_2177_), .B(_2180_), .Y(_2181_) );
OR2X2 OR2X2_1290 ( .A(_2181_), .B(_2176_), .Y(_2182_) );
OR2X2 OR2X2_1291 ( .A(INTERRUPT_flag_bF_buf14_bF_buf0), .B(REGs_USR_REGS_5__9_), .Y(_2183_) );
OR2X2 OR2X2_1292 ( .A(REGs_FIRQ_REGS_5__9_), .B(_1568__bF_buf12), .Y(_2184_) );
AND2X2 AND2X2_1520 ( .A(_2184_), .B(_2183_), .Y(_2185_) );
AND2X2 AND2X2_1521 ( .A(_2185_), .B(_1705__bF_buf1), .Y(_2186_) );
OR2X2 OR2X2_1293 ( .A(INTERRUPT_flag_bF_buf13_bF_buf1), .B(REGs_USR_REGS_4__9_), .Y(_2187_) );
OR2X2 OR2X2_1294 ( .A(REGs_FIRQ_REGS_4__9_), .B(_1568__bF_buf5), .Y(_2188_) );
AND2X2 AND2X2_1522 ( .A(_2188_), .B(_2187_), .Y(_2189_) );
AND2X2 AND2X2_1523 ( .A(_2189_), .B(_1710__bF_buf0), .Y(_2190_) );
OR2X2 OR2X2_1295 ( .A(_2190_), .B(_2186_), .Y(_2191_) );
OR2X2 OR2X2_1296 ( .A(INTERRUPT_flag_bF_buf12_bF_buf1), .B(REGs_USR_REGS_6__9_), .Y(_2192_) );
OR2X2 OR2X2_1297 ( .A(REGs_FIRQ_REGS_6__9_), .B(_1568__bF_buf8), .Y(_2193_) );
AND2X2 AND2X2_1524 ( .A(_2193_), .B(_2192_), .Y(_2194_) );
AND2X2 AND2X2_1525 ( .A(_2194_), .B(_1716__bF_buf2), .Y(_2195_) );
OR2X2 OR2X2_1298 ( .A(INTERRUPT_flag_bF_buf11_bF_buf0), .B(REGs_USR_REGS_7__9_), .Y(_2196_) );
OR2X2 OR2X2_1299 ( .A(REGs_FIRQ_REGS_7__9_), .B(_1568__bF_buf8), .Y(_2197_) );
AND2X2 AND2X2_1526 ( .A(_2197_), .B(_2196_), .Y(_2198_) );
AND2X2 AND2X2_1527 ( .A(_2198_), .B(_1721__bF_buf4), .Y(_2199_) );
OR2X2 OR2X2_1300 ( .A(_2199_), .B(_2195_), .Y(_2200_) );
OR2X2 OR2X2_1301 ( .A(_2191_), .B(_2200_), .Y(_2201_) );
OR2X2 OR2X2_1302 ( .A(INTERRUPT_flag_bF_buf10_bF_buf0), .B(REGs_USR_REGS_0__9_), .Y(_2202_) );
OR2X2 OR2X2_1303 ( .A(REGs_FIRQ_REGS_0__9_), .B(_1568__bF_buf7), .Y(_2203_) );
AND2X2 AND2X2_1528 ( .A(_2203_), .B(_2202_), .Y(_2204_) );
AND2X2 AND2X2_1529 ( .A(_1730__bF_buf1), .B(_2204_), .Y(_2205_) );
OR2X2 OR2X2_1304 ( .A(INTERRUPT_flag_bF_buf9_bF_buf3), .B(REGs_USR_REGS_1__9_), .Y(_2206_) );
OR2X2 OR2X2_1305 ( .A(REGs_FIRQ_REGS_1__9_), .B(_1568__bF_buf3), .Y(_2207_) );
AND2X2 AND2X2_1530 ( .A(_2207_), .B(_2206_), .Y(_2208_) );
AND2X2 AND2X2_1531 ( .A(_1735__bF_buf3), .B(_2208_), .Y(_2209_) );
OR2X2 OR2X2_1306 ( .A(_2205_), .B(_2209_), .Y(_2210_) );
OR2X2 OR2X2_1307 ( .A(INTERRUPT_flag_bF_buf8_bF_buf1), .B(REGs_USR_REGS_3__9_), .Y(_2211_) );
OR2X2 OR2X2_1308 ( .A(REGs_FIRQ_REGS_3__9_), .B(_1568__bF_buf7), .Y(_2212_) );
AND2X2 AND2X2_1532 ( .A(_2212_), .B(_2211_), .Y(_2213_) );
AND2X2 AND2X2_1533 ( .A(_2213_), .B(_1741__bF_buf4), .Y(_2214_) );
OR2X2 OR2X2_1309 ( .A(INTERRUPT_flag_bF_buf7_bF_buf1), .B(REGs_USR_REGS_2__9_), .Y(_2215_) );
OR2X2 OR2X2_1310 ( .A(REGs_FIRQ_REGS_2__9_), .B(_1568__bF_buf15_bF_buf0), .Y(_2216_) );
AND2X2 AND2X2_1534 ( .A(_2216_), .B(_2215_), .Y(_2217_) );
AND2X2 AND2X2_1535 ( .A(_1746__bF_buf4), .B(_2217_), .Y(_2218_) );
OR2X2 OR2X2_1311 ( .A(_2214_), .B(_2218_), .Y(_2219_) );
OR2X2 OR2X2_1312 ( .A(_2219_), .B(_2210_), .Y(_2220_) );
OR2X2 OR2X2_1313 ( .A(_2201_), .B(_2220_), .Y(_2221_) );
OR2X2 OR2X2_1314 ( .A(_2182_), .B(_2221_), .Y(REG_B_9_) );
AND2X2 AND2X2_1536 ( .A(_1678__bF_buf2), .B(REGs_REGS_4__10_), .Y(_2222_) );
AND2X2 AND2X2_1537 ( .A(_1682__bF_buf1), .B(REGs_REGS_5__10_), .Y(_2223_) );
OR2X2 OR2X2_1315 ( .A(_2222_), .B(_2223_), .Y(_2224_) );
AND2X2 AND2X2_1538 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__10_), .Y(_2225_) );
AND2X2 AND2X2_1539 ( .A(_1690__bF_buf0), .B(REGs_REGS_7__10_), .Y(_2226_) );
OR2X2 OR2X2_1316 ( .A(_2226_), .B(_2225_), .Y(_2227_) );
OR2X2 OR2X2_1317 ( .A(_2224_), .B(_2227_), .Y(_2228_) );
AND2X2 AND2X2_1540 ( .A(_1695__bF_buf1), .B(gnd), .Y(_2229_) );
AND2X2 AND2X2_1541 ( .A(_1697__bF_buf1), .B(REGs_REGS_3__10_), .Y(_2230_) );
AND2X2 AND2X2_1542 ( .A(_1699__bF_buf1), .B(REGs_REGS_2__10_), .Y(_2231_) );
OR2X2 OR2X2_1318 ( .A(_2230_), .B(_2231_), .Y(_2232_) );
OR2X2 OR2X2_1319 ( .A(_2229_), .B(_2232_), .Y(_2233_) );
OR2X2 OR2X2_1320 ( .A(_2233_), .B(_2228_), .Y(_2234_) );
OR2X2 OR2X2_1321 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_5__10_), .Y(_2235_) );
OR2X2 OR2X2_1322 ( .A(REGs_FIRQ_REGS_5__10_), .B(_1568__bF_buf12), .Y(_2236_) );
AND2X2 AND2X2_1543 ( .A(_2236_), .B(_2235_), .Y(_2237_) );
AND2X2 AND2X2_1544 ( .A(_2237_), .B(_1705__bF_buf1), .Y(_2238_) );
OR2X2 OR2X2_1323 ( .A(INTERRUPT_flag_bF_buf9), .B(REGs_USR_REGS_4__10_), .Y(_2239_) );
OR2X2 OR2X2_1324 ( .A(REGs_FIRQ_REGS_4__10_), .B(_1568__bF_buf8), .Y(_2240_) );
AND2X2 AND2X2_1545 ( .A(_2240_), .B(_2239_), .Y(_2241_) );
AND2X2 AND2X2_1546 ( .A(_2241_), .B(_1710__bF_buf0), .Y(_2242_) );
OR2X2 OR2X2_1325 ( .A(_2242_), .B(_2238_), .Y(_2243_) );
OR2X2 OR2X2_1326 ( .A(INTERRUPT_flag_bF_buf8), .B(REGs_USR_REGS_6__10_), .Y(_2244_) );
OR2X2 OR2X2_1327 ( .A(REGs_FIRQ_REGS_6__10_), .B(_1568__bF_buf8), .Y(_2245_) );
AND2X2 AND2X2_1547 ( .A(_2245_), .B(_2244_), .Y(_2246_) );
AND2X2 AND2X2_1548 ( .A(_2246_), .B(_1716__bF_buf2), .Y(_2247_) );
OR2X2 OR2X2_1328 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_7__10_), .Y(_2248_) );
OR2X2 OR2X2_1329 ( .A(REGs_FIRQ_REGS_7__10_), .B(_1568__bF_buf5), .Y(_2249_) );
AND2X2 AND2X2_1549 ( .A(_2249_), .B(_2248_), .Y(_2250_) );
AND2X2 AND2X2_1550 ( .A(_2250_), .B(_1721__bF_buf4), .Y(_2251_) );
OR2X2 OR2X2_1330 ( .A(_2251_), .B(_2247_), .Y(_2252_) );
OR2X2 OR2X2_1331 ( .A(_2243_), .B(_2252_), .Y(_2253_) );
OR2X2 OR2X2_1332 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_0__10_), .Y(_2254_) );
OR2X2 OR2X2_1333 ( .A(REGs_FIRQ_REGS_0__10_), .B(_1568__bF_buf10), .Y(_2255_) );
AND2X2 AND2X2_1551 ( .A(_2255_), .B(_2254_), .Y(_2256_) );
AND2X2 AND2X2_1552 ( .A(_1730__bF_buf1), .B(_2256_), .Y(_2257_) );
OR2X2 OR2X2_1334 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_1__10_), .Y(_2258_) );
OR2X2 OR2X2_1335 ( .A(REGs_FIRQ_REGS_1__10_), .B(_1568__bF_buf10), .Y(_2259_) );
AND2X2 AND2X2_1553 ( .A(_2259_), .B(_2258_), .Y(_2260_) );
AND2X2 AND2X2_1554 ( .A(_1735__bF_buf3), .B(_2260_), .Y(_2261_) );
OR2X2 OR2X2_1336 ( .A(_2257_), .B(_2261_), .Y(_2262_) );
OR2X2 OR2X2_1337 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_3__10_), .Y(_2263_) );
OR2X2 OR2X2_1338 ( .A(REGs_FIRQ_REGS_3__10_), .B(_1568__bF_buf7), .Y(_2264_) );
AND2X2 AND2X2_1555 ( .A(_2264_), .B(_2263_), .Y(_2265_) );
AND2X2 AND2X2_1556 ( .A(_2265_), .B(_1741__bF_buf2), .Y(_2266_) );
OR2X2 OR2X2_1339 ( .A(INTERRUPT_flag_bF_buf15_bF_buf0), .B(REGs_USR_REGS_2__10_), .Y(_2267_) );
OR2X2 OR2X2_1340 ( .A(REGs_FIRQ_REGS_2__10_), .B(_1568__bF_buf10), .Y(_2268_) );
AND2X2 AND2X2_1557 ( .A(_2268_), .B(_2267_), .Y(_2269_) );
AND2X2 AND2X2_1558 ( .A(_1746__bF_buf2), .B(_2269_), .Y(_2270_) );
OR2X2 OR2X2_1341 ( .A(_2266_), .B(_2270_), .Y(_2271_) );
OR2X2 OR2X2_1342 ( .A(_2271_), .B(_2262_), .Y(_2272_) );
OR2X2 OR2X2_1343 ( .A(_2253_), .B(_2272_), .Y(_2273_) );
OR2X2 OR2X2_1344 ( .A(_2234_), .B(_2273_), .Y(REG_B_10_) );
AND2X2 AND2X2_1559 ( .A(_1678__bF_buf1), .B(REGs_REGS_4__11_), .Y(_2274_) );
AND2X2 AND2X2_1560 ( .A(_1682__bF_buf0), .B(REGs_REGS_5__11_), .Y(_2275_) );
OR2X2 OR2X2_1345 ( .A(_2274_), .B(_2275_), .Y(_2276_) );
AND2X2 AND2X2_1561 ( .A(_1687__bF_buf0), .B(REGs_REGS_6__11_), .Y(_2277_) );
AND2X2 AND2X2_1562 ( .A(_1690__bF_buf1), .B(REGs_REGS_7__11_), .Y(_2278_) );
OR2X2 OR2X2_1346 ( .A(_2278_), .B(_2277_), .Y(_2279_) );
OR2X2 OR2X2_1347 ( .A(_2276_), .B(_2279_), .Y(_2280_) );
AND2X2 AND2X2_1563 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2281_) );
AND2X2 AND2X2_1564 ( .A(_1697__bF_buf2), .B(REGs_REGS_3__11_), .Y(_2282_) );
AND2X2 AND2X2_1565 ( .A(_1699__bF_buf1), .B(REGs_REGS_2__11_), .Y(_2283_) );
OR2X2 OR2X2_1348 ( .A(_2282_), .B(_2283_), .Y(_2284_) );
OR2X2 OR2X2_1349 ( .A(_2281_), .B(_2284_), .Y(_2285_) );
OR2X2 OR2X2_1350 ( .A(_2285_), .B(_2280_), .Y(_2286_) );
OR2X2 OR2X2_1351 ( .A(INTERRUPT_flag_bF_buf14_bF_buf0), .B(REGs_USR_REGS_5__11_), .Y(_2287_) );
OR2X2 OR2X2_1352 ( .A(REGs_FIRQ_REGS_5__11_), .B(_1568__bF_buf5), .Y(_2288_) );
AND2X2 AND2X2_1566 ( .A(_2288_), .B(_2287_), .Y(_2289_) );
AND2X2 AND2X2_1567 ( .A(_2289_), .B(_1705__bF_buf2), .Y(_2290_) );
OR2X2 OR2X2_1353 ( .A(INTERRUPT_flag_bF_buf13_bF_buf2), .B(REGs_USR_REGS_4__11_), .Y(_2291_) );
OR2X2 OR2X2_1354 ( .A(REGs_FIRQ_REGS_4__11_), .B(_1568__bF_buf12), .Y(_2292_) );
AND2X2 AND2X2_1568 ( .A(_2292_), .B(_2291_), .Y(_2293_) );
AND2X2 AND2X2_1569 ( .A(_2293_), .B(_1710__bF_buf1), .Y(_2294_) );
OR2X2 OR2X2_1355 ( .A(_2294_), .B(_2290_), .Y(_2295_) );
OR2X2 OR2X2_1356 ( .A(INTERRUPT_flag_bF_buf12_bF_buf1), .B(REGs_USR_REGS_6__11_), .Y(_2296_) );
OR2X2 OR2X2_1357 ( .A(REGs_FIRQ_REGS_6__11_), .B(_1568__bF_buf12), .Y(_2297_) );
AND2X2 AND2X2_1570 ( .A(_2297_), .B(_2296_), .Y(_2298_) );
AND2X2 AND2X2_1571 ( .A(_2298_), .B(_1716__bF_buf1), .Y(_2299_) );
OR2X2 OR2X2_1358 ( .A(INTERRUPT_flag_bF_buf11_bF_buf2), .B(REGs_USR_REGS_7__11_), .Y(_2300_) );
OR2X2 OR2X2_1359 ( .A(REGs_FIRQ_REGS_7__11_), .B(_1568__bF_buf12), .Y(_2301_) );
AND2X2 AND2X2_1572 ( .A(_2301_), .B(_2300_), .Y(_2302_) );
AND2X2 AND2X2_1573 ( .A(_2302_), .B(_1721__bF_buf1), .Y(_2303_) );
OR2X2 OR2X2_1360 ( .A(_2303_), .B(_2299_), .Y(_2304_) );
OR2X2 OR2X2_1361 ( .A(_2295_), .B(_2304_), .Y(_2305_) );
OR2X2 OR2X2_1362 ( .A(INTERRUPT_flag_bF_buf10_bF_buf1), .B(REGs_USR_REGS_0__11_), .Y(_2306_) );
OR2X2 OR2X2_1363 ( .A(REGs_FIRQ_REGS_0__11_), .B(_1568__bF_buf13), .Y(_2307_) );
AND2X2 AND2X2_1574 ( .A(_2307_), .B(_2306_), .Y(_2308_) );
AND2X2 AND2X2_1575 ( .A(_1730__bF_buf0), .B(_2308_), .Y(_2309_) );
OR2X2 OR2X2_1364 ( .A(INTERRUPT_flag_bF_buf9_bF_buf2), .B(REGs_USR_REGS_1__11_), .Y(_2310_) );
OR2X2 OR2X2_1365 ( .A(REGs_FIRQ_REGS_1__11_), .B(_1568__bF_buf7), .Y(_2311_) );
AND2X2 AND2X2_1576 ( .A(_2311_), .B(_2310_), .Y(_2312_) );
AND2X2 AND2X2_1577 ( .A(_1735__bF_buf2), .B(_2312_), .Y(_2313_) );
OR2X2 OR2X2_1366 ( .A(_2309_), .B(_2313_), .Y(_2314_) );
OR2X2 OR2X2_1367 ( .A(INTERRUPT_flag_bF_buf8_bF_buf2), .B(REGs_USR_REGS_3__11_), .Y(_2315_) );
OR2X2 OR2X2_1368 ( .A(REGs_FIRQ_REGS_3__11_), .B(_1568__bF_buf7), .Y(_2316_) );
AND2X2 AND2X2_1578 ( .A(_2316_), .B(_2315_), .Y(_2317_) );
AND2X2 AND2X2_1579 ( .A(_2317_), .B(_1741__bF_buf4), .Y(_2318_) );
OR2X2 OR2X2_1369 ( .A(INTERRUPT_flag_bF_buf7_bF_buf2), .B(REGs_USR_REGS_2__11_), .Y(_2319_) );
OR2X2 OR2X2_1370 ( .A(REGs_FIRQ_REGS_2__11_), .B(_1568__bF_buf15_bF_buf2), .Y(_2320_) );
AND2X2 AND2X2_1580 ( .A(_2320_), .B(_2319_), .Y(_2321_) );
AND2X2 AND2X2_1581 ( .A(_1746__bF_buf0), .B(_2321_), .Y(_2322_) );
OR2X2 OR2X2_1371 ( .A(_2318_), .B(_2322_), .Y(_2323_) );
OR2X2 OR2X2_1372 ( .A(_2323_), .B(_2314_), .Y(_2324_) );
OR2X2 OR2X2_1373 ( .A(_2305_), .B(_2324_), .Y(_2325_) );
OR2X2 OR2X2_1374 ( .A(_2286_), .B(_2325_), .Y(REG_B_11_) );
AND2X2 AND2X2_1582 ( .A(_1678__bF_buf0), .B(REGs_REGS_4__12_), .Y(_2326_) );
AND2X2 AND2X2_1583 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__12_), .Y(_2327_) );
OR2X2 OR2X2_1375 ( .A(_2326_), .B(_2327_), .Y(_2328_) );
AND2X2 AND2X2_1584 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__12_), .Y(_2329_) );
AND2X2 AND2X2_1585 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__12_), .Y(_2330_) );
OR2X2 OR2X2_1376 ( .A(_2330_), .B(_2329_), .Y(_2331_) );
OR2X2 OR2X2_1377 ( .A(_2328_), .B(_2331_), .Y(_2332_) );
AND2X2 AND2X2_1586 ( .A(_1695__bF_buf2), .B(gnd), .Y(_2333_) );
AND2X2 AND2X2_1587 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__12_), .Y(_2334_) );
AND2X2 AND2X2_1588 ( .A(_1699__bF_buf2), .B(REGs_REGS_2__12_), .Y(_2335_) );
OR2X2 OR2X2_1378 ( .A(_2334_), .B(_2335_), .Y(_2336_) );
OR2X2 OR2X2_1379 ( .A(_2333_), .B(_2336_), .Y(_2337_) );
OR2X2 OR2X2_1380 ( .A(_2337_), .B(_2332_), .Y(_2338_) );
OR2X2 OR2X2_1381 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_5__12_), .Y(_2339_) );
OR2X2 OR2X2_1382 ( .A(REGs_FIRQ_REGS_5__12_), .B(_1568__bF_buf14), .Y(_2340_) );
AND2X2 AND2X2_1589 ( .A(_2340_), .B(_2339_), .Y(_2341_) );
AND2X2 AND2X2_1590 ( .A(_2341_), .B(_1705__bF_buf4), .Y(_2342_) );
OR2X2 OR2X2_1383 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_4__12_), .Y(_2343_) );
OR2X2 OR2X2_1384 ( .A(REGs_FIRQ_REGS_4__12_), .B(_1568__bF_buf14), .Y(_2344_) );
AND2X2 AND2X2_1591 ( .A(_2344_), .B(_2343_), .Y(_2345_) );
AND2X2 AND2X2_1592 ( .A(_2345_), .B(_1710__bF_buf3), .Y(_2346_) );
OR2X2 OR2X2_1385 ( .A(_2346_), .B(_2342_), .Y(_2347_) );
OR2X2 OR2X2_1386 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_6__12_), .Y(_2348_) );
OR2X2 OR2X2_1387 ( .A(REGs_FIRQ_REGS_6__12_), .B(_1568__bF_buf11), .Y(_2349_) );
AND2X2 AND2X2_1593 ( .A(_2349_), .B(_2348_), .Y(_2350_) );
AND2X2 AND2X2_1594 ( .A(_2350_), .B(_1716__bF_buf4), .Y(_2351_) );
OR2X2 OR2X2_1388 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_7__12_), .Y(_2352_) );
OR2X2 OR2X2_1389 ( .A(REGs_FIRQ_REGS_7__12_), .B(_1568__bF_buf14), .Y(_2353_) );
AND2X2 AND2X2_1595 ( .A(_2353_), .B(_2352_), .Y(_2354_) );
AND2X2 AND2X2_1596 ( .A(_2354_), .B(_1721__bF_buf0), .Y(_2355_) );
OR2X2 OR2X2_1390 ( .A(_2355_), .B(_2351_), .Y(_2356_) );
OR2X2 OR2X2_1391 ( .A(_2347_), .B(_2356_), .Y(_2357_) );
OR2X2 OR2X2_1392 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_0__12_), .Y(_2358_) );
OR2X2 OR2X2_1393 ( .A(REGs_FIRQ_REGS_0__12_), .B(_1568__bF_buf14), .Y(_2359_) );
AND2X2 AND2X2_1597 ( .A(_2359_), .B(_2358_), .Y(_2360_) );
AND2X2 AND2X2_1598 ( .A(_1730__bF_buf3), .B(_2360_), .Y(_2361_) );
OR2X2 OR2X2_1394 ( .A(INTERRUPT_flag_bF_buf10), .B(REGs_USR_REGS_1__12_), .Y(_2362_) );
OR2X2 OR2X2_1395 ( .A(REGs_FIRQ_REGS_1__12_), .B(_1568__bF_buf11), .Y(_2363_) );
AND2X2 AND2X2_1599 ( .A(_2363_), .B(_2362_), .Y(_2364_) );
AND2X2 AND2X2_1600 ( .A(_1735__bF_buf1), .B(_2364_), .Y(_2365_) );
OR2X2 OR2X2_1396 ( .A(_2361_), .B(_2365_), .Y(_2366_) );
OR2X2 OR2X2_1397 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_3__12_), .Y(_2367_) );
OR2X2 OR2X2_1398 ( .A(REGs_FIRQ_REGS_3__12_), .B(_1568__bF_buf11), .Y(_2368_) );
AND2X2 AND2X2_1601 ( .A(_2368_), .B(_2367_), .Y(_2369_) );
AND2X2 AND2X2_1602 ( .A(_2369_), .B(_1741__bF_buf3), .Y(_2370_) );
OR2X2 OR2X2_1399 ( .A(INTERRUPT_flag_bF_buf15_bF_buf1), .B(REGs_USR_REGS_2__12_), .Y(_2371_) );
OR2X2 OR2X2_1400 ( .A(REGs_FIRQ_REGS_2__12_), .B(_1568__bF_buf9), .Y(_2372_) );
AND2X2 AND2X2_1603 ( .A(_2372_), .B(_2371_), .Y(_2373_) );
AND2X2 AND2X2_1604 ( .A(_1746__bF_buf1), .B(_2373_), .Y(_2374_) );
OR2X2 OR2X2_1401 ( .A(_2370_), .B(_2374_), .Y(_2375_) );
OR2X2 OR2X2_1402 ( .A(_2375_), .B(_2366_), .Y(_2376_) );
OR2X2 OR2X2_1403 ( .A(_2357_), .B(_2376_), .Y(_2377_) );
OR2X2 OR2X2_1404 ( .A(_2338_), .B(_2377_), .Y(REG_B_12_) );
AND2X2 AND2X2_1605 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__13_), .Y(_2378_) );
AND2X2 AND2X2_1606 ( .A(_1682__bF_buf2), .B(REGs_REGS_5__13_), .Y(_2379_) );
OR2X2 OR2X2_1405 ( .A(_2378_), .B(_2379_), .Y(_2380_) );
AND2X2 AND2X2_1607 ( .A(_1687__bF_buf1), .B(REGs_REGS_6__13_), .Y(_2381_) );
AND2X2 AND2X2_1608 ( .A(_1690__bF_buf2), .B(REGs_REGS_7__13_), .Y(_2382_) );
OR2X2 OR2X2_1406 ( .A(_2382_), .B(_2381_), .Y(_2383_) );
OR2X2 OR2X2_1407 ( .A(_2380_), .B(_2383_), .Y(_2384_) );
AND2X2 AND2X2_1609 ( .A(_1695__bF_buf4), .B(gnd), .Y(_2385_) );
AND2X2 AND2X2_1610 ( .A(_1697__bF_buf0), .B(REGs_REGS_3__13_), .Y(_2386_) );
AND2X2 AND2X2_1611 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__13_), .Y(_2387_) );
OR2X2 OR2X2_1408 ( .A(_2386_), .B(_2387_), .Y(_2388_) );
OR2X2 OR2X2_1409 ( .A(_2385_), .B(_2388_), .Y(_2389_) );
OR2X2 OR2X2_1410 ( .A(_2389_), .B(_2384_), .Y(_2390_) );
OR2X2 OR2X2_1411 ( .A(INTERRUPT_flag_bF_buf14_bF_buf2), .B(REGs_USR_REGS_5__13_), .Y(_2391_) );
OR2X2 OR2X2_1412 ( .A(REGs_FIRQ_REGS_5__13_), .B(_1568__bF_buf13), .Y(_2392_) );
AND2X2 AND2X2_1612 ( .A(_2392_), .B(_2391_), .Y(_2393_) );
AND2X2 AND2X2_1613 ( .A(_2393_), .B(_1705__bF_buf0), .Y(_2394_) );
OR2X2 OR2X2_1413 ( .A(INTERRUPT_flag_bF_buf13_bF_buf3), .B(REGs_USR_REGS_4__13_), .Y(_2395_) );
OR2X2 OR2X2_1414 ( .A(REGs_FIRQ_REGS_4__13_), .B(_1568__bF_buf13), .Y(_2396_) );
AND2X2 AND2X2_1614 ( .A(_2396_), .B(_2395_), .Y(_2397_) );
AND2X2 AND2X2_1615 ( .A(_2397_), .B(_1710__bF_buf2), .Y(_2398_) );
OR2X2 OR2X2_1415 ( .A(_2398_), .B(_2394_), .Y(_2399_) );
OR2X2 OR2X2_1416 ( .A(INTERRUPT_flag_bF_buf12_bF_buf0), .B(REGs_USR_REGS_6__13_), .Y(_2400_) );
OR2X2 OR2X2_1417 ( .A(REGs_FIRQ_REGS_6__13_), .B(_1568__bF_buf4), .Y(_2401_) );
AND2X2 AND2X2_1616 ( .A(_2401_), .B(_2400_), .Y(_2402_) );
AND2X2 AND2X2_1617 ( .A(_2402_), .B(_1716__bF_buf0), .Y(_2403_) );
OR2X2 OR2X2_1418 ( .A(INTERRUPT_flag_bF_buf11_bF_buf3), .B(REGs_USR_REGS_7__13_), .Y(_2404_) );
OR2X2 OR2X2_1419 ( .A(REGs_FIRQ_REGS_7__13_), .B(_1568__bF_buf13), .Y(_2405_) );
AND2X2 AND2X2_1618 ( .A(_2405_), .B(_2404_), .Y(_2406_) );
AND2X2 AND2X2_1619 ( .A(_2406_), .B(_1721__bF_buf2), .Y(_2407_) );
OR2X2 OR2X2_1420 ( .A(_2407_), .B(_2403_), .Y(_2408_) );
OR2X2 OR2X2_1421 ( .A(_2399_), .B(_2408_), .Y(_2409_) );
OR2X2 OR2X2_1422 ( .A(INTERRUPT_flag_bF_buf10_bF_buf1), .B(REGs_USR_REGS_0__13_), .Y(_2410_) );
OR2X2 OR2X2_1423 ( .A(REGs_FIRQ_REGS_0__13_), .B(_1568__bF_buf4), .Y(_2411_) );
AND2X2 AND2X2_1620 ( .A(_2411_), .B(_2410_), .Y(_2412_) );
AND2X2 AND2X2_1621 ( .A(_1730__bF_buf4), .B(_2412_), .Y(_2413_) );
OR2X2 OR2X2_1424 ( .A(INTERRUPT_flag_bF_buf9_bF_buf0), .B(REGs_USR_REGS_1__13_), .Y(_2414_) );
OR2X2 OR2X2_1425 ( .A(REGs_FIRQ_REGS_1__13_), .B(_1568__bF_buf9), .Y(_2415_) );
AND2X2 AND2X2_1622 ( .A(_2415_), .B(_2414_), .Y(_2416_) );
AND2X2 AND2X2_1623 ( .A(_1735__bF_buf0), .B(_2416_), .Y(_2417_) );
OR2X2 OR2X2_1426 ( .A(_2413_), .B(_2417_), .Y(_2418_) );
OR2X2 OR2X2_1427 ( .A(INTERRUPT_flag_bF_buf8_bF_buf3), .B(REGs_USR_REGS_3__13_), .Y(_2419_) );
OR2X2 OR2X2_1428 ( .A(REGs_FIRQ_REGS_3__13_), .B(_1568__bF_buf2), .Y(_2420_) );
AND2X2 AND2X2_1624 ( .A(_2420_), .B(_2419_), .Y(_2421_) );
AND2X2 AND2X2_1625 ( .A(_2421_), .B(_1741__bF_buf0), .Y(_2422_) );
OR2X2 OR2X2_1429 ( .A(INTERRUPT_flag_bF_buf7_bF_buf3), .B(REGs_USR_REGS_2__13_), .Y(_2423_) );
OR2X2 OR2X2_1430 ( .A(REGs_FIRQ_REGS_2__13_), .B(_1568__bF_buf15_bF_buf3), .Y(_2424_) );
AND2X2 AND2X2_1626 ( .A(_2424_), .B(_2423_), .Y(_2425_) );
AND2X2 AND2X2_1627 ( .A(_1746__bF_buf3), .B(_2425_), .Y(_2426_) );
OR2X2 OR2X2_1431 ( .A(_2422_), .B(_2426_), .Y(_2427_) );
OR2X2 OR2X2_1432 ( .A(_2427_), .B(_2418_), .Y(_2428_) );
OR2X2 OR2X2_1433 ( .A(_2409_), .B(_2428_), .Y(_2429_) );
OR2X2 OR2X2_1434 ( .A(_2390_), .B(_2429_), .Y(REG_B_13_) );
AND2X2 AND2X2_1628 ( .A(_1678__bF_buf2), .B(REGs_REGS_4__14_), .Y(_2430_) );
AND2X2 AND2X2_1629 ( .A(_1682__bF_buf1), .B(REGs_REGS_5__14_), .Y(_2431_) );
OR2X2 OR2X2_1435 ( .A(_2430_), .B(_2431_), .Y(_2432_) );
AND2X2 AND2X2_1630 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__14_), .Y(_2433_) );
AND2X2 AND2X2_1631 ( .A(_1690__bF_buf0), .B(REGs_REGS_7__14_), .Y(_2434_) );
OR2X2 OR2X2_1436 ( .A(_2434_), .B(_2433_), .Y(_2435_) );
OR2X2 OR2X2_1437 ( .A(_2432_), .B(_2435_), .Y(_2436_) );
AND2X2 AND2X2_1632 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2437_) );
AND2X2 AND2X2_1633 ( .A(_1697__bF_buf1), .B(REGs_REGS_3__14_), .Y(_2438_) );
AND2X2 AND2X2_1634 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__14_), .Y(_2439_) );
OR2X2 OR2X2_1438 ( .A(_2438_), .B(_2439_), .Y(_2440_) );
OR2X2 OR2X2_1439 ( .A(_2437_), .B(_2440_), .Y(_2441_) );
OR2X2 OR2X2_1440 ( .A(_2441_), .B(_2436_), .Y(_2442_) );
OR2X2 OR2X2_1441 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_5__14_), .Y(_2443_) );
OR2X2 OR2X2_1442 ( .A(REGs_FIRQ_REGS_5__14_), .B(_1568__bF_buf5), .Y(_2444_) );
AND2X2 AND2X2_1635 ( .A(_2444_), .B(_2443_), .Y(_2445_) );
AND2X2 AND2X2_1636 ( .A(_2445_), .B(_1705__bF_buf1), .Y(_2446_) );
OR2X2 OR2X2_1443 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_4__14_), .Y(_2447_) );
OR2X2 OR2X2_1444 ( .A(REGs_FIRQ_REGS_4__14_), .B(_1568__bF_buf5), .Y(_2448_) );
AND2X2 AND2X2_1637 ( .A(_2448_), .B(_2447_), .Y(_2449_) );
AND2X2 AND2X2_1638 ( .A(_2449_), .B(_1710__bF_buf0), .Y(_2450_) );
OR2X2 OR2X2_1445 ( .A(_2450_), .B(_2446_), .Y(_2451_) );
OR2X2 OR2X2_1446 ( .A(INTERRUPT_flag_bF_buf8), .B(REGs_USR_REGS_6__14_), .Y(_2452_) );
OR2X2 OR2X2_1447 ( .A(REGs_FIRQ_REGS_6__14_), .B(_1568__bF_buf8), .Y(_2453_) );
AND2X2 AND2X2_1639 ( .A(_2453_), .B(_2452_), .Y(_2454_) );
AND2X2 AND2X2_1640 ( .A(_2454_), .B(_1716__bF_buf2), .Y(_2455_) );
OR2X2 OR2X2_1448 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_7__14_), .Y(_2456_) );
OR2X2 OR2X2_1449 ( .A(REGs_FIRQ_REGS_7__14_), .B(_1568__bF_buf5), .Y(_2457_) );
AND2X2 AND2X2_1641 ( .A(_2457_), .B(_2456_), .Y(_2458_) );
AND2X2 AND2X2_1642 ( .A(_2458_), .B(_1721__bF_buf4), .Y(_2459_) );
OR2X2 OR2X2_1450 ( .A(_2459_), .B(_2455_), .Y(_2460_) );
OR2X2 OR2X2_1451 ( .A(_2451_), .B(_2460_), .Y(_2461_) );
OR2X2 OR2X2_1452 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_0__14_), .Y(_2462_) );
OR2X2 OR2X2_1453 ( .A(REGs_FIRQ_REGS_0__14_), .B(_1568__bF_buf10), .Y(_2463_) );
AND2X2 AND2X2_1643 ( .A(_2463_), .B(_2462_), .Y(_2464_) );
AND2X2 AND2X2_1644 ( .A(_1730__bF_buf1), .B(_2464_), .Y(_2465_) );
OR2X2 OR2X2_1454 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_1__14_), .Y(_2466_) );
OR2X2 OR2X2_1455 ( .A(REGs_FIRQ_REGS_1__14_), .B(_1568__bF_buf10), .Y(_2467_) );
AND2X2 AND2X2_1645 ( .A(_2467_), .B(_2466_), .Y(_2468_) );
AND2X2 AND2X2_1646 ( .A(_1735__bF_buf3), .B(_2468_), .Y(_2469_) );
OR2X2 OR2X2_1456 ( .A(_2465_), .B(_2469_), .Y(_2470_) );
OR2X2 OR2X2_1457 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_3__14_), .Y(_2471_) );
OR2X2 OR2X2_1458 ( .A(REGs_FIRQ_REGS_3__14_), .B(_1568__bF_buf10), .Y(_2472_) );
AND2X2 AND2X2_1647 ( .A(_2472_), .B(_2471_), .Y(_2473_) );
AND2X2 AND2X2_1648 ( .A(_2473_), .B(_1741__bF_buf2), .Y(_2474_) );
OR2X2 OR2X2_1459 ( .A(INTERRUPT_flag_bF_buf15_bF_buf0), .B(REGs_USR_REGS_2__14_), .Y(_2475_) );
OR2X2 OR2X2_1460 ( .A(REGs_FIRQ_REGS_2__14_), .B(_1568__bF_buf10), .Y(_2476_) );
AND2X2 AND2X2_1649 ( .A(_2476_), .B(_2475_), .Y(_2477_) );
AND2X2 AND2X2_1650 ( .A(_1746__bF_buf2), .B(_2477_), .Y(_2478_) );
OR2X2 OR2X2_1461 ( .A(_2474_), .B(_2478_), .Y(_2479_) );
OR2X2 OR2X2_1462 ( .A(_2479_), .B(_2470_), .Y(_2480_) );
OR2X2 OR2X2_1463 ( .A(_2461_), .B(_2480_), .Y(_2481_) );
OR2X2 OR2X2_1464 ( .A(_2442_), .B(_2481_), .Y(REG_B_14_) );
AND2X2 AND2X2_1651 ( .A(_1678__bF_buf2), .B(REGs_REGS_4__15_), .Y(_2482_) );
AND2X2 AND2X2_1652 ( .A(_1682__bF_buf1), .B(REGs_REGS_5__15_), .Y(_2483_) );
OR2X2 OR2X2_1465 ( .A(_2482_), .B(_2483_), .Y(_2484_) );
AND2X2 AND2X2_1653 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__15_), .Y(_2485_) );
AND2X2 AND2X2_1654 ( .A(_1690__bF_buf0), .B(REGs_REGS_7__15_), .Y(_2486_) );
OR2X2 OR2X2_1466 ( .A(_2486_), .B(_2485_), .Y(_2487_) );
OR2X2 OR2X2_1467 ( .A(_2484_), .B(_2487_), .Y(_2488_) );
AND2X2 AND2X2_1655 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2489_) );
AND2X2 AND2X2_1656 ( .A(_1697__bF_buf1), .B(REGs_REGS_3__15_), .Y(_2490_) );
AND2X2 AND2X2_1657 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__15_), .Y(_2491_) );
OR2X2 OR2X2_1468 ( .A(_2490_), .B(_2491_), .Y(_2492_) );
OR2X2 OR2X2_1469 ( .A(_2489_), .B(_2492_), .Y(_2493_) );
OR2X2 OR2X2_1470 ( .A(_2493_), .B(_2488_), .Y(_2494_) );
OR2X2 OR2X2_1471 ( .A(INTERRUPT_flag_bF_buf14_bF_buf1), .B(REGs_USR_REGS_5__15_), .Y(_2495_) );
OR2X2 OR2X2_1472 ( .A(REGs_FIRQ_REGS_5__15_), .B(_1568__bF_buf12), .Y(_2496_) );
AND2X2 AND2X2_1658 ( .A(_2496_), .B(_2495_), .Y(_2497_) );
AND2X2 AND2X2_1659 ( .A(_2497_), .B(_1705__bF_buf1), .Y(_2498_) );
OR2X2 OR2X2_1473 ( .A(INTERRUPT_flag_bF_buf13_bF_buf2), .B(REGs_USR_REGS_4__15_), .Y(_2499_) );
OR2X2 OR2X2_1474 ( .A(REGs_FIRQ_REGS_4__15_), .B(_1568__bF_buf12), .Y(_2500_) );
AND2X2 AND2X2_1660 ( .A(_2500_), .B(_2499_), .Y(_2501_) );
AND2X2 AND2X2_1661 ( .A(_2501_), .B(_1710__bF_buf0), .Y(_2502_) );
OR2X2 OR2X2_1475 ( .A(_2502_), .B(_2498_), .Y(_2503_) );
OR2X2 OR2X2_1476 ( .A(INTERRUPT_flag_bF_buf12_bF_buf1), .B(REGs_USR_REGS_6__15_), .Y(_2504_) );
OR2X2 OR2X2_1477 ( .A(REGs_FIRQ_REGS_6__15_), .B(_1568__bF_buf12), .Y(_2505_) );
AND2X2 AND2X2_1662 ( .A(_2505_), .B(_2504_), .Y(_2506_) );
AND2X2 AND2X2_1663 ( .A(_2506_), .B(_1716__bF_buf2), .Y(_2507_) );
OR2X2 OR2X2_1478 ( .A(INTERRUPT_flag_bF_buf11_bF_buf2), .B(REGs_USR_REGS_7__15_), .Y(_2508_) );
OR2X2 OR2X2_1479 ( .A(REGs_FIRQ_REGS_7__15_), .B(_1568__bF_buf12), .Y(_2509_) );
AND2X2 AND2X2_1664 ( .A(_2509_), .B(_2508_), .Y(_2510_) );
AND2X2 AND2X2_1665 ( .A(_2510_), .B(_1721__bF_buf4), .Y(_2511_) );
OR2X2 OR2X2_1480 ( .A(_2511_), .B(_2507_), .Y(_2512_) );
OR2X2 OR2X2_1481 ( .A(_2503_), .B(_2512_), .Y(_2513_) );
OR2X2 OR2X2_1482 ( .A(INTERRUPT_flag_bF_buf10_bF_buf0), .B(REGs_USR_REGS_0__15_), .Y(_2514_) );
OR2X2 OR2X2_1483 ( .A(REGs_FIRQ_REGS_0__15_), .B(_1568__bF_buf3), .Y(_2515_) );
AND2X2 AND2X2_1666 ( .A(_2515_), .B(_2514_), .Y(_2516_) );
AND2X2 AND2X2_1667 ( .A(_1730__bF_buf1), .B(_2516_), .Y(_2517_) );
OR2X2 OR2X2_1484 ( .A(INTERRUPT_flag_bF_buf9_bF_buf3), .B(REGs_USR_REGS_1__15_), .Y(_2518_) );
OR2X2 OR2X2_1485 ( .A(REGs_FIRQ_REGS_1__15_), .B(_1568__bF_buf10), .Y(_2519_) );
AND2X2 AND2X2_1668 ( .A(_2519_), .B(_2518_), .Y(_2520_) );
AND2X2 AND2X2_1669 ( .A(_1735__bF_buf3), .B(_2520_), .Y(_2521_) );
OR2X2 OR2X2_1486 ( .A(_2517_), .B(_2521_), .Y(_2522_) );
OR2X2 OR2X2_1487 ( .A(INTERRUPT_flag_bF_buf8_bF_buf1), .B(REGs_USR_REGS_3__15_), .Y(_2523_) );
OR2X2 OR2X2_1488 ( .A(REGs_FIRQ_REGS_3__15_), .B(_1568__bF_buf10), .Y(_2524_) );
AND2X2 AND2X2_1670 ( .A(_2524_), .B(_2523_), .Y(_2525_) );
AND2X2 AND2X2_1671 ( .A(_2525_), .B(_1741__bF_buf2), .Y(_2526_) );
OR2X2 OR2X2_1489 ( .A(INTERRUPT_flag_bF_buf7_bF_buf0), .B(REGs_USR_REGS_2__15_), .Y(_2527_) );
OR2X2 OR2X2_1490 ( .A(REGs_FIRQ_REGS_2__15_), .B(_1568__bF_buf15_bF_buf0), .Y(_2528_) );
AND2X2 AND2X2_1672 ( .A(_2528_), .B(_2527_), .Y(_2529_) );
AND2X2 AND2X2_1673 ( .A(_1746__bF_buf2), .B(_2529_), .Y(_2530_) );
OR2X2 OR2X2_1491 ( .A(_2526_), .B(_2530_), .Y(_2531_) );
OR2X2 OR2X2_1492 ( .A(_2531_), .B(_2522_), .Y(_2532_) );
OR2X2 OR2X2_1493 ( .A(_2513_), .B(_2532_), .Y(_2533_) );
OR2X2 OR2X2_1494 ( .A(_2494_), .B(_2533_), .Y(REG_B_15_) );
AND2X2 AND2X2_1674 ( .A(_1678__bF_buf2), .B(REGs_REGS_4__16_), .Y(_2534_) );
AND2X2 AND2X2_1675 ( .A(_1682__bF_buf1), .B(REGs_REGS_5__16_), .Y(_2535_) );
OR2X2 OR2X2_1495 ( .A(_2534_), .B(_2535_), .Y(_2536_) );
AND2X2 AND2X2_1676 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__16_), .Y(_2537_) );
AND2X2 AND2X2_1677 ( .A(_1690__bF_buf0), .B(REGs_REGS_7__16_), .Y(_2538_) );
OR2X2 OR2X2_1496 ( .A(_2538_), .B(_2537_), .Y(_2539_) );
OR2X2 OR2X2_1497 ( .A(_2536_), .B(_2539_), .Y(_2540_) );
AND2X2 AND2X2_1678 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2541_) );
AND2X2 AND2X2_1679 ( .A(_1697__bF_buf1), .B(REGs_REGS_3__16_), .Y(_2542_) );
AND2X2 AND2X2_1680 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__16_), .Y(_2543_) );
OR2X2 OR2X2_1498 ( .A(_2542_), .B(_2543_), .Y(_2544_) );
OR2X2 OR2X2_1499 ( .A(_2541_), .B(_2544_), .Y(_2545_) );
OR2X2 OR2X2_1500 ( .A(_2545_), .B(_2540_), .Y(_2546_) );
OR2X2 OR2X2_1501 ( .A(INTERRUPT_flag_bF_buf9), .B(REGs_USR_REGS_5__16_), .Y(_2547_) );
OR2X2 OR2X2_1502 ( .A(REGs_FIRQ_REGS_5__16_), .B(_1568__bF_buf12), .Y(_2548_) );
AND2X2 AND2X2_1681 ( .A(_2548_), .B(_2547_), .Y(_2549_) );
AND2X2 AND2X2_1682 ( .A(_2549_), .B(_1705__bF_buf1), .Y(_2550_) );
OR2X2 OR2X2_1503 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_4__16_), .Y(_2551_) );
OR2X2 OR2X2_1504 ( .A(REGs_FIRQ_REGS_4__16_), .B(_1568__bF_buf5), .Y(_2552_) );
AND2X2 AND2X2_1683 ( .A(_2552_), .B(_2551_), .Y(_2553_) );
AND2X2 AND2X2_1684 ( .A(_2553_), .B(_1710__bF_buf0), .Y(_2554_) );
OR2X2 OR2X2_1505 ( .A(_2554_), .B(_2550_), .Y(_2555_) );
OR2X2 OR2X2_1506 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_6__16_), .Y(_2556_) );
OR2X2 OR2X2_1507 ( .A(REGs_FIRQ_REGS_6__16_), .B(_1568__bF_buf8), .Y(_2557_) );
AND2X2 AND2X2_1685 ( .A(_2557_), .B(_2556_), .Y(_2558_) );
AND2X2 AND2X2_1686 ( .A(_2558_), .B(_1716__bF_buf2), .Y(_2559_) );
OR2X2 OR2X2_1508 ( .A(INTERRUPT_flag_bF_buf14), .B(REGs_USR_REGS_7__16_), .Y(_2560_) );
OR2X2 OR2X2_1509 ( .A(REGs_FIRQ_REGS_7__16_), .B(_1568__bF_buf8), .Y(_2561_) );
AND2X2 AND2X2_1687 ( .A(_2561_), .B(_2560_), .Y(_2562_) );
AND2X2 AND2X2_1688 ( .A(_2562_), .B(_1721__bF_buf4), .Y(_2563_) );
OR2X2 OR2X2_1510 ( .A(_2563_), .B(_2559_), .Y(_2564_) );
OR2X2 OR2X2_1511 ( .A(_2555_), .B(_2564_), .Y(_2565_) );
OR2X2 OR2X2_1512 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_0__16_), .Y(_2566_) );
OR2X2 OR2X2_1513 ( .A(REGs_FIRQ_REGS_0__16_), .B(_1568__bF_buf10), .Y(_2567_) );
AND2X2 AND2X2_1689 ( .A(_2567_), .B(_2566_), .Y(_2568_) );
AND2X2 AND2X2_1690 ( .A(_1730__bF_buf1), .B(_2568_), .Y(_2569_) );
OR2X2 OR2X2_1514 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_1__16_), .Y(_2570_) );
OR2X2 OR2X2_1515 ( .A(REGs_FIRQ_REGS_1__16_), .B(_1568__bF_buf10), .Y(_2571_) );
AND2X2 AND2X2_1691 ( .A(_2571_), .B(_2570_), .Y(_2572_) );
AND2X2 AND2X2_1692 ( .A(_1735__bF_buf3), .B(_2572_), .Y(_2573_) );
OR2X2 OR2X2_1516 ( .A(_2569_), .B(_2573_), .Y(_2574_) );
OR2X2 OR2X2_1517 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_3__16_), .Y(_2575_) );
OR2X2 OR2X2_1518 ( .A(REGs_FIRQ_REGS_3__16_), .B(_1568__bF_buf7), .Y(_2576_) );
AND2X2 AND2X2_1693 ( .A(_2576_), .B(_2575_), .Y(_2577_) );
AND2X2 AND2X2_1694 ( .A(_2577_), .B(_1741__bF_buf2), .Y(_2578_) );
OR2X2 OR2X2_1519 ( .A(INTERRUPT_flag_bF_buf15_bF_buf0), .B(REGs_USR_REGS_2__16_), .Y(_2579_) );
OR2X2 OR2X2_1520 ( .A(REGs_FIRQ_REGS_2__16_), .B(_1568__bF_buf10), .Y(_2580_) );
AND2X2 AND2X2_1695 ( .A(_2580_), .B(_2579_), .Y(_2581_) );
AND2X2 AND2X2_1696 ( .A(_1746__bF_buf2), .B(_2581_), .Y(_2582_) );
OR2X2 OR2X2_1521 ( .A(_2578_), .B(_2582_), .Y(_2583_) );
OR2X2 OR2X2_1522 ( .A(_2583_), .B(_2574_), .Y(_2584_) );
OR2X2 OR2X2_1523 ( .A(_2565_), .B(_2584_), .Y(_2585_) );
OR2X2 OR2X2_1524 ( .A(_2546_), .B(_2585_), .Y(REG_B_16_) );
AND2X2 AND2X2_1697 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__17_), .Y(_2586_) );
AND2X2 AND2X2_1698 ( .A(_1682__bF_buf2), .B(REGs_REGS_5__17_), .Y(_2587_) );
OR2X2 OR2X2_1525 ( .A(_2586_), .B(_2587_), .Y(_2588_) );
AND2X2 AND2X2_1699 ( .A(_1687__bF_buf2), .B(REGs_REGS_6__17_), .Y(_2589_) );
AND2X2 AND2X2_1700 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__17_), .Y(_2590_) );
OR2X2 OR2X2_1526 ( .A(_2590_), .B(_2589_), .Y(_2591_) );
OR2X2 OR2X2_1527 ( .A(_2588_), .B(_2591_), .Y(_2592_) );
AND2X2 AND2X2_1701 ( .A(_1695__bF_buf4), .B(gnd), .Y(_2593_) );
AND2X2 AND2X2_1702 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__17_), .Y(_2594_) );
AND2X2 AND2X2_1703 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__17_), .Y(_2595_) );
OR2X2 OR2X2_1528 ( .A(_2594_), .B(_2595_), .Y(_2596_) );
OR2X2 OR2X2_1529 ( .A(_2593_), .B(_2596_), .Y(_2597_) );
OR2X2 OR2X2_1530 ( .A(_2597_), .B(_2592_), .Y(_2598_) );
OR2X2 OR2X2_1531 ( .A(INTERRUPT_flag_bF_buf14_bF_buf3), .B(REGs_USR_REGS_5__17_), .Y(_2599_) );
OR2X2 OR2X2_1532 ( .A(REGs_FIRQ_REGS_5__17_), .B(_1568__bF_buf15), .Y(_2600_) );
AND2X2 AND2X2_1704 ( .A(_2600_), .B(_2599_), .Y(_2601_) );
AND2X2 AND2X2_1705 ( .A(_2601_), .B(_1705__bF_buf3), .Y(_2602_) );
OR2X2 OR2X2_1533 ( .A(INTERRUPT_flag_bF_buf13_bF_buf0), .B(REGs_USR_REGS_4__17_), .Y(_2603_) );
OR2X2 OR2X2_1534 ( .A(REGs_FIRQ_REGS_4__17_), .B(_1568__bF_buf4), .Y(_2604_) );
AND2X2 AND2X2_1706 ( .A(_2604_), .B(_2603_), .Y(_2605_) );
AND2X2 AND2X2_1707 ( .A(_2605_), .B(_1710__bF_buf4), .Y(_2606_) );
OR2X2 OR2X2_1535 ( .A(_2606_), .B(_2602_), .Y(_2607_) );
OR2X2 OR2X2_1536 ( .A(INTERRUPT_flag_bF_buf12_bF_buf0), .B(REGs_USR_REGS_6__17_), .Y(_2608_) );
OR2X2 OR2X2_1537 ( .A(REGs_FIRQ_REGS_6__17_), .B(_1568__bF_buf1), .Y(_2609_) );
AND2X2 AND2X2_1708 ( .A(_2609_), .B(_2608_), .Y(_2610_) );
AND2X2 AND2X2_1709 ( .A(_2610_), .B(_1716__bF_buf3), .Y(_2611_) );
OR2X2 OR2X2_1538 ( .A(INTERRUPT_flag_bF_buf11_bF_buf1), .B(REGs_USR_REGS_7__17_), .Y(_2612_) );
OR2X2 OR2X2_1539 ( .A(REGs_FIRQ_REGS_7__17_), .B(_1568__bF_buf0), .Y(_2613_) );
AND2X2 AND2X2_1710 ( .A(_2613_), .B(_2612_), .Y(_2614_) );
AND2X2 AND2X2_1711 ( .A(_2614_), .B(_1721__bF_buf3), .Y(_2615_) );
OR2X2 OR2X2_1540 ( .A(_2615_), .B(_2611_), .Y(_2616_) );
OR2X2 OR2X2_1541 ( .A(_2607_), .B(_2616_), .Y(_2617_) );
OR2X2 OR2X2_1542 ( .A(INTERRUPT_flag_bF_buf10_bF_buf2), .B(REGs_USR_REGS_0__17_), .Y(_2618_) );
OR2X2 OR2X2_1543 ( .A(REGs_FIRQ_REGS_0__17_), .B(_1568__bF_buf9), .Y(_2619_) );
AND2X2 AND2X2_1712 ( .A(_2619_), .B(_2618_), .Y(_2620_) );
AND2X2 AND2X2_1713 ( .A(_1730__bF_buf4), .B(_2620_), .Y(_2621_) );
OR2X2 OR2X2_1544 ( .A(INTERRUPT_flag_bF_buf9_bF_buf1), .B(REGs_USR_REGS_1__17_), .Y(_2622_) );
OR2X2 OR2X2_1545 ( .A(REGs_FIRQ_REGS_1__17_), .B(_1568__bF_buf9), .Y(_2623_) );
AND2X2 AND2X2_1714 ( .A(_2623_), .B(_2622_), .Y(_2624_) );
AND2X2 AND2X2_1715 ( .A(_1735__bF_buf4), .B(_2624_), .Y(_2625_) );
OR2X2 OR2X2_1546 ( .A(_2621_), .B(_2625_), .Y(_2626_) );
OR2X2 OR2X2_1547 ( .A(INTERRUPT_flag_bF_buf8_bF_buf3), .B(REGs_USR_REGS_3__17_), .Y(_2627_) );
OR2X2 OR2X2_1548 ( .A(REGs_FIRQ_REGS_3__17_), .B(_1568__bF_buf2), .Y(_2628_) );
AND2X2 AND2X2_1716 ( .A(_2628_), .B(_2627_), .Y(_2629_) );
AND2X2 AND2X2_1717 ( .A(_2629_), .B(_1741__bF_buf0), .Y(_2630_) );
OR2X2 OR2X2_1549 ( .A(INTERRUPT_flag_bF_buf7_bF_buf3), .B(REGs_USR_REGS_2__17_), .Y(_2631_) );
OR2X2 OR2X2_1550 ( .A(REGs_FIRQ_REGS_2__17_), .B(_1568__bF_buf15_bF_buf3), .Y(_2632_) );
AND2X2 AND2X2_1718 ( .A(_2632_), .B(_2631_), .Y(_2633_) );
AND2X2 AND2X2_1719 ( .A(_1746__bF_buf3), .B(_2633_), .Y(_2634_) );
OR2X2 OR2X2_1551 ( .A(_2630_), .B(_2634_), .Y(_2635_) );
OR2X2 OR2X2_1552 ( .A(_2635_), .B(_2626_), .Y(_2636_) );
OR2X2 OR2X2_1553 ( .A(_2617_), .B(_2636_), .Y(_2637_) );
OR2X2 OR2X2_1554 ( .A(_2598_), .B(_2637_), .Y(REG_B_17_) );
AND2X2 AND2X2_1720 ( .A(_1678__bF_buf1), .B(REGs_REGS_4__18_), .Y(_2638_) );
AND2X2 AND2X2_1721 ( .A(_1682__bF_buf0), .B(REGs_REGS_5__18_), .Y(_2639_) );
OR2X2 OR2X2_1555 ( .A(_2638_), .B(_2639_), .Y(_2640_) );
AND2X2 AND2X2_1722 ( .A(_1687__bF_buf2), .B(REGs_REGS_6__18_), .Y(_2641_) );
AND2X2 AND2X2_1723 ( .A(_1690__bF_buf1), .B(REGs_REGS_7__18_), .Y(_2642_) );
OR2X2 OR2X2_1556 ( .A(_2642_), .B(_2641_), .Y(_2643_) );
OR2X2 OR2X2_1557 ( .A(_2640_), .B(_2643_), .Y(_2644_) );
AND2X2 AND2X2_1724 ( .A(_1695__bF_buf1), .B(gnd), .Y(_2645_) );
AND2X2 AND2X2_1725 ( .A(_1697__bF_buf2), .B(REGs_REGS_3__18_), .Y(_2646_) );
AND2X2 AND2X2_1726 ( .A(_1699__bF_buf1), .B(REGs_REGS_2__18_), .Y(_2647_) );
OR2X2 OR2X2_1558 ( .A(_2646_), .B(_2647_), .Y(_2648_) );
OR2X2 OR2X2_1559 ( .A(_2645_), .B(_2648_), .Y(_2649_) );
OR2X2 OR2X2_1560 ( .A(_2649_), .B(_2644_), .Y(_2650_) );
OR2X2 OR2X2_1561 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_5__18_), .Y(_2651_) );
OR2X2 OR2X2_1562 ( .A(REGs_FIRQ_REGS_5__18_), .B(_1568__bF_buf5), .Y(_2652_) );
AND2X2 AND2X2_1727 ( .A(_2652_), .B(_2651_), .Y(_2653_) );
AND2X2 AND2X2_1728 ( .A(_2653_), .B(_1705__bF_buf2), .Y(_2654_) );
OR2X2 OR2X2_1563 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_4__18_), .Y(_2655_) );
OR2X2 OR2X2_1564 ( .A(REGs_FIRQ_REGS_4__18_), .B(_1568__bF_buf5), .Y(_2656_) );
AND2X2 AND2X2_1729 ( .A(_2656_), .B(_2655_), .Y(_2657_) );
AND2X2 AND2X2_1730 ( .A(_2657_), .B(_1710__bF_buf1), .Y(_2658_) );
OR2X2 OR2X2_1565 ( .A(_2658_), .B(_2654_), .Y(_2659_) );
OR2X2 OR2X2_1566 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_6__18_), .Y(_2660_) );
OR2X2 OR2X2_1567 ( .A(REGs_FIRQ_REGS_6__18_), .B(_1568__bF_buf8), .Y(_2661_) );
AND2X2 AND2X2_1731 ( .A(_2661_), .B(_2660_), .Y(_2662_) );
AND2X2 AND2X2_1732 ( .A(_2662_), .B(_1716__bF_buf1), .Y(_2663_) );
OR2X2 OR2X2_1568 ( .A(INTERRUPT_flag_bF_buf5), .B(REGs_USR_REGS_7__18_), .Y(_2664_) );
OR2X2 OR2X2_1569 ( .A(REGs_FIRQ_REGS_7__18_), .B(_1568__bF_buf5), .Y(_2665_) );
AND2X2 AND2X2_1733 ( .A(_2665_), .B(_2664_), .Y(_2666_) );
AND2X2 AND2X2_1734 ( .A(_2666_), .B(_1721__bF_buf1), .Y(_2667_) );
OR2X2 OR2X2_1570 ( .A(_2667_), .B(_2663_), .Y(_2668_) );
OR2X2 OR2X2_1571 ( .A(_2659_), .B(_2668_), .Y(_2669_) );
OR2X2 OR2X2_1572 ( .A(INTERRUPT_flag_bF_buf11), .B(REGs_USR_REGS_0__18_), .Y(_2670_) );
OR2X2 OR2X2_1573 ( .A(REGs_FIRQ_REGS_0__18_), .B(_1568__bF_buf3), .Y(_2671_) );
AND2X2 AND2X2_1735 ( .A(_2671_), .B(_2670_), .Y(_2672_) );
AND2X2 AND2X2_1736 ( .A(_1730__bF_buf1), .B(_2672_), .Y(_2673_) );
OR2X2 OR2X2_1574 ( .A(INTERRUPT_flag_bF_buf11), .B(REGs_USR_REGS_1__18_), .Y(_2674_) );
OR2X2 OR2X2_1575 ( .A(REGs_FIRQ_REGS_1__18_), .B(_1568__bF_buf10), .Y(_2675_) );
AND2X2 AND2X2_1737 ( .A(_2675_), .B(_2674_), .Y(_2676_) );
AND2X2 AND2X2_1738 ( .A(_1735__bF_buf3), .B(_2676_), .Y(_2677_) );
OR2X2 OR2X2_1576 ( .A(_2673_), .B(_2677_), .Y(_2678_) );
OR2X2 OR2X2_1577 ( .A(INTERRUPT_flag_bF_buf11), .B(REGs_USR_REGS_3__18_), .Y(_2679_) );
OR2X2 OR2X2_1578 ( .A(REGs_FIRQ_REGS_3__18_), .B(_1568__bF_buf3), .Y(_2680_) );
AND2X2 AND2X2_1739 ( .A(_2680_), .B(_2679_), .Y(_2681_) );
AND2X2 AND2X2_1740 ( .A(_2681_), .B(_1741__bF_buf2), .Y(_2682_) );
OR2X2 OR2X2_1579 ( .A(INTERRUPT_flag_bF_buf15_bF_buf0), .B(REGs_USR_REGS_2__18_), .Y(_2683_) );
OR2X2 OR2X2_1580 ( .A(REGs_FIRQ_REGS_2__18_), .B(_1568__bF_buf10), .Y(_2684_) );
AND2X2 AND2X2_1741 ( .A(_2684_), .B(_2683_), .Y(_2685_) );
AND2X2 AND2X2_1742 ( .A(_1746__bF_buf2), .B(_2685_), .Y(_2686_) );
OR2X2 OR2X2_1581 ( .A(_2682_), .B(_2686_), .Y(_2687_) );
OR2X2 OR2X2_1582 ( .A(_2687_), .B(_2678_), .Y(_2688_) );
OR2X2 OR2X2_1583 ( .A(_2669_), .B(_2688_), .Y(_2689_) );
OR2X2 OR2X2_1584 ( .A(_2650_), .B(_2689_), .Y(REG_B_18_) );
AND2X2 AND2X2_1743 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__19_), .Y(_2690_) );
AND2X2 AND2X2_1744 ( .A(_1682__bF_buf2), .B(REGs_REGS_5__19_), .Y(_2691_) );
OR2X2 OR2X2_1585 ( .A(_2690_), .B(_2691_), .Y(_2692_) );
AND2X2 AND2X2_1745 ( .A(_1687__bF_buf2), .B(REGs_REGS_6__19_), .Y(_2693_) );
AND2X2 AND2X2_1746 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__19_), .Y(_2694_) );
OR2X2 OR2X2_1586 ( .A(_2694_), .B(_2693_), .Y(_2695_) );
OR2X2 OR2X2_1587 ( .A(_2692_), .B(_2695_), .Y(_2696_) );
AND2X2 AND2X2_1747 ( .A(_1695__bF_buf1), .B(gnd), .Y(_2697_) );
AND2X2 AND2X2_1748 ( .A(_1697__bF_buf0), .B(REGs_REGS_3__19_), .Y(_2698_) );
AND2X2 AND2X2_1749 ( .A(_1699__bF_buf1), .B(REGs_REGS_2__19_), .Y(_2699_) );
OR2X2 OR2X2_1588 ( .A(_2698_), .B(_2699_), .Y(_2700_) );
OR2X2 OR2X2_1589 ( .A(_2697_), .B(_2700_), .Y(_2701_) );
OR2X2 OR2X2_1590 ( .A(_2701_), .B(_2696_), .Y(_2702_) );
OR2X2 OR2X2_1591 ( .A(INTERRUPT_flag_bF_buf14_bF_buf2), .B(REGs_USR_REGS_5__19_), .Y(_2703_) );
OR2X2 OR2X2_1592 ( .A(REGs_FIRQ_REGS_5__19_), .B(_1568__bF_buf13), .Y(_2704_) );
AND2X2 AND2X2_1750 ( .A(_2704_), .B(_2703_), .Y(_2705_) );
AND2X2 AND2X2_1751 ( .A(_2705_), .B(_1705__bF_buf0), .Y(_2706_) );
OR2X2 OR2X2_1593 ( .A(INTERRUPT_flag_bF_buf13_bF_buf3), .B(REGs_USR_REGS_4__19_), .Y(_2707_) );
OR2X2 OR2X2_1594 ( .A(REGs_FIRQ_REGS_4__19_), .B(_1568__bF_buf13), .Y(_2708_) );
AND2X2 AND2X2_1752 ( .A(_2708_), .B(_2707_), .Y(_2709_) );
AND2X2 AND2X2_1753 ( .A(_2709_), .B(_1710__bF_buf2), .Y(_2710_) );
OR2X2 OR2X2_1595 ( .A(_2710_), .B(_2706_), .Y(_2711_) );
OR2X2 OR2X2_1596 ( .A(INTERRUPT_flag_bF_buf12_bF_buf3), .B(REGs_USR_REGS_6__19_), .Y(_2712_) );
OR2X2 OR2X2_1597 ( .A(REGs_FIRQ_REGS_6__19_), .B(_1568__bF_buf13), .Y(_2713_) );
AND2X2 AND2X2_1754 ( .A(_2713_), .B(_2712_), .Y(_2714_) );
AND2X2 AND2X2_1755 ( .A(_2714_), .B(_1716__bF_buf0), .Y(_2715_) );
OR2X2 OR2X2_1598 ( .A(INTERRUPT_flag_bF_buf11_bF_buf3), .B(REGs_USR_REGS_7__19_), .Y(_2716_) );
OR2X2 OR2X2_1599 ( .A(REGs_FIRQ_REGS_7__19_), .B(_1568__bF_buf13), .Y(_2717_) );
AND2X2 AND2X2_1756 ( .A(_2717_), .B(_2716_), .Y(_2718_) );
AND2X2 AND2X2_1757 ( .A(_2718_), .B(_1721__bF_buf2), .Y(_2719_) );
OR2X2 OR2X2_1600 ( .A(_2719_), .B(_2715_), .Y(_2720_) );
OR2X2 OR2X2_1601 ( .A(_2711_), .B(_2720_), .Y(_2721_) );
OR2X2 OR2X2_1602 ( .A(INTERRUPT_flag_bF_buf10_bF_buf1), .B(REGs_USR_REGS_0__19_), .Y(_2722_) );
OR2X2 OR2X2_1603 ( .A(REGs_FIRQ_REGS_0__19_), .B(_1568__bF_buf13), .Y(_2723_) );
AND2X2 AND2X2_1758 ( .A(_2723_), .B(_2722_), .Y(_2724_) );
AND2X2 AND2X2_1759 ( .A(_1730__bF_buf2), .B(_2724_), .Y(_2725_) );
OR2X2 OR2X2_1604 ( .A(INTERRUPT_flag_bF_buf9_bF_buf2), .B(REGs_USR_REGS_1__19_), .Y(_2726_) );
OR2X2 OR2X2_1605 ( .A(REGs_FIRQ_REGS_1__19_), .B(_1568__bF_buf6), .Y(_2727_) );
AND2X2 AND2X2_1760 ( .A(_2727_), .B(_2726_), .Y(_2728_) );
AND2X2 AND2X2_1761 ( .A(_1735__bF_buf0), .B(_2728_), .Y(_2729_) );
OR2X2 OR2X2_1606 ( .A(_2725_), .B(_2729_), .Y(_2730_) );
OR2X2 OR2X2_1607 ( .A(INTERRUPT_flag_bF_buf8_bF_buf0), .B(REGs_USR_REGS_3__19_), .Y(_2731_) );
OR2X2 OR2X2_1608 ( .A(REGs_FIRQ_REGS_3__19_), .B(_1568__bF_buf6), .Y(_2732_) );
AND2X2 AND2X2_1762 ( .A(_2732_), .B(_2731_), .Y(_2733_) );
AND2X2 AND2X2_1763 ( .A(_2733_), .B(_1741__bF_buf1), .Y(_2734_) );
OR2X2 OR2X2_1609 ( .A(INTERRUPT_flag_bF_buf7_bF_buf1), .B(REGs_USR_REGS_2__19_), .Y(_2735_) );
OR2X2 OR2X2_1610 ( .A(REGs_FIRQ_REGS_2__19_), .B(_1568__bF_buf15_bF_buf1), .Y(_2736_) );
AND2X2 AND2X2_1764 ( .A(_2736_), .B(_2735_), .Y(_2737_) );
AND2X2 AND2X2_1765 ( .A(_1746__bF_buf4), .B(_2737_), .Y(_2738_) );
OR2X2 OR2X2_1611 ( .A(_2734_), .B(_2738_), .Y(_2739_) );
OR2X2 OR2X2_1612 ( .A(_2739_), .B(_2730_), .Y(_2740_) );
OR2X2 OR2X2_1613 ( .A(_2721_), .B(_2740_), .Y(_2741_) );
OR2X2 OR2X2_1614 ( .A(_2702_), .B(_2741_), .Y(REG_B_19_) );
AND2X2 AND2X2_1766 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__20_), .Y(_2742_) );
AND2X2 AND2X2_1767 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__20_), .Y(_2743_) );
OR2X2 OR2X2_1615 ( .A(_2742_), .B(_2743_), .Y(_2744_) );
AND2X2 AND2X2_1768 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__20_), .Y(_2745_) );
AND2X2 AND2X2_1769 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__20_), .Y(_2746_) );
OR2X2 OR2X2_1616 ( .A(_2746_), .B(_2745_), .Y(_2747_) );
OR2X2 OR2X2_1617 ( .A(_2744_), .B(_2747_), .Y(_2748_) );
AND2X2 AND2X2_1770 ( .A(_1695__bF_buf0), .B(gnd), .Y(_2749_) );
AND2X2 AND2X2_1771 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__20_), .Y(_2750_) );
AND2X2 AND2X2_1772 ( .A(_1699__bF_buf0), .B(REGs_REGS_2__20_), .Y(_2751_) );
OR2X2 OR2X2_1618 ( .A(_2750_), .B(_2751_), .Y(_2752_) );
OR2X2 OR2X2_1619 ( .A(_2749_), .B(_2752_), .Y(_2753_) );
OR2X2 OR2X2_1620 ( .A(_2753_), .B(_2748_), .Y(_2754_) );
OR2X2 OR2X2_1621 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_5__20_), .Y(_2755_) );
OR2X2 OR2X2_1622 ( .A(REGs_FIRQ_REGS_5__20_), .B(_1568__bF_buf1), .Y(_2756_) );
AND2X2 AND2X2_1773 ( .A(_2756_), .B(_2755_), .Y(_2757_) );
AND2X2 AND2X2_1774 ( .A(_2757_), .B(_1705__bF_buf3), .Y(_2758_) );
OR2X2 OR2X2_1623 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_4__20_), .Y(_2759_) );
OR2X2 OR2X2_1624 ( .A(REGs_FIRQ_REGS_4__20_), .B(_1568__bF_buf2), .Y(_2760_) );
AND2X2 AND2X2_1775 ( .A(_2760_), .B(_2759_), .Y(_2761_) );
AND2X2 AND2X2_1776 ( .A(_2761_), .B(_1710__bF_buf4), .Y(_2762_) );
OR2X2 OR2X2_1625 ( .A(_2762_), .B(_2758_), .Y(_2763_) );
OR2X2 OR2X2_1626 ( .A(INTERRUPT_flag_bF_buf7), .B(REGs_USR_REGS_6__20_), .Y(_2764_) );
OR2X2 OR2X2_1627 ( .A(REGs_FIRQ_REGS_6__20_), .B(_1568__bF_buf4), .Y(_2765_) );
AND2X2 AND2X2_1777 ( .A(_2765_), .B(_2764_), .Y(_2766_) );
AND2X2 AND2X2_1778 ( .A(_2766_), .B(_1716__bF_buf3), .Y(_2767_) );
OR2X2 OR2X2_1628 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_7__20_), .Y(_2768_) );
OR2X2 OR2X2_1629 ( .A(REGs_FIRQ_REGS_7__20_), .B(_1568__bF_buf1), .Y(_2769_) );
AND2X2 AND2X2_1779 ( .A(_2769_), .B(_2768_), .Y(_2770_) );
AND2X2 AND2X2_1780 ( .A(_2770_), .B(_1721__bF_buf3), .Y(_2771_) );
OR2X2 OR2X2_1630 ( .A(_2771_), .B(_2767_), .Y(_2772_) );
OR2X2 OR2X2_1631 ( .A(_2763_), .B(_2772_), .Y(_2773_) );
OR2X2 OR2X2_1632 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_0__20_), .Y(_2774_) );
OR2X2 OR2X2_1633 ( .A(REGs_FIRQ_REGS_0__20_), .B(_1568__bF_buf0), .Y(_2775_) );
AND2X2 AND2X2_1781 ( .A(_2775_), .B(_2774_), .Y(_2776_) );
AND2X2 AND2X2_1782 ( .A(_1730__bF_buf4), .B(_2776_), .Y(_2777_) );
OR2X2 OR2X2_1634 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_1__20_), .Y(_2778_) );
OR2X2 OR2X2_1635 ( .A(REGs_FIRQ_REGS_1__20_), .B(_1568__bF_buf9), .Y(_2779_) );
AND2X2 AND2X2_1783 ( .A(_2779_), .B(_2778_), .Y(_2780_) );
AND2X2 AND2X2_1784 ( .A(_1735__bF_buf4), .B(_2780_), .Y(_2781_) );
OR2X2 OR2X2_1636 ( .A(_2777_), .B(_2781_), .Y(_2782_) );
OR2X2 OR2X2_1637 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_3__20_), .Y(_2783_) );
OR2X2 OR2X2_1638 ( .A(REGs_FIRQ_REGS_3__20_), .B(_1568__bF_buf2), .Y(_2784_) );
AND2X2 AND2X2_1785 ( .A(_2784_), .B(_2783_), .Y(_2785_) );
AND2X2 AND2X2_1786 ( .A(_2785_), .B(_1741__bF_buf0), .Y(_2786_) );
OR2X2 OR2X2_1639 ( .A(INTERRUPT_flag_bF_buf15_bF_buf1), .B(REGs_USR_REGS_2__20_), .Y(_2787_) );
OR2X2 OR2X2_1640 ( .A(REGs_FIRQ_REGS_2__20_), .B(_1568__bF_buf2), .Y(_2788_) );
AND2X2 AND2X2_1787 ( .A(_2788_), .B(_2787_), .Y(_2789_) );
AND2X2 AND2X2_1788 ( .A(_1746__bF_buf3), .B(_2789_), .Y(_2790_) );
OR2X2 OR2X2_1641 ( .A(_2786_), .B(_2790_), .Y(_2791_) );
OR2X2 OR2X2_1642 ( .A(_2791_), .B(_2782_), .Y(_2792_) );
OR2X2 OR2X2_1643 ( .A(_2773_), .B(_2792_), .Y(_2793_) );
OR2X2 OR2X2_1644 ( .A(_2754_), .B(_2793_), .Y(REG_B_20_) );
AND2X2 AND2X2_1789 ( .A(_1678__bF_buf1), .B(REGs_REGS_4__21_), .Y(_2794_) );
AND2X2 AND2X2_1790 ( .A(_1682__bF_buf0), .B(REGs_REGS_5__21_), .Y(_2795_) );
OR2X2 OR2X2_1645 ( .A(_2794_), .B(_2795_), .Y(_2796_) );
AND2X2 AND2X2_1791 ( .A(_1687__bF_buf0), .B(REGs_REGS_6__21_), .Y(_2797_) );
AND2X2 AND2X2_1792 ( .A(_1690__bF_buf1), .B(REGs_REGS_7__21_), .Y(_2798_) );
OR2X2 OR2X2_1646 ( .A(_2798_), .B(_2797_), .Y(_2799_) );
OR2X2 OR2X2_1647 ( .A(_2796_), .B(_2799_), .Y(_2800_) );
AND2X2 AND2X2_1793 ( .A(_1695__bF_buf1), .B(gnd), .Y(_2801_) );
AND2X2 AND2X2_1794 ( .A(_1697__bF_buf2), .B(REGs_REGS_3__21_), .Y(_2802_) );
AND2X2 AND2X2_1795 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__21_), .Y(_2803_) );
OR2X2 OR2X2_1648 ( .A(_2802_), .B(_2803_), .Y(_2804_) );
OR2X2 OR2X2_1649 ( .A(_2801_), .B(_2804_), .Y(_2805_) );
OR2X2 OR2X2_1650 ( .A(_2805_), .B(_2800_), .Y(_2806_) );
OR2X2 OR2X2_1651 ( .A(INTERRUPT_flag_bF_buf14_bF_buf2), .B(REGs_USR_REGS_5__21_), .Y(_2807_) );
OR2X2 OR2X2_1652 ( .A(REGs_FIRQ_REGS_5__21_), .B(_1568__bF_buf7), .Y(_2808_) );
AND2X2 AND2X2_1796 ( .A(_2808_), .B(_2807_), .Y(_2809_) );
AND2X2 AND2X2_1797 ( .A(_2809_), .B(_1705__bF_buf0), .Y(_2810_) );
OR2X2 OR2X2_1653 ( .A(INTERRUPT_flag_bF_buf13_bF_buf2), .B(REGs_USR_REGS_4__21_), .Y(_2811_) );
OR2X2 OR2X2_1654 ( .A(REGs_FIRQ_REGS_4__21_), .B(_1568__bF_buf7), .Y(_2812_) );
AND2X2 AND2X2_1798 ( .A(_2812_), .B(_2811_), .Y(_2813_) );
AND2X2 AND2X2_1799 ( .A(_2813_), .B(_1710__bF_buf2), .Y(_2814_) );
OR2X2 OR2X2_1655 ( .A(_2814_), .B(_2810_), .Y(_2815_) );
OR2X2 OR2X2_1656 ( .A(INTERRUPT_flag_bF_buf12_bF_buf3), .B(REGs_USR_REGS_6__21_), .Y(_2816_) );
OR2X2 OR2X2_1657 ( .A(REGs_FIRQ_REGS_6__21_), .B(_1568__bF_buf8), .Y(_2817_) );
AND2X2 AND2X2_1800 ( .A(_2817_), .B(_2816_), .Y(_2818_) );
AND2X2 AND2X2_1801 ( .A(_2818_), .B(_1716__bF_buf0), .Y(_2819_) );
OR2X2 OR2X2_1658 ( .A(INTERRUPT_flag_bF_buf11_bF_buf0), .B(REGs_USR_REGS_7__21_), .Y(_2820_) );
OR2X2 OR2X2_1659 ( .A(REGs_FIRQ_REGS_7__21_), .B(_1568__bF_buf8), .Y(_2821_) );
AND2X2 AND2X2_1802 ( .A(_2821_), .B(_2820_), .Y(_2822_) );
AND2X2 AND2X2_1803 ( .A(_2822_), .B(_1721__bF_buf4), .Y(_2823_) );
OR2X2 OR2X2_1660 ( .A(_2823_), .B(_2819_), .Y(_2824_) );
OR2X2 OR2X2_1661 ( .A(_2815_), .B(_2824_), .Y(_2825_) );
OR2X2 OR2X2_1662 ( .A(INTERRUPT_flag_bF_buf10_bF_buf0), .B(REGs_USR_REGS_0__21_), .Y(_2826_) );
OR2X2 OR2X2_1663 ( .A(REGs_FIRQ_REGS_0__21_), .B(_1568__bF_buf7), .Y(_2827_) );
AND2X2 AND2X2_1804 ( .A(_2827_), .B(_2826_), .Y(_2828_) );
AND2X2 AND2X2_1805 ( .A(_1730__bF_buf0), .B(_2828_), .Y(_2829_) );
OR2X2 OR2X2_1664 ( .A(INTERRUPT_flag_bF_buf9_bF_buf2), .B(REGs_USR_REGS_1__21_), .Y(_2830_) );
OR2X2 OR2X2_1665 ( .A(REGs_FIRQ_REGS_1__21_), .B(_1568__bF_buf3), .Y(_2831_) );
AND2X2 AND2X2_1806 ( .A(_2831_), .B(_2830_), .Y(_2832_) );
AND2X2 AND2X2_1807 ( .A(_1735__bF_buf2), .B(_2832_), .Y(_2833_) );
OR2X2 OR2X2_1666 ( .A(_2829_), .B(_2833_), .Y(_2834_) );
OR2X2 OR2X2_1667 ( .A(INTERRUPT_flag_bF_buf8_bF_buf1), .B(REGs_USR_REGS_3__21_), .Y(_2835_) );
OR2X2 OR2X2_1668 ( .A(REGs_FIRQ_REGS_3__21_), .B(_1568__bF_buf7), .Y(_2836_) );
AND2X2 AND2X2_1808 ( .A(_2836_), .B(_2835_), .Y(_2837_) );
AND2X2 AND2X2_1809 ( .A(_2837_), .B(_1741__bF_buf2), .Y(_2838_) );
OR2X2 OR2X2_1669 ( .A(INTERRUPT_flag_bF_buf7_bF_buf0), .B(REGs_USR_REGS_2__21_), .Y(_2839_) );
OR2X2 OR2X2_1670 ( .A(REGs_FIRQ_REGS_2__21_), .B(_1568__bF_buf15_bF_buf0), .Y(_2840_) );
AND2X2 AND2X2_1810 ( .A(_2840_), .B(_2839_), .Y(_2841_) );
AND2X2 AND2X2_1811 ( .A(_1746__bF_buf2), .B(_2841_), .Y(_2842_) );
OR2X2 OR2X2_1671 ( .A(_2838_), .B(_2842_), .Y(_2843_) );
OR2X2 OR2X2_1672 ( .A(_2843_), .B(_2834_), .Y(_2844_) );
OR2X2 OR2X2_1673 ( .A(_2825_), .B(_2844_), .Y(_2845_) );
OR2X2 OR2X2_1674 ( .A(_2806_), .B(_2845_), .Y(REG_B_21_) );
AND2X2 AND2X2_1812 ( .A(_1678__bF_buf0), .B(REGs_REGS_4__22_), .Y(_2846_) );
AND2X2 AND2X2_1813 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__22_), .Y(_2847_) );
OR2X2 OR2X2_1675 ( .A(_2846_), .B(_2847_), .Y(_2848_) );
AND2X2 AND2X2_1814 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__22_), .Y(_2849_) );
AND2X2 AND2X2_1815 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__22_), .Y(_2850_) );
OR2X2 OR2X2_1676 ( .A(_2850_), .B(_2849_), .Y(_2851_) );
OR2X2 OR2X2_1677 ( .A(_2848_), .B(_2851_), .Y(_2852_) );
AND2X2 AND2X2_1816 ( .A(_1695__bF_buf2), .B(gnd), .Y(_2853_) );
AND2X2 AND2X2_1817 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__22_), .Y(_2854_) );
AND2X2 AND2X2_1818 ( .A(_1699__bF_buf2), .B(REGs_REGS_2__22_), .Y(_2855_) );
OR2X2 OR2X2_1678 ( .A(_2854_), .B(_2855_), .Y(_2856_) );
OR2X2 OR2X2_1679 ( .A(_2853_), .B(_2856_), .Y(_2857_) );
OR2X2 OR2X2_1680 ( .A(_2857_), .B(_2852_), .Y(_2858_) );
OR2X2 OR2X2_1681 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_5__22_), .Y(_2859_) );
OR2X2 OR2X2_1682 ( .A(REGs_FIRQ_REGS_5__22_), .B(_1568__bF_buf0), .Y(_2860_) );
AND2X2 AND2X2_1819 ( .A(_2860_), .B(_2859_), .Y(_2861_) );
AND2X2 AND2X2_1820 ( .A(_2861_), .B(_1705__bF_buf4), .Y(_2862_) );
OR2X2 OR2X2_1683 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_4__22_), .Y(_2863_) );
OR2X2 OR2X2_1684 ( .A(REGs_FIRQ_REGS_4__22_), .B(_1568__bF_buf14), .Y(_2864_) );
AND2X2 AND2X2_1821 ( .A(_2864_), .B(_2863_), .Y(_2865_) );
AND2X2 AND2X2_1822 ( .A(_2865_), .B(_1710__bF_buf3), .Y(_2866_) );
OR2X2 OR2X2_1685 ( .A(_2866_), .B(_2862_), .Y(_2867_) );
OR2X2 OR2X2_1686 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_6__22_), .Y(_2868_) );
OR2X2 OR2X2_1687 ( .A(REGs_FIRQ_REGS_6__22_), .B(_1568__bF_buf11), .Y(_2869_) );
AND2X2 AND2X2_1823 ( .A(_2869_), .B(_2868_), .Y(_2870_) );
AND2X2 AND2X2_1824 ( .A(_2870_), .B(_1716__bF_buf4), .Y(_2871_) );
OR2X2 OR2X2_1688 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_7__22_), .Y(_2872_) );
OR2X2 OR2X2_1689 ( .A(REGs_FIRQ_REGS_7__22_), .B(_1568__bF_buf0), .Y(_2873_) );
AND2X2 AND2X2_1825 ( .A(_2873_), .B(_2872_), .Y(_2874_) );
AND2X2 AND2X2_1826 ( .A(_2874_), .B(_1721__bF_buf0), .Y(_2875_) );
OR2X2 OR2X2_1690 ( .A(_2875_), .B(_2871_), .Y(_2876_) );
OR2X2 OR2X2_1691 ( .A(_2867_), .B(_2876_), .Y(_2877_) );
OR2X2 OR2X2_1692 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_0__22_), .Y(_2878_) );
OR2X2 OR2X2_1693 ( .A(REGs_FIRQ_REGS_0__22_), .B(_1568__bF_buf14), .Y(_2879_) );
AND2X2 AND2X2_1827 ( .A(_2879_), .B(_2878_), .Y(_2880_) );
AND2X2 AND2X2_1828 ( .A(_1730__bF_buf3), .B(_2880_), .Y(_2881_) );
OR2X2 OR2X2_1694 ( .A(INTERRUPT_flag_bF_buf13), .B(REGs_USR_REGS_1__22_), .Y(_2882_) );
OR2X2 OR2X2_1695 ( .A(REGs_FIRQ_REGS_1__22_), .B(_1568__bF_buf11), .Y(_2883_) );
AND2X2 AND2X2_1829 ( .A(_2883_), .B(_2882_), .Y(_2884_) );
AND2X2 AND2X2_1830 ( .A(_1735__bF_buf1), .B(_2884_), .Y(_2885_) );
OR2X2 OR2X2_1696 ( .A(_2881_), .B(_2885_), .Y(_2886_) );
OR2X2 OR2X2_1697 ( .A(INTERRUPT_flag_bF_buf0), .B(REGs_USR_REGS_3__22_), .Y(_2887_) );
OR2X2 OR2X2_1698 ( .A(REGs_FIRQ_REGS_3__22_), .B(_1568__bF_buf11), .Y(_2888_) );
AND2X2 AND2X2_1831 ( .A(_2888_), .B(_2887_), .Y(_2889_) );
AND2X2 AND2X2_1832 ( .A(_2889_), .B(_1741__bF_buf3), .Y(_2890_) );
OR2X2 OR2X2_1699 ( .A(INTERRUPT_flag_bF_buf15_bF_buf2), .B(REGs_USR_REGS_2__22_), .Y(_2891_) );
OR2X2 OR2X2_1700 ( .A(REGs_FIRQ_REGS_2__22_), .B(_1568__bF_buf11), .Y(_2892_) );
AND2X2 AND2X2_1833 ( .A(_2892_), .B(_2891_), .Y(_2893_) );
AND2X2 AND2X2_1834 ( .A(_1746__bF_buf1), .B(_2893_), .Y(_2894_) );
OR2X2 OR2X2_1701 ( .A(_2890_), .B(_2894_), .Y(_2895_) );
OR2X2 OR2X2_1702 ( .A(_2895_), .B(_2886_), .Y(_2896_) );
OR2X2 OR2X2_1703 ( .A(_2877_), .B(_2896_), .Y(_2897_) );
OR2X2 OR2X2_1704 ( .A(_2858_), .B(_2897_), .Y(REG_B_22_) );
AND2X2 AND2X2_1835 ( .A(_1678__bF_buf2), .B(REGs_REGS_4__23_), .Y(_2898_) );
AND2X2 AND2X2_1836 ( .A(_1682__bF_buf1), .B(REGs_REGS_5__23_), .Y(_2899_) );
OR2X2 OR2X2_1705 ( .A(_2898_), .B(_2899_), .Y(_2900_) );
AND2X2 AND2X2_1837 ( .A(_1687__bF_buf3), .B(REGs_REGS_6__23_), .Y(_2901_) );
AND2X2 AND2X2_1838 ( .A(_1690__bF_buf0), .B(REGs_REGS_7__23_), .Y(_2902_) );
OR2X2 OR2X2_1706 ( .A(_2902_), .B(_2901_), .Y(_2903_) );
OR2X2 OR2X2_1707 ( .A(_2900_), .B(_2903_), .Y(_2904_) );
AND2X2 AND2X2_1839 ( .A(_1695__bF_buf3), .B(gnd), .Y(_2905_) );
AND2X2 AND2X2_1840 ( .A(_1697__bF_buf1), .B(REGs_REGS_3__23_), .Y(_2906_) );
AND2X2 AND2X2_1841 ( .A(_1699__bF_buf3), .B(REGs_REGS_2__23_), .Y(_2907_) );
OR2X2 OR2X2_1708 ( .A(_2906_), .B(_2907_), .Y(_2908_) );
OR2X2 OR2X2_1709 ( .A(_2905_), .B(_2908_), .Y(_2909_) );
OR2X2 OR2X2_1710 ( .A(_2909_), .B(_2904_), .Y(_2910_) );
OR2X2 OR2X2_1711 ( .A(INTERRUPT_flag_bF_buf14_bF_buf0), .B(REGs_USR_REGS_5__23_), .Y(_2911_) );
OR2X2 OR2X2_1712 ( .A(REGs_FIRQ_REGS_5__23_), .B(_1568__bF_buf5), .Y(_2912_) );
AND2X2 AND2X2_1842 ( .A(_2912_), .B(_2911_), .Y(_2913_) );
AND2X2 AND2X2_1843 ( .A(_2913_), .B(_1705__bF_buf2), .Y(_2914_) );
OR2X2 OR2X2_1713 ( .A(INTERRUPT_flag_bF_buf13_bF_buf1), .B(REGs_USR_REGS_4__23_), .Y(_2915_) );
OR2X2 OR2X2_1714 ( .A(REGs_FIRQ_REGS_4__23_), .B(_1568__bF_buf5), .Y(_2916_) );
AND2X2 AND2X2_1844 ( .A(_2916_), .B(_2915_), .Y(_2917_) );
AND2X2 AND2X2_1845 ( .A(_2917_), .B(_1710__bF_buf1), .Y(_2918_) );
OR2X2 OR2X2_1715 ( .A(_2918_), .B(_2914_), .Y(_2919_) );
OR2X2 OR2X2_1716 ( .A(INTERRUPT_flag_bF_buf12_bF_buf3), .B(REGs_USR_REGS_6__23_), .Y(_2920_) );
OR2X2 OR2X2_1717 ( .A(REGs_FIRQ_REGS_6__23_), .B(_1568__bF_buf8), .Y(_2921_) );
AND2X2 AND2X2_1846 ( .A(_2921_), .B(_2920_), .Y(_2922_) );
AND2X2 AND2X2_1847 ( .A(_2922_), .B(_1716__bF_buf1), .Y(_2923_) );
OR2X2 OR2X2_1718 ( .A(INTERRUPT_flag_bF_buf11_bF_buf2), .B(REGs_USR_REGS_7__23_), .Y(_2924_) );
OR2X2 OR2X2_1719 ( .A(REGs_FIRQ_REGS_7__23_), .B(_1568__bF_buf8), .Y(_2925_) );
AND2X2 AND2X2_1848 ( .A(_2925_), .B(_2924_), .Y(_2926_) );
AND2X2 AND2X2_1849 ( .A(_2926_), .B(_1721__bF_buf1), .Y(_2927_) );
OR2X2 OR2X2_1720 ( .A(_2927_), .B(_2923_), .Y(_2928_) );
OR2X2 OR2X2_1721 ( .A(_2919_), .B(_2928_), .Y(_2929_) );
OR2X2 OR2X2_1722 ( .A(INTERRUPT_flag_bF_buf10_bF_buf0), .B(REGs_USR_REGS_0__23_), .Y(_2930_) );
OR2X2 OR2X2_1723 ( .A(REGs_FIRQ_REGS_0__23_), .B(_1568__bF_buf7), .Y(_2931_) );
AND2X2 AND2X2_1850 ( .A(_2931_), .B(_2930_), .Y(_2932_) );
AND2X2 AND2X2_1851 ( .A(_1730__bF_buf0), .B(_2932_), .Y(_2933_) );
OR2X2 OR2X2_1724 ( .A(INTERRUPT_flag_bF_buf9_bF_buf3), .B(REGs_USR_REGS_1__23_), .Y(_2934_) );
OR2X2 OR2X2_1725 ( .A(REGs_FIRQ_REGS_1__23_), .B(_1568__bF_buf3), .Y(_2935_) );
AND2X2 AND2X2_1852 ( .A(_2935_), .B(_2934_), .Y(_2936_) );
AND2X2 AND2X2_1853 ( .A(_1735__bF_buf3), .B(_2936_), .Y(_2937_) );
OR2X2 OR2X2_1726 ( .A(_2933_), .B(_2937_), .Y(_2938_) );
OR2X2 OR2X2_1727 ( .A(INTERRUPT_flag_bF_buf8_bF_buf2), .B(REGs_USR_REGS_3__23_), .Y(_2939_) );
OR2X2 OR2X2_1728 ( .A(REGs_FIRQ_REGS_3__23_), .B(_1568__bF_buf3), .Y(_2940_) );
AND2X2 AND2X2_1854 ( .A(_2940_), .B(_2939_), .Y(_2941_) );
AND2X2 AND2X2_1855 ( .A(_2941_), .B(_1741__bF_buf4), .Y(_2942_) );
OR2X2 OR2X2_1729 ( .A(INTERRUPT_flag_bF_buf7_bF_buf0), .B(REGs_USR_REGS_2__23_), .Y(_2943_) );
OR2X2 OR2X2_1730 ( .A(REGs_FIRQ_REGS_2__23_), .B(_1568__bF_buf15_bF_buf0), .Y(_2944_) );
AND2X2 AND2X2_1856 ( .A(_2944_), .B(_2943_), .Y(_2945_) );
AND2X2 AND2X2_1857 ( .A(_1746__bF_buf4), .B(_2945_), .Y(_2946_) );
OR2X2 OR2X2_1731 ( .A(_2942_), .B(_2946_), .Y(_2947_) );
OR2X2 OR2X2_1732 ( .A(_2947_), .B(_2938_), .Y(_2948_) );
OR2X2 OR2X2_1733 ( .A(_2929_), .B(_2948_), .Y(_2949_) );
OR2X2 OR2X2_1734 ( .A(_2910_), .B(_2949_), .Y(REG_B_23_) );
AND2X2 AND2X2_1858 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__24_), .Y(_2950_) );
AND2X2 AND2X2_1859 ( .A(_1682__bF_buf2), .B(REGs_REGS_5__24_), .Y(_2951_) );
OR2X2 OR2X2_1735 ( .A(_2950_), .B(_2951_), .Y(_2952_) );
AND2X2 AND2X2_1860 ( .A(_1687__bF_buf2), .B(REGs_REGS_6__24_), .Y(_2953_) );
AND2X2 AND2X2_1861 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__24_), .Y(_2954_) );
OR2X2 OR2X2_1736 ( .A(_2954_), .B(_2953_), .Y(_2955_) );
OR2X2 OR2X2_1737 ( .A(_2952_), .B(_2955_), .Y(_2956_) );
AND2X2 AND2X2_1862 ( .A(_1695__bF_buf4), .B(gnd), .Y(_2957_) );
AND2X2 AND2X2_1863 ( .A(_1697__bF_buf0), .B(REGs_REGS_3__24_), .Y(_2958_) );
AND2X2 AND2X2_1864 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__24_), .Y(_2959_) );
OR2X2 OR2X2_1738 ( .A(_2958_), .B(_2959_), .Y(_2960_) );
OR2X2 OR2X2_1739 ( .A(_2957_), .B(_2960_), .Y(_2961_) );
OR2X2 OR2X2_1740 ( .A(_2961_), .B(_2956_), .Y(_2962_) );
OR2X2 OR2X2_1741 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_5__24_), .Y(_2963_) );
OR2X2 OR2X2_1742 ( .A(REGs_FIRQ_REGS_5__24_), .B(_1568__bF_buf4), .Y(_2964_) );
AND2X2 AND2X2_1865 ( .A(_2964_), .B(_2963_), .Y(_2965_) );
AND2X2 AND2X2_1866 ( .A(_2965_), .B(_1705__bF_buf3), .Y(_2966_) );
OR2X2 OR2X2_1743 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_4__24_), .Y(_2967_) );
OR2X2 OR2X2_1744 ( .A(REGs_FIRQ_REGS_4__24_), .B(_1568__bF_buf2), .Y(_2968_) );
AND2X2 AND2X2_1867 ( .A(_2968_), .B(_2967_), .Y(_2969_) );
AND2X2 AND2X2_1868 ( .A(_2969_), .B(_1710__bF_buf4), .Y(_2970_) );
OR2X2 OR2X2_1745 ( .A(_2970_), .B(_2966_), .Y(_2971_) );
OR2X2 OR2X2_1746 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_6__24_), .Y(_2972_) );
OR2X2 OR2X2_1747 ( .A(REGs_FIRQ_REGS_6__24_), .B(_1568__bF_buf13), .Y(_2973_) );
AND2X2 AND2X2_1869 ( .A(_2973_), .B(_2972_), .Y(_2974_) );
AND2X2 AND2X2_1870 ( .A(_2974_), .B(_1716__bF_buf0), .Y(_2975_) );
OR2X2 OR2X2_1748 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_7__24_), .Y(_2976_) );
OR2X2 OR2X2_1749 ( .A(REGs_FIRQ_REGS_7__24_), .B(_1568__bF_buf4), .Y(_2977_) );
AND2X2 AND2X2_1871 ( .A(_2977_), .B(_2976_), .Y(_2978_) );
AND2X2 AND2X2_1872 ( .A(_2978_), .B(_1721__bF_buf2), .Y(_2979_) );
OR2X2 OR2X2_1750 ( .A(_2979_), .B(_2975_), .Y(_2980_) );
OR2X2 OR2X2_1751 ( .A(_2971_), .B(_2980_), .Y(_2981_) );
OR2X2 OR2X2_1752 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_0__24_), .Y(_2982_) );
OR2X2 OR2X2_1753 ( .A(REGs_FIRQ_REGS_0__24_), .B(_1568__bF_buf4), .Y(_2983_) );
AND2X2 AND2X2_1873 ( .A(_2983_), .B(_2982_), .Y(_2984_) );
AND2X2 AND2X2_1874 ( .A(_1730__bF_buf2), .B(_2984_), .Y(_2985_) );
OR2X2 OR2X2_1754 ( .A(INTERRUPT_flag_bF_buf2), .B(REGs_USR_REGS_1__24_), .Y(_2986_) );
OR2X2 OR2X2_1755 ( .A(REGs_FIRQ_REGS_1__24_), .B(_1568__bF_buf4), .Y(_2987_) );
AND2X2 AND2X2_1875 ( .A(_2987_), .B(_2986_), .Y(_2988_) );
AND2X2 AND2X2_1876 ( .A(_1735__bF_buf0), .B(_2988_), .Y(_2989_) );
OR2X2 OR2X2_1756 ( .A(_2985_), .B(_2989_), .Y(_2990_) );
OR2X2 OR2X2_1757 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_3__24_), .Y(_2991_) );
OR2X2 OR2X2_1758 ( .A(REGs_FIRQ_REGS_3__24_), .B(_1568__bF_buf6), .Y(_2992_) );
AND2X2 AND2X2_1877 ( .A(_2992_), .B(_2991_), .Y(_2993_) );
AND2X2 AND2X2_1878 ( .A(_2993_), .B(_1741__bF_buf1), .Y(_2994_) );
OR2X2 OR2X2_1759 ( .A(INTERRUPT_flag_bF_buf15_bF_buf3), .B(REGs_USR_REGS_2__24_), .Y(_2995_) );
OR2X2 OR2X2_1760 ( .A(REGs_FIRQ_REGS_2__24_), .B(_1568__bF_buf2), .Y(_2996_) );
AND2X2 AND2X2_1879 ( .A(_2996_), .B(_2995_), .Y(_2997_) );
AND2X2 AND2X2_1880 ( .A(_1746__bF_buf0), .B(_2997_), .Y(_2998_) );
OR2X2 OR2X2_1761 ( .A(_2994_), .B(_2998_), .Y(_2999_) );
OR2X2 OR2X2_1762 ( .A(_2999_), .B(_2990_), .Y(_3000_) );
OR2X2 OR2X2_1763 ( .A(_2981_), .B(_3000_), .Y(_3001_) );
OR2X2 OR2X2_1764 ( .A(_2962_), .B(_3001_), .Y(REG_B_24_) );
AND2X2 AND2X2_1881 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__25_), .Y(_3002_) );
AND2X2 AND2X2_1882 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__25_), .Y(_3003_) );
OR2X2 OR2X2_1765 ( .A(_3002_), .B(_3003_), .Y(_3004_) );
AND2X2 AND2X2_1883 ( .A(_1687__bF_buf1), .B(REGs_REGS_6__25_), .Y(_3005_) );
AND2X2 AND2X2_1884 ( .A(_1690__bF_buf2), .B(REGs_REGS_7__25_), .Y(_3006_) );
OR2X2 OR2X2_1766 ( .A(_3006_), .B(_3005_), .Y(_3007_) );
OR2X2 OR2X2_1767 ( .A(_3004_), .B(_3007_), .Y(_3008_) );
AND2X2 AND2X2_1885 ( .A(_1695__bF_buf0), .B(gnd), .Y(_3009_) );
AND2X2 AND2X2_1886 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__25_), .Y(_3010_) );
AND2X2 AND2X2_1887 ( .A(_1699__bF_buf0), .B(REGs_REGS_2__25_), .Y(_3011_) );
OR2X2 OR2X2_1768 ( .A(_3010_), .B(_3011_), .Y(_3012_) );
OR2X2 OR2X2_1769 ( .A(_3009_), .B(_3012_), .Y(_3013_) );
OR2X2 OR2X2_1770 ( .A(_3013_), .B(_3008_), .Y(_3014_) );
OR2X2 OR2X2_1771 ( .A(INTERRUPT_flag_bF_buf14_bF_buf0), .B(REGs_USR_REGS_5__25_), .Y(_3015_) );
OR2X2 OR2X2_1772 ( .A(REGs_FIRQ_REGS_5__25_), .B(_1568__bF_buf13), .Y(_3016_) );
AND2X2 AND2X2_1888 ( .A(_3016_), .B(_3015_), .Y(_3017_) );
AND2X2 AND2X2_1889 ( .A(_3017_), .B(_1705__bF_buf3), .Y(_3018_) );
OR2X2 OR2X2_1773 ( .A(INTERRUPT_flag_bF_buf13_bF_buf3), .B(REGs_USR_REGS_4__25_), .Y(_3019_) );
OR2X2 OR2X2_1774 ( .A(REGs_FIRQ_REGS_4__25_), .B(_1568__bF_buf2), .Y(_3020_) );
AND2X2 AND2X2_1890 ( .A(_3020_), .B(_3019_), .Y(_3021_) );
AND2X2 AND2X2_1891 ( .A(_3021_), .B(_1710__bF_buf4), .Y(_3022_) );
OR2X2 OR2X2_1775 ( .A(_3022_), .B(_3018_), .Y(_3023_) );
OR2X2 OR2X2_1776 ( .A(INTERRUPT_flag_bF_buf12_bF_buf0), .B(REGs_USR_REGS_6__25_), .Y(_3024_) );
OR2X2 OR2X2_1777 ( .A(REGs_FIRQ_REGS_6__25_), .B(_1568__bF_buf4), .Y(_3025_) );
AND2X2 AND2X2_1892 ( .A(_3025_), .B(_3024_), .Y(_3026_) );
AND2X2 AND2X2_1893 ( .A(_3026_), .B(_1716__bF_buf3), .Y(_3027_) );
OR2X2 OR2X2_1778 ( .A(INTERRUPT_flag_bF_buf11_bF_buf3), .B(REGs_USR_REGS_7__25_), .Y(_3028_) );
OR2X2 OR2X2_1779 ( .A(REGs_FIRQ_REGS_7__25_), .B(_1568__bF_buf4), .Y(_3029_) );
AND2X2 AND2X2_1894 ( .A(_3029_), .B(_3028_), .Y(_3030_) );
AND2X2 AND2X2_1895 ( .A(_3030_), .B(_1721__bF_buf3), .Y(_3031_) );
OR2X2 OR2X2_1780 ( .A(_3031_), .B(_3027_), .Y(_3032_) );
OR2X2 OR2X2_1781 ( .A(_3023_), .B(_3032_), .Y(_3033_) );
OR2X2 OR2X2_1782 ( .A(INTERRUPT_flag_bF_buf10_bF_buf2), .B(REGs_USR_REGS_0__25_), .Y(_3034_) );
OR2X2 OR2X2_1783 ( .A(REGs_FIRQ_REGS_0__25_), .B(_1568__bF_buf9), .Y(_3035_) );
AND2X2 AND2X2_1896 ( .A(_3035_), .B(_3034_), .Y(_3036_) );
AND2X2 AND2X2_1897 ( .A(_1730__bF_buf4), .B(_3036_), .Y(_3037_) );
OR2X2 OR2X2_1784 ( .A(INTERRUPT_flag_bF_buf9_bF_buf1), .B(REGs_USR_REGS_1__25_), .Y(_3038_) );
OR2X2 OR2X2_1785 ( .A(REGs_FIRQ_REGS_1__25_), .B(_1568__bF_buf2), .Y(_3039_) );
AND2X2 AND2X2_1898 ( .A(_3039_), .B(_3038_), .Y(_3040_) );
AND2X2 AND2X2_1899 ( .A(_1735__bF_buf4), .B(_3040_), .Y(_3041_) );
OR2X2 OR2X2_1786 ( .A(_3037_), .B(_3041_), .Y(_3042_) );
OR2X2 OR2X2_1787 ( .A(INTERRUPT_flag_bF_buf8_bF_buf3), .B(REGs_USR_REGS_3__25_), .Y(_3043_) );
OR2X2 OR2X2_1788 ( .A(REGs_FIRQ_REGS_3__25_), .B(_1568__bF_buf2), .Y(_3044_) );
AND2X2 AND2X2_1900 ( .A(_3044_), .B(_3043_), .Y(_3045_) );
AND2X2 AND2X2_1901 ( .A(_3045_), .B(_1741__bF_buf0), .Y(_3046_) );
OR2X2 OR2X2_1789 ( .A(INTERRUPT_flag_bF_buf7_bF_buf3), .B(REGs_USR_REGS_2__25_), .Y(_3047_) );
OR2X2 OR2X2_1790 ( .A(REGs_FIRQ_REGS_2__25_), .B(_1568__bF_buf15_bF_buf3), .Y(_3048_) );
AND2X2 AND2X2_1902 ( .A(_3048_), .B(_3047_), .Y(_3049_) );
AND2X2 AND2X2_1903 ( .A(_1746__bF_buf3), .B(_3049_), .Y(_3050_) );
OR2X2 OR2X2_1791 ( .A(_3046_), .B(_3050_), .Y(_3051_) );
OR2X2 OR2X2_1792 ( .A(_3051_), .B(_3042_), .Y(_3052_) );
OR2X2 OR2X2_1793 ( .A(_3033_), .B(_3052_), .Y(_3053_) );
OR2X2 OR2X2_1794 ( .A(_3014_), .B(_3053_), .Y(REG_B_25_) );
AND2X2 AND2X2_1904 ( .A(_1678__bF_buf0), .B(REGs_REGS_4__26_), .Y(_3054_) );
AND2X2 AND2X2_1905 ( .A(_1682__bF_buf3), .B(REGs_REGS_5__26_), .Y(_3055_) );
OR2X2 OR2X2_1795 ( .A(_3054_), .B(_3055_), .Y(_3056_) );
AND2X2 AND2X2_1906 ( .A(_1687__bF_buf4), .B(REGs_REGS_6__26_), .Y(_3057_) );
AND2X2 AND2X2_1907 ( .A(_1690__bF_buf3), .B(REGs_REGS_7__26_), .Y(_3058_) );
OR2X2 OR2X2_1796 ( .A(_3058_), .B(_3057_), .Y(_3059_) );
OR2X2 OR2X2_1797 ( .A(_3056_), .B(_3059_), .Y(_3060_) );
AND2X2 AND2X2_1908 ( .A(_1695__bF_buf2), .B(gnd), .Y(_3061_) );
AND2X2 AND2X2_1909 ( .A(_1697__bF_buf4), .B(REGs_REGS_3__26_), .Y(_3062_) );
AND2X2 AND2X2_1910 ( .A(_1699__bF_buf2), .B(REGs_REGS_2__26_), .Y(_3063_) );
OR2X2 OR2X2_1798 ( .A(_3062_), .B(_3063_), .Y(_3064_) );
OR2X2 OR2X2_1799 ( .A(_3061_), .B(_3064_), .Y(_3065_) );
OR2X2 OR2X2_1800 ( .A(_3065_), .B(_3060_), .Y(_3066_) );
OR2X2 OR2X2_1801 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_5__26_), .Y(_3067_) );
OR2X2 OR2X2_1802 ( .A(REGs_FIRQ_REGS_5__26_), .B(_1568__bF_buf0), .Y(_3068_) );
AND2X2 AND2X2_1911 ( .A(_3068_), .B(_3067_), .Y(_3069_) );
AND2X2 AND2X2_1912 ( .A(_3069_), .B(_1705__bF_buf4), .Y(_3070_) );
OR2X2 OR2X2_1803 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_4__26_), .Y(_3071_) );
OR2X2 OR2X2_1804 ( .A(REGs_FIRQ_REGS_4__26_), .B(_1568__bF_buf11), .Y(_3072_) );
AND2X2 AND2X2_1913 ( .A(_3072_), .B(_3071_), .Y(_3073_) );
AND2X2 AND2X2_1914 ( .A(_3073_), .B(_1710__bF_buf3), .Y(_3074_) );
OR2X2 OR2X2_1805 ( .A(_3074_), .B(_3070_), .Y(_3075_) );
OR2X2 OR2X2_1806 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_6__26_), .Y(_3076_) );
OR2X2 OR2X2_1807 ( .A(REGs_FIRQ_REGS_6__26_), .B(_1568__bF_buf11), .Y(_3077_) );
AND2X2 AND2X2_1915 ( .A(_3077_), .B(_3076_), .Y(_3078_) );
AND2X2 AND2X2_1916 ( .A(_3078_), .B(_1716__bF_buf4), .Y(_3079_) );
OR2X2 OR2X2_1808 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_7__26_), .Y(_3080_) );
OR2X2 OR2X2_1809 ( .A(REGs_FIRQ_REGS_7__26_), .B(_1568__bF_buf1), .Y(_3081_) );
AND2X2 AND2X2_1917 ( .A(_3081_), .B(_3080_), .Y(_3082_) );
AND2X2 AND2X2_1918 ( .A(_3082_), .B(_1721__bF_buf3), .Y(_3083_) );
OR2X2 OR2X2_1810 ( .A(_3083_), .B(_3079_), .Y(_3084_) );
OR2X2 OR2X2_1811 ( .A(_3075_), .B(_3084_), .Y(_3085_) );
OR2X2 OR2X2_1812 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_0__26_), .Y(_3086_) );
OR2X2 OR2X2_1813 ( .A(REGs_FIRQ_REGS_0__26_), .B(_1568__bF_buf9), .Y(_3087_) );
AND2X2 AND2X2_1919 ( .A(_3087_), .B(_3086_), .Y(_3088_) );
AND2X2 AND2X2_1920 ( .A(_1730__bF_buf3), .B(_3088_), .Y(_3089_) );
OR2X2 OR2X2_1814 ( .A(INTERRUPT_flag_bF_buf10), .B(REGs_USR_REGS_1__26_), .Y(_3090_) );
OR2X2 OR2X2_1815 ( .A(REGs_FIRQ_REGS_1__26_), .B(_1568__bF_buf11), .Y(_3091_) );
AND2X2 AND2X2_1921 ( .A(_3091_), .B(_3090_), .Y(_3092_) );
AND2X2 AND2X2_1922 ( .A(_1735__bF_buf4), .B(_3092_), .Y(_3093_) );
OR2X2 OR2X2_1816 ( .A(_3089_), .B(_3093_), .Y(_3094_) );
OR2X2 OR2X2_1817 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_3__26_), .Y(_3095_) );
OR2X2 OR2X2_1818 ( .A(REGs_FIRQ_REGS_3__26_), .B(_1568__bF_buf9), .Y(_3096_) );
AND2X2 AND2X2_1923 ( .A(_3096_), .B(_3095_), .Y(_3097_) );
AND2X2 AND2X2_1924 ( .A(_3097_), .B(_1741__bF_buf3), .Y(_3098_) );
OR2X2 OR2X2_1819 ( .A(INTERRUPT_flag_bF_buf15_bF_buf2), .B(REGs_USR_REGS_2__26_), .Y(_3099_) );
OR2X2 OR2X2_1820 ( .A(REGs_FIRQ_REGS_2__26_), .B(_1568__bF_buf9), .Y(_3100_) );
AND2X2 AND2X2_1925 ( .A(_3100_), .B(_3099_), .Y(_3101_) );
AND2X2 AND2X2_1926 ( .A(_1746__bF_buf1), .B(_3101_), .Y(_3102_) );
OR2X2 OR2X2_1821 ( .A(_3098_), .B(_3102_), .Y(_3103_) );
OR2X2 OR2X2_1822 ( .A(_3103_), .B(_3094_), .Y(_3104_) );
OR2X2 OR2X2_1823 ( .A(_3085_), .B(_3104_), .Y(_3105_) );
OR2X2 OR2X2_1824 ( .A(_3066_), .B(_3105_), .Y(REG_B_26_) );
AND2X2 AND2X2_1927 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__27_), .Y(_3106_) );
AND2X2 AND2X2_1928 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__27_), .Y(_3107_) );
OR2X2 OR2X2_1825 ( .A(_3106_), .B(_3107_), .Y(_3108_) );
AND2X2 AND2X2_1929 ( .A(_1687__bF_buf1), .B(REGs_REGS_6__27_), .Y(_3109_) );
AND2X2 AND2X2_1930 ( .A(_1690__bF_buf2), .B(REGs_REGS_7__27_), .Y(_3110_) );
OR2X2 OR2X2_1826 ( .A(_3110_), .B(_3109_), .Y(_3111_) );
OR2X2 OR2X2_1827 ( .A(_3108_), .B(_3111_), .Y(_3112_) );
AND2X2 AND2X2_1931 ( .A(_1695__bF_buf0), .B(gnd), .Y(_3113_) );
AND2X2 AND2X2_1932 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__27_), .Y(_3114_) );
AND2X2 AND2X2_1933 ( .A(_1699__bF_buf0), .B(REGs_REGS_2__27_), .Y(_3115_) );
OR2X2 OR2X2_1828 ( .A(_3114_), .B(_3115_), .Y(_3116_) );
OR2X2 OR2X2_1829 ( .A(_3113_), .B(_3116_), .Y(_3117_) );
OR2X2 OR2X2_1830 ( .A(_3117_), .B(_3112_), .Y(_3118_) );
OR2X2 OR2X2_1831 ( .A(INTERRUPT_flag_bF_buf14_bF_buf3), .B(REGs_USR_REGS_5__27_), .Y(_3119_) );
OR2X2 OR2X2_1832 ( .A(REGs_FIRQ_REGS_5__27_), .B(_1568__bF_buf0), .Y(_3120_) );
AND2X2 AND2X2_1934 ( .A(_3120_), .B(_3119_), .Y(_3121_) );
AND2X2 AND2X2_1935 ( .A(_3121_), .B(_1705__bF_buf3), .Y(_3122_) );
OR2X2 OR2X2_1833 ( .A(INTERRUPT_flag_bF_buf13_bF_buf0), .B(REGs_USR_REGS_4__27_), .Y(_3123_) );
OR2X2 OR2X2_1834 ( .A(REGs_FIRQ_REGS_4__27_), .B(_1568__bF_buf1), .Y(_3124_) );
AND2X2 AND2X2_1936 ( .A(_3124_), .B(_3123_), .Y(_3125_) );
AND2X2 AND2X2_1937 ( .A(_3125_), .B(_1710__bF_buf4), .Y(_3126_) );
OR2X2 OR2X2_1835 ( .A(_3126_), .B(_3122_), .Y(_3127_) );
OR2X2 OR2X2_1836 ( .A(INTERRUPT_flag_bF_buf12_bF_buf2), .B(REGs_USR_REGS_6__27_), .Y(_3128_) );
OR2X2 OR2X2_1837 ( .A(REGs_FIRQ_REGS_6__27_), .B(_1568__bF_buf11), .Y(_3129_) );
AND2X2 AND2X2_1938 ( .A(_3129_), .B(_3128_), .Y(_3130_) );
AND2X2 AND2X2_1939 ( .A(_3130_), .B(_1716__bF_buf3), .Y(_3131_) );
OR2X2 OR2X2_1838 ( .A(INTERRUPT_flag_bF_buf11_bF_buf1), .B(REGs_USR_REGS_7__27_), .Y(_3132_) );
OR2X2 OR2X2_1839 ( .A(REGs_FIRQ_REGS_7__27_), .B(_1568__bF_buf0), .Y(_3133_) );
AND2X2 AND2X2_1940 ( .A(_3133_), .B(_3132_), .Y(_3134_) );
AND2X2 AND2X2_1941 ( .A(_3134_), .B(_1721__bF_buf3), .Y(_3135_) );
OR2X2 OR2X2_1840 ( .A(_3135_), .B(_3131_), .Y(_3136_) );
OR2X2 OR2X2_1841 ( .A(_3127_), .B(_3136_), .Y(_3137_) );
OR2X2 OR2X2_1842 ( .A(INTERRUPT_flag_bF_buf10_bF_buf2), .B(REGs_USR_REGS_0__27_), .Y(_3138_) );
OR2X2 OR2X2_1843 ( .A(REGs_FIRQ_REGS_0__27_), .B(_1568__bF_buf9), .Y(_3139_) );
AND2X2 AND2X2_1942 ( .A(_3139_), .B(_3138_), .Y(_3140_) );
AND2X2 AND2X2_1943 ( .A(_1730__bF_buf4), .B(_3140_), .Y(_3141_) );
OR2X2 OR2X2_1844 ( .A(INTERRUPT_flag_bF_buf9_bF_buf1), .B(REGs_USR_REGS_1__27_), .Y(_3142_) );
OR2X2 OR2X2_1845 ( .A(REGs_FIRQ_REGS_1__27_), .B(_1568__bF_buf9), .Y(_3143_) );
AND2X2 AND2X2_1944 ( .A(_3143_), .B(_3142_), .Y(_3144_) );
AND2X2 AND2X2_1945 ( .A(_1735__bF_buf4), .B(_3144_), .Y(_3145_) );
OR2X2 OR2X2_1846 ( .A(_3141_), .B(_3145_), .Y(_3146_) );
OR2X2 OR2X2_1847 ( .A(INTERRUPT_flag_bF_buf8_bF_buf3), .B(REGs_USR_REGS_3__27_), .Y(_3147_) );
OR2X2 OR2X2_1848 ( .A(REGs_FIRQ_REGS_3__27_), .B(_1568__bF_buf2), .Y(_3148_) );
AND2X2 AND2X2_1946 ( .A(_3148_), .B(_3147_), .Y(_3149_) );
AND2X2 AND2X2_1947 ( .A(_3149_), .B(_1741__bF_buf0), .Y(_3150_) );
OR2X2 OR2X2_1849 ( .A(INTERRUPT_flag_bF_buf7_bF_buf3), .B(REGs_USR_REGS_2__27_), .Y(_3151_) );
OR2X2 OR2X2_1850 ( .A(REGs_FIRQ_REGS_2__27_), .B(_1568__bF_buf15_bF_buf3), .Y(_3152_) );
AND2X2 AND2X2_1948 ( .A(_3152_), .B(_3151_), .Y(_3153_) );
AND2X2 AND2X2_1949 ( .A(_1746__bF_buf3), .B(_3153_), .Y(_3154_) );
OR2X2 OR2X2_1851 ( .A(_3150_), .B(_3154_), .Y(_3155_) );
OR2X2 OR2X2_1852 ( .A(_3155_), .B(_3146_), .Y(_3156_) );
OR2X2 OR2X2_1853 ( .A(_3137_), .B(_3156_), .Y(_3157_) );
OR2X2 OR2X2_1854 ( .A(_3118_), .B(_3157_), .Y(REG_B_27_) );
AND2X2 AND2X2_1950 ( .A(_1678__bF_buf1), .B(REGs_REGS_4__28_), .Y(_3158_) );
AND2X2 AND2X2_1951 ( .A(_1682__bF_buf0), .B(REGs_REGS_5__28_), .Y(_3159_) );
OR2X2 OR2X2_1855 ( .A(_3158_), .B(_3159_), .Y(_3160_) );
AND2X2 AND2X2_1952 ( .A(_1687__bF_buf0), .B(REGs_REGS_6__28_), .Y(_3161_) );
AND2X2 AND2X2_1953 ( .A(_1690__bF_buf1), .B(REGs_REGS_7__28_), .Y(_3162_) );
OR2X2 OR2X2_1856 ( .A(_3162_), .B(_3161_), .Y(_3163_) );
OR2X2 OR2X2_1857 ( .A(_3160_), .B(_3163_), .Y(_3164_) );
AND2X2 AND2X2_1954 ( .A(_1695__bF_buf1), .B(gnd), .Y(_3165_) );
AND2X2 AND2X2_1955 ( .A(_1697__bF_buf2), .B(REGs_REGS_3__28_), .Y(_3166_) );
AND2X2 AND2X2_1956 ( .A(_1699__bF_buf1), .B(REGs_REGS_2__28_), .Y(_3167_) );
OR2X2 OR2X2_1858 ( .A(_3166_), .B(_3167_), .Y(_3168_) );
OR2X2 OR2X2_1859 ( .A(_3165_), .B(_3168_), .Y(_3169_) );
OR2X2 OR2X2_1860 ( .A(_3169_), .B(_3164_), .Y(_3170_) );
OR2X2 OR2X2_1861 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_5__28_), .Y(_3171_) );
OR2X2 OR2X2_1862 ( .A(REGs_FIRQ_REGS_5__28_), .B(_1568__bF_buf12), .Y(_3172_) );
AND2X2 AND2X2_1957 ( .A(_3172_), .B(_3171_), .Y(_3173_) );
AND2X2 AND2X2_1958 ( .A(_3173_), .B(_1705__bF_buf2), .Y(_3174_) );
OR2X2 OR2X2_1863 ( .A(INTERRUPT_flag_bF_buf14), .B(REGs_USR_REGS_4__28_), .Y(_3175_) );
OR2X2 OR2X2_1864 ( .A(REGs_FIRQ_REGS_4__28_), .B(_1568__bF_buf8), .Y(_3176_) );
AND2X2 AND2X2_1959 ( .A(_3176_), .B(_3175_), .Y(_3177_) );
AND2X2 AND2X2_1960 ( .A(_3177_), .B(_1710__bF_buf1), .Y(_3178_) );
OR2X2 OR2X2_1865 ( .A(_3178_), .B(_3174_), .Y(_3179_) );
OR2X2 OR2X2_1866 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_6__28_), .Y(_3180_) );
OR2X2 OR2X2_1867 ( .A(REGs_FIRQ_REGS_6__28_), .B(_1568__bF_buf8), .Y(_3181_) );
AND2X2 AND2X2_1961 ( .A(_3181_), .B(_3180_), .Y(_3182_) );
AND2X2 AND2X2_1962 ( .A(_3182_), .B(_1716__bF_buf1), .Y(_3183_) );
OR2X2 OR2X2_1868 ( .A(INTERRUPT_flag_bF_buf8), .B(REGs_USR_REGS_7__28_), .Y(_3184_) );
OR2X2 OR2X2_1869 ( .A(REGs_FIRQ_REGS_7__28_), .B(_1568__bF_buf8), .Y(_3185_) );
AND2X2 AND2X2_1963 ( .A(_3185_), .B(_3184_), .Y(_3186_) );
AND2X2 AND2X2_1964 ( .A(_3186_), .B(_1721__bF_buf1), .Y(_3187_) );
OR2X2 OR2X2_1870 ( .A(_3187_), .B(_3183_), .Y(_3188_) );
OR2X2 OR2X2_1871 ( .A(_3179_), .B(_3188_), .Y(_3189_) );
OR2X2 OR2X2_1872 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_0__28_), .Y(_3190_) );
OR2X2 OR2X2_1873 ( .A(REGs_FIRQ_REGS_0__28_), .B(_1568__bF_buf3), .Y(_3191_) );
AND2X2 AND2X2_1965 ( .A(_3191_), .B(_3190_), .Y(_3192_) );
AND2X2 AND2X2_1966 ( .A(_1730__bF_buf0), .B(_3192_), .Y(_3193_) );
OR2X2 OR2X2_1874 ( .A(INTERRUPT_flag_bF_buf4), .B(REGs_USR_REGS_1__28_), .Y(_3194_) );
OR2X2 OR2X2_1875 ( .A(REGs_FIRQ_REGS_1__28_), .B(_1568__bF_buf7), .Y(_3195_) );
AND2X2 AND2X2_1967 ( .A(_3195_), .B(_3194_), .Y(_3196_) );
AND2X2 AND2X2_1968 ( .A(_1735__bF_buf2), .B(_3196_), .Y(_3197_) );
OR2X2 OR2X2_1876 ( .A(_3193_), .B(_3197_), .Y(_3198_) );
OR2X2 OR2X2_1877 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_3__28_), .Y(_3199_) );
OR2X2 OR2X2_1878 ( .A(REGs_FIRQ_REGS_3__28_), .B(_1568__bF_buf3), .Y(_3200_) );
AND2X2 AND2X2_1969 ( .A(_3200_), .B(_3199_), .Y(_3201_) );
AND2X2 AND2X2_1970 ( .A(_3201_), .B(_1741__bF_buf4), .Y(_3202_) );
OR2X2 OR2X2_1879 ( .A(INTERRUPT_flag_bF_buf15_bF_buf3), .B(REGs_USR_REGS_2__28_), .Y(_3203_) );
OR2X2 OR2X2_1880 ( .A(REGs_FIRQ_REGS_2__28_), .B(_1568__bF_buf6), .Y(_3204_) );
AND2X2 AND2X2_1971 ( .A(_3204_), .B(_3203_), .Y(_3205_) );
AND2X2 AND2X2_1972 ( .A(_1746__bF_buf4), .B(_3205_), .Y(_3206_) );
OR2X2 OR2X2_1881 ( .A(_3202_), .B(_3206_), .Y(_3207_) );
OR2X2 OR2X2_1882 ( .A(_3207_), .B(_3198_), .Y(_3208_) );
OR2X2 OR2X2_1883 ( .A(_3189_), .B(_3208_), .Y(_3209_) );
OR2X2 OR2X2_1884 ( .A(_3170_), .B(_3209_), .Y(REG_B_28_) );
AND2X2 AND2X2_1973 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__29_), .Y(_3210_) );
AND2X2 AND2X2_1974 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__29_), .Y(_3211_) );
OR2X2 OR2X2_1885 ( .A(_3210_), .B(_3211_), .Y(_3212_) );
AND2X2 AND2X2_1975 ( .A(_1687__bF_buf2), .B(REGs_REGS_6__29_), .Y(_3213_) );
AND2X2 AND2X2_1976 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__29_), .Y(_3214_) );
OR2X2 OR2X2_1886 ( .A(_3214_), .B(_3213_), .Y(_3215_) );
OR2X2 OR2X2_1887 ( .A(_3212_), .B(_3215_), .Y(_3216_) );
AND2X2 AND2X2_1977 ( .A(_1695__bF_buf4), .B(gnd), .Y(_3217_) );
AND2X2 AND2X2_1978 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__29_), .Y(_3218_) );
AND2X2 AND2X2_1979 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__29_), .Y(_3219_) );
OR2X2 OR2X2_1888 ( .A(_3218_), .B(_3219_), .Y(_3220_) );
OR2X2 OR2X2_1889 ( .A(_3217_), .B(_3220_), .Y(_3221_) );
OR2X2 OR2X2_1890 ( .A(_3221_), .B(_3216_), .Y(_3222_) );
OR2X2 OR2X2_1891 ( .A(INTERRUPT_flag_bF_buf14_bF_buf2), .B(REGs_USR_REGS_5__29_), .Y(_3223_) );
OR2X2 OR2X2_1892 ( .A(REGs_FIRQ_REGS_5__29_), .B(_1568__bF_buf13), .Y(_3224_) );
AND2X2 AND2X2_1980 ( .A(_3224_), .B(_3223_), .Y(_3225_) );
AND2X2 AND2X2_1981 ( .A(_3225_), .B(_1705__bF_buf0), .Y(_3226_) );
OR2X2 OR2X2_1893 ( .A(INTERRUPT_flag_bF_buf13_bF_buf3), .B(REGs_USR_REGS_4__29_), .Y(_3227_) );
OR2X2 OR2X2_1894 ( .A(REGs_FIRQ_REGS_4__29_), .B(_1568__bF_buf6), .Y(_3228_) );
AND2X2 AND2X2_1982 ( .A(_3228_), .B(_3227_), .Y(_3229_) );
AND2X2 AND2X2_1983 ( .A(_3229_), .B(_1710__bF_buf2), .Y(_3230_) );
OR2X2 OR2X2_1895 ( .A(_3230_), .B(_3226_), .Y(_3231_) );
OR2X2 OR2X2_1896 ( .A(INTERRUPT_flag_bF_buf12_bF_buf0), .B(REGs_USR_REGS_6__29_), .Y(_3232_) );
OR2X2 OR2X2_1897 ( .A(REGs_FIRQ_REGS_6__29_), .B(_1568__bF_buf4), .Y(_3233_) );
AND2X2 AND2X2_1984 ( .A(_3233_), .B(_3232_), .Y(_3234_) );
AND2X2 AND2X2_1985 ( .A(_3234_), .B(_1716__bF_buf3), .Y(_3235_) );
OR2X2 OR2X2_1898 ( .A(INTERRUPT_flag_bF_buf11_bF_buf3), .B(REGs_USR_REGS_7__29_), .Y(_3236_) );
OR2X2 OR2X2_1899 ( .A(REGs_FIRQ_REGS_7__29_), .B(_1568__bF_buf13), .Y(_3237_) );
AND2X2 AND2X2_1986 ( .A(_3237_), .B(_3236_), .Y(_3238_) );
AND2X2 AND2X2_1987 ( .A(_3238_), .B(_1721__bF_buf2), .Y(_3239_) );
OR2X2 OR2X2_1900 ( .A(_3239_), .B(_3235_), .Y(_3240_) );
OR2X2 OR2X2_1901 ( .A(_3231_), .B(_3240_), .Y(_3241_) );
OR2X2 OR2X2_1902 ( .A(INTERRUPT_flag_bF_buf10_bF_buf3), .B(REGs_USR_REGS_0__29_), .Y(_3242_) );
OR2X2 OR2X2_1903 ( .A(REGs_FIRQ_REGS_0__29_), .B(_1568__bF_buf6), .Y(_3243_) );
AND2X2 AND2X2_1988 ( .A(_3243_), .B(_3242_), .Y(_3244_) );
AND2X2 AND2X2_1989 ( .A(_1730__bF_buf2), .B(_3244_), .Y(_3245_) );
OR2X2 OR2X2_1904 ( .A(INTERRUPT_flag_bF_buf9_bF_buf2), .B(REGs_USR_REGS_1__29_), .Y(_3246_) );
OR2X2 OR2X2_1905 ( .A(REGs_FIRQ_REGS_1__29_), .B(_1568__bF_buf4), .Y(_3247_) );
AND2X2 AND2X2_1990 ( .A(_3247_), .B(_3246_), .Y(_3248_) );
AND2X2 AND2X2_1991 ( .A(_1735__bF_buf0), .B(_3248_), .Y(_3249_) );
OR2X2 OR2X2_1906 ( .A(_3245_), .B(_3249_), .Y(_3250_) );
OR2X2 OR2X2_1907 ( .A(INTERRUPT_flag_bF_buf8_bF_buf0), .B(REGs_USR_REGS_3__29_), .Y(_3251_) );
OR2X2 OR2X2_1908 ( .A(REGs_FIRQ_REGS_3__29_), .B(_1568__bF_buf6), .Y(_3252_) );
AND2X2 AND2X2_1992 ( .A(_3252_), .B(_3251_), .Y(_3253_) );
AND2X2 AND2X2_1993 ( .A(_3253_), .B(_1741__bF_buf1), .Y(_3254_) );
OR2X2 OR2X2_1909 ( .A(INTERRUPT_flag_bF_buf7_bF_buf2), .B(REGs_USR_REGS_2__29_), .Y(_3255_) );
OR2X2 OR2X2_1910 ( .A(REGs_FIRQ_REGS_2__29_), .B(_1568__bF_buf15_bF_buf2), .Y(_3256_) );
AND2X2 AND2X2_1994 ( .A(_3256_), .B(_3255_), .Y(_3257_) );
AND2X2 AND2X2_1995 ( .A(_1746__bF_buf0), .B(_3257_), .Y(_3258_) );
OR2X2 OR2X2_1911 ( .A(_3254_), .B(_3258_), .Y(_3259_) );
OR2X2 OR2X2_1912 ( .A(_3259_), .B(_3250_), .Y(_3260_) );
OR2X2 OR2X2_1913 ( .A(_3241_), .B(_3260_), .Y(_3261_) );
OR2X2 OR2X2_1914 ( .A(_3222_), .B(_3261_), .Y(REG_B_29_) );
AND2X2 AND2X2_1996 ( .A(_1678__bF_buf3), .B(REGs_REGS_4__30_), .Y(_3262_) );
AND2X2 AND2X2_1997 ( .A(_1682__bF_buf4), .B(REGs_REGS_5__30_), .Y(_3263_) );
OR2X2 OR2X2_1915 ( .A(_3262_), .B(_3263_), .Y(_3264_) );
AND2X2 AND2X2_1998 ( .A(_1687__bF_buf1), .B(REGs_REGS_6__30_), .Y(_3265_) );
AND2X2 AND2X2_1999 ( .A(_1690__bF_buf2), .B(REGs_REGS_7__30_), .Y(_3266_) );
OR2X2 OR2X2_1916 ( .A(_3266_), .B(_3265_), .Y(_3267_) );
OR2X2 OR2X2_1917 ( .A(_3264_), .B(_3267_), .Y(_3268_) );
AND2X2 AND2X2_2000 ( .A(_1695__bF_buf0), .B(gnd), .Y(_3269_) );
AND2X2 AND2X2_2001 ( .A(_1697__bF_buf3), .B(REGs_REGS_3__30_), .Y(_3270_) );
AND2X2 AND2X2_2002 ( .A(_1699__bF_buf0), .B(REGs_REGS_2__30_), .Y(_3271_) );
OR2X2 OR2X2_1918 ( .A(_3270_), .B(_3271_), .Y(_3272_) );
OR2X2 OR2X2_1919 ( .A(_3269_), .B(_3272_), .Y(_3273_) );
OR2X2 OR2X2_1920 ( .A(_3273_), .B(_3268_), .Y(_3274_) );
OR2X2 OR2X2_1921 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_5__30_), .Y(_3275_) );
OR2X2 OR2X2_1922 ( .A(REGs_FIRQ_REGS_5__30_), .B(_1568__bF_buf0), .Y(_3276_) );
AND2X2 AND2X2_2003 ( .A(_3276_), .B(_3275_), .Y(_3277_) );
AND2X2 AND2X2_2004 ( .A(_3277_), .B(_1705__bF_buf3), .Y(_3278_) );
OR2X2 OR2X2_1923 ( .A(INTERRUPT_flag_bF_buf7), .B(REGs_USR_REGS_4__30_), .Y(_3279_) );
OR2X2 OR2X2_1924 ( .A(REGs_FIRQ_REGS_4__30_), .B(_1568__bF_buf1), .Y(_3280_) );
AND2X2 AND2X2_2005 ( .A(_3280_), .B(_3279_), .Y(_3281_) );
AND2X2 AND2X2_2006 ( .A(_3281_), .B(_1710__bF_buf4), .Y(_3282_) );
OR2X2 OR2X2_1925 ( .A(_3282_), .B(_3278_), .Y(_3283_) );
OR2X2 OR2X2_1926 ( .A(INTERRUPT_flag_bF_buf6), .B(REGs_USR_REGS_6__30_), .Y(_3284_) );
OR2X2 OR2X2_1927 ( .A(REGs_FIRQ_REGS_6__30_), .B(_1568__bF_buf9), .Y(_3285_) );
AND2X2 AND2X2_2007 ( .A(_3285_), .B(_3284_), .Y(_3286_) );
AND2X2 AND2X2_2008 ( .A(_3286_), .B(_1716__bF_buf3), .Y(_3287_) );
OR2X2 OR2X2_1928 ( .A(INTERRUPT_flag_bF_buf3), .B(REGs_USR_REGS_7__30_), .Y(_3288_) );
OR2X2 OR2X2_1929 ( .A(REGs_FIRQ_REGS_7__30_), .B(_1568__bF_buf1), .Y(_3289_) );
AND2X2 AND2X2_2009 ( .A(_3289_), .B(_3288_), .Y(_3290_) );
AND2X2 AND2X2_2010 ( .A(_3290_), .B(_1721__bF_buf3), .Y(_3291_) );
OR2X2 OR2X2_1930 ( .A(_3291_), .B(_3287_), .Y(_3292_) );
OR2X2 OR2X2_1931 ( .A(_3283_), .B(_3292_), .Y(_3293_) );
OR2X2 OR2X2_1932 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_0__30_), .Y(_3294_) );
OR2X2 OR2X2_1933 ( .A(REGs_FIRQ_REGS_0__30_), .B(_1568__bF_buf0), .Y(_3295_) );
AND2X2 AND2X2_2011 ( .A(_3295_), .B(_3294_), .Y(_3296_) );
AND2X2 AND2X2_2012 ( .A(_1730__bF_buf4), .B(_3296_), .Y(_3297_) );
OR2X2 OR2X2_1934 ( .A(INTERRUPT_flag_bF_buf7), .B(REGs_USR_REGS_1__30_), .Y(_3298_) );
OR2X2 OR2X2_1935 ( .A(REGs_FIRQ_REGS_1__30_), .B(_1568__bF_buf1), .Y(_3299_) );
AND2X2 AND2X2_2013 ( .A(_3299_), .B(_3298_), .Y(_3300_) );
AND2X2 AND2X2_2014 ( .A(_1735__bF_buf4), .B(_3300_), .Y(_3301_) );
OR2X2 OR2X2_1936 ( .A(_3297_), .B(_3301_), .Y(_3302_) );
OR2X2 OR2X2_1937 ( .A(INTERRUPT_flag_bF_buf1), .B(REGs_USR_REGS_3__30_), .Y(_3303_) );
OR2X2 OR2X2_1938 ( .A(REGs_FIRQ_REGS_3__30_), .B(_1568__bF_buf1), .Y(_3304_) );
AND2X2 AND2X2_2015 ( .A(_3304_), .B(_3303_), .Y(_3305_) );
AND2X2 AND2X2_2016 ( .A(_3305_), .B(_1741__bF_buf1), .Y(_3306_) );
OR2X2 OR2X2_1939 ( .A(INTERRUPT_flag_bF_buf15_bF_buf1), .B(REGs_USR_REGS_2__30_), .Y(_3307_) );
OR2X2 OR2X2_1940 ( .A(REGs_FIRQ_REGS_2__30_), .B(_1568__bF_buf1), .Y(_3308_) );
AND2X2 AND2X2_2017 ( .A(_3308_), .B(_3307_), .Y(_3309_) );
AND2X2 AND2X2_2018 ( .A(_1746__bF_buf3), .B(_3309_), .Y(_3310_) );
OR2X2 OR2X2_1941 ( .A(_3306_), .B(_3310_), .Y(_3311_) );
OR2X2 OR2X2_1942 ( .A(_3311_), .B(_3302_), .Y(_3312_) );
OR2X2 OR2X2_1943 ( .A(_3293_), .B(_3312_), .Y(_3313_) );
OR2X2 OR2X2_1944 ( .A(_3274_), .B(_3313_), .Y(REG_B_30_) );
AND2X2 AND2X2_2019 ( .A(_1678__bF_buf4), .B(REGs_REGS_4__31_), .Y(_3314_) );
AND2X2 AND2X2_2020 ( .A(_1682__bF_buf2), .B(REGs_REGS_5__31_), .Y(_3315_) );
OR2X2 OR2X2_1945 ( .A(_3314_), .B(_3315_), .Y(_3316_) );
AND2X2 AND2X2_2021 ( .A(_1687__bF_buf2), .B(REGs_REGS_6__31_), .Y(_3317_) );
AND2X2 AND2X2_2022 ( .A(_1690__bF_buf4), .B(REGs_REGS_7__31_), .Y(_3318_) );
OR2X2 OR2X2_1946 ( .A(_3318_), .B(_3317_), .Y(_3319_) );
OR2X2 OR2X2_1947 ( .A(_3316_), .B(_3319_), .Y(_3320_) );
AND2X2 AND2X2_2023 ( .A(_1695__bF_buf4), .B(gnd), .Y(_3321_) );
AND2X2 AND2X2_2024 ( .A(_1697__bF_buf0), .B(REGs_REGS_3__31_), .Y(_3322_) );
AND2X2 AND2X2_2025 ( .A(_1699__bF_buf4), .B(REGs_REGS_2__31_), .Y(_3323_) );
OR2X2 OR2X2_1948 ( .A(_3322_), .B(_3323_), .Y(_3324_) );
OR2X2 OR2X2_1949 ( .A(_3321_), .B(_3324_), .Y(_3325_) );
OR2X2 OR2X2_1950 ( .A(_3325_), .B(_3320_), .Y(_3326_) );
OR2X2 OR2X2_1951 ( .A(INTERRUPT_flag_bF_buf14_bF_buf1), .B(REGs_USR_REGS_5__31_), .Y(_3327_) );
OR2X2 OR2X2_1952 ( .A(REGs_FIRQ_REGS_5__31_), .B(_1568__bF_buf12), .Y(_3328_) );
AND2X2 AND2X2_2026 ( .A(_3328_), .B(_3327_), .Y(_3329_) );
AND2X2 AND2X2_2027 ( .A(_3329_), .B(_1705__bF_buf2), .Y(_3330_) );
OR2X2 OR2X2_1953 ( .A(INTERRUPT_flag_bF_buf13_bF_buf2), .B(REGs_USR_REGS_4__31_), .Y(_3331_) );
OR2X2 OR2X2_1954 ( .A(REGs_FIRQ_REGS_4__31_), .B(_1568__bF_buf12), .Y(_3332_) );
AND2X2 AND2X2_2028 ( .A(_3332_), .B(_3331_), .Y(_3333_) );
AND2X2 AND2X2_2029 ( .A(_3333_), .B(_1710__bF_buf1), .Y(_3334_) );
OR2X2 OR2X2_1955 ( .A(_3334_), .B(_3330_), .Y(_3335_) );
OR2X2 OR2X2_1956 ( .A(INTERRUPT_flag_bF_buf12_bF_buf3), .B(REGs_USR_REGS_6__31_), .Y(_3336_) );
OR2X2 OR2X2_1957 ( .A(REGs_FIRQ_REGS_6__31_), .B(_1568__bF_buf3), .Y(_3337_) );
AND2X2 AND2X2_2030 ( .A(_3337_), .B(_3336_), .Y(_3338_) );
AND2X2 AND2X2_2031 ( .A(_3338_), .B(_1716__bF_buf1), .Y(_3339_) );
OR2X2 OR2X2_1958 ( .A(INTERRUPT_flag_bF_buf11_bF_buf0), .B(REGs_USR_REGS_7__31_), .Y(_3340_) );
OR2X2 OR2X2_1959 ( .A(REGs_FIRQ_REGS_7__31_), .B(_1568__bF_buf3), .Y(_3341_) );
AND2X2 AND2X2_2032 ( .A(_3341_), .B(_3340_), .Y(_3342_) );
AND2X2 AND2X2_2033 ( .A(_3342_), .B(_1721__bF_buf1), .Y(_3343_) );
OR2X2 OR2X2_1960 ( .A(_3343_), .B(_3339_), .Y(_3344_) );
OR2X2 OR2X2_1961 ( .A(_3335_), .B(_3344_), .Y(_3345_) );
OR2X2 OR2X2_1962 ( .A(INTERRUPT_flag_bF_buf10_bF_buf1), .B(REGs_USR_REGS_0__31_), .Y(_3346_) );
OR2X2 OR2X2_1963 ( .A(REGs_FIRQ_REGS_0__31_), .B(_1568__bF_buf4), .Y(_3347_) );
AND2X2 AND2X2_2034 ( .A(_3347_), .B(_3346_), .Y(_3348_) );
AND2X2 AND2X2_2035 ( .A(_1730__bF_buf2), .B(_3348_), .Y(_3349_) );
OR2X2 OR2X2_1964 ( .A(INTERRUPT_flag_bF_buf9_bF_buf0), .B(REGs_USR_REGS_1__31_), .Y(_3350_) );
OR2X2 OR2X2_1965 ( .A(REGs_FIRQ_REGS_1__31_), .B(_1568__bF_buf4), .Y(_3351_) );
AND2X2 AND2X2_2036 ( .A(_3351_), .B(_3350_), .Y(_3352_) );
AND2X2 AND2X2_2037 ( .A(_1735__bF_buf0), .B(_3352_), .Y(_3353_) );
OR2X2 OR2X2_1966 ( .A(_3349_), .B(_3353_), .Y(_3354_) );
OR2X2 OR2X2_1967 ( .A(INTERRUPT_flag_bF_buf8_bF_buf0), .B(REGs_USR_REGS_3__31_), .Y(_3355_) );
OR2X2 OR2X2_1968 ( .A(REGs_FIRQ_REGS_3__31_), .B(_1568__bF_buf6), .Y(_3356_) );
AND2X2 AND2X2_2038 ( .A(_3356_), .B(_3355_), .Y(_3357_) );
AND2X2 AND2X2_2039 ( .A(_3357_), .B(_1741__bF_buf1), .Y(_3358_) );
OR2X2 OR2X2_1969 ( .A(INTERRUPT_flag_bF_buf7_bF_buf2), .B(REGs_USR_REGS_2__31_), .Y(_3359_) );
OR2X2 OR2X2_1970 ( .A(REGs_FIRQ_REGS_2__31_), .B(_1568__bF_buf15_bF_buf2), .Y(_3360_) );
AND2X2 AND2X2_2040 ( .A(_3360_), .B(_3359_), .Y(_3361_) );
AND2X2 AND2X2_2041 ( .A(_1746__bF_buf0), .B(_3361_), .Y(_3362_) );
OR2X2 OR2X2_1971 ( .A(_3358_), .B(_3362_), .Y(_3363_) );
OR2X2 OR2X2_1972 ( .A(_3363_), .B(_3354_), .Y(_3364_) );
OR2X2 OR2X2_1973 ( .A(_3345_), .B(_3364_), .Y(_3365_) );
OR2X2 OR2X2_1974 ( .A(_3326_), .B(_3365_), .Y(REG_B_31_) );
INVX1 INVX1_327 ( .A(CORE_REG_RF1_3_), .Y(_3366_) );
AND2X2 AND2X2_2042 ( .A(_3366_), .B(CORE_REG_RF1_2_), .Y(_3367_) );
NOR2X1 NOR2X1_177 ( .A(CORE_REG_RF1_1_), .B(CORE_REG_RF1_0_), .Y(_3368_) );
AND2X2 AND2X2_2043 ( .A(_3367_), .B(_3368_), .Y(_3369_) );
AND2X2 AND2X2_2044 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__0_), .Y(_3370_) );
INVX1 INVX1_328 ( .A(CORE_REG_RF1_1_), .Y(_3371_) );
AND2X2 AND2X2_2045 ( .A(_3371_), .B(CORE_REG_RF1_0_), .Y(_3372_) );
AND2X2 AND2X2_2046 ( .A(_3367_), .B(_3372_), .Y(_3373_) );
AND2X2 AND2X2_2047 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__0_), .Y(_3374_) );
OR2X2 OR2X2_1975 ( .A(_3370_), .B(_3374_), .Y(_3375_) );
INVX1 INVX1_329 ( .A(CORE_REG_RF1_0_), .Y(_3376_) );
AND2X2 AND2X2_2048 ( .A(_3376_), .B(CORE_REG_RF1_1_), .Y(_3377_) );
AND2X2 AND2X2_2049 ( .A(_3367_), .B(_3377_), .Y(_3378_) );
AND2X2 AND2X2_2050 ( .A(_3378__bF_buf1), .B(REGs_REGS_6__0_), .Y(_3379_) );
AND2X2 AND2X2_2051 ( .A(CORE_REG_RF1_1_), .B(CORE_REG_RF1_0_), .Y(_3380_) );
AND2X2 AND2X2_2052 ( .A(_3367_), .B(_3380_), .Y(_3381_) );
AND2X2 AND2X2_2053 ( .A(_3381__bF_buf0), .B(REGs_REGS_7__0_), .Y(_3382_) );
OR2X2 OR2X2_1976 ( .A(_3382_), .B(_3379_), .Y(_3383_) );
OR2X2 OR2X2_1977 ( .A(_3375_), .B(_3383_), .Y(_3384_) );
NOR2X1 NOR2X1_178 ( .A(CORE_REG_RF1_3_), .B(CORE_REG_RF1_2_), .Y(_3385_) );
AND2X2 AND2X2_2054 ( .A(_3372_), .B(_3385_), .Y(_3386_) );
AND2X2 AND2X2_2055 ( .A(_3386__bF_buf1), .B(PC_ADDR_stack_1__0_), .Y(_3387_) );
AND2X2 AND2X2_2056 ( .A(_3385_), .B(_3380_), .Y(_3388_) );
AND2X2 AND2X2_2057 ( .A(_3388__bF_buf0), .B(REGs_REGS_3__0_), .Y(_3389_) );
AND2X2 AND2X2_2058 ( .A(_3377_), .B(_3385_), .Y(_3390_) );
AND2X2 AND2X2_2059 ( .A(_3390__bF_buf2), .B(REGs_REGS_2__0_), .Y(_3391_) );
OR2X2 OR2X2_1978 ( .A(_3389_), .B(_3391_), .Y(_3392_) );
OR2X2 OR2X2_1979 ( .A(_3387_), .B(_3392_), .Y(_3393_) );
OR2X2 OR2X2_1980 ( .A(_3393_), .B(_3384_), .Y(_3394_) );
AND2X2 AND2X2_2060 ( .A(CORE_REG_RF1_3_), .B(CORE_REG_RF1_2_), .Y(_3395_) );
AND2X2 AND2X2_2061 ( .A(_3372_), .B(_3395_), .Y(_3396_) );
AND2X2 AND2X2_2062 ( .A(_1708_), .B(_3396__bF_buf4), .Y(_3397_) );
AND2X2 AND2X2_2063 ( .A(_3368_), .B(_3395_), .Y(_3398_) );
AND2X2 AND2X2_2064 ( .A(_1713_), .B(_3398__bF_buf2), .Y(_3399_) );
OR2X2 OR2X2_1981 ( .A(_3399_), .B(_3397_), .Y(_3400_) );
AND2X2 AND2X2_2065 ( .A(_3377_), .B(_3395_), .Y(_3401_) );
AND2X2 AND2X2_2066 ( .A(_1719_), .B(_3401__bF_buf2), .Y(_3402_) );
AND2X2 AND2X2_2067 ( .A(_3380_), .B(_3395_), .Y(_3403_) );
AND2X2 AND2X2_2068 ( .A(_1724_), .B(_3403__bF_buf0), .Y(_3404_) );
OR2X2 OR2X2_1982 ( .A(_3404_), .B(_3402_), .Y(_3405_) );
OR2X2 OR2X2_1983 ( .A(_3400_), .B(_3405_), .Y(_3406_) );
INVX1 INVX1_330 ( .A(CORE_REG_RF1_2_), .Y(_3407_) );
AND2X2 AND2X2_2069 ( .A(_3407_), .B(CORE_REG_RF1_3_), .Y(_3408_) );
AND2X2 AND2X2_2070 ( .A(_3408_), .B(_3368_), .Y(_3409_) );
AND2X2 AND2X2_2071 ( .A(_3409__bF_buf0), .B(_1733_), .Y(_3410_) );
AND2X2 AND2X2_2072 ( .A(_3372_), .B(_3408_), .Y(_3411_) );
AND2X2 AND2X2_2073 ( .A(_3411__bF_buf4), .B(_1738_), .Y(_3412_) );
OR2X2 OR2X2_1984 ( .A(_3410_), .B(_3412_), .Y(_3413_) );
AND2X2 AND2X2_2074 ( .A(_3408_), .B(_3380_), .Y(_3414_) );
AND2X2 AND2X2_2075 ( .A(_1744_), .B(_3414__bF_buf0), .Y(_3415_) );
AND2X2 AND2X2_2076 ( .A(_3408_), .B(_3377_), .Y(_3416_) );
AND2X2 AND2X2_2077 ( .A(_3416__bF_buf1), .B(_1749_), .Y(_3417_) );
OR2X2 OR2X2_1985 ( .A(_3415_), .B(_3417_), .Y(_3418_) );
OR2X2 OR2X2_1986 ( .A(_3418_), .B(_3413_), .Y(_3419_) );
OR2X2 OR2X2_1987 ( .A(_3406_), .B(_3419_), .Y(_3420_) );
OR2X2 OR2X2_1988 ( .A(_3394_), .B(_3420_), .Y(REG_A_0_) );
AND2X2 AND2X2_2078 ( .A(_3369__bF_buf0), .B(REGs_REGS_4__1_), .Y(_3421_) );
AND2X2 AND2X2_2079 ( .A(_3373__bF_buf3), .B(REGs_REGS_5__1_), .Y(_3422_) );
OR2X2 OR2X2_1989 ( .A(_3421_), .B(_3422_), .Y(_3423_) );
AND2X2 AND2X2_2080 ( .A(_3378__bF_buf1), .B(REGs_REGS_6__1_), .Y(_3424_) );
AND2X2 AND2X2_2081 ( .A(_3381__bF_buf0), .B(REGs_REGS_7__1_), .Y(_3425_) );
OR2X2 OR2X2_1990 ( .A(_3425_), .B(_3424_), .Y(_3426_) );
OR2X2 OR2X2_1991 ( .A(_3423_), .B(_3426_), .Y(_3427_) );
AND2X2 AND2X2_2082 ( .A(_3386__bF_buf1), .B(PC_ADDR_stack_1__1_), .Y(_3428_) );
AND2X2 AND2X2_2083 ( .A(_3388__bF_buf0), .B(REGs_REGS_3__1_), .Y(_3429_) );
AND2X2 AND2X2_2084 ( .A(_3390__bF_buf2), .B(REGs_REGS_2__1_), .Y(_3430_) );
OR2X2 OR2X2_1992 ( .A(_3429_), .B(_3430_), .Y(_3431_) );
OR2X2 OR2X2_1993 ( .A(_3428_), .B(_3431_), .Y(_3432_) );
OR2X2 OR2X2_1994 ( .A(_3432_), .B(_3427_), .Y(_3433_) );
AND2X2 AND2X2_2085 ( .A(_1769_), .B(_3396__bF_buf0), .Y(_3434_) );
AND2X2 AND2X2_2086 ( .A(_1773_), .B(_3398__bF_buf4), .Y(_3435_) );
OR2X2 OR2X2_1995 ( .A(_3435_), .B(_3434_), .Y(_3436_) );
AND2X2 AND2X2_2087 ( .A(_1778_), .B(_3401__bF_buf4), .Y(_3437_) );
AND2X2 AND2X2_2088 ( .A(_1782_), .B(_3403__bF_buf1), .Y(_3438_) );
OR2X2 OR2X2_1996 ( .A(_3438_), .B(_3437_), .Y(_3439_) );
OR2X2 OR2X2_1997 ( .A(_3436_), .B(_3439_), .Y(_3440_) );
AND2X2 AND2X2_2089 ( .A(_3409__bF_buf2), .B(_1788_), .Y(_3441_) );
AND2X2 AND2X2_2090 ( .A(_3411__bF_buf1), .B(_1792_), .Y(_3442_) );
OR2X2 OR2X2_1998 ( .A(_3441_), .B(_3442_), .Y(_3443_) );
AND2X2 AND2X2_2091 ( .A(_1797_), .B(_3414__bF_buf2), .Y(_3444_) );
AND2X2 AND2X2_2092 ( .A(_3416__bF_buf2), .B(_1801_), .Y(_3445_) );
OR2X2 OR2X2_1999 ( .A(_3444_), .B(_3445_), .Y(_3446_) );
OR2X2 OR2X2_2000 ( .A(_3446_), .B(_3443_), .Y(_3447_) );
OR2X2 OR2X2_2001 ( .A(_3440_), .B(_3447_), .Y(_3448_) );
OR2X2 OR2X2_2002 ( .A(_3433_), .B(_3448_), .Y(REG_A_1_) );
AND2X2 AND2X2_2093 ( .A(_3369__bF_buf3), .B(REGs_REGS_4__2_), .Y(_3449_) );
AND2X2 AND2X2_2094 ( .A(_3373__bF_buf0), .B(REGs_REGS_5__2_), .Y(_3450_) );
OR2X2 OR2X2_2003 ( .A(_3449_), .B(_3450_), .Y(_3451_) );
AND2X2 AND2X2_2095 ( .A(_3378__bF_buf2), .B(REGs_REGS_6__2_), .Y(_3452_) );
AND2X2 AND2X2_2096 ( .A(_3381__bF_buf2), .B(REGs_REGS_7__2_), .Y(_3453_) );
OR2X2 OR2X2_2004 ( .A(_3453_), .B(_3452_), .Y(_3454_) );
OR2X2 OR2X2_2005 ( .A(_3451_), .B(_3454_), .Y(_3455_) );
AND2X2 AND2X2_2097 ( .A(_3386__bF_buf2), .B(PC_ADDR_stack_1__2_), .Y(_3456_) );
AND2X2 AND2X2_2098 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__2_), .Y(_3457_) );
AND2X2 AND2X2_2099 ( .A(_3390__bF_buf3), .B(REGs_REGS_2__2_), .Y(_3458_) );
OR2X2 OR2X2_2006 ( .A(_3457_), .B(_3458_), .Y(_3459_) );
OR2X2 OR2X2_2007 ( .A(_3456_), .B(_3459_), .Y(_3460_) );
OR2X2 OR2X2_2008 ( .A(_3460_), .B(_3455_), .Y(_3461_) );
AND2X2 AND2X2_2100 ( .A(_1821_), .B(_3396__bF_buf2), .Y(_3462_) );
AND2X2 AND2X2_2101 ( .A(_1825_), .B(_3398__bF_buf3), .Y(_3463_) );
OR2X2 OR2X2_2009 ( .A(_3463_), .B(_3462_), .Y(_3464_) );
AND2X2 AND2X2_2102 ( .A(_1830_), .B(_3401__bF_buf3), .Y(_3465_) );
AND2X2 AND2X2_2103 ( .A(_1834_), .B(_3403__bF_buf2), .Y(_3466_) );
OR2X2 OR2X2_2010 ( .A(_3466_), .B(_3465_), .Y(_3467_) );
OR2X2 OR2X2_2011 ( .A(_3464_), .B(_3467_), .Y(_3468_) );
AND2X2 AND2X2_2104 ( .A(_3409__bF_buf1), .B(_1840_), .Y(_3469_) );
AND2X2 AND2X2_2105 ( .A(_3411__bF_buf4), .B(_1844_), .Y(_3470_) );
OR2X2 OR2X2_2012 ( .A(_3469_), .B(_3470_), .Y(_3471_) );
AND2X2 AND2X2_2106 ( .A(_1849_), .B(_3414__bF_buf3), .Y(_3472_) );
AND2X2 AND2X2_2107 ( .A(_3416__bF_buf1), .B(_1853_), .Y(_3473_) );
OR2X2 OR2X2_2013 ( .A(_3472_), .B(_3473_), .Y(_3474_) );
OR2X2 OR2X2_2014 ( .A(_3474_), .B(_3471_), .Y(_3475_) );
OR2X2 OR2X2_2015 ( .A(_3468_), .B(_3475_), .Y(_3476_) );
OR2X2 OR2X2_2016 ( .A(_3461_), .B(_3476_), .Y(REG_A_2_) );
AND2X2 AND2X2_2108 ( .A(_3369__bF_buf4), .B(REGs_REGS_4__3_), .Y(_3477_) );
AND2X2 AND2X2_2109 ( .A(_3373__bF_buf0), .B(REGs_REGS_5__3_), .Y(_3478_) );
OR2X2 OR2X2_2017 ( .A(_3477_), .B(_3478_), .Y(_3479_) );
AND2X2 AND2X2_2110 ( .A(_3378__bF_buf2), .B(REGs_REGS_6__3_), .Y(_3480_) );
AND2X2 AND2X2_2111 ( .A(_3381__bF_buf2), .B(REGs_REGS_7__3_), .Y(_3481_) );
OR2X2 OR2X2_2018 ( .A(_3481_), .B(_3480_), .Y(_3482_) );
OR2X2 OR2X2_2019 ( .A(_3479_), .B(_3482_), .Y(_3483_) );
AND2X2 AND2X2_2112 ( .A(_3386__bF_buf2), .B(PC_ADDR_stack_1__3_), .Y(_3484_) );
AND2X2 AND2X2_2113 ( .A(_3388__bF_buf3), .B(REGs_REGS_3__3_), .Y(_3485_) );
endmodule
