magic
tech scmos
magscale 1 4
timestamp 1516238463
<< metal1 >>
rect 1608 3937 1619 3943
rect 2024 3937 2035 3943
rect 3336 3937 3347 3943
rect 3400 3937 3411 3943
rect 509 3897 520 3903
rect 1725 3897 1736 3903
rect 1933 3897 1971 3903
rect 61 3877 72 3883
rect 189 3877 200 3883
rect 589 3877 627 3883
rect 696 3877 707 3883
rect 797 3877 808 3883
rect 1117 3877 1155 3883
rect 1933 3883 1939 3897
rect 2076 3897 2088 3903
rect 2076 3892 2084 3897
rect 2365 3897 2376 3903
rect 2653 3897 2664 3903
rect 3016 3897 3027 3903
rect 3741 3897 3763 3903
rect 3805 3897 3816 3903
rect 1901 3877 1939 3883
rect 2776 3877 2787 3883
rect 2936 3877 2947 3883
rect 3757 3883 3763 3897
rect 3949 3897 3960 3903
rect 3464 3877 3491 3883
rect 3757 3877 3768 3883
rect 3949 3877 3976 3883
rect 4621 3877 4632 3883
rect 5965 3877 5976 3883
rect 984 3837 1011 3843
rect 109 3737 120 3743
rect 301 3737 312 3743
rect 445 3737 483 3743
rect 669 3737 707 3743
rect 888 3737 899 3743
rect 1389 3737 1400 3743
rect 1517 3737 1528 3743
rect 1645 3737 1656 3743
rect 3240 3737 3267 3743
rect 3629 3737 3651 3743
rect 2525 3717 2536 3723
rect 2797 3717 2824 3723
rect 3544 3717 3555 3723
rect 3629 3723 3635 3737
rect 4408 3737 4419 3743
rect 4765 3737 4776 3743
rect 5005 3737 5075 3743
rect 5277 3737 5288 3743
rect 5357 3737 5395 3743
rect 5485 3737 5496 3743
rect 5661 3737 5699 3743
rect 3613 3717 3635 3723
rect 4056 3717 4083 3723
rect 200 3677 211 3683
rect 1288 3677 1299 3683
rect 3176 3677 3187 3683
rect 3032 3637 3059 3643
rect 1069 3503 1075 3523
rect 2808 3517 2819 3523
rect 1052 3497 1075 3503
rect 1052 3492 1060 3497
rect 1112 3497 1123 3503
rect 2285 3497 2296 3503
rect 2941 3497 2968 3503
rect 3565 3503 3571 3523
rect 3549 3497 3571 3503
rect 3672 3497 3683 3503
rect 4024 3497 4083 3503
rect 4856 3497 4867 3503
rect 5064 3497 5091 3503
rect 445 3477 467 3483
rect 765 3477 787 3483
rect 1053 3477 1064 3483
rect 1213 3477 1224 3483
rect 2509 3477 2520 3483
rect 2680 3477 2691 3483
rect 3053 3477 3075 3483
rect 3789 3477 3811 3483
rect 4280 3477 4291 3483
rect 5037 3477 5064 3483
rect 5565 3477 5576 3483
rect 893 3437 920 3443
rect 2984 3437 3011 3443
rect 3981 3377 4019 3383
rect 2957 3357 2984 3363
rect 3981 3363 3987 3377
rect 3965 3357 3987 3363
rect 5021 3357 5032 3363
rect 520 3337 531 3343
rect 584 3337 595 3343
rect 765 3337 776 3343
rect 1597 3337 1619 3343
rect 2349 3337 2371 3343
rect 2941 3337 2979 3343
rect 3053 3337 3075 3343
rect 3101 3337 3139 3343
rect 1917 3317 1960 3323
rect 2973 3323 2979 3337
rect 3288 3337 3299 3343
rect 3325 3337 3352 3343
rect 3821 3337 3832 3343
rect 4493 3337 4504 3343
rect 4621 3337 4632 3343
rect 2973 3317 3011 3323
rect 5277 3317 5288 3323
rect 1608 3297 1619 3303
rect 3912 3277 3923 3283
rect 920 3237 947 3243
rect 584 3117 595 3123
rect 1048 3117 1059 3123
rect 1112 3117 1123 3123
rect 2797 3117 2808 3123
rect 797 3097 835 3103
rect 2008 3097 2020 3103
rect 2012 3092 2020 3097
rect 2909 3103 2915 3123
rect 4920 3117 4931 3123
rect 2893 3097 2915 3103
rect 3512 3097 3523 3103
rect 3581 3097 3592 3103
rect 3928 3097 3939 3103
rect 3992 3097 4036 3103
rect 4028 3092 4036 3097
rect 5325 3097 5347 3103
rect 253 3077 275 3083
rect 392 3077 419 3083
rect 1773 3077 1795 3083
rect 2573 3077 2595 3083
rect 2845 3077 2856 3083
rect 4472 3077 4483 3083
rect 5037 3077 5091 3083
rect 5117 3077 5128 3083
rect 5288 3077 5299 3083
rect 5373 3077 5411 3083
rect 5581 3077 5592 3083
rect 2488 2957 2499 2963
rect 1016 2937 1027 2943
rect 1480 2937 1491 2943
rect 1944 2937 1971 2943
rect 2333 2937 2360 2943
rect 2765 2937 2776 2943
rect 4109 2937 4120 2943
rect 4765 2937 4787 2943
rect 3469 2917 3480 2923
rect 3565 2917 3576 2923
rect 4984 2917 4995 2923
rect 573 2897 584 2903
rect 3144 2877 3155 2883
rect 3272 2877 3283 2883
rect 893 2837 904 2843
rect 1256 2697 1268 2703
rect 1260 2692 1268 2697
rect 1976 2697 2003 2703
rect 2988 2697 3016 2703
rect 2988 2692 2996 2697
rect 3148 2697 3160 2703
rect 3148 2692 3156 2697
rect 3197 2703 3203 2723
rect 3197 2697 3219 2703
rect 3773 2703 3779 2723
rect 3756 2697 3779 2703
rect 3756 2692 3764 2697
rect 3996 2697 4024 2703
rect 3996 2692 4004 2697
rect 4200 2697 4211 2703
rect 5661 2697 5684 2703
rect 5676 2692 5684 2697
rect 5981 2697 5992 2703
rect 125 2677 147 2683
rect 445 2677 467 2683
rect 1053 2677 1075 2683
rect 1741 2677 1752 2683
rect 2797 2677 2819 2683
rect 2861 2677 2899 2683
rect 2861 2657 2867 2677
rect 4685 2677 4696 2683
rect 4813 2677 4851 2683
rect 4941 2677 4952 2683
rect 5021 2677 5048 2683
rect 5181 2677 5203 2683
rect 5917 2677 5955 2683
rect 3224 2657 3235 2663
rect 1949 2637 1976 2643
rect 3032 2637 3043 2643
rect 5048 2637 5075 2643
rect 2957 2577 2995 2583
rect 1549 2557 1571 2563
rect 2989 2563 2995 2577
rect 2989 2557 3011 2563
rect 408 2537 419 2543
rect 621 2537 659 2543
rect 1101 2537 1112 2543
rect 1213 2537 1240 2543
rect 1677 2537 1699 2543
rect 1800 2537 1827 2543
rect 2445 2537 2456 2543
rect 2813 2537 2851 2543
rect 4093 2537 4104 2543
rect 4429 2537 4440 2543
rect 4760 2537 4787 2543
rect 5805 2537 5832 2543
rect 2104 2517 2115 2523
rect 4253 2517 4264 2523
rect 4328 2517 4339 2523
rect 5048 2517 5075 2523
rect 5517 2517 5528 2523
rect 4317 2497 4339 2503
rect 5128 2497 5139 2503
rect 5949 2437 5960 2443
rect 4008 2337 4035 2343
rect 904 2317 947 2323
rect 1192 2317 1203 2323
rect 1965 2317 2008 2323
rect 2061 2317 2072 2323
rect 456 2297 468 2303
rect 460 2292 468 2297
rect 701 2297 712 2303
rect 892 2297 904 2303
rect 892 2292 900 2297
rect 1821 2297 1832 2303
rect 1912 2297 1924 2303
rect 1916 2292 1924 2297
rect 2589 2297 2600 2303
rect 3080 2297 3091 2303
rect 3208 2297 3219 2303
rect 3576 2297 3588 2303
rect 3580 2292 3588 2297
rect 4076 2297 4088 2303
rect 4076 2292 4084 2297
rect 4397 2297 4408 2303
rect 301 2277 312 2283
rect 749 2277 787 2283
rect 781 2268 787 2277
rect 1245 2277 1267 2283
rect 1293 2277 1304 2283
rect 1784 2277 1795 2283
rect 2573 2277 2627 2283
rect 3309 2277 3331 2283
rect 3853 2277 3875 2283
rect 4333 2277 4387 2283
rect 4397 2277 4403 2297
rect 4456 2297 4468 2303
rect 4460 2292 4468 2297
rect 5708 2297 5720 2303
rect 5708 2292 5716 2297
rect 5880 2297 5892 2303
rect 5884 2292 5892 2297
rect 4573 2277 4584 2283
rect 4685 2277 4696 2283
rect 4765 2277 4792 2283
rect 4877 2277 4888 2283
rect 5064 2277 5075 2283
rect 1320 2257 1331 2263
rect 3000 2237 3011 2243
rect 280 2137 307 2143
rect 461 2137 499 2143
rect 781 2137 792 2143
rect 952 2137 979 2143
rect 1773 2137 1795 2143
rect 1896 2137 1939 2143
rect 1965 2137 2019 2143
rect 2280 2137 2291 2143
rect 2317 2137 2339 2143
rect 2568 2137 2579 2143
rect 2744 2137 2787 2143
rect 4221 2137 4232 2143
rect 4621 2137 4648 2143
rect 4744 2137 4755 2143
rect 5197 2137 5219 2143
rect 2541 2117 2563 2123
rect 3837 2117 3848 2123
rect 3960 2117 4019 2123
rect 4328 2117 4339 2123
rect 4408 2117 4419 2123
rect 5000 2117 5032 2123
rect 5213 2123 5219 2137
rect 5805 2137 5816 2143
rect 5213 2117 5224 2123
rect 5837 2123 5843 2143
rect 5832 2117 5843 2123
rect 1656 2097 1667 2103
rect 2061 2097 2072 2103
rect 4781 2097 4803 2103
rect 29 1917 40 1923
rect 1240 1917 1251 1923
rect 1496 1917 1507 1923
rect 3485 1917 3496 1923
rect 189 1897 227 1903
rect 301 1897 339 1903
rect 776 1897 787 1903
rect 940 1897 968 1903
rect 940 1892 948 1897
rect 2973 1897 2984 1903
rect 3181 1897 3208 1903
rect 4301 1897 4323 1903
rect 61 1877 99 1883
rect 232 1877 243 1883
rect 317 1877 328 1883
rect 392 1877 403 1883
rect 685 1877 712 1883
rect 1037 1877 1048 1883
rect 2077 1877 2115 1883
rect 2077 1868 2083 1877
rect 2920 1877 2931 1883
rect 3448 1877 3459 1883
rect 4301 1877 4307 1897
rect 5336 1897 5347 1903
rect 4909 1877 4931 1883
rect 4957 1877 4968 1883
rect 5533 1877 5544 1883
rect 5741 1877 5752 1883
rect 3432 1857 3443 1863
rect 3656 1857 3667 1863
rect 3997 1857 4008 1863
rect 968 1837 995 1843
rect 1837 1777 1848 1783
rect 4040 1777 4067 1783
rect 5933 1777 5944 1783
rect 109 1743 115 1763
rect 2989 1757 3016 1763
rect 3576 1757 3587 1763
rect 3704 1757 3715 1763
rect 77 1737 115 1743
rect 141 1737 179 1743
rect 1933 1737 1987 1743
rect 2184 1737 2195 1743
rect 2285 1737 2307 1743
rect 3592 1737 3603 1743
rect 4109 1737 4120 1743
rect 4413 1737 4424 1743
rect 4493 1737 4515 1743
rect 4541 1737 4552 1743
rect 5528 1737 5555 1743
rect 45 1717 67 1723
rect 45 1708 51 1717
rect 1165 1717 1176 1723
rect 3100 1723 3108 1728
rect 3085 1717 3108 1723
rect 3452 1723 3460 1728
rect 3448 1717 3460 1723
rect 4205 1717 4216 1723
rect 5037 1717 5080 1723
rect 5192 1717 5203 1723
rect 3016 1697 3043 1703
rect 652 1683 660 1688
rect 605 1677 660 1683
rect 1837 1677 1864 1683
rect 2845 1537 2867 1543
rect 1400 1517 1411 1523
rect 2136 1517 2147 1523
rect 2861 1517 2867 1537
rect 3128 1537 3155 1543
rect 204 1503 212 1506
rect 189 1497 212 1503
rect 797 1497 808 1503
rect 1149 1497 1187 1503
rect 1452 1497 1464 1503
rect 1452 1492 1460 1497
rect 1629 1497 1656 1503
rect 1965 1497 1976 1503
rect 2072 1497 2083 1503
rect 2744 1497 2755 1503
rect 3005 1503 3011 1523
rect 3400 1517 3411 1523
rect 3544 1517 3555 1523
rect 3688 1517 3699 1523
rect 2941 1497 3011 1503
rect 3021 1497 3032 1503
rect 4024 1497 4051 1503
rect 509 1477 563 1483
rect 765 1477 776 1483
rect 984 1477 1011 1483
rect 1581 1477 1592 1483
rect 2781 1477 2808 1483
rect 3085 1477 3096 1483
rect 3485 1477 3496 1483
rect 3981 1477 4008 1483
rect 4520 1477 4531 1483
rect 4557 1477 4568 1483
rect 4637 1477 4675 1483
rect 5165 1477 5203 1483
rect 5389 1477 5411 1483
rect 5773 1477 5784 1483
rect 5928 1477 5939 1483
rect 3144 1457 3155 1463
rect 4237 1437 4248 1443
rect 5032 1437 5059 1443
rect 4040 1377 4051 1383
rect 637 1357 659 1363
rect 1117 1337 1128 1343
rect 1837 1343 1843 1352
rect 1720 1337 1731 1343
rect 1821 1337 1843 1343
rect 1960 1337 2003 1343
rect 2536 1337 2547 1343
rect 2573 1337 2595 1343
rect 93 1317 116 1323
rect 108 1314 116 1317
rect 3101 1337 3112 1343
rect 3389 1343 3395 1363
rect 3357 1337 3395 1343
rect 4600 1337 4611 1343
rect 4749 1337 4760 1343
rect 5016 1337 5075 1343
rect 5485 1343 5491 1363
rect 5464 1337 5491 1343
rect 5645 1337 5656 1343
rect 808 1317 819 1323
rect 2893 1317 2915 1323
rect 3384 1317 3395 1323
rect 3624 1317 3635 1323
rect 3656 1317 3667 1323
rect 1080 1297 1091 1303
rect 1933 1297 1944 1303
rect 3661 1297 3667 1317
rect 4892 1323 4900 1328
rect 4892 1317 4904 1323
rect 5916 1323 5924 1328
rect 5916 1317 5960 1323
rect 648 1277 659 1283
rect 1357 1277 1384 1283
rect 1357 1257 1363 1277
rect 2296 1277 2307 1283
rect 1000 1237 1027 1243
rect 3997 1237 4024 1243
rect 780 1137 792 1143
rect 780 1132 788 1137
rect 1389 1137 1400 1143
rect 4712 1137 4723 1143
rect 5192 1137 5203 1143
rect 1917 1117 1960 1123
rect 2152 1117 2163 1123
rect 2344 1117 2355 1123
rect 2904 1117 2915 1123
rect 4264 1117 4275 1123
rect 5256 1117 5267 1123
rect 204 1103 212 1106
rect 189 1097 212 1103
rect 952 1097 979 1103
rect 1213 1097 1251 1103
rect 1672 1097 1684 1103
rect 1676 1092 1684 1097
rect 1864 1097 1891 1103
rect 1928 1097 1987 1103
rect 2024 1097 2035 1103
rect 2076 1097 2099 1103
rect 2076 1092 2084 1097
rect 2412 1103 2420 1108
rect 2397 1097 2420 1103
rect 744 1077 755 1083
rect 1149 1077 1187 1083
rect 1197 1077 1208 1083
rect 1149 1057 1155 1077
rect 1512 1077 1523 1083
rect 2397 1077 2403 1097
rect 3533 1097 3571 1103
rect 5308 1097 5331 1103
rect 5308 1092 5316 1097
rect 3000 1077 3011 1083
rect 3405 1077 3416 1083
rect 3517 1077 3528 1083
rect 3992 1077 4019 1083
rect 4317 1077 4328 1083
rect 4317 1057 4323 1077
rect 5021 1077 5048 1083
rect 5357 1077 5368 1083
rect 5501 1077 5523 1083
rect 5741 1077 5752 1083
rect 893 1037 904 1043
rect 5048 1037 5075 1043
rect 2989 977 3016 983
rect 1597 957 1635 963
rect 189 917 212 923
rect 204 914 212 917
rect 920 937 963 943
rect 1533 937 1544 943
rect 1976 937 2003 943
rect 2109 937 2131 943
rect 2584 937 2595 943
rect 3096 937 3107 943
rect 3325 943 3331 963
rect 3997 957 4040 963
rect 5917 957 5928 963
rect 3272 937 3283 943
rect 3293 937 3331 943
rect 3640 937 3651 943
rect 3741 937 3763 943
rect 4093 937 4115 943
rect 4296 937 4307 943
rect 4888 937 4899 943
rect 4973 937 5011 943
rect 780 923 788 928
rect 765 917 788 923
rect 920 917 947 923
rect 2748 923 2756 928
rect 2748 917 2760 923
rect 3117 917 3155 923
rect 701 897 712 903
rect 1949 897 1976 903
rect 3149 897 3155 917
rect 3613 917 3635 923
rect 5005 923 5011 937
rect 5661 937 5683 943
rect 5736 937 5747 943
rect 5005 917 5043 923
rect 5596 923 5604 928
rect 5596 917 5619 923
rect 5480 877 5491 883
rect 3992 777 4019 783
rect 2141 737 2216 743
rect 701 717 712 723
rect 1053 697 1091 703
rect 1133 697 1171 703
rect 1325 697 1347 703
rect 1496 697 1507 703
rect 1581 697 1619 703
rect 1724 697 1736 703
rect 1724 692 1732 697
rect 1773 703 1779 723
rect 2189 717 2200 723
rect 2621 717 2659 723
rect 3208 717 3219 723
rect 1773 697 1811 703
rect 2301 697 2339 703
rect 3245 697 3283 703
rect 3400 697 3411 703
rect 1037 677 1048 683
rect 1288 677 1299 683
rect 1469 677 1480 683
rect 1912 677 1923 683
rect 2461 677 2483 683
rect 3101 677 3112 683
rect 2941 657 2968 663
rect 3101 657 3107 677
rect 3288 677 3299 683
rect 3645 677 3667 683
rect 5165 677 5176 683
rect 5229 677 5240 683
rect 5485 677 5496 683
rect 5629 677 5651 683
rect 5021 657 5043 663
rect 5181 657 5203 663
rect 920 637 947 643
rect 5037 643 5043 657
rect 5037 637 5075 643
rect 3992 577 4019 583
rect 845 537 856 543
rect 1437 543 1443 563
rect 1640 556 1644 564
rect 1437 537 1475 543
rect 1485 537 1496 543
rect 1864 537 1875 543
rect 2701 543 2707 563
rect 3112 556 3116 564
rect 2632 537 2659 543
rect 2669 537 2707 543
rect 2797 537 2808 543
rect 2925 537 2979 543
rect 684 523 692 528
rect 440 517 451 523
rect 669 517 692 523
rect 861 517 899 523
rect 1117 517 1128 523
rect 1501 517 1539 523
rect 2941 517 2952 523
rect 2973 523 2979 537
rect 3160 537 3171 543
rect 3309 537 3320 543
rect 3565 537 3576 543
rect 3709 543 3715 552
rect 3709 537 3747 543
rect 3949 537 3960 543
rect 4365 537 4403 543
rect 4877 537 4931 543
rect 5549 537 5571 543
rect 5661 537 5672 543
rect 5917 537 5976 543
rect 2973 517 2995 523
rect 5016 517 5059 523
rect 733 497 744 503
rect 2269 497 2291 503
rect 3096 497 3107 503
rect 5240 477 5251 483
rect 584 336 586 344
rect 1037 317 1048 323
rect 1837 317 1848 323
rect 3080 317 3091 323
rect 4088 317 4099 323
rect 4152 317 4163 323
rect 2444 303 2452 306
rect 2429 297 2452 303
rect 3000 297 3027 303
rect 3132 297 3144 303
rect 3132 292 3140 297
rect 3997 297 4035 303
rect 2749 277 2771 283
rect 2765 257 2771 277
rect 3133 277 3155 283
rect 3149 257 3155 277
rect 3997 283 4003 297
rect 4888 297 4915 303
rect 5016 297 5043 303
rect 3981 277 4003 283
rect 4189 277 4200 283
rect 4861 277 4899 283
rect 5405 277 5427 283
rect 2973 237 2984 243
rect 1912 177 1923 183
rect 5032 177 5059 183
rect 5608 157 5619 163
rect 941 137 979 143
rect 429 117 452 123
rect 444 114 452 117
rect 941 123 947 137
rect 2989 137 3027 143
rect 925 117 947 123
rect 1101 117 1124 123
rect 1116 114 1124 117
rect 1676 117 1699 123
rect 1676 114 1684 117
rect 1869 117 1896 123
rect 2556 117 2579 123
rect 2556 114 2564 117
rect 3021 123 3027 137
rect 4013 137 4051 143
rect 2940 117 2963 123
rect 3021 117 3043 123
rect 2940 114 2948 117
rect 3229 117 3240 123
rect 3516 117 3539 123
rect 3516 114 3524 117
rect 3757 117 3780 123
rect 3772 114 3780 117
rect 4013 123 4019 137
rect 5229 137 5251 143
rect 3997 117 4019 123
rect 4120 117 4131 123
rect 4428 117 4451 123
rect 4428 114 4436 117
rect 5624 137 5635 143
rect 5661 137 5699 143
rect 4844 117 4867 123
rect 4844 114 4852 117
<< m2contact >>
rect 925 4002 961 4018
rect 2973 4002 3009 4018
rect 5021 4002 5057 4018
rect 5848 3972 5864 3988
rect 1592 3932 1608 3948
rect 2008 3932 2024 3948
rect 3320 3932 3336 3948
rect 3384 3932 3400 3948
rect 5128 3932 5144 3948
rect 5000 3912 5016 3928
rect 216 3892 232 3908
rect 296 3892 312 3908
rect 344 3892 360 3908
rect 392 3892 424 3908
rect 440 3892 456 3908
rect 488 3892 504 3908
rect 520 3892 552 3908
rect 584 3892 600 3908
rect 664 3892 680 3908
rect 824 3892 840 3908
rect 888 3892 904 3908
rect 936 3892 968 3908
rect 1144 3892 1160 3908
rect 1192 3892 1224 3908
rect 1240 3892 1256 3908
rect 1272 3892 1288 3908
rect 1384 3892 1400 3908
rect 1416 3892 1432 3908
rect 1576 3892 1608 3908
rect 1736 3892 1752 3908
rect 40 3876 56 3892
rect 88 3888 104 3892
rect 72 3876 104 3888
rect 168 3876 184 3892
rect 72 3872 88 3876
rect 200 3872 216 3888
rect 312 3872 328 3888
rect 632 3876 648 3892
rect 680 3872 696 3888
rect 776 3876 792 3892
rect 1032 3888 1048 3892
rect 808 3872 824 3888
rect 1032 3876 1064 3888
rect 1096 3876 1112 3892
rect 1448 3888 1464 3892
rect 1512 3888 1528 3892
rect 1640 3888 1656 3892
rect 1832 3888 1848 3892
rect 1048 3872 1064 3876
rect 1224 3872 1240 3888
rect 1320 3872 1336 3888
rect 1400 3872 1416 3888
rect 1448 3876 1480 3888
rect 1512 3876 1544 3888
rect 1640 3876 1672 3888
rect 1464 3872 1480 3876
rect 1528 3872 1544 3876
rect 1656 3872 1672 3876
rect 1768 3872 1784 3888
rect 1832 3876 1864 3888
rect 2056 3892 2072 3908
rect 2088 3892 2136 3908
rect 2152 3892 2184 3908
rect 2200 3892 2216 3908
rect 2248 3892 2280 3908
rect 2296 3892 2312 3908
rect 2344 3892 2360 3908
rect 2376 3892 2408 3908
rect 2440 3892 2472 3908
rect 2520 3892 2536 3908
rect 2584 3892 2600 3908
rect 2664 3892 2696 3908
rect 2728 3892 2760 3908
rect 2776 3892 2792 3908
rect 2824 3892 2856 3908
rect 2904 3892 2920 3908
rect 2968 3892 2984 3908
rect 3000 3892 3016 3908
rect 3080 3892 3096 3908
rect 3176 3892 3192 3908
rect 3304 3892 3320 3908
rect 3432 3892 3448 3908
rect 3480 3892 3496 3908
rect 3528 3892 3560 3908
rect 3576 3892 3592 3908
rect 3624 3892 3656 3908
rect 3672 3892 3688 3908
rect 3720 3892 3736 3908
rect 1992 3888 2008 3892
rect 3368 3888 3384 3892
rect 1992 3876 2024 3888
rect 1848 3872 1864 3876
rect 2008 3872 2024 3876
rect 2200 3872 2216 3888
rect 2296 3872 2312 3888
rect 2392 3872 2408 3888
rect 2760 3872 2776 3888
rect 2920 3872 2936 3888
rect 3048 3872 3064 3888
rect 3192 3872 3208 3888
rect 3240 3872 3256 3888
rect 3320 3872 3336 3888
rect 3368 3876 3400 3888
rect 3384 3872 3400 3876
rect 3448 3872 3464 3888
rect 3816 3892 3832 3908
rect 3880 3892 3912 3908
rect 3960 3892 3976 3908
rect 4008 3892 4040 3908
rect 4072 3892 4088 3908
rect 4104 3892 4136 3908
rect 4168 3892 4184 3908
rect 4200 3892 4232 3908
rect 4264 3892 4280 3908
rect 4296 3892 4328 3908
rect 4360 3892 4376 3908
rect 4488 3892 4504 3908
rect 4552 3892 4568 3908
rect 4648 3892 4664 3908
rect 4680 3892 4696 3908
rect 4872 3892 4888 3908
rect 4952 3892 4984 3908
rect 5064 3892 5080 3908
rect 5160 3892 5176 3908
rect 5288 3892 5304 3908
rect 5352 3892 5368 3908
rect 5400 3892 5416 3908
rect 5432 3892 5448 3908
rect 5608 3892 5624 3908
rect 5816 3892 5832 3908
rect 4424 3888 4440 3892
rect 4744 3888 4760 3892
rect 4808 3888 4824 3892
rect 5224 3888 5240 3892
rect 5544 3888 5560 3892
rect 5672 3888 5688 3892
rect 5736 3888 5752 3892
rect 3768 3872 3784 3888
rect 3976 3872 3992 3888
rect 4072 3872 4088 3888
rect 4264 3872 4280 3888
rect 4360 3872 4376 3888
rect 4424 3876 4456 3888
rect 4440 3872 4456 3876
rect 4504 3872 4520 3888
rect 4568 3872 4584 3888
rect 4632 3872 4648 3888
rect 4696 3872 4712 3888
rect 4744 3876 4776 3888
rect 4808 3876 4840 3888
rect 4760 3872 4776 3876
rect 4824 3872 4840 3876
rect 4888 3872 4904 3888
rect 4920 3872 4936 3888
rect 5176 3872 5192 3888
rect 5224 3876 5256 3888
rect 5240 3872 5256 3876
rect 5304 3872 5320 3888
rect 5368 3872 5400 3888
rect 5480 3872 5496 3888
rect 5544 3876 5576 3888
rect 5560 3872 5576 3876
rect 5624 3872 5640 3888
rect 5672 3876 5704 3888
rect 5736 3876 5768 3888
rect 5688 3872 5704 3876
rect 5752 3872 5768 3876
rect 5800 3872 5816 3888
rect 5864 3872 5880 3888
rect 5976 3872 5992 3888
rect 360 3852 376 3868
rect 680 3852 696 3868
rect 1176 3852 1192 3868
rect 1336 3852 1352 3868
rect 1912 3852 1928 3868
rect 2872 3852 2888 3868
rect 3256 3852 3272 3868
rect 3592 3852 3608 3868
rect 4632 3852 4648 3868
rect 5496 3852 5512 3868
rect 8 3832 24 3848
rect 120 3832 152 3848
rect 248 3832 280 3848
rect 456 3832 472 3848
rect 552 3832 568 3848
rect 728 3832 760 3848
rect 856 3832 872 3848
rect 904 3832 920 3848
rect 968 3832 984 3848
rect 1064 3832 1080 3848
rect 1288 3832 1304 3848
rect 1352 3832 1368 3848
rect 1480 3832 1496 3848
rect 1544 3832 1560 3848
rect 1688 3832 1704 3848
rect 1800 3832 1816 3848
rect 1864 3832 1880 3848
rect 2488 3832 2504 3848
rect 2552 3832 2568 3848
rect 2616 3832 2632 3848
rect 2696 3832 2712 3848
rect 3112 3832 3128 3848
rect 3144 3832 3160 3848
rect 3208 3832 3224 3848
rect 3272 3832 3288 3848
rect 3688 3832 3704 3848
rect 3848 3832 3864 3848
rect 4152 3832 4168 3848
rect 4392 3832 4408 3848
rect 4456 3832 4472 3848
rect 4520 3832 4536 3848
rect 4584 3832 4600 3848
rect 4712 3832 4728 3848
rect 4776 3832 4792 3848
rect 4840 3832 4856 3848
rect 5096 3832 5112 3848
rect 5192 3832 5208 3848
rect 5256 3832 5272 3848
rect 5320 3832 5336 3848
rect 5448 3832 5464 3848
rect 5512 3832 5528 3848
rect 5576 3832 5592 3848
rect 5640 3832 5656 3848
rect 5704 3832 5720 3848
rect 5912 3832 5928 3848
rect 1933 3802 1969 3818
rect 3981 3802 4017 3818
rect 392 3772 408 3788
rect 744 3772 760 3788
rect 1544 3772 1560 3788
rect 1800 3772 1816 3788
rect 1864 3772 1880 3788
rect 2024 3772 2040 3788
rect 2680 3772 2696 3788
rect 2776 3772 2792 3788
rect 3112 3772 3128 3788
rect 3800 3772 3816 3788
rect 4184 3772 4200 3788
rect 4280 3772 4296 3788
rect 4472 3772 4488 3788
rect 4536 3772 4552 3788
rect 5384 3772 5400 3788
rect 5432 3772 5448 3788
rect 5656 3772 5672 3788
rect 5736 3772 5752 3788
rect 5800 3772 5816 3788
rect 8 3752 24 3768
rect 120 3752 136 3768
rect 248 3752 264 3768
rect 312 3752 328 3768
rect 504 3752 520 3768
rect 616 3752 632 3768
rect 680 3752 696 3768
rect 856 3752 872 3768
rect 1208 3752 1224 3768
rect 1336 3752 1352 3768
rect 1400 3752 1416 3768
rect 1528 3752 1544 3768
rect 1656 3752 1672 3768
rect 1784 3752 1800 3768
rect 2008 3752 2024 3768
rect 3096 3752 3112 3768
rect 4264 3752 4280 3768
rect 4392 3752 4408 3768
rect 4456 3752 4472 3768
rect 4776 3752 4792 3768
rect 4840 3752 4856 3768
rect 4984 3752 5000 3768
rect 5048 3752 5064 3768
rect 5160 3752 5176 3768
rect 5224 3752 5240 3768
rect 5288 3752 5304 3768
rect 5496 3752 5512 3768
rect 5608 3752 5624 3768
rect 5816 3752 5832 3768
rect 24 3732 40 3748
rect 120 3732 136 3748
rect 168 3728 184 3744
rect 232 3732 248 3748
rect 312 3732 328 3748
rect 376 3732 392 3748
rect 424 3728 440 3744
rect 552 3732 568 3748
rect 632 3732 648 3748
rect 792 3744 808 3748
rect 776 3732 808 3744
rect 840 3732 856 3748
rect 872 3732 888 3748
rect 1192 3732 1208 3748
rect 1320 3732 1336 3748
rect 1400 3732 1416 3748
rect 776 3728 792 3732
rect 1448 3728 1464 3744
rect 1528 3732 1544 3748
rect 1592 3732 1608 3748
rect 1656 3732 1672 3748
rect 1768 3732 1784 3748
rect 1848 3732 1864 3748
rect 1912 3732 1928 3748
rect 1960 3732 1976 3748
rect 1992 3732 2008 3748
rect 2072 3732 2088 3748
rect 2136 3732 2152 3748
rect 3080 3732 3096 3748
rect 3160 3732 3176 3748
rect 3224 3732 3240 3748
rect 136 3712 152 3728
rect 184 3712 200 3728
rect 328 3712 344 3728
rect 360 3712 376 3728
rect 472 3712 488 3728
rect 520 3712 552 3728
rect 568 3712 584 3728
rect 600 3712 616 3728
rect 888 3712 904 3728
rect 936 3712 968 3728
rect 1016 3712 1048 3728
rect 1064 3712 1096 3728
rect 1128 3712 1144 3728
rect 1256 3712 1288 3728
rect 1416 3712 1432 3728
rect 1464 3712 1480 3728
rect 1576 3712 1592 3728
rect 1672 3712 1688 3728
rect 1704 3712 1736 3728
rect 1832 3712 1848 3728
rect 1896 3712 1912 3728
rect 2056 3712 2072 3728
rect 2088 3712 2104 3728
rect 2120 3712 2136 3728
rect 2168 3712 2184 3728
rect 2216 3712 2248 3728
rect 2264 3712 2280 3728
rect 2312 3712 2344 3728
rect 2360 3712 2376 3728
rect 2408 3712 2440 3728
rect 2456 3712 2472 3728
rect 2504 3712 2520 3728
rect 2536 3712 2568 3728
rect 2600 3712 2664 3728
rect 2696 3712 2712 3728
rect 2728 3712 2760 3728
rect 2824 3712 2856 3728
rect 2888 3712 2920 3728
rect 2936 3712 2952 3728
rect 2984 3712 3016 3728
rect 3144 3712 3160 3728
rect 3208 3712 3224 3728
rect 3256 3712 3272 3728
rect 3304 3712 3336 3728
rect 3352 3712 3368 3728
rect 3400 3712 3432 3728
rect 3448 3712 3464 3728
rect 3496 3712 3544 3728
rect 3592 3712 3608 3728
rect 4200 3732 4216 3748
rect 4248 3732 4264 3748
rect 4328 3732 4344 3748
rect 4376 3732 4408 3748
rect 4440 3732 4456 3748
rect 4520 3732 4536 3748
rect 4584 3732 4600 3748
rect 4776 3732 4792 3748
rect 4824 3732 4840 3748
rect 4904 3732 4920 3748
rect 5144 3732 5160 3748
rect 5208 3732 5224 3748
rect 5288 3732 5304 3748
rect 5496 3732 5528 3748
rect 5592 3732 5608 3748
rect 5752 3732 5768 3748
rect 5832 3732 5848 3748
rect 3672 3712 3720 3728
rect 3752 3712 3768 3728
rect 3832 3712 3848 3728
rect 3864 3712 3880 3728
rect 3912 3712 3976 3728
rect 4008 3712 4024 3728
rect 4040 3712 4056 3728
rect 4088 3712 4104 3728
rect 4136 3712 4152 3728
rect 4312 3712 4328 3728
rect 4504 3712 4520 3728
rect 4568 3712 4584 3728
rect 4648 3712 4664 3728
rect 4712 3712 4728 3728
rect 4888 3712 4904 3728
rect 4920 3712 4936 3728
rect 5304 3712 5320 3728
rect 5336 3712 5352 3728
rect 5416 3712 5432 3728
rect 5464 3712 5480 3728
rect 5624 3712 5640 3728
rect 5704 3712 5720 3728
rect 5768 3712 5784 3728
rect 5880 3712 5896 3728
rect 1144 3692 1160 3708
rect 3368 3692 3384 3708
rect 3640 3692 3656 3708
rect 184 3672 200 3688
rect 1112 3672 1128 3688
rect 1272 3672 1288 3688
rect 3160 3672 3176 3688
rect 3880 3672 3896 3688
rect 4856 3672 4872 3688
rect 1160 3652 1176 3668
rect 4120 3652 4136 3668
rect 56 3632 88 3648
rect 264 3632 280 3648
rect 728 3632 744 3648
rect 808 3632 824 3648
rect 1128 3632 1144 3648
rect 1224 3632 1240 3648
rect 1352 3632 1368 3648
rect 1480 3632 1496 3648
rect 1608 3632 1624 3648
rect 1736 3632 1752 3648
rect 2184 3632 2200 3648
rect 2280 3632 2296 3648
rect 2376 3632 2392 3648
rect 2472 3632 2488 3648
rect 2568 3632 2584 3648
rect 2856 3632 2872 3648
rect 2952 3632 2968 3648
rect 3016 3632 3032 3648
rect 3464 3632 3480 3648
rect 3560 3632 3576 3648
rect 3736 3632 3752 3648
rect 3800 3632 3816 3648
rect 3992 3632 4008 3648
rect 4216 3632 4232 3648
rect 4344 3632 4360 3648
rect 4616 3632 4632 3648
rect 4680 3632 4696 3648
rect 4728 3632 4744 3648
rect 4792 3632 4808 3648
rect 4952 3632 4968 3648
rect 5096 3632 5128 3648
rect 5176 3632 5192 3648
rect 5240 3632 5256 3648
rect 5384 3632 5400 3648
rect 5544 3632 5576 3648
rect 5656 3632 5672 3648
rect 5864 3632 5880 3648
rect 5912 3632 5928 3648
rect 925 3602 961 3618
rect 2973 3602 3009 3618
rect 5021 3602 5057 3618
rect 2744 3572 2760 3588
rect 3736 3572 3752 3588
rect 4088 3572 4104 3588
rect 1448 3552 1464 3568
rect 2616 3552 2632 3568
rect 3560 3532 3576 3548
rect 40 3492 56 3508
rect 72 3492 88 3508
rect 168 3492 184 3508
rect 264 3492 280 3508
rect 328 3492 344 3508
rect 424 3492 440 3508
rect 456 3492 472 3508
rect 552 3492 568 3508
rect 616 3492 632 3508
rect 664 3492 680 3508
rect 744 3492 760 3508
rect 840 3492 872 3508
rect 1032 3492 1048 3508
rect 2792 3512 2808 3528
rect 1096 3492 1112 3508
rect 1144 3492 1160 3508
rect 1272 3492 1288 3508
rect 1336 3492 1352 3508
rect 1480 3492 1496 3508
rect 1528 3492 1592 3508
rect 1656 3492 1672 3508
rect 1784 3492 1800 3508
rect 1864 3492 1880 3508
rect 1912 3492 1928 3508
rect 1976 3492 2008 3508
rect 2040 3492 2056 3508
rect 2104 3492 2136 3508
rect 2168 3492 2184 3508
rect 2216 3492 2232 3508
rect 2264 3492 2280 3508
rect 2296 3492 2344 3508
rect 2360 3492 2392 3508
rect 2424 3492 2440 3508
rect 2488 3492 2504 3508
rect 2536 3492 2552 3508
rect 2584 3492 2616 3508
rect 2648 3492 2664 3508
rect 2696 3492 2712 3508
rect 2776 3492 2792 3508
rect 2840 3492 2856 3508
rect 2872 3492 2904 3508
rect 2968 3492 2984 3508
rect 3032 3492 3048 3508
rect 3064 3492 3096 3508
rect 3112 3492 3128 3508
rect 3224 3492 3240 3508
rect 3256 3492 3272 3508
rect 3288 3492 3304 3508
rect 3320 3492 3336 3508
rect 3352 3492 3368 3508
rect 3480 3492 3496 3508
rect 4728 3512 4744 3528
rect 4808 3512 4824 3528
rect 5864 3512 5880 3528
rect 3656 3492 3672 3508
rect 3784 3492 3800 3508
rect 3816 3492 3832 3508
rect 3896 3492 3960 3508
rect 3992 3492 4024 3508
rect 4120 3492 4152 3508
rect 4200 3492 4216 3508
rect 4376 3492 4392 3508
rect 4408 3492 4424 3508
rect 4440 3492 4456 3508
rect 4488 3492 4504 3508
rect 4552 3492 4568 3508
rect 4696 3492 4712 3508
rect 4760 3492 4776 3508
rect 4840 3492 4856 3508
rect 5016 3492 5032 3508
rect 5048 3492 5064 3508
rect 5112 3492 5144 3508
rect 5336 3492 5368 3508
rect 5544 3492 5560 3508
rect 5592 3492 5608 3508
rect 5704 3492 5736 3508
rect 5800 3492 5816 3508
rect 5832 3492 5848 3508
rect 5928 3492 5944 3508
rect 56 3472 72 3488
rect 88 3476 104 3492
rect 232 3488 248 3492
rect 184 3472 200 3488
rect 232 3476 264 3488
rect 280 3476 296 3492
rect 344 3476 360 3492
rect 472 3476 488 3492
rect 1720 3488 1736 3492
rect 248 3472 264 3476
rect 568 3472 584 3488
rect 632 3472 664 3488
rect 808 3472 840 3488
rect 936 3472 952 3488
rect 968 3472 984 3488
rect 1064 3472 1080 3488
rect 1096 3472 1112 3488
rect 1160 3472 1176 3488
rect 1224 3472 1240 3488
rect 1288 3472 1304 3488
rect 1352 3472 1368 3488
rect 1400 3472 1416 3488
rect 1672 3472 1688 3488
rect 1720 3476 1752 3488
rect 1736 3472 1752 3476
rect 1800 3472 1816 3488
rect 1848 3476 1864 3492
rect 1928 3472 1944 3488
rect 2184 3472 2200 3488
rect 2440 3472 2456 3488
rect 2520 3472 2536 3488
rect 2664 3472 2680 3488
rect 2792 3472 2808 3488
rect 2856 3472 2872 3488
rect 3160 3472 3176 3488
rect 3240 3472 3256 3488
rect 3304 3472 3320 3488
rect 3368 3472 3384 3488
rect 3416 3472 3432 3488
rect 3496 3472 3512 3488
rect 3592 3472 3608 3488
rect 3768 3476 3784 3492
rect 3992 3472 4008 3488
rect 4184 3476 4200 3492
rect 4248 3488 4264 3492
rect 5176 3488 5192 3492
rect 5304 3488 5320 3492
rect 5672 3488 5688 3492
rect 4248 3476 4280 3488
rect 4264 3472 4280 3476
rect 4312 3472 4328 3488
rect 4392 3472 4408 3488
rect 4456 3472 4488 3488
rect 4536 3472 4552 3488
rect 4632 3472 4648 3488
rect 4712 3472 4728 3488
rect 4776 3472 4792 3488
rect 4952 3472 4968 3488
rect 5064 3472 5080 3488
rect 5176 3476 5208 3488
rect 5192 3472 5208 3476
rect 5240 3472 5256 3488
rect 5304 3476 5336 3488
rect 5320 3472 5336 3476
rect 5400 3472 5416 3488
rect 5496 3472 5512 3488
rect 5576 3472 5592 3488
rect 5672 3476 5704 3488
rect 5688 3472 5704 3476
rect 5816 3472 5832 3488
rect 5944 3472 5960 3488
rect 824 3452 840 3468
rect 984 3452 1000 3468
rect 1080 3452 1096 3468
rect 1224 3452 1240 3468
rect 1416 3452 1432 3468
rect 2920 3452 2936 3468
rect 3176 3452 3192 3468
rect 3432 3452 3448 3468
rect 3512 3452 3528 3468
rect 4328 3452 4344 3468
rect 4648 3452 4664 3468
rect 4968 3452 4984 3468
rect 5256 3452 5272 3468
rect 8 3432 24 3448
rect 120 3432 152 3448
rect 200 3432 216 3448
rect 312 3432 328 3448
rect 376 3432 408 3448
rect 504 3432 536 3448
rect 584 3432 600 3448
rect 696 3432 728 3448
rect 920 3432 936 3448
rect 1000 3432 1016 3448
rect 1176 3432 1192 3448
rect 1240 3432 1256 3448
rect 1304 3432 1320 3448
rect 1368 3432 1384 3448
rect 1496 3432 1512 3448
rect 1608 3432 1640 3448
rect 1688 3432 1704 3448
rect 1752 3432 1768 3448
rect 1816 3432 1832 3448
rect 1880 3432 1896 3448
rect 2024 3432 2040 3448
rect 2072 3432 2088 3448
rect 2136 3432 2152 3448
rect 2232 3432 2248 3448
rect 2392 3432 2408 3448
rect 2456 3432 2472 3448
rect 2552 3432 2568 3448
rect 2728 3432 2744 3448
rect 2968 3432 2984 3448
rect 3128 3432 3144 3448
rect 3192 3432 3208 3448
rect 3384 3432 3400 3448
rect 3448 3432 3464 3448
rect 3528 3432 3544 3448
rect 3560 3432 3576 3448
rect 3624 3432 3640 3448
rect 3704 3432 3720 3448
rect 3848 3432 3880 3448
rect 4152 3432 4168 3448
rect 4216 3432 4232 3448
rect 4344 3432 4360 3448
rect 4520 3432 4536 3448
rect 4584 3432 4616 3448
rect 4664 3432 4680 3448
rect 4888 3432 4904 3448
rect 4920 3432 4936 3448
rect 4984 3432 5000 3448
rect 5144 3432 5160 3448
rect 5208 3432 5224 3448
rect 5272 3432 5288 3448
rect 5384 3432 5400 3448
rect 5448 3432 5464 3448
rect 5512 3432 5528 3448
rect 5624 3432 5656 3448
rect 5752 3432 5784 3448
rect 5896 3432 5912 3448
rect 1933 3402 1969 3418
rect 3981 3402 4017 3418
rect 328 3372 344 3388
rect 440 3372 456 3388
rect 712 3372 728 3388
rect 1192 3372 1208 3388
rect 1752 3372 1768 3388
rect 1976 3372 1992 3388
rect 2120 3372 2136 3388
rect 2600 3372 2616 3388
rect 2776 3372 2792 3388
rect 2872 3372 2888 3388
rect 3208 3372 3224 3388
rect 8 3352 24 3368
rect 136 3352 152 3368
rect 248 3352 264 3368
rect 312 3352 328 3368
rect 504 3352 520 3368
rect 568 3352 584 3368
rect 632 3352 648 3368
rect 696 3352 712 3368
rect 888 3352 904 3368
rect 984 3352 1000 3368
rect 1048 3352 1064 3368
rect 1400 3352 1416 3368
rect 1656 3352 1688 3368
rect 1720 3352 1736 3368
rect 1848 3352 1864 3368
rect 2072 3352 2088 3368
rect 2184 3352 2200 3368
rect 2408 3352 2424 3368
rect 2472 3352 2488 3368
rect 2536 3352 2552 3368
rect 2696 3352 2712 3368
rect 2760 3352 2776 3368
rect 2984 3352 3000 3368
rect 3112 3352 3128 3368
rect 3144 3352 3160 3368
rect 3272 3352 3288 3368
rect 3336 3352 3352 3368
rect 3480 3352 3496 3368
rect 3832 3352 3848 3368
rect 4072 3372 4088 3388
rect 4264 3372 4280 3388
rect 4776 3372 4792 3388
rect 4840 3372 4856 3388
rect 5336 3372 5352 3388
rect 5480 3372 5496 3388
rect 5832 3372 5848 3388
rect 4184 3352 4200 3368
rect 4248 3352 4264 3368
rect 4456 3352 4472 3368
rect 4504 3352 4520 3368
rect 4632 3352 4648 3368
rect 4760 3352 4776 3368
rect 5032 3352 5048 3368
rect 5176 3352 5192 3368
rect 5400 3352 5416 3368
rect 5464 3352 5480 3368
rect 5608 3352 5624 3368
rect 5784 3352 5800 3368
rect 24 3332 40 3348
rect 120 3332 136 3348
rect 152 3332 168 3348
rect 232 3332 248 3348
rect 296 3332 312 3348
rect 392 3332 408 3348
rect 488 3332 520 3348
rect 552 3332 584 3348
rect 616 3332 632 3348
rect 680 3332 696 3348
rect 776 3344 792 3348
rect 776 3332 808 3344
rect 872 3332 888 3348
rect 968 3332 984 3348
rect 1032 3332 1048 3348
rect 1112 3344 1144 3348
rect 1096 3332 1144 3344
rect 1240 3332 1256 3348
rect 1384 3332 1400 3348
rect 1464 3332 1480 3348
rect 1640 3332 1656 3348
rect 1704 3332 1720 3348
rect 1832 3332 1848 3348
rect 2056 3332 2072 3348
rect 2088 3332 2104 3348
rect 2168 3332 2184 3348
rect 2216 3332 2232 3348
rect 792 3328 808 3332
rect 1096 3328 1112 3332
rect 2328 3328 2344 3344
rect 2392 3332 2408 3348
rect 2456 3332 2472 3348
rect 2520 3332 2536 3348
rect 2680 3332 2696 3348
rect 2744 3332 2760 3348
rect 2824 3344 2840 3348
rect 2808 3332 2840 3344
rect 2808 3328 2824 3332
rect 72 3312 88 3328
rect 104 3312 120 3328
rect 360 3312 392 3328
rect 408 3312 424 3328
rect 744 3312 760 3328
rect 824 3312 840 3328
rect 1064 3312 1080 3328
rect 1144 3312 1160 3328
rect 1176 3312 1192 3328
rect 1224 3312 1240 3328
rect 1272 3312 1288 3328
rect 1320 3312 1352 3328
rect 1416 3312 1432 3328
rect 1448 3312 1464 3328
rect 1528 3312 1560 3328
rect 1576 3312 1592 3328
rect 1784 3312 1800 3328
rect 1960 3312 1976 3328
rect 2008 3312 2024 3328
rect 2216 3312 2232 3328
rect 2264 3312 2296 3328
rect 2552 3312 2584 3328
rect 2616 3312 2632 3328
rect 2840 3312 2856 3328
rect 3160 3332 3176 3348
rect 3256 3332 3288 3348
rect 3352 3332 3384 3348
rect 3832 3332 3848 3348
rect 3944 3332 3960 3348
rect 4056 3332 4072 3348
rect 4120 3344 4136 3348
rect 4104 3332 4136 3344
rect 4168 3332 4184 3348
rect 4232 3332 4248 3348
rect 4440 3332 4456 3348
rect 4504 3332 4520 3348
rect 4568 3332 4584 3348
rect 4632 3332 4648 3348
rect 4696 3332 4712 3348
rect 4744 3332 4760 3348
rect 4824 3332 4840 3348
rect 4888 3332 4920 3348
rect 5000 3332 5016 3348
rect 5064 3344 5080 3348
rect 5064 3332 5096 3344
rect 5160 3332 5176 3348
rect 5384 3332 5400 3348
rect 5448 3332 5464 3348
rect 5528 3332 5544 3348
rect 5592 3332 5608 3348
rect 5624 3332 5640 3348
rect 5688 3332 5704 3348
rect 5768 3332 5784 3348
rect 4104 3328 4120 3332
rect 5080 3328 5096 3332
rect 3032 3312 3048 3328
rect 3176 3312 3192 3328
rect 3368 3312 3384 3328
rect 3416 3312 3464 3328
rect 3512 3312 3528 3328
rect 3560 3312 3592 3328
rect 3608 3312 3624 3328
rect 3656 3312 3720 3328
rect 3752 3312 3768 3328
rect 3848 3312 3864 3328
rect 3880 3312 3912 3328
rect 4040 3312 4056 3328
rect 4296 3312 4344 3328
rect 4360 3312 4392 3328
rect 4424 3312 4440 3328
rect 4520 3312 4536 3328
rect 4552 3312 4568 3328
rect 4648 3312 4664 3328
rect 4680 3312 4696 3328
rect 4808 3312 4824 3328
rect 4872 3312 4888 3328
rect 4920 3312 4936 3328
rect 4952 3312 4984 3328
rect 5112 3312 5128 3328
rect 5208 3312 5224 3328
rect 5256 3312 5272 3328
rect 5288 3312 5320 3328
rect 5512 3312 5528 3328
rect 5576 3312 5592 3328
rect 5720 3312 5736 3328
rect 5800 3312 5816 3328
rect 5864 3312 5896 3328
rect 5928 3312 5960 3328
rect 1592 3292 1608 3308
rect 2120 3292 2136 3308
rect 4584 3292 4600 3308
rect 1496 3272 1512 3288
rect 3128 3272 3144 3288
rect 3528 3272 3544 3288
rect 3896 3272 3912 3288
rect 840 3252 856 3268
rect 2296 3252 2312 3268
rect 3448 3252 3464 3268
rect 3624 3252 3640 3268
rect 56 3232 72 3248
rect 184 3232 216 3248
rect 264 3232 280 3248
rect 456 3232 472 3248
rect 648 3232 664 3248
rect 904 3232 920 3248
rect 1000 3232 1016 3248
rect 1304 3232 1320 3248
rect 1352 3232 1368 3248
rect 1800 3232 1816 3248
rect 1880 3232 1896 3248
rect 2024 3232 2040 3248
rect 2136 3232 2152 3248
rect 2424 3232 2440 3248
rect 2488 3232 2504 3248
rect 2648 3232 2664 3248
rect 2712 3232 2728 3248
rect 2904 3232 2920 3248
rect 3224 3232 3240 3248
rect 3736 3232 3752 3248
rect 3784 3232 3800 3248
rect 4136 3232 4152 3248
rect 4200 3232 4216 3248
rect 4392 3232 4408 3248
rect 4712 3232 4728 3248
rect 5128 3232 5144 3248
rect 5224 3232 5240 3248
rect 5352 3232 5368 3248
rect 5416 3232 5432 3248
rect 5544 3232 5560 3248
rect 5656 3232 5672 3248
rect 5736 3232 5752 3248
rect 5896 3232 5912 3248
rect 925 3202 961 3218
rect 2973 3202 3009 3218
rect 5021 3202 5057 3218
rect 3016 3172 3032 3188
rect 3768 3172 3784 3188
rect 4984 3172 5000 3188
rect 5320 3172 5336 3188
rect 4664 3152 4680 3168
rect 2904 3132 2920 3148
rect 4632 3132 4648 3148
rect 568 3112 584 3128
rect 808 3112 824 3128
rect 1032 3112 1048 3128
rect 1096 3112 1112 3128
rect 2520 3112 2536 3128
rect 2808 3112 2824 3128
rect 56 3092 88 3108
rect 184 3092 200 3108
rect 280 3092 296 3108
rect 328 3092 344 3108
rect 440 3092 456 3108
rect 488 3092 520 3108
rect 552 3092 568 3108
rect 632 3092 648 3108
rect 744 3092 760 3108
rect 888 3092 920 3108
rect 1016 3092 1032 3108
rect 1144 3092 1192 3108
rect 1208 3092 1224 3108
rect 1320 3092 1336 3108
rect 1368 3092 1400 3108
rect 1448 3092 1464 3108
rect 1496 3092 1512 3108
rect 1544 3092 1560 3108
rect 1592 3092 1624 3108
rect 1640 3092 1656 3108
rect 1672 3092 1688 3108
rect 1880 3092 1912 3108
rect 1944 3092 1960 3108
rect 1992 3092 2008 3108
rect 2024 3092 2040 3108
rect 2104 3092 2120 3108
rect 2232 3092 2264 3108
rect 2296 3092 2312 3108
rect 2376 3092 2392 3108
rect 2488 3092 2520 3108
rect 2552 3092 2568 3108
rect 2584 3092 2616 3108
rect 2680 3092 2696 3108
rect 3208 3112 3224 3128
rect 3448 3112 3464 3128
rect 4344 3112 4360 3128
rect 4600 3112 4616 3128
rect 4648 3112 4664 3128
rect 4904 3112 4920 3128
rect 2984 3092 3000 3108
rect 3048 3092 3064 3108
rect 3080 3092 3112 3108
rect 3144 3092 3160 3108
rect 3176 3092 3192 3108
rect 3240 3092 3272 3108
rect 3336 3092 3352 3108
rect 3400 3092 3416 3108
rect 3480 3092 3512 3108
rect 3560 3092 3576 3108
rect 3592 3092 3624 3108
rect 3656 3092 3672 3108
rect 3720 3092 3736 3108
rect 3864 3092 3880 3108
rect 3912 3092 3928 3108
rect 3976 3092 3992 3108
rect 4120 3092 4152 3108
rect 4184 3092 4200 3108
rect 4312 3092 4328 3108
rect 4440 3092 4456 3108
rect 4536 3092 4552 3108
rect 4568 3092 4584 3108
rect 4616 3092 4632 3108
rect 4696 3092 4712 3108
rect 4760 3092 4792 3108
rect 4888 3092 4904 3108
rect 4952 3092 4968 3108
rect 5016 3092 5032 3108
rect 5144 3092 5160 3108
rect 5176 3092 5192 3108
rect 5208 3092 5224 3108
rect 5240 3092 5272 3108
rect 5416 3092 5432 3108
rect 5496 3092 5512 3108
rect 5560 3092 5576 3108
rect 5608 3092 5624 3108
rect 5704 3092 5720 3108
rect 5736 3092 5752 3108
rect 5800 3092 5816 3108
rect 40 3076 56 3092
rect 88 3076 104 3092
rect 168 3076 184 3092
rect 216 3072 232 3088
rect 360 3072 392 3088
rect 568 3072 584 3088
rect 616 3076 632 3092
rect 1080 3088 1096 3092
rect 664 3072 680 3088
rect 760 3072 792 3088
rect 840 3072 856 3088
rect 1032 3072 1048 3088
rect 1080 3076 1112 3088
rect 1096 3072 1112 3076
rect 1224 3072 1256 3088
rect 1272 3072 1288 3088
rect 1512 3072 1544 3088
rect 1656 3072 1672 3088
rect 1736 3072 1752 3088
rect 1800 3076 1816 3092
rect 2168 3088 2184 3092
rect 1960 3072 1976 3088
rect 2120 3072 2136 3088
rect 2168 3076 2200 3088
rect 2184 3072 2200 3076
rect 2312 3072 2328 3088
rect 2360 3072 2376 3088
rect 2424 3072 2440 3088
rect 2696 3072 2712 3088
rect 2744 3072 2760 3088
rect 2856 3072 2872 3088
rect 2936 3072 2952 3088
rect 3160 3072 3176 3088
rect 3352 3072 3368 3088
rect 3416 3072 3432 3088
rect 3736 3072 3768 3088
rect 3832 3072 3848 3088
rect 3960 3072 3976 3088
rect 4040 3076 4056 3092
rect 5864 3088 5880 3092
rect 4200 3072 4216 3088
rect 4248 3072 4264 3088
rect 4328 3072 4344 3088
rect 4376 3072 4392 3088
rect 4456 3072 4472 3088
rect 4504 3072 4520 3088
rect 4584 3072 4600 3088
rect 4712 3072 4728 3088
rect 4824 3072 4840 3088
rect 4904 3072 4920 3088
rect 4968 3072 4984 3088
rect 5128 3072 5144 3088
rect 5192 3072 5208 3088
rect 5272 3072 5288 3088
rect 5512 3072 5528 3088
rect 5592 3072 5608 3088
rect 5672 3072 5688 3088
rect 5720 3072 5736 3088
rect 5784 3072 5800 3088
rect 5848 3076 5880 3088
rect 5848 3072 5864 3076
rect 5928 3072 5944 3088
rect 200 3052 216 3068
rect 376 3052 408 3068
rect 648 3052 664 3068
rect 872 3052 888 3068
rect 1288 3052 1304 3068
rect 1720 3052 1736 3068
rect 2328 3052 2344 3068
rect 2440 3052 2456 3068
rect 2760 3052 2792 3068
rect 2856 3052 2872 3068
rect 2920 3052 2936 3068
rect 3848 3052 3864 3068
rect 4216 3052 4232 3068
rect 4264 3052 4280 3068
rect 4392 3052 4408 3068
rect 4520 3052 4536 3068
rect 4840 3052 4856 3068
rect 5128 3052 5144 3068
rect 5272 3052 5288 3068
rect 5912 3052 5928 3068
rect 8 3032 24 3048
rect 120 3032 152 3048
rect 312 3032 328 3048
rect 456 3032 472 3048
rect 520 3032 536 3048
rect 696 3032 728 3048
rect 856 3032 872 3048
rect 936 3032 952 3048
rect 984 3032 1000 3048
rect 1336 3032 1352 3048
rect 1416 3032 1432 3048
rect 1464 3032 1480 3048
rect 1576 3032 1592 3048
rect 1704 3032 1720 3048
rect 1832 3032 1864 3048
rect 1912 3032 1928 3048
rect 2056 3032 2088 3048
rect 2136 3032 2152 3048
rect 2200 3032 2216 3048
rect 2264 3032 2280 3048
rect 2344 3032 2360 3048
rect 2392 3032 2408 3048
rect 2456 3032 2472 3048
rect 2632 3032 2664 3048
rect 2712 3032 2728 3048
rect 2808 3032 2824 3048
rect 2872 3032 2888 3048
rect 3016 3032 3032 3048
rect 3112 3032 3128 3048
rect 3288 3032 3320 3048
rect 3368 3032 3384 3048
rect 3528 3032 3544 3048
rect 3640 3032 3656 3048
rect 3688 3032 3704 3048
rect 3800 3032 3816 3048
rect 3896 3032 3912 3048
rect 4072 3032 4104 3048
rect 4152 3032 4168 3048
rect 4280 3032 4296 3048
rect 4408 3032 4424 3048
rect 4728 3032 4744 3048
rect 4792 3032 4808 3048
rect 4856 3032 4872 3048
rect 5320 3032 5336 3048
rect 5368 3032 5384 3048
rect 5448 3032 5480 3048
rect 5528 3032 5544 3048
rect 5640 3032 5656 3048
rect 5768 3032 5784 3048
rect 5832 3032 5848 3048
rect 5896 3032 5912 3048
rect 5960 3032 5976 3048
rect 1933 3002 1969 3018
rect 3981 3002 4017 3018
rect 56 2972 72 2988
rect 328 2972 344 2988
rect 504 2972 520 2988
rect 632 2972 648 2988
rect 776 2972 792 2988
rect 1608 2972 1624 2988
rect 1672 2972 1688 2988
rect 2280 2972 2296 2988
rect 2488 2972 2504 2988
rect 2856 2972 2872 2988
rect 3080 2972 3096 2988
rect 3208 2972 3224 2988
rect 3720 2972 3736 2988
rect 4024 2972 4040 2988
rect 4648 2972 4664 2988
rect 4840 2972 4856 2988
rect 4904 2972 4920 2988
rect 5144 2972 5160 2988
rect 5288 2972 5304 2988
rect 5544 2972 5560 2988
rect 5720 2972 5736 2988
rect 120 2952 136 2968
rect 184 2952 200 2968
rect 248 2952 264 2968
rect 392 2952 408 2968
rect 456 2952 472 2968
rect 520 2952 536 2968
rect 648 2952 664 2968
rect 712 2952 728 2968
rect 840 2952 856 2968
rect 952 2952 968 2968
rect 1000 2952 1016 2968
rect 1048 2952 1064 2968
rect 1112 2952 1128 2968
rect 1176 2952 1192 2968
rect 1336 2952 1368 2968
rect 1464 2952 1480 2968
rect 1592 2952 1608 2968
rect 1784 2952 1800 2968
rect 1864 2952 1880 2968
rect 2072 2952 2088 2968
rect 2136 2952 2152 2968
rect 2200 2952 2216 2968
rect 2264 2952 2280 2968
rect 2344 2952 2360 2968
rect 2472 2952 2488 2968
rect 2584 2952 2600 2968
rect 2648 2952 2664 2968
rect 2776 2952 2792 2968
rect 2840 2952 2856 2968
rect 2920 2952 2936 2968
rect 3064 2952 3080 2968
rect 3320 2952 3336 2968
rect 3384 2952 3400 2968
rect 3640 2952 3656 2968
rect 3704 2952 3720 2968
rect 3960 2952 3976 2968
rect 4120 2952 4136 2968
rect 4200 2952 4216 2968
rect 4632 2952 4648 2968
rect 4824 2952 4840 2968
rect 5224 2952 5240 2968
rect 5304 2952 5320 2968
rect 5416 2952 5432 2968
rect 5528 2952 5544 2968
rect 5608 2952 5624 2968
rect 5736 2952 5752 2968
rect 5800 2952 5816 2968
rect 104 2932 120 2948
rect 168 2932 184 2948
rect 232 2932 248 2948
rect 312 2932 328 2948
rect 376 2932 392 2948
rect 408 2932 424 2948
rect 472 2932 488 2948
rect 536 2932 552 2948
rect 584 2932 600 2948
rect 664 2932 680 2948
rect 728 2932 744 2948
rect 824 2932 840 2948
rect 856 2932 872 2948
rect 1000 2932 1016 2948
rect 1096 2932 1112 2948
rect 1160 2932 1176 2948
rect 1320 2932 1336 2948
rect 1368 2932 1384 2948
rect 1448 2932 1480 2948
rect 1576 2932 1592 2948
rect 1656 2944 1672 2948
rect 1640 2932 1672 2944
rect 1720 2932 1736 2948
rect 1768 2932 1784 2948
rect 1848 2932 1864 2948
rect 1880 2932 1896 2948
rect 1928 2932 1944 2948
rect 2056 2932 2072 2948
rect 2120 2932 2136 2948
rect 2184 2932 2200 2948
rect 2248 2932 2264 2948
rect 2360 2932 2376 2948
rect 2488 2932 2504 2948
rect 2568 2932 2584 2948
rect 2632 2932 2648 2948
rect 2776 2932 2792 2948
rect 2824 2932 2840 2948
rect 2904 2944 2920 2948
rect 2888 2932 2920 2944
rect 2936 2932 2952 2948
rect 3048 2932 3064 2948
rect 3128 2932 3144 2948
rect 3192 2932 3208 2948
rect 3256 2932 3272 2948
rect 3304 2932 3320 2948
rect 3368 2932 3384 2948
rect 3464 2932 3480 2948
rect 3560 2932 3576 2948
rect 3624 2932 3640 2948
rect 3688 2932 3704 2948
rect 3768 2932 3784 2948
rect 3848 2932 3864 2948
rect 3944 2932 3960 2948
rect 4120 2932 4136 2948
rect 4184 2932 4200 2948
rect 4216 2932 4232 2948
rect 4312 2932 4328 2948
rect 4344 2932 4360 2948
rect 4472 2932 4488 2948
rect 4616 2932 4632 2948
rect 4696 2932 4712 2948
rect 4808 2932 4824 2948
rect 4952 2932 4968 2948
rect 4984 2932 5000 2948
rect 5096 2932 5112 2948
rect 5160 2932 5176 2948
rect 5240 2932 5256 2948
rect 5432 2932 5448 2948
rect 5512 2932 5528 2948
rect 5592 2944 5608 2948
rect 5576 2932 5608 2944
rect 5624 2932 5640 2948
rect 5752 2932 5768 2948
rect 5816 2932 5832 2948
rect 5864 2932 5880 2948
rect 1640 2928 1656 2932
rect 2888 2928 2904 2932
rect 5576 2928 5592 2932
rect 8 2912 40 2928
rect 264 2912 280 2928
rect 296 2912 312 2928
rect 360 2912 376 2928
rect 600 2912 616 2928
rect 808 2912 824 2928
rect 984 2912 1000 2928
rect 1192 2912 1224 2928
rect 1256 2912 1272 2928
rect 1416 2912 1432 2928
rect 1496 2912 1512 2928
rect 1704 2912 1720 2928
rect 1816 2912 1848 2928
rect 1976 2912 1992 2928
rect 2008 2912 2024 2928
rect 2312 2912 2328 2928
rect 2472 2912 2488 2928
rect 2664 2912 2696 2928
rect 2712 2912 2728 2928
rect 3112 2912 3128 2928
rect 3176 2912 3192 2928
rect 3240 2912 3256 2928
rect 3400 2912 3432 2928
rect 3480 2912 3528 2928
rect 3576 2912 3592 2928
rect 3752 2912 3768 2928
rect 3800 2912 3816 2928
rect 3864 2912 3880 2928
rect 3896 2912 3912 2928
rect 4056 2912 4072 2928
rect 4136 2912 4152 2928
rect 4168 2912 4184 2928
rect 4264 2912 4280 2928
rect 4296 2912 4312 2928
rect 4344 2912 4360 2928
rect 4392 2912 4424 2928
rect 4456 2912 4472 2928
rect 4488 2912 4520 2928
rect 4552 2912 4568 2928
rect 4680 2912 4696 2928
rect 4712 2912 4728 2928
rect 4744 2912 4760 2928
rect 4872 2912 4904 2928
rect 4936 2912 4952 2928
rect 4968 2912 4984 2928
rect 5032 2912 5064 2928
rect 5112 2912 5128 2928
rect 5176 2912 5192 2928
rect 5208 2912 5224 2928
rect 5320 2912 5352 2928
rect 5384 2912 5400 2928
rect 5672 2912 5704 2928
rect 5880 2912 5896 2928
rect 584 2892 600 2908
rect 1508 2892 1524 2908
rect 1528 2892 1544 2908
rect 1800 2892 1816 2908
rect 2792 2892 2808 2908
rect 3784 2892 3800 2908
rect 3128 2872 3144 2888
rect 3256 2872 3272 2888
rect 3816 2872 3832 2888
rect 4584 2872 4600 2888
rect 2600 2852 2616 2868
rect 2968 2852 2984 2868
rect 3592 2852 3608 2868
rect 72 2832 88 2848
rect 136 2832 152 2848
rect 200 2832 216 2848
rect 440 2832 456 2848
rect 696 2832 712 2848
rect 760 2832 776 2848
rect 904 2832 920 2848
rect 1064 2832 1080 2848
rect 1128 2832 1144 2848
rect 1240 2832 1256 2848
rect 1288 2832 1304 2848
rect 1400 2832 1416 2848
rect 1544 2832 1560 2848
rect 1736 2832 1752 2848
rect 1912 2832 1928 2848
rect 2024 2832 2040 2848
rect 2088 2832 2104 2848
rect 2152 2832 2168 2848
rect 2216 2832 2232 2848
rect 2392 2832 2408 2848
rect 2536 2832 2552 2848
rect 2728 2832 2744 2848
rect 3016 2832 3032 2848
rect 3336 2832 3352 2848
rect 3656 2832 3672 2848
rect 3832 2832 3848 2848
rect 3912 2832 3928 2848
rect 4072 2832 4088 2848
rect 4248 2832 4264 2848
rect 4424 2832 4440 2848
rect 4520 2832 4536 2848
rect 5272 2832 5288 2848
rect 5368 2832 5384 2848
rect 5464 2832 5496 2848
rect 5656 2832 5672 2848
rect 5784 2832 5800 2848
rect 5848 2832 5864 2848
rect 5912 2832 5928 2848
rect 925 2802 961 2818
rect 2973 2802 3009 2818
rect 5021 2802 5057 2818
rect 968 2772 984 2788
rect 1224 2772 1240 2788
rect 2392 2772 2408 2788
rect 2744 2772 2760 2788
rect 3320 2772 3336 2788
rect 3944 2772 3960 2788
rect 4088 2772 4104 2788
rect 5368 2772 5384 2788
rect 1672 2752 1688 2768
rect 3192 2732 3208 2748
rect 3768 2732 3784 2748
rect 2888 2712 2904 2728
rect 2936 2712 2952 2728
rect 24 2692 40 2708
rect 56 2692 72 2708
rect 152 2692 168 2708
rect 232 2692 248 2708
rect 296 2692 328 2708
rect 344 2692 360 2708
rect 424 2692 440 2708
rect 456 2692 488 2708
rect 520 2692 552 2708
rect 616 2692 648 2708
rect 696 2692 744 2708
rect 808 2692 856 2708
rect 936 2692 952 2708
rect 1080 2692 1096 2708
rect 1128 2692 1144 2708
rect 1160 2692 1176 2708
rect 1192 2692 1208 2708
rect 1240 2692 1256 2708
rect 1272 2692 1288 2708
rect 1352 2692 1384 2708
rect 1416 2692 1464 2708
rect 1544 2692 1592 2708
rect 1640 2692 1656 2708
rect 1800 2692 1832 2708
rect 1960 2692 1976 2708
rect 2024 2692 2056 2708
rect 2184 2692 2200 2708
rect 2280 2692 2296 2708
rect 2328 2692 2376 2708
rect 2488 2692 2504 2708
rect 2552 2692 2584 2708
rect 2680 2692 2696 2708
rect 2712 2692 2728 2708
rect 2776 2692 2792 2708
rect 2920 2692 2936 2708
rect 3016 2692 3032 2708
rect 3064 2692 3080 2708
rect 3128 2692 3144 2708
rect 3160 2692 3176 2708
rect 3272 2692 3288 2708
rect 3352 2692 3368 2708
rect 3416 2692 3464 2708
rect 3640 2692 3656 2708
rect 3736 2692 3752 2708
rect 3816 2692 3848 2708
rect 3880 2692 3896 2708
rect 3976 2692 3992 2708
rect 4024 2692 4072 2708
rect 4104 2692 4120 2708
rect 4184 2692 4200 2708
rect 4296 2692 4312 2708
rect 4360 2692 4392 2708
rect 4424 2692 4440 2708
rect 4488 2692 4504 2708
rect 4536 2692 4552 2708
rect 4600 2692 4616 2708
rect 4712 2692 4728 2708
rect 4744 2692 4760 2708
rect 4776 2692 4792 2708
rect 4840 2692 4872 2708
rect 5000 2692 5016 2708
rect 5128 2692 5144 2708
rect 5160 2692 5176 2708
rect 5192 2692 5224 2708
rect 5288 2692 5304 2708
rect 5336 2692 5352 2708
rect 5416 2692 5448 2708
rect 5480 2692 5496 2708
rect 5592 2692 5608 2708
rect 5640 2692 5656 2708
rect 5688 2692 5704 2708
rect 5752 2692 5768 2708
rect 5864 2692 5880 2708
rect 5896 2692 5912 2708
rect 5992 2692 6008 2708
rect 8 2672 24 2688
rect 88 2672 104 2688
rect 248 2672 264 2688
rect 328 2672 344 2688
rect 680 2676 696 2692
rect 872 2672 888 2688
rect 1016 2672 1032 2688
rect 1176 2672 1192 2688
rect 1592 2672 1608 2688
rect 1752 2672 1768 2688
rect 1864 2672 1880 2688
rect 1912 2672 1928 2688
rect 2072 2672 2088 2688
rect 2136 2672 2152 2688
rect 2200 2676 2216 2692
rect 2456 2672 2472 2688
rect 2520 2672 2536 2688
rect 2632 2672 2648 2688
rect 2664 2672 2680 2688
rect 2728 2672 2744 2688
rect 2840 2672 2856 2688
rect 72 2652 88 2668
rect 1000 2652 1016 2668
rect 1624 2652 1640 2668
rect 1752 2652 1768 2668
rect 1880 2652 1912 2668
rect 2056 2652 2072 2668
rect 2120 2652 2136 2668
rect 2248 2652 2264 2668
rect 2472 2652 2488 2668
rect 2536 2652 2552 2668
rect 2616 2652 2632 2668
rect 2968 2676 2984 2692
rect 3544 2688 3560 2692
rect 5544 2688 5560 2692
rect 3080 2672 3096 2688
rect 3160 2672 3176 2688
rect 3256 2672 3272 2688
rect 3368 2672 3384 2688
rect 3480 2672 3496 2688
rect 3544 2676 3592 2688
rect 3560 2672 3592 2676
rect 3608 2672 3624 2688
rect 3672 2672 3688 2688
rect 3800 2672 3816 2688
rect 4312 2672 4328 2688
rect 4440 2672 4456 2688
rect 4504 2672 4536 2688
rect 4584 2672 4600 2688
rect 4696 2672 4712 2688
rect 4760 2672 4776 2688
rect 4952 2672 4968 2688
rect 5048 2672 5064 2688
rect 5096 2672 5112 2688
rect 5304 2672 5336 2688
rect 5496 2672 5512 2688
rect 5544 2676 5576 2688
rect 5560 2672 5576 2676
rect 5672 2672 5688 2688
rect 5736 2672 5752 2688
rect 5816 2672 5832 2688
rect 3208 2652 3224 2668
rect 3240 2652 3256 2668
rect 3624 2652 3640 2668
rect 3688 2652 3704 2668
rect 4696 2652 4712 2668
rect 4824 2652 4840 2668
rect 4952 2652 4968 2668
rect 5112 2652 5128 2668
rect 5800 2652 5816 2668
rect 184 2632 216 2648
rect 264 2632 280 2648
rect 376 2632 408 2648
rect 504 2632 520 2648
rect 568 2632 600 2648
rect 648 2632 664 2648
rect 760 2632 792 2648
rect 1112 2632 1128 2648
rect 1304 2632 1336 2648
rect 1384 2632 1400 2648
rect 1480 2632 1496 2648
rect 1512 2632 1528 2648
rect 1608 2632 1624 2648
rect 1704 2632 1720 2648
rect 1768 2632 1784 2648
rect 1832 2632 1848 2648
rect 1976 2632 1992 2648
rect 2104 2632 2120 2648
rect 2168 2632 2184 2648
rect 2232 2632 2248 2648
rect 2264 2632 2280 2648
rect 2296 2632 2312 2648
rect 2424 2632 2440 2648
rect 2600 2632 2616 2648
rect 3016 2632 3032 2648
rect 3096 2632 3112 2648
rect 3192 2632 3208 2648
rect 3304 2632 3320 2648
rect 3384 2632 3400 2648
rect 3512 2632 3528 2648
rect 3704 2632 3720 2648
rect 3768 2632 3784 2648
rect 3864 2632 3880 2648
rect 3912 2632 3928 2648
rect 4152 2632 4168 2648
rect 4232 2632 4248 2648
rect 4264 2632 4280 2648
rect 4328 2632 4344 2648
rect 4392 2632 4408 2648
rect 4456 2632 4472 2648
rect 4568 2632 4584 2648
rect 4632 2632 4664 2648
rect 4888 2632 4920 2648
rect 4968 2632 4984 2648
rect 5032 2632 5048 2648
rect 5240 2632 5272 2648
rect 5384 2632 5400 2648
rect 5448 2632 5464 2648
rect 5512 2632 5528 2648
rect 5608 2632 5624 2648
rect 5720 2632 5736 2648
rect 5784 2632 5800 2648
rect 5848 2632 5864 2648
rect 5944 2632 5960 2648
rect 1933 2602 1969 2618
rect 3981 2602 4017 2618
rect 104 2572 120 2588
rect 472 2572 488 2588
rect 824 2572 840 2588
rect 1288 2572 1304 2588
rect 1624 2572 1640 2588
rect 40 2552 56 2568
rect 184 2552 200 2568
rect 264 2552 280 2568
rect 328 2552 344 2568
rect 392 2552 408 2568
rect 504 2552 520 2568
rect 568 2552 584 2568
rect 632 2552 648 2568
rect 808 2552 824 2568
rect 936 2552 952 2568
rect 984 2552 1000 2568
rect 1032 2552 1048 2568
rect 1112 2552 1128 2568
rect 1224 2552 1240 2568
rect 1304 2552 1320 2568
rect 1480 2552 1512 2568
rect 1736 2552 1752 2568
rect 1800 2552 1816 2568
rect 1880 2552 1896 2568
rect 1976 2552 1992 2568
rect 2120 2552 2152 2568
rect 2200 2552 2216 2568
rect 2312 2552 2328 2568
rect 2392 2552 2408 2568
rect 2456 2552 2472 2568
rect 2520 2552 2536 2568
rect 2760 2552 2776 2568
rect 2824 2552 2840 2568
rect 2888 2552 2904 2568
rect 3864 2572 3880 2588
rect 4584 2572 4600 2588
rect 4824 2572 4840 2588
rect 5272 2572 5288 2588
rect 5384 2572 5400 2588
rect 5656 2572 5672 2588
rect 5720 2572 5736 2588
rect 3160 2552 3176 2568
rect 3240 2552 3256 2568
rect 3304 2552 3320 2568
rect 3416 2552 3432 2568
rect 3528 2552 3544 2568
rect 3592 2552 3624 2568
rect 3848 2552 3864 2568
rect 4104 2552 4120 2568
rect 4376 2552 4392 2568
rect 4440 2552 4456 2568
rect 4568 2552 4584 2568
rect 4760 2552 4776 2568
rect 4888 2552 4904 2568
rect 4952 2552 4984 2568
rect 5240 2552 5256 2568
rect 5368 2552 5384 2568
rect 5832 2552 5848 2568
rect 5896 2552 5912 2568
rect 168 2532 184 2548
rect 248 2544 264 2548
rect 232 2532 264 2544
rect 280 2532 296 2548
rect 344 2532 360 2548
rect 392 2532 408 2548
rect 488 2532 504 2548
rect 520 2532 536 2548
rect 584 2532 600 2548
rect 792 2532 808 2548
rect 872 2544 888 2548
rect 856 2532 888 2544
rect 920 2532 936 2548
rect 1000 2532 1016 2548
rect 1112 2532 1144 2548
rect 1176 2532 1192 2548
rect 1240 2532 1256 2548
rect 1320 2532 1336 2548
rect 1416 2544 1432 2548
rect 1400 2532 1432 2544
rect 1464 2532 1480 2548
rect 1512 2532 1528 2548
rect 1576 2532 1592 2548
rect 1720 2532 1736 2548
rect 1784 2532 1800 2548
rect 1896 2532 1912 2548
rect 1992 2532 2008 2548
rect 2040 2532 2056 2548
rect 2184 2532 2200 2548
rect 2216 2532 2232 2548
rect 2296 2532 2312 2548
rect 2408 2532 2424 2548
rect 2456 2532 2488 2548
rect 2536 2532 2552 2548
rect 2632 2532 2648 2548
rect 2744 2532 2760 2548
rect 2872 2532 2888 2548
rect 2904 2532 2920 2548
rect 3016 2532 3032 2548
rect 3112 2532 3128 2548
rect 3224 2532 3240 2548
rect 3288 2532 3304 2548
rect 3432 2532 3448 2548
rect 3512 2532 3528 2548
rect 3576 2532 3592 2548
rect 3624 2532 3640 2548
rect 3736 2532 3752 2548
rect 3832 2532 3848 2548
rect 3912 2532 3928 2548
rect 4104 2532 4120 2548
rect 4280 2532 4296 2548
rect 4360 2532 4376 2548
rect 4440 2532 4456 2548
rect 4504 2532 4520 2548
rect 4552 2532 4568 2548
rect 4632 2544 4664 2548
rect 4632 2532 4680 2544
rect 4744 2532 4760 2548
rect 4872 2532 4888 2548
rect 4936 2532 4952 2548
rect 4984 2532 5000 2548
rect 5112 2532 5128 2548
rect 5176 2532 5192 2548
rect 5224 2532 5240 2548
rect 5352 2532 5368 2548
rect 232 2528 248 2532
rect 856 2528 872 2532
rect 1400 2528 1416 2532
rect 4664 2528 4680 2532
rect 5416 2528 5432 2544
rect 5832 2532 5864 2548
rect 5912 2532 5928 2548
rect 8 2512 24 2528
rect 72 2512 88 2528
rect 200 2512 216 2528
rect 696 2512 712 2528
rect 728 2512 760 2528
rect 888 2512 904 2528
rect 1048 2512 1064 2528
rect 1080 2512 1096 2528
rect 1256 2512 1272 2528
rect 1368 2512 1384 2528
rect 1656 2512 1672 2528
rect 1832 2512 1848 2528
rect 1864 2512 1880 2528
rect 2056 2512 2072 2528
rect 2088 2512 2104 2528
rect 2168 2512 2184 2528
rect 2328 2512 2344 2528
rect 2616 2512 2632 2528
rect 2664 2512 2680 2528
rect 2920 2512 2936 2528
rect 3096 2512 3112 2528
rect 3144 2512 3160 2528
rect 3192 2512 3208 2528
rect 3256 2512 3272 2528
rect 3336 2512 3352 2528
rect 3384 2512 3416 2528
rect 3704 2512 3720 2528
rect 3752 2512 3768 2528
rect 3784 2512 3800 2528
rect 3896 2512 3912 2528
rect 3944 2512 3960 2528
rect 3992 2512 4024 2528
rect 4120 2512 4136 2528
rect 4152 2512 4216 2528
rect 4264 2512 4280 2528
rect 4312 2512 4328 2528
rect 4456 2512 4472 2528
rect 4488 2512 4504 2528
rect 4616 2512 4632 2528
rect 4792 2512 4808 2528
rect 5032 2512 5048 2528
rect 5096 2512 5112 2528
rect 5160 2512 5176 2528
rect 5304 2512 5320 2528
rect 5432 2512 5480 2528
rect 5528 2512 5576 2528
rect 5608 2512 5624 2528
rect 5688 2512 5704 2528
rect 5752 2512 5784 2528
rect 2068 2492 2084 2508
rect 2088 2492 2104 2508
rect 2136 2492 2152 2508
rect 2584 2492 2600 2508
rect 2604 2492 2620 2508
rect 2648 2492 2664 2508
rect 3128 2492 3144 2508
rect 3720 2492 3736 2508
rect 5112 2492 5128 2508
rect 2024 2472 2040 2488
rect 2680 2472 2696 2488
rect 3160 2472 3176 2488
rect 3656 2472 3672 2488
rect 3688 2472 3704 2488
rect 2664 2452 2680 2468
rect 5016 2452 5032 2468
rect 136 2432 152 2448
rect 312 2432 328 2448
rect 376 2432 392 2448
rect 440 2432 456 2448
rect 552 2432 568 2448
rect 680 2432 696 2448
rect 760 2432 776 2448
rect 1160 2432 1176 2448
rect 1352 2432 1368 2448
rect 1432 2432 1448 2448
rect 1608 2432 1624 2448
rect 1688 2432 1704 2448
rect 1752 2432 1768 2448
rect 1928 2432 1944 2448
rect 2248 2432 2280 2448
rect 2360 2432 2376 2448
rect 2504 2432 2520 2448
rect 2568 2432 2584 2448
rect 2712 2432 2728 2448
rect 2776 2432 2792 2448
rect 3048 2432 3080 2448
rect 3352 2432 3368 2448
rect 3464 2432 3496 2448
rect 3544 2432 3560 2448
rect 3704 2432 3720 2448
rect 3800 2432 3816 2448
rect 3976 2432 3992 2448
rect 4056 2432 4072 2448
rect 4216 2432 4232 2448
rect 4296 2432 4312 2448
rect 4392 2432 4408 2448
rect 4520 2432 4536 2448
rect 4696 2432 4728 2448
rect 4840 2432 4856 2448
rect 4904 2432 4920 2448
rect 5192 2432 5208 2448
rect 5320 2432 5336 2448
rect 5480 2432 5496 2448
rect 5592 2432 5608 2448
rect 5880 2432 5896 2448
rect 5960 2432 5976 2448
rect 925 2402 961 2418
rect 2973 2402 3009 2418
rect 5021 2402 5057 2418
rect 424 2372 440 2388
rect 1848 2372 1864 2388
rect 3752 2372 3768 2388
rect 5304 2372 5320 2388
rect 5928 2372 5944 2388
rect 1608 2332 1624 2348
rect 2600 2332 2616 2348
rect 3992 2332 4008 2348
rect 888 2312 904 2328
rect 1176 2312 1192 2328
rect 2008 2312 2024 2328
rect 2072 2312 2088 2328
rect 2776 2312 2792 2328
rect 3112 2312 3128 2328
rect 3240 2312 3256 2328
rect 4248 2312 4264 2328
rect 4360 2312 4376 2328
rect 4440 2312 4456 2328
rect 40 2292 72 2308
rect 104 2292 136 2308
rect 168 2292 200 2308
rect 328 2292 344 2308
rect 360 2292 408 2308
rect 440 2292 456 2308
rect 472 2292 488 2308
rect 520 2292 536 2308
rect 600 2292 616 2308
rect 712 2292 728 2308
rect 872 2292 888 2308
rect 904 2292 920 2308
rect 1000 2292 1016 2308
rect 1160 2292 1176 2308
rect 1224 2292 1240 2308
rect 1384 2292 1400 2308
rect 1496 2292 1512 2308
rect 1560 2292 1592 2308
rect 1704 2292 1736 2308
rect 1752 2292 1768 2308
rect 1832 2292 1848 2308
rect 1896 2292 1912 2308
rect 2024 2292 2040 2308
rect 2088 2292 2104 2308
rect 2248 2292 2264 2308
rect 2280 2292 2296 2308
rect 2344 2292 2360 2308
rect 2456 2292 2488 2308
rect 2504 2292 2536 2308
rect 2600 2292 2616 2308
rect 2664 2292 2680 2308
rect 2712 2292 2744 2308
rect 2824 2292 2840 2308
rect 3032 2292 3080 2308
rect 3144 2292 3160 2308
rect 3192 2292 3208 2308
rect 3224 2292 3240 2308
rect 3336 2292 3352 2308
rect 3368 2292 3400 2308
rect 3464 2292 3480 2308
rect 3512 2292 3528 2308
rect 3560 2292 3576 2308
rect 3592 2292 3608 2308
rect 3704 2292 3736 2308
rect 3768 2292 3784 2308
rect 3928 2292 3944 2308
rect 4056 2292 4072 2308
rect 4088 2292 4120 2308
rect 4152 2292 4184 2308
rect 4344 2292 4360 2308
rect 216 2272 232 2288
rect 312 2272 328 2288
rect 552 2272 568 2288
rect 584 2272 600 2288
rect 664 2272 680 2288
rect 792 2272 808 2288
rect 968 2272 984 2288
rect 1080 2272 1096 2288
rect 1176 2272 1192 2288
rect 1304 2272 1320 2288
rect 1336 2272 1352 2288
rect 1464 2272 1480 2288
rect 1528 2272 1544 2288
rect 1672 2272 1688 2288
rect 1768 2272 1784 2288
rect 1832 2272 1848 2288
rect 1928 2276 1944 2292
rect 2008 2272 2024 2288
rect 2072 2272 2088 2288
rect 2152 2272 2168 2288
rect 2216 2272 2232 2288
rect 2264 2272 2280 2288
rect 2328 2272 2344 2288
rect 2408 2272 2424 2288
rect 2536 2272 2568 2288
rect 2632 2272 2664 2288
rect 2808 2276 2824 2292
rect 2840 2272 2856 2288
rect 2872 2272 2888 2288
rect 2936 2272 2952 2288
rect 3064 2272 3080 2288
rect 3112 2272 3144 2288
rect 3192 2272 3208 2288
rect 3272 2272 3288 2288
rect 3416 2272 3432 2288
rect 3448 2272 3464 2288
rect 3672 2272 3688 2288
rect 3816 2272 3832 2288
rect 3880 2276 3896 2292
rect 4200 2272 4216 2288
rect 4280 2272 4296 2288
rect 4408 2292 4424 2308
rect 4440 2292 4456 2308
rect 4472 2292 4488 2308
rect 4552 2292 4568 2308
rect 4600 2292 4616 2308
rect 4712 2292 4728 2308
rect 4744 2292 4760 2308
rect 4776 2292 4792 2308
rect 4840 2292 4856 2308
rect 4904 2292 4920 2308
rect 4936 2292 4952 2308
rect 5000 2292 5016 2308
rect 5160 2292 5176 2308
rect 5224 2292 5256 2308
rect 5448 2292 5464 2308
rect 5496 2292 5544 2308
rect 5608 2292 5624 2308
rect 5688 2292 5704 2308
rect 5720 2292 5752 2308
rect 5784 2292 5832 2308
rect 5864 2292 5880 2308
rect 5896 2292 5912 2308
rect 4408 2272 4424 2288
rect 4584 2272 4600 2288
rect 4696 2272 4712 2288
rect 4792 2272 4808 2288
rect 4888 2272 4904 2288
rect 4952 2272 4968 2288
rect 5016 2272 5032 2288
rect 5048 2272 5064 2288
rect 5096 2272 5112 2288
rect 5176 2272 5192 2288
rect 5272 2272 5288 2288
rect 5320 2272 5336 2288
rect 5416 2272 5432 2288
rect 5560 2272 5576 2288
rect 5592 2272 5608 2288
rect 200 2252 216 2268
rect 264 2252 280 2268
rect 312 2252 328 2268
rect 568 2252 584 2268
rect 648 2252 664 2268
rect 776 2252 792 2268
rect 984 2252 1000 2268
rect 1064 2252 1080 2268
rect 1304 2252 1320 2268
rect 1416 2252 1432 2268
rect 1448 2252 1464 2268
rect 1512 2252 1528 2268
rect 1688 2252 1704 2268
rect 1768 2252 1784 2268
rect 2136 2252 2152 2268
rect 2200 2252 2216 2268
rect 2392 2252 2408 2268
rect 2888 2252 2904 2268
rect 2952 2252 2968 2268
rect 3256 2252 3272 2268
rect 3432 2252 3448 2268
rect 3688 2252 3704 2268
rect 3800 2252 3816 2268
rect 4184 2252 4200 2268
rect 4296 2252 4312 2268
rect 4696 2252 4712 2268
rect 4824 2252 4840 2268
rect 4888 2252 4904 2268
rect 5112 2252 5128 2268
rect 5256 2252 5272 2268
rect 8 2232 24 2248
rect 72 2232 88 2248
rect 136 2232 152 2248
rect 248 2232 264 2248
rect 504 2232 520 2248
rect 632 2232 648 2248
rect 824 2232 856 2248
rect 1032 2232 1048 2248
rect 1112 2232 1144 2248
rect 1368 2232 1384 2248
rect 1640 2232 1656 2248
rect 2120 2232 2136 2248
rect 2184 2232 2200 2248
rect 2312 2232 2328 2248
rect 2376 2232 2392 2248
rect 2440 2232 2456 2248
rect 2696 2232 2712 2248
rect 2760 2232 2776 2248
rect 2904 2232 2920 2248
rect 2984 2232 3000 2248
rect 3176 2232 3192 2248
rect 3496 2232 3512 2248
rect 3544 2232 3560 2248
rect 3624 2232 3656 2248
rect 3912 2232 3928 2248
rect 3960 2232 3976 2248
rect 4120 2232 4136 2248
rect 4232 2232 4248 2248
rect 4264 2232 4280 2248
rect 4312 2232 4328 2248
rect 4424 2232 4440 2248
rect 4504 2232 4536 2248
rect 4632 2232 4664 2248
rect 4808 2232 4824 2248
rect 4968 2232 4984 2248
rect 5128 2232 5144 2248
rect 5192 2232 5208 2248
rect 5368 2232 5384 2248
rect 5464 2232 5480 2248
rect 5640 2232 5672 2248
rect 5752 2232 5768 2248
rect 5848 2232 5864 2248
rect 1933 2202 1969 2218
rect 3981 2202 4017 2218
rect 728 2172 744 2188
rect 840 2172 856 2188
rect 1208 2172 1224 2188
rect 1336 2172 1352 2188
rect 1720 2172 1736 2188
rect 2120 2172 2136 2188
rect 2376 2172 2392 2188
rect 2536 2172 2552 2188
rect 2888 2172 2904 2188
rect 3064 2172 3080 2188
rect 3096 2172 3112 2188
rect 3192 2172 3208 2188
rect 3256 2172 3272 2188
rect 4904 2172 4920 2188
rect 5144 2172 5160 2188
rect 5304 2172 5320 2188
rect 5560 2172 5576 2188
rect 5880 2172 5896 2188
rect 8 2152 24 2168
rect 280 2152 296 2168
rect 408 2152 424 2168
rect 472 2152 488 2168
rect 536 2152 552 2168
rect 648 2152 664 2168
rect 792 2152 808 2168
rect 856 2152 872 2168
rect 952 2152 968 2168
rect 1080 2152 1096 2168
rect 1192 2152 1208 2168
rect 1272 2152 1288 2168
rect 1400 2152 1416 2168
rect 1464 2152 1480 2168
rect 1528 2152 1544 2168
rect 1704 2152 1720 2168
rect 1832 2152 1848 2168
rect 1896 2152 1928 2168
rect 2136 2152 2152 2168
rect 2264 2152 2280 2168
rect 2392 2152 2408 2168
rect 2520 2152 2536 2168
rect 2744 2152 2776 2168
rect 2872 2152 2888 2168
rect 3080 2152 3096 2168
rect 3208 2152 3224 2168
rect 3464 2152 3480 2168
rect 3752 2152 3768 2168
rect 4232 2152 4248 2168
rect 4568 2152 4584 2168
rect 4632 2152 4648 2168
rect 4696 2152 4712 2168
rect 4840 2152 4856 2168
rect 5416 2152 5432 2168
rect 5544 2152 5560 2168
rect 5672 2152 5688 2168
rect 232 2132 248 2148
rect 264 2132 280 2148
rect 424 2132 440 2148
rect 552 2132 568 2148
rect 600 2132 616 2148
rect 632 2132 648 2148
rect 712 2144 728 2148
rect 696 2132 728 2144
rect 696 2128 712 2132
rect 760 2128 776 2144
rect 792 2132 824 2148
rect 872 2132 888 2148
rect 936 2132 952 2148
rect 1016 2144 1032 2148
rect 1016 2132 1048 2144
rect 1096 2132 1112 2148
rect 1144 2132 1160 2148
rect 1176 2132 1192 2148
rect 1288 2132 1304 2148
rect 1384 2144 1400 2148
rect 1368 2132 1400 2144
rect 1416 2132 1432 2148
rect 1480 2132 1496 2148
rect 1512 2132 1528 2148
rect 1544 2132 1560 2148
rect 1640 2132 1656 2148
rect 1688 2132 1704 2148
rect 1816 2132 1832 2148
rect 1880 2132 1896 2148
rect 2072 2132 2088 2148
rect 2152 2132 2168 2148
rect 2200 2132 2216 2148
rect 2264 2132 2280 2148
rect 2408 2132 2424 2148
rect 2456 2132 2472 2148
rect 2504 2132 2520 2148
rect 2552 2132 2568 2148
rect 2600 2132 2616 2148
rect 2696 2132 2712 2148
rect 2728 2132 2744 2148
rect 2856 2132 2872 2148
rect 2936 2132 2952 2148
rect 2984 2132 3000 2148
rect 3144 2132 3160 2148
rect 3176 2132 3192 2148
rect 3352 2132 3368 2148
rect 3416 2132 3432 2148
rect 3448 2132 3464 2148
rect 3480 2132 3496 2148
rect 3592 2132 3608 2148
rect 3736 2132 3752 2148
rect 4232 2132 4248 2148
rect 4552 2132 4568 2148
rect 4584 2132 4600 2148
rect 4648 2132 4664 2148
rect 4728 2132 4744 2148
rect 4824 2132 4840 2148
rect 4856 2132 4872 2148
rect 1032 2128 1048 2132
rect 1368 2128 1384 2132
rect 5176 2128 5192 2144
rect 72 2112 88 2128
rect 136 2112 152 2128
rect 200 2112 216 2128
rect 376 2112 392 2128
rect 664 2112 680 2128
rect 1240 2112 1272 2128
rect 1592 2112 1608 2128
rect 1624 2112 1640 2128
rect 1752 2112 1768 2128
rect 2024 2112 2040 2128
rect 2088 2112 2104 2128
rect 2216 2112 2232 2128
rect 2248 2112 2264 2128
rect 2344 2112 2360 2128
rect 2488 2112 2504 2128
rect 2616 2112 2632 2128
rect 2648 2112 2664 2128
rect 2808 2112 2824 2128
rect 2920 2112 2936 2128
rect 3000 2112 3016 2128
rect 3048 2112 3064 2128
rect 3128 2112 3144 2128
rect 3160 2112 3176 2128
rect 3224 2112 3240 2128
rect 3320 2112 3336 2128
rect 3368 2112 3384 2128
rect 3400 2112 3416 2128
rect 3496 2112 3512 2128
rect 3576 2112 3592 2128
rect 3608 2112 3640 2128
rect 3672 2112 3688 2128
rect 3768 2112 3800 2128
rect 3848 2112 3896 2128
rect 3928 2112 3960 2128
rect 4056 2112 4120 2128
rect 4152 2112 4168 2128
rect 4280 2112 4296 2128
rect 4312 2112 4328 2128
rect 4376 2112 4408 2128
rect 4424 2112 4440 2128
rect 4472 2112 4488 2128
rect 4536 2112 4552 2128
rect 4680 2112 4696 2128
rect 4728 2112 4744 2128
rect 4872 2112 4888 2128
rect 4920 2112 4952 2128
rect 4984 2112 5000 2128
rect 5032 2112 5080 2128
rect 5096 2112 5128 2128
rect 5224 2132 5240 2148
rect 5400 2132 5416 2148
rect 5432 2132 5448 2148
rect 5528 2132 5544 2148
rect 5608 2132 5624 2148
rect 5656 2132 5672 2148
rect 5784 2132 5800 2148
rect 5816 2132 5832 2148
rect 5224 2112 5240 2128
rect 5272 2112 5304 2128
rect 5336 2112 5368 2128
rect 5448 2112 5464 2128
rect 5480 2112 5496 2128
rect 5592 2112 5608 2128
rect 5688 2112 5720 2128
rect 5752 2112 5768 2128
rect 5816 2112 5832 2128
rect 5928 2132 5944 2148
rect 88 2092 104 2108
rect 152 2092 168 2108
rect 216 2092 232 2108
rect 264 2092 280 2108
rect 392 2092 408 2108
rect 1640 2092 1656 2108
rect 2072 2092 2088 2108
rect 2456 2092 2472 2108
rect 2632 2092 2648 2108
rect 2888 2092 2904 2108
rect 3336 2092 3352 2108
rect 3544 2092 3560 2108
rect 4296 2092 4312 2108
rect 4760 2092 4776 2108
rect 5496 2092 5512 2108
rect 56 2072 72 2088
rect 120 2072 136 2088
rect 184 2072 200 2088
rect 360 2072 376 2088
rect 1848 2072 1864 2088
rect 2664 2072 2680 2088
rect 3304 2072 3320 2088
rect 3704 2072 3720 2088
rect 4264 2072 4280 2088
rect 4968 2072 4984 2088
rect 5368 2072 5384 2088
rect 5816 2072 5832 2088
rect 3288 2052 3304 2068
rect 4184 2052 4200 2068
rect 4248 2052 4264 2068
rect 4360 2052 4376 2068
rect 24 2032 40 2048
rect 72 2032 88 2048
rect 136 2032 152 2048
rect 200 2032 216 2048
rect 248 2032 264 2048
rect 328 2032 344 2048
rect 376 2032 392 2048
rect 520 2032 536 2048
rect 584 2032 600 2048
rect 904 2032 920 2048
rect 1000 2032 1016 2048
rect 1064 2032 1080 2048
rect 1128 2032 1144 2048
rect 1320 2032 1336 2048
rect 1448 2032 1464 2048
rect 1576 2032 1592 2048
rect 2184 2032 2200 2048
rect 2440 2032 2456 2048
rect 2568 2032 2584 2048
rect 2680 2032 2696 2048
rect 2824 2032 2840 2048
rect 3032 2032 3048 2048
rect 3528 2032 3544 2048
rect 3656 2032 3672 2048
rect 3816 2032 3832 2048
rect 3912 2032 3928 2048
rect 4024 2032 4040 2048
rect 4136 2032 4152 2048
rect 4456 2032 4472 2048
rect 4504 2032 4520 2048
rect 4712 2032 4728 2048
rect 4792 2032 4808 2048
rect 5624 2032 5640 2048
rect 5736 2032 5752 2048
rect 925 2002 961 2018
rect 2973 2002 3009 2018
rect 5021 2002 5057 2018
rect 1832 1972 1848 1988
rect 1864 1972 1880 1988
rect 2408 1972 2424 1988
rect 2664 1972 2680 1988
rect 3288 1972 3304 1988
rect 4040 1972 4056 1988
rect 5800 1972 5816 1988
rect 1720 1952 1736 1968
rect 3880 1952 3896 1968
rect 3944 1952 3960 1968
rect 488 1932 504 1948
rect 1704 1932 1720 1948
rect 2024 1932 2040 1948
rect 2648 1932 2664 1948
rect 2888 1932 2904 1948
rect 3656 1932 3672 1948
rect 40 1912 56 1928
rect 72 1912 88 1928
rect 200 1912 216 1928
rect 280 1912 296 1928
rect 456 1912 472 1928
rect 712 1912 728 1928
rect 808 1912 824 1928
rect 888 1912 904 1928
rect 1224 1912 1240 1928
rect 1480 1912 1496 1928
rect 1736 1912 1752 1928
rect 1848 1912 1864 1928
rect 2376 1912 2392 1928
rect 2680 1912 2696 1928
rect 3192 1912 3208 1928
rect 3496 1912 3512 1928
rect 3624 1912 3640 1928
rect 4248 1912 4264 1928
rect 104 1892 120 1908
rect 168 1892 184 1908
rect 408 1892 424 1908
rect 472 1892 488 1908
rect 504 1892 552 1908
rect 600 1892 616 1908
rect 760 1892 776 1908
rect 792 1892 808 1908
rect 824 1892 856 1908
rect 920 1892 936 1908
rect 968 1892 984 1908
rect 1016 1892 1032 1908
rect 1096 1892 1112 1908
rect 1128 1892 1144 1908
rect 1208 1892 1224 1908
rect 1272 1892 1320 1908
rect 1352 1892 1368 1908
rect 1384 1892 1400 1908
rect 1432 1892 1448 1908
rect 1464 1892 1480 1908
rect 1544 1892 1592 1908
rect 1624 1892 1640 1908
rect 1656 1892 1688 1908
rect 1720 1892 1736 1908
rect 1752 1892 1768 1908
rect 1896 1892 1912 1908
rect 2136 1892 2152 1908
rect 2216 1892 2248 1908
rect 2264 1892 2280 1908
rect 2296 1892 2312 1908
rect 2328 1892 2360 1908
rect 2440 1892 2472 1908
rect 2504 1892 2520 1908
rect 2536 1892 2552 1908
rect 2584 1892 2600 1908
rect 2664 1892 2680 1908
rect 2696 1892 2728 1908
rect 2824 1892 2840 1908
rect 2936 1892 2952 1908
rect 2984 1892 3000 1908
rect 3160 1892 3176 1908
rect 3208 1892 3224 1908
rect 3256 1892 3272 1908
rect 3304 1892 3320 1908
rect 3512 1892 3528 1908
rect 3592 1892 3624 1908
rect 3640 1892 3656 1908
rect 3688 1892 3704 1908
rect 3784 1892 3800 1908
rect 3832 1892 3848 1908
rect 4184 1892 4200 1908
rect 4264 1892 4296 1908
rect 40 1872 56 1888
rect 152 1872 168 1888
rect 216 1872 232 1888
rect 328 1872 360 1888
rect 376 1872 392 1888
rect 584 1872 600 1888
rect 648 1872 664 1888
rect 712 1872 728 1888
rect 744 1872 776 1888
rect 1048 1872 1080 1888
rect 1112 1872 1128 1888
rect 1224 1872 1240 1888
rect 1320 1876 1336 1892
rect 1368 1872 1384 1888
rect 1480 1872 1496 1888
rect 1528 1876 1544 1892
rect 1768 1876 1784 1892
rect 1816 1872 1832 1888
rect 1912 1872 1928 1888
rect 1992 1872 2008 1888
rect 2056 1872 2072 1888
rect 2168 1872 2184 1888
rect 2200 1872 2216 1888
rect 2280 1872 2296 1888
rect 2424 1872 2440 1888
rect 2552 1872 2584 1888
rect 2792 1872 2808 1888
rect 2840 1872 2856 1888
rect 2904 1872 2920 1888
rect 3016 1872 3032 1888
rect 3048 1872 3064 1888
rect 3112 1872 3128 1888
rect 3144 1872 3160 1888
rect 3400 1872 3416 1888
rect 3432 1872 3448 1888
rect 3496 1872 3512 1888
rect 3704 1876 3720 1892
rect 3800 1872 3832 1888
rect 3912 1872 3928 1888
rect 3976 1872 3992 1888
rect 4056 1872 4088 1888
rect 4168 1872 4184 1888
rect 4216 1872 4232 1888
rect 4360 1892 4376 1908
rect 4472 1892 4520 1908
rect 4536 1892 4552 1908
rect 4600 1892 4616 1908
rect 4648 1892 4664 1908
rect 4696 1892 4728 1908
rect 4744 1892 4760 1908
rect 4824 1892 4840 1908
rect 4888 1892 4904 1908
rect 5016 1892 5032 1908
rect 5080 1892 5112 1908
rect 5144 1892 5160 1908
rect 5240 1892 5272 1908
rect 5304 1892 5336 1908
rect 5368 1892 5384 1908
rect 5416 1892 5432 1908
rect 5464 1892 5496 1908
rect 5528 1892 5544 1908
rect 5640 1892 5656 1908
rect 5720 1892 5736 1908
rect 5768 1892 5784 1908
rect 5848 1892 5864 1908
rect 5880 1892 5912 1908
rect 4344 1876 4360 1892
rect 5592 1888 5608 1892
rect 4376 1872 4392 1888
rect 4408 1872 4424 1888
rect 4552 1872 4568 1888
rect 4616 1872 4632 1888
rect 4728 1872 4744 1888
rect 4840 1872 4856 1888
rect 4968 1872 4984 1888
rect 5032 1872 5048 1888
rect 5208 1872 5224 1888
rect 5384 1872 5416 1888
rect 5544 1872 5560 1888
rect 5592 1876 5640 1888
rect 5608 1872 5640 1876
rect 5752 1872 5768 1888
rect 5864 1872 5880 1888
rect 8 1852 24 1868
rect 264 1852 280 1868
rect 376 1852 392 1868
rect 696 1852 712 1868
rect 1960 1852 1976 1868
rect 2008 1852 2024 1868
rect 2072 1852 2088 1868
rect 2152 1852 2168 1868
rect 2808 1852 2824 1868
rect 2872 1852 2888 1868
rect 2904 1852 2920 1868
rect 3064 1852 3080 1868
rect 3128 1852 3144 1868
rect 3224 1852 3240 1868
rect 3272 1852 3288 1868
rect 3368 1852 3384 1868
rect 3416 1852 3432 1868
rect 3640 1852 3656 1868
rect 3928 1852 3944 1868
rect 4008 1852 4024 1868
rect 4232 1852 4248 1868
rect 4424 1852 4440 1868
rect 4968 1852 4984 1868
rect 5224 1852 5240 1868
rect 136 1832 152 1848
rect 248 1832 264 1848
rect 360 1832 376 1848
rect 440 1832 456 1848
rect 568 1832 584 1848
rect 632 1832 648 1848
rect 728 1832 744 1848
rect 872 1832 888 1848
rect 952 1832 968 1848
rect 1160 1832 1192 1848
rect 1416 1832 1432 1848
rect 1608 1832 1624 1848
rect 1800 1832 1816 1848
rect 2408 1832 2424 1848
rect 2488 1832 2504 1848
rect 2616 1832 2632 1848
rect 2744 1832 2776 1848
rect 2856 1832 2872 1848
rect 3080 1832 3096 1848
rect 3336 1832 3352 1848
rect 3544 1832 3576 1848
rect 3736 1832 3768 1848
rect 3864 1832 3880 1848
rect 4120 1832 4136 1848
rect 4440 1832 4456 1848
rect 4568 1832 4584 1848
rect 4680 1832 4696 1848
rect 4776 1832 4808 1848
rect 4856 1832 4872 1848
rect 4984 1832 5000 1848
rect 5128 1832 5144 1848
rect 5176 1832 5192 1848
rect 5288 1832 5304 1848
rect 5448 1832 5464 1848
rect 5560 1832 5576 1848
rect 5672 1832 5704 1848
rect 5816 1832 5832 1848
rect 5928 1832 5944 1848
rect 1933 1802 1969 1818
rect 3981 1802 4017 1818
rect 568 1772 584 1788
rect 824 1772 840 1788
rect 1000 1772 1016 1788
rect 1224 1772 1240 1788
rect 1288 1772 1304 1788
rect 1352 1772 1384 1788
rect 1848 1772 1864 1788
rect 1880 1772 1896 1788
rect 2344 1772 2360 1788
rect 2456 1772 2472 1788
rect 2792 1772 2808 1788
rect 2968 1772 2984 1788
rect 3144 1772 3160 1788
rect 3896 1772 3912 1788
rect 4024 1772 4040 1788
rect 4200 1772 4216 1788
rect 4360 1772 4376 1788
rect 5944 1772 5960 1788
rect 88 1752 104 1768
rect 8 1732 24 1748
rect 184 1752 216 1768
rect 344 1752 360 1768
rect 392 1752 408 1768
rect 456 1752 472 1768
rect 1096 1752 1112 1768
rect 1544 1752 1560 1768
rect 1608 1752 1624 1768
rect 2024 1752 2040 1768
rect 2088 1752 2104 1768
rect 2168 1752 2184 1768
rect 2232 1752 2248 1768
rect 2408 1752 2424 1768
rect 2520 1752 2536 1768
rect 3016 1752 3032 1768
rect 3208 1752 3224 1768
rect 3272 1752 3288 1768
rect 3400 1752 3416 1768
rect 3432 1752 3448 1768
rect 3560 1752 3576 1768
rect 3688 1752 3704 1768
rect 3816 1752 3832 1768
rect 3880 1752 3896 1768
rect 4312 1752 4328 1768
rect 4424 1752 4440 1768
rect 4552 1752 4568 1768
rect 4728 1752 4744 1768
rect 4776 1752 4792 1768
rect 4936 1752 4952 1768
rect 5128 1752 5144 1768
rect 5512 1752 5528 1768
rect 5688 1752 5704 1768
rect 5816 1752 5832 1768
rect 120 1732 136 1748
rect 216 1732 232 1748
rect 408 1732 424 1748
rect 472 1732 488 1748
rect 520 1732 536 1748
rect 680 1732 696 1748
rect 760 1732 776 1748
rect 808 1732 824 1748
rect 856 1728 872 1744
rect 888 1732 904 1748
rect 936 1732 952 1748
rect 1048 1732 1064 1748
rect 1080 1732 1096 1748
rect 1128 1728 1144 1744
rect 1176 1732 1192 1748
rect 1240 1732 1256 1748
rect 1320 1728 1336 1744
rect 1528 1732 1544 1748
rect 1592 1732 1608 1748
rect 1640 1732 1656 1748
rect 1672 1732 1688 1748
rect 1752 1732 1768 1748
rect 1800 1732 1816 1748
rect 1912 1728 1928 1744
rect 2008 1732 2024 1748
rect 2072 1732 2088 1748
rect 2104 1732 2120 1748
rect 2168 1732 2184 1748
rect 2248 1732 2264 1748
rect 2392 1732 2408 1748
rect 2552 1732 2568 1748
rect 2600 1732 2616 1748
rect 2632 1732 2648 1748
rect 2664 1732 2680 1748
rect 2744 1732 2760 1748
rect 2856 1732 2872 1748
rect 2904 1728 2920 1744
rect 2952 1732 2968 1748
rect 3160 1732 3176 1748
rect 3192 1732 3208 1748
rect 3256 1732 3272 1748
rect 3304 1728 3320 1744
rect 3384 1732 3400 1748
rect 3544 1732 3560 1748
rect 3576 1732 3592 1748
rect 3672 1732 3688 1748
rect 3720 1732 3736 1748
rect 3768 1732 3784 1748
rect 3800 1732 3816 1748
rect 3864 1732 3880 1748
rect 3944 1744 3960 1748
rect 3928 1732 3960 1744
rect 4008 1732 4024 1748
rect 4120 1732 4136 1748
rect 4184 1732 4200 1748
rect 4328 1732 4344 1748
rect 4424 1732 4440 1748
rect 4552 1732 4568 1748
rect 4616 1732 4632 1748
rect 4760 1732 4776 1748
rect 4920 1732 4936 1748
rect 5192 1732 5208 1748
rect 5496 1732 5528 1748
rect 5624 1732 5640 1748
rect 5704 1732 5720 1748
rect 5768 1732 5784 1748
rect 5832 1732 5848 1748
rect 5880 1732 5896 1748
rect 3928 1728 3944 1732
rect 24 1712 40 1728
rect 152 1712 168 1728
rect 248 1712 296 1728
rect 360 1712 376 1728
rect 536 1712 552 1728
rect 616 1712 632 1728
rect 728 1712 744 1728
rect 776 1712 792 1728
rect 872 1712 888 1728
rect 904 1712 920 1728
rect 1032 1712 1048 1728
rect 1112 1712 1128 1728
rect 1176 1712 1208 1728
rect 1256 1712 1272 1728
rect 1304 1712 1320 1728
rect 1400 1712 1448 1728
rect 1464 1712 1496 1728
rect 1560 1712 1576 1728
rect 1656 1712 1672 1728
rect 1688 1712 1704 1728
rect 1768 1712 1784 1728
rect 1848 1712 1864 1728
rect 2120 1712 2136 1728
rect 2152 1712 2168 1728
rect 2216 1712 2232 1728
rect 2312 1712 2328 1728
rect 2424 1712 2440 1728
rect 2488 1712 2504 1728
rect 2584 1712 2600 1728
rect 2648 1712 2664 1728
rect 2680 1712 2712 1728
rect 2760 1712 2776 1728
rect 2840 1712 2856 1728
rect 2872 1712 2888 1728
rect 2920 1712 2952 1728
rect 3048 1712 3064 1728
rect 3112 1712 3128 1728
rect 3288 1712 3304 1728
rect 3432 1712 3448 1728
rect 3464 1712 3480 1728
rect 3512 1712 3528 1728
rect 3960 1712 3976 1728
rect 3992 1712 4008 1728
rect 4088 1712 4104 1728
rect 4136 1712 4152 1728
rect 4216 1712 4248 1728
rect 4280 1712 4312 1728
rect 4440 1712 4456 1728
rect 4472 1712 4488 1728
rect 4568 1712 4584 1728
rect 4600 1712 4616 1728
rect 4632 1712 4664 1728
rect 4696 1712 4712 1728
rect 4792 1712 4824 1728
rect 4856 1712 4872 1728
rect 4968 1712 4984 1728
rect 5016 1712 5032 1728
rect 5080 1712 5112 1728
rect 5144 1712 5192 1728
rect 5240 1712 5272 1728
rect 5288 1712 5304 1728
rect 5336 1712 5368 1728
rect 5384 1712 5400 1728
rect 5432 1712 5464 1728
rect 5544 1712 5560 1728
rect 5592 1712 5624 1728
rect 5640 1712 5656 1728
rect 5672 1712 5688 1728
rect 5800 1712 5816 1728
rect 5896 1712 5912 1728
rect 40 1692 56 1708
rect 312 1692 328 1708
rect 376 1692 392 1708
rect 440 1692 456 1708
rect 600 1692 616 1708
rect 632 1692 648 1708
rect 744 1692 760 1708
rect 808 1692 824 1708
rect 936 1692 952 1708
rect 1224 1692 1240 1708
rect 1288 1692 1304 1708
rect 1624 1692 1640 1708
rect 1800 1692 1816 1708
rect 1832 1692 1848 1708
rect 1864 1692 1880 1708
rect 2552 1692 2568 1708
rect 2616 1692 2632 1708
rect 2808 1692 2824 1708
rect 2828 1692 2844 1708
rect 3000 1692 3016 1708
rect 3352 1692 3368 1708
rect 3640 1692 3656 1708
rect 4376 1692 4392 1708
rect 344 1672 360 1688
rect 712 1672 728 1688
rect 1864 1672 1880 1688
rect 2040 1672 2056 1688
rect 3064 1672 3080 1688
rect 4264 1672 4280 1688
rect 1720 1652 1736 1668
rect 3224 1652 3240 1668
rect 168 1632 184 1648
rect 504 1632 520 1648
rect 616 1632 632 1648
rect 664 1632 680 1648
rect 728 1632 744 1648
rect 1496 1632 1512 1648
rect 2360 1632 2376 1648
rect 2728 1632 2744 1648
rect 3336 1632 3352 1648
rect 3416 1632 3432 1648
rect 3496 1632 3512 1648
rect 3624 1632 3640 1648
rect 3752 1632 3768 1648
rect 3832 1632 3848 1648
rect 4168 1632 4184 1648
rect 4680 1632 4696 1648
rect 4840 1632 4856 1648
rect 4888 1632 4904 1648
rect 5000 1632 5016 1648
rect 5304 1632 5320 1648
rect 5400 1632 5416 1648
rect 5464 1632 5480 1648
rect 5736 1632 5752 1648
rect 5864 1632 5880 1648
rect 925 1602 961 1618
rect 2973 1602 3009 1618
rect 5021 1602 5057 1618
rect 56 1572 72 1588
rect 584 1572 600 1588
rect 1208 1572 1224 1588
rect 1672 1572 1688 1588
rect 1784 1572 1800 1588
rect 1864 1572 1880 1588
rect 2264 1572 2280 1588
rect 2392 1572 2408 1588
rect 2504 1572 2520 1588
rect 2552 1572 2568 1588
rect 2712 1572 2728 1588
rect 2872 1572 2888 1588
rect 8 1552 24 1568
rect 3592 1552 3608 1568
rect 600 1532 616 1548
rect 1224 1532 1240 1548
rect 1336 1532 1352 1548
rect 2232 1532 2248 1548
rect 2408 1532 2424 1548
rect 2520 1532 2536 1548
rect 2568 1532 2584 1548
rect 424 1512 440 1528
rect 536 1512 552 1528
rect 632 1512 648 1528
rect 1048 1512 1064 1528
rect 1160 1512 1176 1528
rect 1256 1512 1272 1528
rect 1320 1512 1336 1528
rect 1384 1512 1400 1528
rect 1528 1512 1544 1528
rect 1640 1512 1656 1528
rect 2040 1512 2056 1528
rect 2120 1512 2136 1528
rect 2200 1512 2216 1528
rect 2360 1512 2392 1528
rect 2440 1512 2472 1528
rect 2488 1512 2504 1528
rect 2600 1512 2616 1528
rect 2644 1512 2660 1528
rect 2664 1512 2680 1528
rect 2888 1532 2904 1548
rect 3112 1532 3128 1548
rect 4232 1532 4248 1548
rect 4744 1532 4760 1548
rect 2952 1512 2968 1528
rect 40 1492 56 1508
rect 88 1492 104 1508
rect 136 1492 152 1508
rect 328 1490 344 1506
rect 392 1492 408 1508
rect 440 1492 456 1508
rect 520 1492 536 1508
rect 616 1492 632 1508
rect 664 1492 680 1508
rect 712 1492 728 1508
rect 744 1492 760 1508
rect 776 1492 792 1508
rect 808 1492 824 1508
rect 840 1492 856 1508
rect 984 1492 1000 1508
rect 1064 1492 1080 1508
rect 1240 1492 1256 1508
rect 1288 1492 1320 1508
rect 1432 1492 1448 1508
rect 1464 1492 1480 1508
rect 1512 1492 1576 1508
rect 1608 1492 1624 1508
rect 1656 1492 1672 1508
rect 1704 1492 1720 1508
rect 1736 1492 1752 1508
rect 1896 1492 1928 1508
rect 1976 1492 1992 1508
rect 2008 1492 2024 1508
rect 2056 1492 2072 1508
rect 2104 1492 2120 1508
rect 2184 1492 2200 1508
rect 2216 1492 2232 1508
rect 2392 1492 2408 1508
rect 2504 1492 2520 1508
rect 2584 1492 2600 1508
rect 2632 1492 2648 1508
rect 2680 1492 2696 1508
rect 2728 1492 2744 1508
rect 2840 1492 2856 1508
rect 2872 1492 2888 1508
rect 3112 1512 3128 1528
rect 3176 1512 3192 1528
rect 3224 1512 3240 1528
rect 3272 1512 3288 1528
rect 3384 1512 3400 1528
rect 3448 1512 3464 1528
rect 3496 1512 3512 1528
rect 3528 1512 3544 1528
rect 3672 1512 3688 1528
rect 4104 1512 4120 1528
rect 4264 1512 4280 1528
rect 4344 1512 4360 1528
rect 4392 1512 4408 1528
rect 3032 1492 3048 1508
rect 3096 1492 3112 1508
rect 3128 1492 3144 1508
rect 3288 1492 3320 1508
rect 3368 1492 3384 1508
rect 3656 1492 3672 1508
rect 3720 1492 3752 1508
rect 3816 1492 3848 1508
rect 3912 1492 3928 1508
rect 4008 1492 4024 1508
rect 4168 1492 4184 1508
rect 4248 1492 4264 1508
rect 4296 1492 4312 1508
rect 4456 1492 4472 1508
rect 4584 1492 4600 1508
rect 4616 1492 4632 1508
rect 4664 1492 4680 1508
rect 4712 1492 4744 1508
rect 4776 1492 4792 1508
rect 4808 1492 4840 1508
rect 4872 1492 4888 1508
rect 5080 1492 5112 1508
rect 5144 1492 5160 1508
rect 5192 1492 5208 1508
rect 5240 1492 5304 1508
rect 5368 1492 5384 1508
rect 5400 1492 5432 1508
rect 5528 1492 5544 1508
rect 5640 1492 5656 1508
rect 5704 1492 5720 1508
rect 5800 1492 5816 1508
rect 5880 1492 5912 1508
rect 1368 1488 1384 1492
rect 104 1472 120 1488
rect 152 1472 168 1488
rect 264 1472 280 1488
rect 360 1472 376 1488
rect 456 1472 472 1488
rect 568 1472 584 1488
rect 648 1472 664 1488
rect 776 1472 792 1488
rect 824 1472 840 1488
rect 904 1472 920 1488
rect 968 1472 984 1488
rect 1080 1472 1096 1488
rect 1128 1472 1144 1488
rect 1192 1472 1208 1488
rect 1272 1472 1288 1488
rect 1368 1476 1400 1488
rect 1384 1472 1400 1476
rect 1592 1472 1608 1488
rect 1720 1472 1736 1488
rect 1816 1472 1832 1488
rect 1928 1476 1944 1492
rect 2120 1472 2136 1488
rect 2168 1476 2184 1492
rect 2296 1472 2312 1488
rect 2328 1472 2344 1488
rect 2472 1472 2488 1488
rect 2616 1472 2632 1488
rect 2808 1472 2824 1488
rect 2920 1472 2936 1488
rect 3032 1472 3048 1488
rect 3096 1472 3112 1488
rect 3208 1472 3224 1488
rect 3256 1472 3272 1488
rect 3320 1472 3336 1488
rect 3384 1472 3400 1488
rect 3432 1472 3448 1488
rect 3496 1472 3512 1488
rect 3528 1472 3544 1488
rect 3576 1472 3592 1488
rect 3608 1472 3624 1488
rect 3672 1472 3688 1488
rect 3784 1472 3800 1488
rect 3928 1472 3944 1488
rect 4008 1472 4024 1488
rect 4072 1472 4088 1488
rect 4136 1472 4152 1488
rect 4280 1472 4296 1488
rect 4376 1472 4392 1488
rect 4424 1472 4440 1488
rect 4488 1472 4520 1488
rect 4568 1472 4584 1488
rect 4792 1472 4808 1488
rect 4904 1472 4920 1488
rect 5000 1472 5016 1488
rect 5480 1472 5496 1488
rect 5544 1476 5560 1492
rect 5608 1472 5624 1488
rect 5752 1476 5768 1492
rect 5784 1472 5800 1488
rect 5912 1472 5928 1488
rect 5960 1472 5976 1488
rect 408 1452 424 1468
rect 472 1452 488 1468
rect 808 1452 824 1468
rect 888 1452 904 1468
rect 936 1452 952 1468
rect 1032 1452 1048 1468
rect 1096 1452 1112 1468
rect 1832 1452 1848 1468
rect 2232 1452 2248 1468
rect 2312 1452 2328 1468
rect 2808 1452 2824 1468
rect 3048 1452 3064 1468
rect 3128 1452 3144 1468
rect 3192 1452 3208 1468
rect 3416 1452 3432 1468
rect 3512 1452 3528 1468
rect 3800 1452 3816 1468
rect 3944 1452 3960 1468
rect 3992 1452 4008 1468
rect 4088 1452 4104 1468
rect 4152 1452 4168 1468
rect 4200 1452 4216 1468
rect 4440 1452 4456 1468
rect 4504 1452 4520 1468
rect 4568 1452 4584 1468
rect 4856 1452 4872 1468
rect 5464 1452 5480 1468
rect 5912 1452 5928 1468
rect 488 1432 504 1448
rect 696 1432 712 1448
rect 872 1432 888 1448
rect 1016 1432 1032 1448
rect 1112 1432 1128 1448
rect 1480 1432 1496 1448
rect 1768 1432 1784 1448
rect 2344 1432 2360 1448
rect 2776 1432 2792 1448
rect 3064 1432 3080 1448
rect 3224 1432 3240 1448
rect 3336 1432 3352 1448
rect 3448 1432 3464 1448
rect 3544 1432 3560 1448
rect 3624 1432 3640 1448
rect 3752 1432 3768 1448
rect 3864 1432 3896 1448
rect 4184 1432 4200 1448
rect 4248 1432 4264 1448
rect 4328 1432 4360 1448
rect 4952 1432 4968 1448
rect 5016 1432 5032 1448
rect 5112 1432 5128 1448
rect 5320 1432 5352 1448
rect 5448 1432 5464 1448
rect 5512 1432 5528 1448
rect 5576 1432 5592 1448
rect 5672 1432 5688 1448
rect 5720 1432 5736 1448
rect 5832 1432 5864 1448
rect 1933 1402 1969 1418
rect 3981 1402 4017 1418
rect 296 1372 312 1388
rect 1432 1372 1448 1388
rect 1624 1372 1640 1388
rect 1672 1372 1688 1388
rect 1720 1372 1736 1388
rect 1992 1372 2008 1388
rect 2040 1372 2056 1388
rect 2232 1372 2248 1388
rect 2632 1372 2664 1388
rect 2728 1372 2744 1388
rect 2792 1372 2808 1388
rect 2888 1372 2904 1388
rect 2936 1372 2952 1388
rect 3480 1372 3496 1388
rect 4024 1372 4040 1388
rect 4840 1372 4856 1388
rect 5352 1372 5368 1388
rect 5528 1372 5544 1388
rect 5752 1372 5768 1388
rect 488 1352 504 1368
rect 552 1352 568 1368
rect 696 1352 712 1368
rect 760 1352 776 1368
rect 792 1352 808 1368
rect 1128 1352 1144 1368
rect 1448 1352 1464 1368
rect 1688 1352 1704 1368
rect 1832 1352 1848 1368
rect 2344 1352 2360 1368
rect 2408 1352 2424 1368
rect 2520 1352 2536 1368
rect 2776 1352 2792 1368
rect 2808 1352 2824 1368
rect 3048 1352 3080 1368
rect 3112 1352 3128 1368
rect 3224 1352 3256 1368
rect 3304 1352 3320 1368
rect 8 1332 24 1348
rect 56 1332 72 1348
rect 264 1332 280 1348
rect 504 1332 520 1348
rect 568 1332 584 1348
rect 680 1332 696 1348
rect 744 1332 760 1348
rect 856 1332 888 1348
rect 968 1332 984 1348
rect 1064 1332 1080 1348
rect 1128 1332 1144 1348
rect 1192 1344 1208 1348
rect 1176 1332 1208 1344
rect 1304 1332 1320 1348
rect 1464 1332 1480 1348
rect 1656 1332 1672 1348
rect 1704 1332 1720 1348
rect 1848 1332 1864 1348
rect 1880 1332 1896 1348
rect 1928 1332 1960 1348
rect 2088 1332 2104 1348
rect 2280 1332 2296 1348
rect 2328 1332 2344 1348
rect 2360 1332 2376 1348
rect 2392 1332 2408 1348
rect 2488 1332 2536 1348
rect 40 1312 56 1328
rect 232 1314 248 1330
rect 360 1312 376 1328
rect 424 1314 440 1330
rect 1176 1328 1192 1332
rect 2600 1328 2616 1344
rect 2696 1332 2728 1348
rect 2824 1332 2840 1348
rect 2872 1332 2888 1348
rect 3032 1332 3048 1348
rect 3112 1332 3128 1348
rect 3176 1332 3192 1348
rect 3208 1332 3224 1348
rect 3288 1332 3304 1348
rect 3496 1352 3512 1368
rect 3528 1352 3544 1368
rect 3592 1352 3624 1368
rect 3880 1352 3896 1368
rect 4216 1352 4232 1368
rect 4328 1352 4344 1368
rect 4440 1352 4456 1368
rect 4504 1352 4520 1368
rect 4584 1352 4600 1368
rect 4760 1352 4776 1368
rect 4824 1352 4840 1368
rect 5144 1352 5160 1368
rect 5272 1352 5288 1368
rect 5336 1352 5352 1368
rect 3416 1332 3432 1348
rect 3464 1332 3480 1348
rect 3512 1332 3528 1348
rect 3560 1332 3576 1348
rect 3672 1332 3704 1348
rect 3736 1332 3752 1348
rect 3896 1332 3912 1348
rect 3944 1332 3960 1348
rect 4088 1332 4120 1348
rect 4200 1332 4216 1348
rect 4248 1332 4264 1348
rect 4312 1332 4328 1348
rect 4376 1332 4392 1348
rect 4424 1332 4440 1348
rect 4456 1332 4472 1348
rect 4488 1332 4504 1348
rect 4584 1332 4600 1348
rect 4728 1332 4744 1348
rect 4760 1332 4776 1348
rect 4808 1332 4824 1348
rect 4904 1332 4920 1348
rect 5000 1332 5016 1348
rect 5080 1332 5096 1348
rect 5128 1332 5144 1348
rect 5160 1332 5176 1348
rect 5256 1332 5272 1348
rect 5320 1332 5336 1348
rect 5384 1328 5400 1344
rect 5448 1332 5464 1348
rect 5656 1352 5672 1368
rect 5848 1352 5864 1368
rect 5496 1332 5512 1348
rect 5544 1332 5560 1348
rect 5656 1332 5672 1348
rect 5704 1328 5720 1344
rect 5832 1332 5848 1348
rect 5896 1328 5912 1344
rect 616 1312 632 1328
rect 792 1312 808 1328
rect 840 1312 856 1328
rect 904 1312 920 1328
rect 1048 1312 1064 1328
rect 1144 1312 1160 1328
rect 1224 1312 1240 1328
rect 1352 1312 1368 1328
rect 1384 1312 1416 1328
rect 1496 1312 1528 1328
rect 1544 1312 1560 1328
rect 1576 1312 1608 1328
rect 1640 1312 1656 1328
rect 1752 1312 1784 1328
rect 1800 1312 1816 1328
rect 1864 1312 1880 1328
rect 1896 1312 1912 1328
rect 2024 1312 2040 1328
rect 2072 1312 2088 1328
rect 2152 1312 2168 1328
rect 2216 1312 2232 1328
rect 2264 1312 2280 1328
rect 2424 1312 2440 1328
rect 2680 1312 2696 1328
rect 2760 1312 2776 1328
rect 3128 1312 3144 1328
rect 3160 1312 3176 1328
rect 3192 1312 3208 1328
rect 3320 1312 3336 1328
rect 3368 1312 3384 1328
rect 3432 1312 3464 1328
rect 3544 1312 3560 1328
rect 3608 1312 3624 1328
rect 3640 1312 3656 1328
rect 1064 1292 1080 1308
rect 1208 1292 1224 1308
rect 1368 1292 1384 1308
rect 1560 1292 1576 1308
rect 1944 1292 1960 1308
rect 2744 1292 2760 1308
rect 3768 1312 3784 1328
rect 3816 1312 3832 1328
rect 3848 1312 3880 1328
rect 3928 1312 3944 1328
rect 3960 1312 3976 1328
rect 4072 1312 4088 1328
rect 4264 1312 4280 1328
rect 4360 1312 4376 1328
rect 4520 1312 4552 1328
rect 4568 1312 4584 1328
rect 4696 1312 4728 1328
rect 4872 1312 4888 1328
rect 4904 1312 4920 1328
rect 5176 1312 5192 1328
rect 5208 1312 5240 1328
rect 5400 1312 5432 1328
rect 5560 1312 5576 1328
rect 5592 1312 5608 1328
rect 5672 1312 5688 1328
rect 5720 1312 5736 1328
rect 5784 1312 5800 1328
rect 5960 1312 5976 1328
rect 3752 1292 3768 1308
rect 4280 1292 4296 1308
rect 4344 1292 4360 1308
rect 4392 1292 4408 1308
rect 5048 1292 5064 1308
rect 632 1272 648 1288
rect 1240 1272 1256 1288
rect 1272 1272 1288 1288
rect 1336 1272 1352 1288
rect 1384 1272 1400 1288
rect 1528 1272 1544 1288
rect 2280 1272 2296 1288
rect 2776 1272 2792 1288
rect 3704 1272 3720 1288
rect 3784 1272 3800 1288
rect 4776 1272 4792 1288
rect 5800 1252 5816 1268
rect 536 1232 552 1248
rect 600 1232 616 1248
rect 712 1232 728 1248
rect 776 1232 792 1248
rect 984 1232 1000 1248
rect 1224 1232 1240 1248
rect 1288 1232 1304 1248
rect 2120 1232 2136 1248
rect 2184 1232 2200 1248
rect 2456 1232 2472 1248
rect 2856 1232 2872 1248
rect 2936 1232 2952 1248
rect 3000 1232 3016 1248
rect 3256 1232 3272 1248
rect 3352 1232 3368 1248
rect 3592 1232 3608 1248
rect 3720 1232 3736 1248
rect 3768 1232 3784 1248
rect 4024 1232 4040 1248
rect 4152 1232 4168 1248
rect 4216 1232 4232 1248
rect 4632 1232 4648 1248
rect 4664 1232 4680 1248
rect 4952 1232 4968 1248
rect 5096 1232 5112 1248
rect 5288 1232 5304 1248
rect 5608 1232 5624 1248
rect 5864 1232 5880 1248
rect 925 1202 961 1218
rect 2973 1202 3009 1218
rect 5021 1202 5057 1218
rect 2264 1172 2280 1188
rect 2424 1172 2440 1188
rect 2568 1172 2584 1188
rect 3096 1172 3112 1188
rect 3160 1172 3176 1188
rect 4136 1172 4152 1188
rect 104 1152 120 1168
rect 2472 1152 2488 1168
rect 8 1132 24 1148
rect 424 1132 440 1148
rect 792 1132 808 1148
rect 888 1132 904 1148
rect 1400 1132 1416 1148
rect 2440 1132 2456 1148
rect 2552 1132 2568 1148
rect 3144 1132 3160 1148
rect 4200 1132 4216 1148
rect 4696 1132 4712 1148
rect 5176 1132 5192 1148
rect 760 1112 776 1128
rect 824 1112 840 1128
rect 920 1112 936 1128
rect 1256 1112 1272 1128
rect 1416 1112 1432 1128
rect 1828 1112 1844 1128
rect 1848 1112 1864 1128
rect 1960 1112 1976 1128
rect 2136 1112 2152 1128
rect 2172 1112 2188 1128
rect 2308 1112 2324 1128
rect 2328 1112 2344 1128
rect 2364 1112 2380 1128
rect 2408 1112 2424 1128
rect 2584 1112 2600 1128
rect 2664 1112 2680 1128
rect 2792 1112 2808 1128
rect 2888 1112 2904 1128
rect 3048 1112 3064 1128
rect 3176 1112 3192 1128
rect 3352 1112 3368 1128
rect 3464 1112 3480 1128
rect 3576 1112 3592 1128
rect 3720 1112 3736 1128
rect 4248 1112 4264 1128
rect 4456 1112 4472 1128
rect 4792 1112 4808 1128
rect 5240 1112 5256 1128
rect 40 1092 56 1108
rect 88 1092 104 1108
rect 136 1092 152 1108
rect 328 1090 344 1106
rect 392 1092 408 1108
rect 552 1090 568 1106
rect 632 1092 648 1108
rect 904 1092 920 1108
rect 936 1092 952 1108
rect 1000 1092 1048 1108
rect 1064 1092 1080 1108
rect 1304 1092 1336 1108
rect 1480 1092 1496 1108
rect 1544 1092 1560 1108
rect 1656 1092 1672 1108
rect 1752 1092 1768 1108
rect 1816 1092 1832 1108
rect 1848 1092 1864 1108
rect 1912 1092 1928 1108
rect 1992 1092 2024 1108
rect 2056 1092 2072 1108
rect 2120 1092 2136 1108
rect 2184 1092 2200 1108
rect 2296 1092 2312 1108
rect 2376 1092 2392 1108
rect 56 1072 72 1088
rect 152 1072 168 1088
rect 360 1072 376 1088
rect 584 1072 600 1088
rect 616 1072 632 1088
rect 680 1072 696 1088
rect 712 1072 744 1088
rect 856 1072 872 1088
rect 1080 1072 1096 1088
rect 1128 1072 1144 1088
rect 408 1052 424 1068
rect 728 1052 744 1068
rect 792 1052 808 1068
rect 840 1052 856 1068
rect 1208 1072 1240 1088
rect 1352 1072 1368 1088
rect 1496 1072 1512 1088
rect 1560 1072 1576 1088
rect 1656 1072 1672 1088
rect 1688 1076 1704 1092
rect 1736 1072 1752 1088
rect 1800 1072 1816 1088
rect 1864 1072 1880 1088
rect 2008 1072 2024 1088
rect 2136 1072 2152 1088
rect 2200 1072 2216 1088
rect 2232 1072 2248 1088
rect 2280 1072 2296 1088
rect 2424 1092 2440 1108
rect 2568 1092 2584 1108
rect 2600 1092 2632 1108
rect 2680 1092 2712 1108
rect 2760 1092 2792 1108
rect 2872 1092 2888 1108
rect 2936 1092 2968 1108
rect 3016 1092 3032 1108
rect 3064 1092 3080 1108
rect 3160 1092 3176 1108
rect 3192 1092 3208 1108
rect 3272 1092 3288 1108
rect 3336 1092 3352 1108
rect 3416 1092 3432 1108
rect 3656 1092 3688 1108
rect 3880 1092 3912 1108
rect 3944 1092 3976 1108
rect 4104 1092 4120 1108
rect 4232 1092 4248 1108
rect 4344 1092 4360 1108
rect 4552 1092 4568 1108
rect 4616 1092 4632 1108
rect 4680 1092 4696 1108
rect 4824 1092 4840 1108
rect 4872 1092 4888 1108
rect 5000 1092 5016 1108
rect 5160 1092 5176 1108
rect 5224 1092 5240 1108
rect 5288 1092 5304 1108
rect 5368 1092 5384 1108
rect 5416 1092 5432 1108
rect 5480 1092 5496 1108
rect 5512 1092 5544 1108
rect 5608 1092 5640 1108
rect 5672 1092 5688 1108
rect 5704 1092 5720 1108
rect 5800 1092 5816 1108
rect 5896 1092 5912 1108
rect 4744 1088 4760 1092
rect 2504 1072 2520 1088
rect 2712 1072 2728 1088
rect 2824 1072 2840 1088
rect 2888 1072 2904 1088
rect 2984 1072 3000 1088
rect 3208 1072 3224 1088
rect 3256 1072 3272 1088
rect 3320 1072 3336 1088
rect 3416 1072 3464 1088
rect 3528 1072 3560 1088
rect 3592 1072 3608 1088
rect 3624 1072 3640 1088
rect 3752 1072 3768 1088
rect 3816 1072 3832 1088
rect 3976 1072 3992 1088
rect 4040 1072 4056 1088
rect 4120 1072 4136 1088
rect 4168 1072 4184 1088
rect 4248 1072 4264 1088
rect 4296 1072 4312 1088
rect 1160 1052 1176 1068
rect 1336 1052 1352 1068
rect 1400 1052 1416 1068
rect 2216 1052 2232 1068
rect 2520 1052 2536 1068
rect 3240 1052 3256 1068
rect 3368 1052 3384 1068
rect 3480 1052 3496 1068
rect 3640 1052 3656 1068
rect 3768 1052 3800 1068
rect 3832 1052 3848 1068
rect 4056 1052 4072 1068
rect 4184 1052 4200 1068
rect 4328 1072 4344 1088
rect 4392 1072 4408 1088
rect 4424 1072 4440 1088
rect 4488 1072 4504 1088
rect 4568 1072 4584 1088
rect 4632 1072 4648 1088
rect 4696 1072 4712 1088
rect 4744 1076 4776 1088
rect 4760 1072 4776 1076
rect 4888 1072 4904 1088
rect 4936 1072 4952 1088
rect 5048 1072 5064 1088
rect 5096 1072 5112 1088
rect 5176 1072 5192 1088
rect 5240 1072 5256 1088
rect 5368 1072 5384 1088
rect 5432 1072 5448 1088
rect 5688 1072 5704 1088
rect 5752 1072 5768 1088
rect 5816 1072 5832 1088
rect 5864 1072 5880 1088
rect 5912 1076 5928 1092
rect 4440 1052 4456 1068
rect 4504 1052 4520 1068
rect 4952 1052 4968 1068
rect 5112 1052 5128 1068
rect 5320 1052 5336 1068
rect 5752 1052 5768 1068
rect 5880 1052 5896 1068
rect 664 1032 680 1048
rect 808 1032 824 1048
rect 904 1032 920 1048
rect 1096 1032 1112 1048
rect 1272 1032 1288 1048
rect 1448 1032 1464 1048
rect 1608 1032 1624 1048
rect 1720 1032 1736 1048
rect 1784 1032 1800 1048
rect 1912 1032 1928 1048
rect 2648 1032 2664 1048
rect 2728 1032 2744 1048
rect 2792 1032 2808 1048
rect 2840 1032 2856 1048
rect 3048 1032 3064 1048
rect 3224 1032 3240 1048
rect 3304 1032 3320 1048
rect 3384 1032 3400 1048
rect 3496 1032 3512 1048
rect 3704 1032 3720 1048
rect 3848 1032 3864 1048
rect 3912 1032 3928 1048
rect 4072 1032 4088 1048
rect 4376 1032 4392 1048
rect 4520 1032 4536 1048
rect 4584 1032 4600 1048
rect 4648 1032 4664 1048
rect 4840 1032 4856 1048
rect 4904 1032 4920 1048
rect 4968 1032 4984 1048
rect 5032 1032 5048 1048
rect 5128 1032 5144 1048
rect 5384 1032 5400 1048
rect 5448 1032 5464 1048
rect 5560 1032 5592 1048
rect 5640 1032 5656 1048
rect 5768 1032 5784 1048
rect 5832 1032 5848 1048
rect 5944 1032 5960 1048
rect 1933 1002 1969 1018
rect 3981 1002 4017 1018
rect 424 972 440 988
rect 1048 972 1064 988
rect 1464 972 1496 988
rect 1576 972 1592 988
rect 2040 972 2056 988
rect 2168 972 2184 988
rect 2232 972 2248 988
rect 2376 972 2392 988
rect 2696 972 2712 988
rect 2792 972 2824 988
rect 3016 972 3032 988
rect 3448 972 3464 988
rect 3688 972 3704 988
rect 4152 972 4168 988
rect 4232 972 4248 988
rect 4808 972 4824 988
rect 5176 972 5192 988
rect 5544 972 5560 988
rect 5864 972 5880 988
rect 56 952 72 968
rect 408 952 424 968
rect 632 952 648 968
rect 888 952 904 968
rect 968 952 1000 968
rect 1352 952 1368 968
rect 1640 952 1656 968
rect 1768 952 1784 968
rect 1832 952 1848 968
rect 1912 952 1928 968
rect 2296 952 2312 968
rect 2488 952 2504 968
rect 2888 952 2904 968
rect 3080 952 3096 968
rect 3208 952 3224 968
rect 3304 952 3320 968
rect 8 932 24 948
rect 104 932 120 948
rect 152 932 168 948
rect 360 932 376 948
rect 584 932 600 948
rect 648 932 664 948
rect 712 944 728 948
rect 712 932 744 944
rect 40 912 56 928
rect 88 912 104 928
rect 136 912 152 928
rect 328 914 344 930
rect 392 912 408 928
rect 552 914 568 930
rect 728 928 744 932
rect 792 928 808 944
rect 872 932 888 948
rect 904 932 920 948
rect 1000 932 1016 948
rect 1096 932 1112 948
rect 1208 932 1224 948
rect 1272 944 1288 948
rect 1256 932 1288 944
rect 1368 932 1384 948
rect 1544 932 1576 948
rect 1752 932 1768 948
rect 1784 932 1800 948
rect 1848 932 1864 948
rect 1880 932 1896 948
rect 1960 932 1976 948
rect 1256 928 1272 932
rect 2008 928 2024 944
rect 2056 932 2072 948
rect 2280 932 2296 948
rect 2408 928 2424 944
rect 2440 932 2456 948
rect 2472 932 2488 948
rect 2568 932 2584 948
rect 2632 932 2648 948
rect 2760 932 2776 948
rect 2936 932 2952 948
rect 3064 932 3096 948
rect 3176 932 3192 948
rect 3256 932 3272 948
rect 3384 952 3400 968
rect 3560 952 3576 968
rect 3672 952 3688 968
rect 3800 952 3816 968
rect 3864 952 3880 968
rect 3928 952 3944 968
rect 4040 952 4056 968
rect 4216 952 4232 968
rect 4344 952 4360 968
rect 4408 952 4424 968
rect 4472 952 4488 968
rect 4536 952 4552 968
rect 4600 952 4616 968
rect 4936 952 4952 968
rect 4984 952 5000 968
rect 5144 952 5160 968
rect 5272 952 5288 968
rect 5336 952 5352 968
rect 5528 952 5544 968
rect 5720 952 5736 968
rect 5784 952 5800 968
rect 5928 952 5944 968
rect 3336 932 3352 948
rect 3400 932 3416 948
rect 3496 932 3528 948
rect 3576 932 3592 948
rect 3624 932 3640 948
rect 3784 932 3800 948
rect 3848 932 3864 948
rect 3912 932 3928 948
rect 3976 932 3992 948
rect 4056 932 4072 948
rect 4200 932 4216 948
rect 4280 944 4296 948
rect 4264 932 4296 944
rect 4328 932 4344 948
rect 4392 932 4408 948
rect 4456 932 4472 948
rect 4520 932 4536 948
rect 4584 932 4600 948
rect 4664 932 4680 948
rect 4792 932 4808 948
rect 4856 932 4888 948
rect 4264 928 4280 932
rect 616 912 632 928
rect 664 912 680 928
rect 904 912 920 928
rect 1128 912 1144 928
rect 1304 912 1320 928
rect 1400 912 1448 928
rect 1512 912 1528 928
rect 1544 912 1560 928
rect 1608 912 1624 928
rect 1672 912 1688 928
rect 1928 912 1944 928
rect 2072 912 2088 928
rect 2136 912 2152 928
rect 2184 912 2216 928
rect 2248 912 2264 928
rect 2360 912 2376 928
rect 2424 912 2440 928
rect 2520 912 2536 928
rect 2616 912 2632 928
rect 2648 912 2664 928
rect 2728 912 2744 928
rect 2760 912 2776 928
rect 2840 912 2872 928
rect 2904 912 2920 928
rect 2952 912 2968 928
rect 3032 912 3048 928
rect 712 892 728 908
rect 1112 892 1128 908
rect 1176 892 1192 908
rect 1288 892 1304 908
rect 1656 892 1672 908
rect 1976 892 1992 908
rect 2104 892 2120 908
rect 2328 892 2344 908
rect 2504 892 2520 908
rect 2792 892 2808 908
rect 2920 892 2936 908
rect 3160 912 3176 928
rect 3224 912 3240 928
rect 3256 912 3272 928
rect 3480 912 3496 928
rect 3528 912 3544 928
rect 3720 912 3736 928
rect 4120 912 4136 928
rect 4616 912 4632 928
rect 4648 912 4664 928
rect 4680 912 4696 928
rect 4712 912 4744 928
rect 4776 912 4792 928
rect 4840 912 4856 928
rect 4920 912 4936 928
rect 5080 932 5096 948
rect 5128 932 5144 948
rect 5224 932 5240 948
rect 5256 932 5272 948
rect 5320 932 5336 948
rect 5400 932 5416 948
rect 5464 932 5480 948
rect 5512 932 5528 948
rect 5576 928 5592 944
rect 5704 932 5736 948
rect 5768 932 5784 948
rect 5896 932 5912 948
rect 5064 912 5080 928
rect 5208 912 5224 928
rect 5384 912 5400 928
rect 5416 912 5432 928
rect 5448 912 5464 928
rect 5640 912 5656 928
rect 5800 912 5816 928
rect 5832 912 5864 928
rect 3240 892 3256 908
rect 3544 892 3560 908
rect 3944 892 3960 908
rect 1144 872 1160 888
rect 1320 872 1336 888
rect 1688 872 1704 888
rect 1720 872 1736 888
rect 1912 872 1928 888
rect 2536 872 2552 888
rect 2888 872 2904 888
rect 3128 872 3144 888
rect 3208 872 3224 888
rect 4744 872 4760 888
rect 5464 872 5480 888
rect 2520 852 2536 868
rect 824 832 856 848
rect 1128 832 1144 848
rect 1192 832 1208 848
rect 1224 832 1240 848
rect 1304 832 1320 848
rect 1672 832 1688 848
rect 1736 832 1752 848
rect 1816 832 1832 848
rect 2680 832 2696 848
rect 3368 832 3384 848
rect 3432 832 3448 848
rect 3672 832 3688 848
rect 3816 832 3832 848
rect 3880 832 3896 848
rect 4168 832 4184 848
rect 4360 832 4376 848
rect 4424 832 4440 848
rect 4488 832 4504 848
rect 4552 832 4568 848
rect 5096 832 5112 848
rect 5176 832 5192 848
rect 5288 832 5304 848
rect 5352 832 5368 848
rect 925 802 961 818
rect 2973 802 3009 818
rect 5021 802 5057 818
rect 520 772 536 788
rect 1400 772 1416 788
rect 2088 772 2104 788
rect 2152 772 2168 788
rect 2408 772 2424 788
rect 2696 772 2712 788
rect 2840 772 2856 788
rect 2888 772 2904 788
rect 3000 772 3016 788
rect 3048 772 3064 788
rect 3352 772 3368 788
rect 3432 772 3448 788
rect 3976 772 3992 788
rect 4072 772 4088 788
rect 4504 772 4520 788
rect 4584 772 4600 788
rect 5480 772 5496 788
rect 5944 772 5960 788
rect 1528 752 1544 768
rect 4392 752 4408 768
rect 4776 752 4792 768
rect 5128 752 5144 768
rect 8 732 24 748
rect 328 732 344 748
rect 1224 732 1240 748
rect 1384 732 1400 748
rect 1784 732 1800 748
rect 1848 732 1864 748
rect 2072 732 2088 748
rect 2216 732 2232 748
rect 2360 732 2376 748
rect 2600 732 2616 748
rect 2856 732 2872 748
rect 3016 732 3032 748
rect 3144 732 3160 748
rect 3176 732 3192 748
rect 4904 732 4920 748
rect 712 712 728 728
rect 1096 712 1112 728
rect 1144 712 1160 728
rect 1240 712 1256 728
rect 1336 712 1352 728
rect 1416 712 1432 728
rect 1592 712 1608 728
rect 40 692 56 708
rect 88 692 104 708
rect 232 690 248 706
rect 296 692 312 708
rect 456 690 472 706
rect 552 692 568 708
rect 600 692 616 708
rect 648 692 680 708
rect 728 692 744 708
rect 968 692 984 708
rect 1400 692 1416 708
rect 1432 692 1448 708
rect 1480 692 1496 708
rect 1704 692 1720 708
rect 1736 692 1768 708
rect 1880 712 1896 728
rect 2104 712 2120 728
rect 2168 712 2184 728
rect 2200 712 2216 728
rect 2312 712 2328 728
rect 2376 712 2392 728
rect 2824 712 2840 728
rect 2984 712 3000 728
rect 3128 712 3144 728
rect 3192 712 3208 728
rect 3224 712 3240 728
rect 3912 712 3928 728
rect 4200 712 4216 728
rect 4520 712 4536 728
rect 1864 692 1880 708
rect 1896 692 1912 708
rect 2024 692 2056 708
rect 2088 692 2104 708
rect 2152 692 2168 708
rect 2200 692 2216 708
rect 2440 692 2456 708
rect 2536 692 2552 708
rect 2728 692 2744 708
rect 2792 692 2824 708
rect 2840 692 2856 708
rect 3000 692 3016 708
rect 3176 692 3192 708
rect 3384 692 3400 708
rect 3464 692 3480 708
rect 3624 692 3640 708
rect 3752 692 3784 708
rect 3848 692 3864 708
rect 3880 692 3912 708
rect 4136 692 4152 708
rect 4232 692 4280 708
rect 4328 692 4344 708
rect 4360 692 4376 708
rect 4424 692 4456 708
rect 4616 692 4648 708
rect 4840 692 4856 708
rect 4936 692 4984 708
rect 5096 692 5112 708
rect 5256 692 5272 708
rect 5288 692 5320 708
rect 5448 692 5464 708
rect 5544 692 5576 708
rect 5608 692 5624 708
rect 5640 692 5672 708
rect 5800 692 5816 708
rect 5896 692 5928 708
rect 5960 692 5976 708
rect 4744 688 4760 692
rect 4808 688 4824 692
rect 5416 688 5432 692
rect 5736 688 5752 692
rect 56 672 72 688
rect 264 672 280 688
rect 440 672 456 688
rect 584 672 600 688
rect 712 672 728 688
rect 776 672 792 688
rect 808 672 824 688
rect 872 672 888 688
rect 984 672 1000 688
rect 1048 672 1080 688
rect 1112 672 1128 688
rect 1176 672 1192 688
rect 1256 672 1288 688
rect 1352 672 1368 688
rect 1480 672 1496 688
rect 1560 672 1576 688
rect 1624 672 1640 688
rect 1736 672 1752 688
rect 1816 672 1832 688
rect 1896 672 1912 688
rect 2280 672 2296 688
rect 2344 672 2360 688
rect 2392 672 2408 688
rect 2504 672 2520 688
rect 2568 672 2584 688
rect 2632 672 2648 688
rect 2680 672 2696 688
rect 2744 672 2760 688
rect 2920 672 2936 688
rect 3080 672 3096 688
rect 312 652 328 668
rect 536 652 552 668
rect 568 652 584 668
rect 824 652 840 668
rect 888 652 904 668
rect 1000 652 1016 668
rect 1208 652 1224 668
rect 1656 652 1672 668
rect 1848 652 1864 668
rect 1944 652 1960 668
rect 2216 652 2232 668
rect 2248 652 2264 668
rect 2520 652 2536 668
rect 2584 652 2600 668
rect 2968 652 2984 668
rect 3112 672 3128 688
rect 3256 672 3288 688
rect 3496 672 3512 688
rect 3528 672 3544 688
rect 3560 672 3576 688
rect 3688 672 3704 688
rect 3800 672 3816 688
rect 3944 672 3960 688
rect 4040 672 4056 688
rect 4104 672 4120 688
rect 4168 672 4184 688
rect 4296 672 4312 688
rect 4376 672 4392 688
rect 4472 672 4488 688
rect 4552 672 4568 688
rect 4648 672 4664 688
rect 4680 672 4696 688
rect 4744 676 4776 688
rect 4808 676 4840 688
rect 4760 672 4776 676
rect 4824 672 4840 676
rect 5000 672 5016 688
rect 5112 672 5128 688
rect 5176 672 5192 688
rect 5240 672 5256 688
rect 5320 672 5336 688
rect 5352 672 5368 688
rect 5416 676 5448 688
rect 5432 672 5448 676
rect 5496 672 5512 688
rect 5736 676 5768 688
rect 5752 672 5768 676
rect 5816 672 5832 688
rect 5848 672 5864 688
rect 3320 652 3336 668
rect 3512 652 3528 668
rect 3576 652 3592 668
rect 3704 652 3720 668
rect 3784 652 3800 668
rect 3960 652 3976 668
rect 4056 652 4072 668
rect 4120 652 4136 668
rect 4184 652 4200 668
rect 4312 652 4328 668
rect 4456 652 4472 668
rect 4568 652 4584 668
rect 4696 652 4712 668
rect 104 632 120 648
rect 632 632 648 648
rect 760 632 776 648
rect 840 632 856 648
rect 904 632 920 648
rect 1016 632 1032 648
rect 1192 632 1208 648
rect 1288 632 1304 648
rect 1640 632 1656 648
rect 1672 632 1688 648
rect 1928 632 1944 648
rect 1992 632 2008 648
rect 2264 632 2280 648
rect 2648 632 2664 648
rect 2760 632 2776 648
rect 3176 632 3192 648
rect 3304 632 3320 648
rect 3592 632 3608 648
rect 3720 632 3736 648
rect 3832 632 3848 648
rect 4712 632 4728 648
rect 4872 632 4888 648
rect 5240 652 5256 668
rect 5368 652 5384 668
rect 5832 652 5848 668
rect 5880 652 5896 668
rect 5384 632 5400 648
rect 5512 632 5528 648
rect 5576 632 5592 648
rect 5688 632 5720 648
rect 5768 632 5784 648
rect 1933 602 1969 618
rect 3981 602 4017 618
rect 824 572 840 588
rect 1032 572 1048 588
rect 1080 572 1096 588
rect 1352 572 1368 588
rect 1736 572 1752 588
rect 1992 572 2008 588
rect 2584 572 2600 588
rect 2760 572 2776 588
rect 2904 572 2920 588
rect 3240 572 3256 588
rect 3432 572 3448 588
rect 3976 572 3992 588
rect 4072 572 4088 588
rect 4312 572 4328 588
rect 4456 572 4472 588
rect 4568 572 4600 588
rect 4712 572 4728 588
rect 4984 572 5000 588
rect 5112 572 5128 588
rect 5176 572 5192 588
rect 5336 572 5352 588
rect 5432 572 5448 588
rect 5496 572 5512 588
rect 5880 572 5896 588
rect 312 552 328 568
rect 536 552 552 568
rect 568 552 584 568
rect 600 552 616 568
rect 808 552 824 568
rect 1160 552 1176 568
rect 1256 552 1272 568
rect 8 532 24 548
rect 56 532 72 548
rect 264 532 280 548
rect 488 532 504 548
rect 584 532 600 548
rect 616 544 632 548
rect 616 532 648 544
rect 744 532 760 548
rect 856 532 888 548
rect 1016 532 1032 548
rect 1240 532 1256 548
rect 1272 532 1288 548
rect 1416 532 1432 548
rect 1448 552 1464 568
rect 1624 552 1640 568
rect 1720 552 1736 568
rect 1896 552 1912 568
rect 1944 552 1960 568
rect 2056 552 2072 568
rect 2088 552 2104 568
rect 2200 552 2216 568
rect 2536 552 2552 568
rect 2616 552 2632 568
rect 2680 552 2696 568
rect 1496 532 1528 548
rect 1656 532 1688 548
rect 1752 532 1768 548
rect 1848 532 1864 548
rect 1880 532 1896 548
rect 1928 532 1944 548
rect 2104 532 2120 548
rect 2184 532 2200 548
rect 2296 532 2312 548
rect 2328 532 2344 548
rect 2408 532 2424 548
rect 2552 532 2568 548
rect 2616 532 2632 548
rect 2808 552 2824 568
rect 2888 552 2904 568
rect 3096 552 3112 568
rect 3320 552 3336 568
rect 3512 552 3528 568
rect 3576 552 3592 568
rect 3704 552 3720 568
rect 3832 552 3864 568
rect 4120 552 4152 568
rect 4184 552 4200 568
rect 4232 552 4248 568
rect 4264 552 4280 568
rect 4376 552 4392 568
rect 4440 552 4456 568
rect 4632 552 4648 568
rect 4696 552 4712 568
rect 4888 552 4904 568
rect 4936 552 4952 568
rect 5288 552 5304 568
rect 5416 552 5432 568
rect 5608 552 5624 568
rect 5672 552 5688 568
rect 5864 552 5880 568
rect 5928 552 5944 568
rect 2712 532 2728 548
rect 2808 532 2824 548
rect 2872 532 2888 548
rect 632 528 648 532
rect 40 512 56 528
rect 88 512 104 528
rect 216 512 232 528
rect 424 512 440 528
rect 696 512 712 528
rect 760 512 776 528
rect 968 512 984 528
rect 1128 512 1144 528
rect 1224 512 1240 528
rect 1320 512 1336 528
rect 1576 512 1592 528
rect 1768 512 1784 528
rect 1800 512 1816 528
rect 2024 512 2056 528
rect 2232 512 2248 528
rect 2312 512 2328 528
rect 2344 512 2360 528
rect 2376 512 2408 528
rect 2424 512 2440 528
rect 2456 512 2472 528
rect 2488 512 2504 528
rect 2520 512 2536 528
rect 2632 512 2648 528
rect 2824 512 2840 528
rect 2856 512 2872 528
rect 2952 512 2968 528
rect 3064 532 3096 548
rect 3128 532 3160 548
rect 3320 532 3336 548
rect 3368 528 3384 544
rect 3496 532 3512 548
rect 3576 532 3592 548
rect 3640 544 3656 548
rect 3624 532 3656 544
rect 3688 532 3704 548
rect 3784 532 3800 548
rect 3816 532 3832 548
rect 3864 532 3880 548
rect 3960 532 3976 548
rect 4104 532 4120 548
rect 4168 532 4184 548
rect 4280 532 4296 548
rect 4424 532 4440 548
rect 4504 532 4520 548
rect 4616 532 4632 548
rect 4680 532 4696 548
rect 4760 532 4776 548
rect 4840 532 4856 548
rect 5096 532 5112 548
rect 5224 532 5240 548
rect 5272 532 5288 548
rect 5400 532 5416 548
rect 5592 532 5608 548
rect 5672 532 5688 548
rect 5736 532 5768 548
rect 5848 532 5864 548
rect 5976 532 5992 548
rect 3624 528 3640 532
rect 3016 512 3032 528
rect 3192 512 3224 528
rect 3336 512 3352 528
rect 3384 512 3416 528
rect 3592 512 3608 528
rect 3768 512 3784 528
rect 3912 512 3928 528
rect 4040 512 4072 528
rect 4200 512 4216 528
rect 4328 512 4344 528
rect 4488 512 4504 528
rect 4520 512 4552 528
rect 4744 512 4760 528
rect 4776 512 4792 528
rect 4808 512 4840 528
rect 4904 512 4920 528
rect 4952 512 4968 528
rect 5000 512 5016 528
rect 5080 512 5096 528
rect 5144 512 5176 528
rect 5208 512 5224 528
rect 5304 512 5320 528
rect 5368 512 5384 528
rect 5464 512 5496 528
rect 5528 512 5544 528
rect 5688 512 5704 528
rect 5720 512 5736 528
rect 5768 512 5784 528
rect 552 492 568 508
rect 744 492 760 508
rect 904 492 920 508
rect 952 492 968 508
rect 1544 492 1576 508
rect 1624 492 1640 508
rect 1704 492 1720 508
rect 1784 492 1800 508
rect 2216 492 2232 508
rect 2472 492 2488 508
rect 3032 492 3064 508
rect 3080 492 3096 508
rect 3656 492 3672 508
rect 4648 492 4664 508
rect 984 472 1000 488
rect 1048 472 1064 488
rect 1592 472 1608 488
rect 1816 472 1832 488
rect 1848 472 1864 488
rect 2248 472 2264 488
rect 2504 472 2520 488
rect 3000 472 3016 488
rect 5224 472 5240 488
rect 968 452 984 468
rect 1576 452 1592 468
rect 1688 452 1704 468
rect 1800 452 1816 468
rect 104 432 120 448
rect 296 432 312 448
rect 328 432 344 448
rect 520 432 536 448
rect 792 432 808 448
rect 1192 432 1208 448
rect 1304 432 1320 448
rect 1384 432 1400 448
rect 2072 432 2088 448
rect 2136 432 2168 448
rect 2600 432 2616 448
rect 2744 432 2760 448
rect 3272 432 3288 448
rect 3464 432 3480 448
rect 3528 432 3544 448
rect 3896 432 3912 448
rect 5560 432 5576 448
rect 5624 432 5640 448
rect 5800 432 5832 448
rect 925 402 961 418
rect 2973 402 3009 418
rect 5021 402 5057 418
rect 1432 372 1448 388
rect 1672 372 1688 388
rect 1896 372 1928 388
rect 2040 372 2056 388
rect 3928 372 3944 388
rect 4280 372 4296 388
rect 4856 372 4872 388
rect 4968 372 4984 388
rect 5160 372 5176 388
rect 5912 372 5928 388
rect 5976 372 5992 388
rect 8 332 24 348
rect 568 332 584 348
rect 1736 332 1752 348
rect 2024 332 2040 348
rect 3352 332 3368 348
rect 5112 332 5128 348
rect 1048 312 1064 328
rect 1768 312 1784 328
rect 1848 312 1864 328
rect 2056 312 2072 328
rect 2632 312 2648 328
rect 3064 312 3080 328
rect 3368 312 3384 328
rect 3528 312 3544 328
rect 4072 312 4088 328
rect 4136 312 4152 328
rect 4760 312 4776 328
rect 4920 312 4936 328
rect 5144 312 5160 328
rect 5320 312 5336 328
rect 40 292 56 308
rect 88 292 104 308
rect 216 292 232 308
rect 328 292 344 308
rect 456 292 472 308
rect 664 290 680 306
rect 728 292 744 308
rect 808 290 824 306
rect 1000 292 1016 308
rect 1064 292 1080 308
rect 1096 292 1112 308
rect 1128 292 1144 308
rect 1160 292 1192 308
rect 1208 292 1224 308
rect 1352 292 1368 308
rect 1464 292 1480 308
rect 1496 292 1512 308
rect 1528 292 1544 308
rect 1592 292 1608 308
rect 1624 292 1656 308
rect 1704 292 1736 308
rect 1752 292 1768 308
rect 1848 292 1880 308
rect 2040 292 2056 308
rect 2120 290 2136 306
rect 2328 292 2344 308
rect 2360 292 2376 308
rect 2552 292 2568 308
rect 2744 292 2760 308
rect 2776 292 2792 308
rect 2664 288 2680 292
rect 56 272 72 288
rect 264 272 280 288
rect 440 272 456 288
rect 504 272 520 288
rect 600 272 616 288
rect 696 272 712 288
rect 840 272 856 288
rect 984 272 1000 288
rect 1048 272 1064 288
rect 1112 272 1128 288
rect 1224 272 1240 288
rect 1400 272 1416 288
rect 1480 272 1496 288
rect 1544 272 1560 288
rect 1800 272 1816 288
rect 1944 272 1960 288
rect 2280 272 2296 288
rect 2376 272 2392 288
rect 2600 272 2616 288
rect 2664 276 2696 288
rect 2728 276 2744 292
rect 2840 290 2856 306
rect 2984 292 3000 308
rect 3048 292 3064 308
rect 3112 292 3128 308
rect 3144 292 3176 308
rect 3224 290 3240 306
rect 3400 292 3416 308
rect 3432 292 3448 308
rect 3496 292 3512 308
rect 3592 290 3608 306
rect 3784 290 3800 306
rect 3960 292 3976 308
rect 2680 272 2696 276
rect 744 252 760 268
rect 1576 252 1592 268
rect 1784 252 1800 268
rect 1960 252 1976 268
rect 2120 252 2136 268
rect 2264 252 2280 268
rect 3064 272 3080 288
rect 2840 252 2856 268
rect 3256 272 3272 288
rect 3416 272 3432 288
rect 3560 272 3576 288
rect 3752 272 3768 288
rect 4056 292 4072 308
rect 4120 292 4136 308
rect 4216 292 4232 308
rect 4248 292 4264 308
rect 4488 292 4504 308
rect 4552 290 4568 306
rect 4696 292 4728 308
rect 4824 292 4840 308
rect 4872 292 4888 308
rect 4936 292 4952 308
rect 5000 292 5016 308
rect 5128 292 5144 308
rect 5240 292 5256 308
rect 5288 292 5304 308
rect 5384 292 5400 308
rect 5416 292 5448 308
rect 5496 292 5512 308
rect 5576 292 5592 308
rect 5688 292 5704 308
rect 5736 292 5752 308
rect 5816 292 5832 308
rect 5864 292 5896 308
rect 5944 292 5960 308
rect 5192 288 5208 292
rect 5624 288 5640 292
rect 4072 272 4088 288
rect 4136 272 4152 288
rect 4200 272 4216 288
rect 4264 272 4280 288
rect 4312 272 4328 288
rect 4344 272 4360 288
rect 4376 272 4392 288
rect 4408 272 4424 288
rect 4440 272 4456 288
rect 4520 272 4536 288
rect 4792 272 4808 288
rect 5192 276 5240 288
rect 5208 272 5240 276
rect 5480 272 5496 288
rect 5592 276 5640 288
rect 5592 272 5624 276
rect 5672 272 5688 288
rect 5752 276 5768 292
rect 5800 272 5816 288
rect 5928 272 5944 288
rect 3480 252 3496 268
rect 3512 252 3528 268
rect 4200 252 4216 268
rect 4328 252 4344 268
rect 4392 252 4408 268
rect 4456 252 4488 268
rect 4808 252 4824 268
rect 5112 252 5128 268
rect 104 232 120 248
rect 296 232 312 248
rect 344 232 360 248
rect 536 232 552 248
rect 936 232 952 248
rect 1240 232 1256 248
rect 1560 232 1576 248
rect 2248 232 2264 248
rect 2312 232 2328 248
rect 2392 232 2408 248
rect 2696 232 2712 248
rect 2984 232 3000 248
rect 3464 232 3480 248
rect 3720 232 3736 248
rect 3912 232 3928 248
rect 4680 232 4696 248
rect 4744 232 4760 248
rect 4920 232 4936 248
rect 5064 232 5080 248
rect 5272 232 5288 248
rect 5352 232 5368 248
rect 5464 232 5480 248
rect 5528 232 5560 248
rect 5656 232 5672 248
rect 5720 232 5736 248
rect 5784 232 5800 248
rect 5848 232 5864 248
rect 1933 202 1969 218
rect 3981 202 4017 218
rect 744 172 760 188
rect 808 172 824 188
rect 1896 172 1912 188
rect 2664 172 2680 188
rect 3192 172 3208 188
rect 3272 172 3288 188
rect 4088 172 4104 188
rect 5016 172 5032 188
rect 5112 172 5128 188
rect 5176 172 5192 188
rect 5240 172 5256 188
rect 5480 172 5496 188
rect 5896 172 5912 188
rect 5976 172 5992 188
rect 72 154 88 170
rect 872 152 888 168
rect 1416 152 1432 168
rect 2120 152 2136 168
rect 2344 152 2360 168
rect 2728 152 2744 168
rect 3304 152 3320 168
rect 4104 152 4120 168
rect 4216 152 4232 168
rect 4632 152 4648 168
rect 4952 152 4968 168
rect 5160 152 5176 168
rect 5288 152 5304 168
rect 5320 152 5336 168
rect 5464 152 5480 168
rect 5592 152 5608 168
rect 5672 152 5688 168
rect 5720 152 5736 168
rect 5784 152 5800 168
rect 5848 152 5864 168
rect 8 132 24 148
rect 56 132 72 148
rect 136 132 152 148
rect 296 132 312 148
rect 392 132 408 148
rect 600 132 616 148
rect 664 132 680 148
rect 40 112 56 128
rect 88 112 120 128
rect 152 112 168 128
rect 232 112 248 128
rect 280 112 296 128
rect 328 112 344 128
rect 376 112 392 128
rect 568 114 584 130
rect 632 112 648 128
rect 680 112 696 128
rect 776 112 792 128
rect 840 112 872 128
rect 1064 132 1080 148
rect 1272 132 1288 148
rect 1336 132 1352 148
rect 1448 132 1464 148
rect 1512 132 1528 148
rect 1720 132 1736 148
rect 1832 132 1848 148
rect 2072 132 2088 148
rect 2136 132 2152 148
rect 2280 132 2296 148
rect 2360 132 2376 148
rect 2392 132 2408 148
rect 2600 132 2616 148
rect 2712 132 2728 148
rect 2776 132 2792 148
rect 2840 132 2856 148
rect 1000 112 1016 128
rect 1048 112 1064 128
rect 1240 114 1256 130
rect 1304 112 1320 128
rect 1352 112 1368 128
rect 1400 112 1416 128
rect 1480 112 1496 128
rect 1560 112 1576 128
rect 1736 112 1752 128
rect 1784 112 1800 128
rect 1896 112 1912 128
rect 2040 114 2056 130
rect 2104 112 2120 128
rect 2152 112 2168 128
rect 2184 112 2200 128
rect 2232 112 2264 128
rect 2296 112 2312 128
rect 2440 112 2456 128
rect 2616 112 2632 128
rect 2696 112 2712 128
rect 2744 112 2760 128
rect 2808 114 2824 130
rect 3112 132 3128 148
rect 3352 132 3368 148
rect 3560 132 3576 148
rect 3720 132 3736 148
rect 3864 132 3880 148
rect 3080 112 3096 128
rect 3128 112 3144 128
rect 3240 112 3256 128
rect 3320 112 3336 128
rect 3384 114 3400 130
rect 3576 112 3592 128
rect 3624 112 3640 128
rect 3672 112 3688 128
rect 3896 114 3912 130
rect 4152 132 4168 148
rect 4264 132 4280 148
rect 4472 132 4488 148
rect 4584 132 4600 148
rect 4680 132 4696 148
rect 4888 132 4904 148
rect 4968 132 4984 148
rect 5144 132 5160 148
rect 5272 132 5288 148
rect 5336 132 5352 148
rect 5400 144 5416 148
rect 5384 132 5416 144
rect 5448 132 5464 148
rect 4072 112 4088 128
rect 4104 112 4120 128
rect 4168 112 4184 128
rect 4232 112 4248 128
rect 4296 114 4312 130
rect 4488 112 4504 128
rect 4568 112 4584 128
rect 4616 112 4632 128
rect 4648 112 4664 128
rect 4712 114 4728 130
rect 5384 128 5400 132
rect 5512 128 5528 144
rect 5576 132 5592 148
rect 5608 132 5624 148
rect 5736 132 5752 148
rect 5768 132 5784 148
rect 5832 132 5848 148
rect 5928 144 5944 148
rect 5928 132 5960 144
rect 5944 128 5960 132
rect 4904 112 4920 128
rect 5000 112 5016 128
rect 5080 112 5112 128
rect 5208 112 5224 128
rect 5352 112 5368 128
rect 5416 112 5432 128
rect 5528 112 5560 128
rect 5864 112 5880 128
rect 5800 92 5816 108
rect 184 32 216 48
rect 248 32 264 48
rect 344 32 360 48
rect 712 32 728 48
rect 888 32 904 48
rect 1016 32 1032 48
rect 1384 32 1400 48
rect 1768 32 1784 48
rect 1816 32 1832 48
rect 2200 32 2216 48
rect 2328 32 2344 48
rect 2648 32 2664 48
rect 3064 32 3080 48
rect 3160 32 3176 48
rect 3608 32 3624 48
rect 3656 32 3672 48
rect 3704 32 3720 48
rect 3960 32 3976 48
rect 4200 32 4216 48
rect 4520 32 4552 48
rect 4936 32 4952 48
rect 925 2 961 18
rect 2973 2 3009 18
rect 5021 2 5057 18
<< metal2 >>
rect 349 3908 355 3912
rect 397 3908 403 4012
rect 445 3908 451 4063
rect 493 4028 499 4063
rect 13 3788 19 3832
rect 29 3763 35 3792
rect 45 3768 51 3876
rect 77 3868 83 3872
rect 24 3757 35 3763
rect 93 3708 99 3876
rect 125 3768 131 3832
rect 141 3808 147 3832
rect 173 3808 179 3876
rect 205 3848 211 3872
rect 221 3768 227 3892
rect 253 3783 259 3832
rect 237 3777 259 3783
rect 173 3744 179 3752
rect 237 3748 243 3777
rect 269 3763 275 3832
rect 301 3808 307 3892
rect 413 3868 419 3892
rect 445 3888 451 3892
rect 317 3768 323 3772
rect 264 3757 275 3763
rect 136 3737 147 3743
rect 141 3728 147 3737
rect 328 3737 339 3743
rect 333 3728 339 3737
rect 365 3728 371 3792
rect 381 3748 387 3812
rect 429 3744 435 3752
rect 477 3728 483 4012
rect 893 3988 899 4063
rect 541 3908 547 3912
rect 893 3908 899 3972
rect 1197 3968 1203 4063
rect 525 3868 531 3892
rect 669 3883 675 3892
rect 669 3877 680 3883
rect 509 3748 515 3752
rect 541 3728 547 3852
rect 557 3828 563 3832
rect 637 3828 643 3876
rect 685 3848 691 3852
rect 637 3768 643 3812
rect 605 3728 611 3732
rect 45 3508 51 3512
rect 61 3508 67 3632
rect 77 3508 83 3632
rect 173 3508 179 3512
rect 189 3508 195 3672
rect 189 3488 195 3492
rect 93 3468 99 3476
rect 253 3488 259 3652
rect 269 3508 275 3632
rect 429 3508 435 3512
rect 461 3508 467 3532
rect 477 3528 483 3712
rect 525 3628 531 3712
rect 573 3708 579 3712
rect 573 3588 579 3692
rect 621 3528 627 3752
rect 733 3688 739 3832
rect 781 3808 787 3876
rect 813 3848 819 3872
rect 829 3828 835 3892
rect 941 3888 947 3892
rect 957 3868 963 3892
rect 1053 3888 1059 3912
rect 1149 3908 1155 3952
rect 1485 3943 1491 4063
rect 2109 4008 2115 4063
rect 1485 3937 1507 3943
rect 749 3768 755 3772
rect 829 3768 835 3812
rect 861 3803 867 3832
rect 845 3797 867 3803
rect 781 3744 787 3752
rect 845 3748 851 3797
rect 861 3768 867 3772
rect 877 3728 883 3732
rect 957 3728 963 3852
rect 973 3788 979 3832
rect 1037 3808 1043 3876
rect 1069 3768 1075 3832
rect 1101 3828 1107 3876
rect 1181 3868 1187 3872
rect 1213 3868 1219 3892
rect 893 3708 899 3712
rect 744 3637 755 3643
rect 621 3508 627 3512
rect 13 3368 19 3432
rect 77 3328 83 3332
rect 109 3328 115 3452
rect 237 3448 243 3476
rect 637 3488 643 3552
rect 749 3508 755 3637
rect 285 3448 291 3476
rect 349 3468 355 3476
rect 477 3448 483 3476
rect 669 3448 675 3492
rect 829 3488 835 3672
rect 845 3568 851 3632
rect 845 3508 851 3552
rect 125 3403 131 3432
rect 141 3423 147 3432
rect 141 3417 163 3423
rect 125 3397 147 3403
rect 125 3348 131 3372
rect 141 3368 147 3397
rect 157 3348 163 3417
rect 205 3348 211 3432
rect 253 3368 259 3392
rect 317 3383 323 3432
rect 301 3377 323 3383
rect 301 3348 307 3377
rect 333 3363 339 3372
rect 381 3368 387 3432
rect 397 3408 403 3432
rect 509 3383 515 3432
rect 493 3377 515 3383
rect 328 3357 339 3363
rect 397 3348 403 3372
rect 493 3348 499 3377
rect 525 3363 531 3432
rect 589 3408 595 3432
rect 520 3357 531 3363
rect 557 3348 563 3392
rect 621 3348 627 3412
rect 637 3368 643 3372
rect 381 3328 387 3332
rect 365 3288 371 3312
rect 72 3237 83 3243
rect 61 3108 67 3212
rect 77 3108 83 3237
rect 189 3108 195 3232
rect 269 3088 275 3232
rect 365 3088 371 3112
rect 381 3088 387 3312
rect 413 3288 419 3312
rect 13 2988 19 3032
rect 45 3028 51 3076
rect 93 3068 99 3076
rect 13 2928 19 2932
rect 29 2928 35 3012
rect 125 2988 131 3032
rect 61 2968 67 2972
rect 13 2688 19 2912
rect 29 2568 35 2692
rect 77 2683 83 2832
rect 93 2688 99 2972
rect 141 2968 147 3032
rect 173 3028 179 3076
rect 397 3068 403 3272
rect 509 3108 515 3332
rect 573 3228 579 3332
rect 493 3088 499 3092
rect 573 3088 579 3112
rect 493 3068 499 3072
rect 189 2968 195 2992
rect 173 2948 179 2952
rect 109 2928 115 2932
rect 205 2888 211 3052
rect 381 3048 387 3052
rect 317 2988 323 3032
rect 381 3028 387 3032
rect 333 2988 339 2992
rect 237 2948 243 2972
rect 253 2948 259 2952
rect 317 2948 323 2952
rect 381 2948 387 2992
rect 461 2983 467 3032
rect 461 2977 483 2983
rect 397 2948 403 2952
rect 413 2948 419 2972
rect 461 2948 467 2952
rect 477 2948 483 2977
rect 301 2888 307 2912
rect 125 2837 136 2843
rect 61 2677 83 2683
rect 45 2308 51 2352
rect 61 2308 67 2677
rect 77 2528 83 2592
rect 109 2588 115 2712
rect 109 2308 115 2352
rect 125 2308 131 2837
rect 157 2368 163 2692
rect 205 2668 211 2832
rect 237 2728 243 2872
rect 237 2708 243 2712
rect 301 2708 307 2732
rect 317 2708 323 2932
rect 493 2923 499 3052
rect 509 2988 515 2992
rect 525 2983 531 3032
rect 589 2988 595 3212
rect 637 3108 643 3152
rect 653 3108 659 3232
rect 669 3088 675 3392
rect 701 3383 707 3432
rect 717 3408 723 3432
rect 685 3377 707 3383
rect 685 3348 691 3377
rect 717 3363 723 3372
rect 712 3357 723 3363
rect 781 3348 787 3352
rect 797 3344 803 3452
rect 813 3348 819 3472
rect 861 3388 867 3492
rect 973 3488 979 3752
rect 1021 3628 1027 3712
rect 1069 3688 1075 3712
rect 1101 3708 1107 3812
rect 1133 3728 1139 3852
rect 1149 3708 1155 3752
rect 1197 3748 1203 3812
rect 1245 3808 1251 3892
rect 1277 3888 1283 3892
rect 1325 3888 1331 3892
rect 1389 3888 1395 3892
rect 1341 3868 1347 3872
rect 1405 3848 1411 3872
rect 1293 3828 1299 3832
rect 1357 3808 1363 3832
rect 1245 3788 1251 3792
rect 1213 3768 1219 3772
rect 1037 3528 1043 3552
rect 1037 3508 1043 3512
rect 989 3468 995 3492
rect 925 3408 931 3432
rect 877 3328 883 3332
rect 893 3328 899 3352
rect 973 3348 979 3392
rect 1005 3363 1011 3432
rect 1069 3408 1075 3472
rect 1101 3468 1107 3472
rect 1000 3357 1011 3363
rect 1053 3348 1059 3352
rect 749 3288 755 3312
rect 621 3068 627 3072
rect 653 3048 659 3052
rect 749 3048 755 3092
rect 765 3088 771 3172
rect 781 3088 787 3272
rect 813 3128 819 3292
rect 1053 3288 1059 3332
rect 1085 3248 1091 3452
rect 1133 3348 1139 3632
rect 1165 3488 1171 3512
rect 1229 3488 1235 3632
rect 1245 3508 1251 3772
rect 1405 3768 1411 3792
rect 1261 3568 1267 3712
rect 1341 3688 1347 3752
rect 1453 3748 1459 3872
rect 1485 3808 1491 3832
rect 1416 3737 1427 3743
rect 1421 3728 1427 3737
rect 1469 3708 1475 3712
rect 1277 3508 1283 3672
rect 1357 3548 1363 3632
rect 1501 3623 1507 3937
rect 1517 3828 1523 3876
rect 1549 3803 1555 3832
rect 1549 3797 1571 3803
rect 1485 3617 1507 3623
rect 1405 3488 1411 3532
rect 1485 3508 1491 3617
rect 1293 3468 1299 3472
rect 1229 3448 1235 3452
rect 1197 3388 1203 3412
rect 1245 3348 1251 3432
rect 1341 3408 1347 3472
rect 1421 3468 1427 3492
rect 1016 3237 1027 3243
rect 845 3088 851 3232
rect 909 3228 915 3232
rect 893 3108 899 3112
rect 1021 3108 1027 3237
rect 1149 3128 1155 3312
rect 1165 3188 1171 3332
rect 1277 3328 1283 3392
rect 1341 3328 1347 3392
rect 1325 3308 1331 3312
rect 525 2977 547 2983
rect 525 2948 531 2952
rect 541 2948 547 2977
rect 589 2948 595 2972
rect 605 2928 611 3032
rect 477 2917 499 2923
rect 365 2868 371 2912
rect 173 2548 179 2652
rect 189 2588 195 2632
rect 205 2563 211 2632
rect 269 2583 275 2632
rect 269 2577 291 2583
rect 200 2557 211 2563
rect 205 2528 211 2532
rect 173 2308 179 2432
rect 221 2288 227 2572
rect 237 2544 243 2552
rect 253 2548 259 2572
rect 269 2548 275 2552
rect 285 2548 291 2577
rect 349 2548 355 2572
rect 365 2568 371 2852
rect 429 2708 435 2712
rect 461 2708 467 2812
rect 477 2708 483 2917
rect 381 2543 387 2632
rect 397 2568 403 2632
rect 477 2588 483 2652
rect 493 2548 499 2712
rect 525 2708 531 2832
rect 605 2748 611 2912
rect 605 2688 611 2732
rect 621 2728 627 3032
rect 701 3028 707 3032
rect 717 2983 723 3032
rect 717 2977 739 2983
rect 637 2963 643 2972
rect 637 2957 648 2963
rect 701 2957 712 2963
rect 669 2948 675 2952
rect 701 2908 707 2957
rect 733 2948 739 2977
rect 781 2968 787 2972
rect 829 2948 835 3032
rect 845 2968 851 2992
rect 861 2948 867 3032
rect 909 3028 915 3092
rect 1037 3088 1043 3112
rect 1101 3108 1107 3112
rect 1149 3108 1155 3112
rect 1165 3108 1171 3172
rect 1293 3108 1299 3112
rect 1085 3068 1091 3076
rect 621 2708 627 2712
rect 637 2708 643 2772
rect 701 2708 707 2832
rect 717 2708 723 2912
rect 813 2868 819 2912
rect 733 2708 739 2752
rect 829 2708 835 2932
rect 813 2688 819 2692
rect 685 2648 691 2676
rect 845 2668 851 2692
rect 509 2583 515 2632
rect 573 2628 579 2632
rect 509 2577 531 2583
rect 525 2548 531 2577
rect 589 2568 595 2632
rect 653 2563 659 2632
rect 648 2557 659 2563
rect 381 2537 392 2543
rect 573 2508 579 2552
rect 701 2528 707 2532
rect 317 2428 323 2432
rect 365 2308 371 2372
rect 381 2348 387 2412
rect 381 2308 387 2332
rect 397 2308 403 2312
rect 445 2308 451 2432
rect 477 2308 483 2352
rect 333 2283 339 2292
rect 397 2288 403 2292
rect 557 2288 563 2432
rect 653 2388 659 2472
rect 589 2288 595 2292
rect 328 2277 339 2283
rect 557 2268 563 2272
rect 653 2268 659 2372
rect 669 2288 675 2492
rect 733 2488 739 2512
rect 765 2463 771 2632
rect 781 2543 787 2632
rect 829 2563 835 2572
rect 861 2568 867 2912
rect 877 2688 883 3012
rect 941 2848 947 3032
rect 957 2948 963 2952
rect 824 2557 835 2563
rect 781 2537 792 2543
rect 861 2544 867 2552
rect 765 2457 787 2463
rect 13 2208 19 2232
rect 77 2228 83 2232
rect 141 2188 147 2232
rect 77 2128 83 2152
rect 141 2128 147 2152
rect 205 2128 211 2132
rect 29 1883 35 2032
rect 29 1877 40 1883
rect 61 1868 67 2072
rect 13 1748 19 1792
rect 93 1788 99 2092
rect 189 2088 195 2112
rect 253 2108 259 2232
rect 285 2148 291 2152
rect 269 2108 275 2132
rect 317 2128 323 2252
rect 429 2148 435 2212
rect 509 2188 515 2232
rect 573 2208 579 2252
rect 637 2228 643 2232
rect 541 2168 547 2192
rect 669 2163 675 2272
rect 664 2157 675 2163
rect 381 2128 387 2132
rect 477 2128 483 2152
rect 653 2128 659 2152
rect 669 2128 675 2132
rect 269 2088 275 2092
rect 109 1908 115 2032
rect 205 2028 211 2032
rect 173 1908 179 1912
rect 205 1908 211 1912
rect 221 1888 227 2032
rect 253 1928 259 2032
rect 333 1888 339 1892
rect 349 1888 355 2012
rect 381 1888 387 2032
rect 141 1828 147 1832
rect 253 1808 259 1832
rect 157 1728 163 1772
rect 189 1728 195 1752
rect 61 1588 67 1592
rect 173 1568 179 1632
rect 189 1548 195 1712
rect 221 1628 227 1732
rect 269 1588 275 1712
rect 333 1668 339 1872
rect 397 1788 403 2092
rect 413 1908 419 2032
rect 509 2023 515 2092
rect 685 2068 691 2432
rect 781 2283 787 2457
rect 781 2277 792 2283
rect 717 2148 723 2232
rect 733 2168 739 2172
rect 781 2168 787 2252
rect 797 2168 803 2212
rect 813 2148 819 2492
rect 893 2368 899 2512
rect 877 2317 888 2323
rect 877 2308 883 2317
rect 909 2308 915 2832
rect 973 2788 979 3052
rect 989 2943 995 3032
rect 1117 2968 1123 3092
rect 1213 3088 1219 3092
rect 1181 3008 1187 3072
rect 1181 2968 1187 2992
rect 989 2937 1000 2943
rect 1197 2928 1203 3052
rect 1213 2928 1219 2972
rect 1229 2948 1235 3072
rect 1293 3068 1299 3092
rect 1309 2928 1315 3232
rect 1325 3108 1331 3232
rect 1357 3048 1363 3232
rect 1373 3168 1379 3432
rect 1421 3388 1427 3452
rect 1416 3357 1427 3363
rect 1421 3328 1427 3357
rect 1453 3288 1459 3312
rect 1469 3248 1475 3332
rect 1485 3328 1491 3492
rect 1501 3348 1507 3432
rect 1485 3168 1491 3312
rect 1373 3108 1379 3132
rect 1485 3128 1491 3152
rect 1453 3108 1459 3112
rect 1517 3088 1523 3792
rect 1549 3763 1555 3772
rect 1544 3757 1555 3763
rect 1565 3743 1571 3797
rect 1581 3748 1587 3892
rect 1661 3888 1667 3892
rect 1645 3828 1651 3876
rect 1741 3848 1747 3892
rect 1544 3737 1571 3743
rect 1597 3708 1603 3732
rect 1645 3728 1651 3812
rect 1661 3768 1667 3812
rect 1693 3768 1699 3832
rect 1805 3828 1811 3832
rect 1805 3763 1811 3772
rect 1800 3757 1811 3763
rect 1773 3748 1779 3752
rect 1837 3748 1843 3872
rect 1917 3868 1923 3932
rect 2093 3908 2099 3912
rect 2109 3908 2115 3992
rect 2205 3988 2211 4063
rect 2253 4028 2259 4063
rect 2157 3908 2163 3912
rect 2205 3908 2211 3972
rect 1869 3808 1875 3832
rect 1869 3768 1875 3772
rect 1997 3768 2003 3876
rect 2029 3763 2035 3772
rect 2024 3757 2035 3763
rect 1672 3737 1683 3743
rect 1677 3728 1683 3737
rect 1837 3728 1843 3732
rect 1853 3728 1859 3732
rect 1901 3728 1907 3752
rect 1917 3728 1923 3732
rect 1997 3728 2003 3732
rect 2061 3728 2067 3892
rect 2125 3788 2131 3792
rect 2125 3728 2131 3772
rect 1533 3508 1539 3552
rect 1549 3508 1555 3632
rect 1565 3528 1571 3612
rect 1613 3548 1619 3632
rect 1565 3508 1571 3512
rect 1709 3508 1715 3712
rect 1581 3488 1587 3492
rect 1805 3488 1811 3512
rect 1837 3488 1843 3712
rect 1869 3528 1875 3552
rect 1869 3508 1875 3512
rect 1901 3508 1907 3712
rect 2061 3668 2067 3712
rect 2125 3708 2131 3712
rect 2141 3683 2147 3732
rect 2125 3677 2147 3683
rect 2045 3508 2051 3532
rect 2109 3508 2115 3652
rect 2125 3608 2131 3677
rect 2157 3648 2163 3892
rect 2221 3728 2227 4012
rect 2253 3908 2259 3992
rect 2397 3928 2403 4063
rect 2605 4057 2627 4063
rect 2301 3908 2307 3912
rect 2349 3908 2355 3912
rect 2397 3908 2403 3912
rect 2445 3908 2451 3932
rect 2237 3728 2243 3892
rect 2253 3888 2259 3892
rect 2317 3728 2323 3732
rect 2269 3708 2275 3712
rect 2333 3708 2339 3712
rect 2125 3508 2131 3592
rect 2173 3508 2179 3692
rect 2333 3668 2339 3692
rect 2349 3668 2355 3892
rect 2365 3748 2371 3772
rect 2365 3728 2371 3732
rect 2429 3728 2435 3812
rect 2445 3748 2451 3892
rect 2493 3808 2499 3832
rect 2509 3728 2515 3952
rect 2525 3908 2531 3912
rect 2541 3728 2547 3892
rect 2557 3768 2563 3832
rect 2573 3723 2579 3952
rect 2589 3908 2595 3912
rect 2605 3728 2611 4057
rect 2749 4028 2755 4063
rect 2621 3828 2627 3832
rect 2637 3728 2643 3892
rect 2653 3728 2659 3972
rect 2669 3848 2675 3892
rect 2685 3888 2691 3892
rect 2733 3888 2739 3892
rect 2781 3888 2787 3892
rect 2797 3888 2803 4063
rect 2829 3908 2835 4063
rect 2877 3988 2883 4063
rect 2925 4028 2931 4063
rect 2957 4057 2979 4063
rect 2749 3877 2760 3883
rect 2717 3863 2723 3872
rect 2749 3863 2755 3877
rect 2717 3857 2755 3863
rect 2701 3788 2707 3832
rect 2685 3768 2691 3772
rect 2829 3728 2835 3892
rect 2877 3888 2883 3972
rect 2909 3888 2915 3892
rect 2925 3888 2931 3892
rect 2957 3888 2963 4057
rect 2973 3888 2979 3892
rect 2845 3728 2851 3872
rect 2973 3788 2979 3872
rect 3005 3848 3011 3892
rect 2909 3728 2915 3752
rect 3005 3728 3011 3752
rect 3021 3728 3027 4063
rect 3085 3908 3091 3912
rect 3053 3888 3059 3892
rect 3117 3828 3123 3832
rect 2568 3717 2579 3723
rect 2189 3628 2195 3632
rect 2285 3588 2291 3632
rect 1677 3468 1683 3472
rect 1741 3468 1747 3472
rect 1933 3468 1939 3472
rect 1741 3448 1747 3452
rect 1549 3328 1555 3332
rect 1581 3328 1587 3392
rect 1613 3348 1619 3432
rect 1629 3428 1635 3432
rect 1661 3368 1667 3412
rect 1693 3343 1699 3432
rect 1757 3428 1763 3432
rect 1725 3368 1731 3412
rect 1757 3388 1763 3392
rect 1693 3337 1704 3343
rect 1821 3343 1827 3432
rect 1885 3368 1891 3432
rect 1981 3388 1987 3492
rect 2189 3488 2195 3512
rect 2221 3508 2227 3572
rect 2317 3508 2323 3592
rect 2381 3548 2387 3632
rect 2413 3608 2419 3712
rect 2429 3708 2435 3712
rect 2365 3508 2371 3512
rect 2429 3508 2435 3692
rect 2509 3648 2515 3712
rect 2477 3608 2483 3632
rect 2493 3543 2499 3592
rect 2477 3537 2499 3543
rect 2029 3428 2035 3432
rect 1821 3337 1832 3343
rect 1533 3088 1539 3132
rect 1597 3108 1603 3232
rect 1613 3108 1619 3112
rect 1661 3088 1667 3132
rect 1885 3128 1891 3232
rect 1885 3108 1891 3112
rect 1901 3108 1907 3112
rect 1341 2988 1347 3032
rect 1421 3008 1427 3032
rect 1469 2968 1475 3032
rect 1325 2928 1331 2932
rect 989 2868 995 2912
rect 925 2548 931 2732
rect 941 2668 947 2692
rect 1021 2688 1027 2832
rect 1005 2668 1011 2672
rect 941 2568 947 2612
rect 1069 2588 1075 2832
rect 1133 2788 1139 2832
rect 1085 2648 1091 2692
rect 1133 2688 1139 2692
rect 1117 2568 1123 2632
rect 1165 2628 1171 2692
rect 1181 2688 1187 2712
rect 1245 2708 1251 2832
rect 1293 2768 1299 2832
rect 1341 2788 1347 2952
rect 1373 2948 1379 2952
rect 1469 2948 1475 2952
rect 1453 2928 1459 2932
rect 1533 2908 1539 3052
rect 1581 2948 1587 3032
rect 1645 2988 1651 2992
rect 1613 2963 1619 2972
rect 1608 2957 1619 2963
rect 1645 2944 1651 2972
rect 1661 2948 1667 3012
rect 1677 3008 1683 3092
rect 1741 3088 1747 3092
rect 1949 3088 1955 3092
rect 1965 3088 1971 3212
rect 1997 3208 2003 3412
rect 2077 3368 2083 3432
rect 2141 3368 2147 3432
rect 2189 3368 2195 3372
rect 2061 3348 2067 3352
rect 2173 3348 2179 3352
rect 2221 3348 2227 3432
rect 2013 3208 2019 3312
rect 2221 3308 2227 3312
rect 2125 3288 2131 3292
rect 2237 3283 2243 3432
rect 2285 3328 2291 3412
rect 2301 3388 2307 3492
rect 2365 3488 2371 3492
rect 2333 3344 2339 3372
rect 2397 3363 2403 3432
rect 2397 3357 2408 3363
rect 2461 3348 2467 3432
rect 2477 3368 2483 3537
rect 2541 3508 2547 3572
rect 2557 3548 2563 3712
rect 2573 3568 2579 3632
rect 2605 3543 2611 3712
rect 2653 3708 2659 3712
rect 2701 3708 2707 3712
rect 2605 3537 2627 3543
rect 2541 3488 2547 3492
rect 2525 3468 2531 3472
rect 2573 3428 2579 3532
rect 2589 3488 2595 3492
rect 2541 3368 2547 3392
rect 2573 3343 2579 3412
rect 2605 3388 2611 3472
rect 2557 3337 2579 3343
rect 2397 3288 2403 3332
rect 2557 3328 2563 3337
rect 2573 3308 2579 3312
rect 2221 3277 2243 3283
rect 1997 3108 2003 3192
rect 2029 3128 2035 3232
rect 1805 3068 1811 3076
rect 1709 3057 1720 3063
rect 1709 3048 1715 3057
rect 1677 2968 1683 2972
rect 1725 2948 1731 2992
rect 1341 2768 1347 2772
rect 1357 2708 1363 2752
rect 1373 2728 1379 2792
rect 1373 2708 1379 2712
rect 1437 2708 1443 2832
rect 1533 2768 1539 2892
rect 1533 2703 1539 2752
rect 1549 2748 1555 2832
rect 1565 2708 1571 2832
rect 1581 2708 1587 2892
rect 1533 2697 1544 2703
rect 1197 2668 1203 2692
rect 989 2508 995 2552
rect 1133 2548 1139 2552
rect 1229 2548 1235 2552
rect 1245 2548 1251 2672
rect 1053 2528 1059 2532
rect 1085 2488 1091 2512
rect 829 2088 835 2232
rect 845 2228 851 2232
rect 845 2188 851 2192
rect 877 2148 883 2252
rect 941 2148 947 2352
rect 973 2288 979 2392
rect 989 2208 995 2252
rect 1021 2148 1027 2452
rect 1117 2328 1123 2532
rect 1261 2528 1267 2532
rect 1165 2388 1171 2432
rect 1277 2388 1283 2692
rect 1309 2588 1315 2632
rect 1293 2563 1299 2572
rect 1293 2557 1304 2563
rect 1325 2548 1331 2632
rect 1357 2368 1363 2432
rect 1085 2288 1091 2312
rect 1181 2303 1187 2312
rect 1176 2297 1187 2303
rect 1197 2283 1203 2312
rect 1192 2277 1203 2283
rect 1213 2297 1224 2303
rect 1037 2228 1043 2232
rect 1069 2168 1075 2252
rect 1101 2148 1107 2232
rect 1117 2168 1123 2232
rect 589 2028 595 2032
rect 509 2017 531 2023
rect 365 1728 371 1732
rect 349 1688 355 1712
rect 381 1708 387 1772
rect 429 1763 435 1832
rect 461 1788 467 1912
rect 477 1908 483 1912
rect 525 1908 531 2017
rect 717 1928 723 1932
rect 509 1888 515 1892
rect 429 1757 456 1763
rect 397 1748 403 1752
rect 477 1748 483 1792
rect 541 1768 547 1892
rect 605 1888 611 1892
rect 701 1868 707 1892
rect 717 1888 723 1912
rect 765 1908 771 1912
rect 749 1888 755 1892
rect 637 1848 643 1852
rect 557 1837 568 1843
rect 525 1748 531 1752
rect 413 1728 419 1732
rect 541 1708 547 1712
rect 429 1528 435 1532
rect 45 1488 51 1492
rect 141 1388 147 1492
rect 157 1488 163 1492
rect 461 1488 467 1652
rect 509 1548 515 1632
rect 541 1528 547 1552
rect 269 1348 275 1472
rect 13 1328 19 1332
rect 61 1323 67 1332
rect 56 1317 67 1323
rect 365 1328 371 1472
rect 413 1388 419 1452
rect 13 1128 19 1132
rect 93 1108 99 1132
rect 56 1097 67 1103
rect 61 1088 67 1097
rect 152 1097 163 1103
rect 157 1088 163 1097
rect 365 1088 371 1312
rect 429 1168 435 1314
rect 13 928 19 932
rect 109 923 115 932
rect 141 928 147 972
rect 365 948 371 1072
rect 157 928 163 932
rect 104 917 115 923
rect 461 908 467 1472
rect 493 1368 499 1432
rect 557 1408 563 1837
rect 573 1788 579 1812
rect 621 1728 627 1732
rect 605 1708 611 1712
rect 637 1668 643 1692
rect 717 1688 723 1872
rect 733 1768 739 1832
rect 749 1723 755 1872
rect 765 1748 771 1872
rect 813 1828 819 1912
rect 829 1908 835 2012
rect 909 1948 915 2032
rect 1005 1988 1011 2032
rect 845 1908 851 1912
rect 973 1908 979 1912
rect 877 1788 883 1832
rect 1005 1808 1011 1952
rect 1021 1908 1027 1992
rect 1069 1903 1075 2032
rect 1101 1908 1107 2112
rect 1133 2108 1139 2232
rect 1197 2168 1203 2192
rect 1213 2188 1219 2297
rect 1277 2168 1283 2212
rect 1293 2148 1299 2332
rect 1309 2288 1315 2332
rect 1357 2283 1363 2352
rect 1389 2328 1395 2632
rect 1405 2548 1411 2632
rect 1421 2548 1427 2612
rect 1453 2608 1459 2692
rect 1597 2688 1603 2892
rect 1709 2768 1715 2912
rect 1629 2648 1635 2652
rect 1517 2568 1523 2632
rect 1613 2588 1619 2632
rect 1645 2588 1651 2692
rect 1469 2528 1475 2532
rect 1501 2508 1507 2552
rect 1533 2543 1539 2552
rect 1581 2548 1587 2572
rect 1629 2568 1635 2572
rect 1528 2537 1539 2543
rect 1661 2528 1667 2632
rect 1352 2277 1363 2283
rect 1309 2208 1315 2252
rect 1341 2188 1347 2252
rect 1384 2237 1395 2243
rect 1133 1908 1139 1932
rect 1053 1897 1075 1903
rect 1053 1888 1059 1897
rect 1229 1888 1235 1912
rect 1005 1788 1011 1792
rect 1085 1748 1091 1872
rect 1117 1828 1123 1872
rect 744 1717 755 1723
rect 749 1668 755 1692
rect 573 1488 579 1652
rect 621 1628 627 1632
rect 605 1548 611 1612
rect 509 1348 515 1392
rect 605 1308 611 1532
rect 621 1508 627 1592
rect 669 1588 675 1632
rect 765 1568 771 1732
rect 781 1728 787 1732
rect 877 1708 883 1712
rect 813 1688 819 1692
rect 893 1568 899 1732
rect 909 1728 915 1732
rect 941 1688 947 1692
rect 621 1428 627 1492
rect 637 1408 643 1512
rect 749 1508 755 1512
rect 717 1488 723 1492
rect 781 1468 787 1472
rect 701 1348 707 1352
rect 525 788 531 1152
rect 557 1106 563 1212
rect 605 1168 611 1232
rect 637 1108 643 1272
rect 701 1237 712 1243
rect 589 948 595 1072
rect 621 968 627 1072
rect 653 948 659 1232
rect 701 1068 707 1237
rect 733 1108 739 1412
rect 749 1348 755 1432
rect 765 1368 771 1412
rect 829 1348 835 1472
rect 845 1408 851 1492
rect 909 1488 915 1492
rect 973 1488 979 1632
rect 1037 1628 1043 1712
rect 1085 1608 1091 1732
rect 1053 1528 1059 1532
rect 1101 1508 1107 1752
rect 1117 1588 1123 1712
rect 1165 1648 1171 1832
rect 1181 1768 1187 1832
rect 1245 1783 1251 2112
rect 1261 2108 1267 2112
rect 1277 1908 1283 1932
rect 1293 1908 1299 2072
rect 1309 1908 1315 2152
rect 1373 2144 1379 2152
rect 1389 2148 1395 2237
rect 1405 2168 1411 2192
rect 1437 2148 1443 2432
rect 1501 2368 1507 2492
rect 1469 2288 1475 2352
rect 1533 2348 1539 2432
rect 1613 2428 1619 2432
rect 1661 2348 1667 2512
rect 1533 2288 1539 2332
rect 1453 2228 1459 2252
rect 1517 2228 1523 2252
rect 1469 2168 1475 2212
rect 1533 2168 1539 2212
rect 1517 2148 1523 2152
rect 1549 2148 1555 2272
rect 1581 2128 1587 2292
rect 1661 2288 1667 2332
rect 1677 2288 1683 2452
rect 1693 2348 1699 2432
rect 1709 2408 1715 2632
rect 1725 2628 1731 2852
rect 1757 2688 1763 3032
rect 1853 2968 1859 3032
rect 1869 2988 1875 3072
rect 2029 3068 2035 3092
rect 1869 2968 1875 2972
rect 1853 2948 1859 2952
rect 1885 2948 1891 3012
rect 1773 2928 1779 2932
rect 1917 2928 1923 3032
rect 1933 2948 1939 2972
rect 1981 2928 1987 3052
rect 2061 3008 2067 3032
rect 2077 2983 2083 3032
rect 2061 2977 2083 2983
rect 2061 2948 2067 2977
rect 2093 2963 2099 3252
rect 2109 3088 2115 3092
rect 2125 3088 2131 3112
rect 2141 3023 2147 3032
rect 2088 2957 2099 2963
rect 2125 3017 2147 3023
rect 2125 2948 2131 3017
rect 2205 3008 2211 3032
rect 2141 2968 2147 2992
rect 2221 2988 2227 3277
rect 2365 3268 2371 3272
rect 2253 3108 2259 3112
rect 2333 3068 2339 3092
rect 2365 3088 2371 3252
rect 2429 3188 2435 3232
rect 2381 3088 2387 3092
rect 2429 3088 2435 3112
rect 2456 3057 2467 3063
rect 2461 3048 2467 3057
rect 2269 2983 2275 3032
rect 2253 2977 2275 2983
rect 2253 2948 2259 2977
rect 2349 2983 2355 3032
rect 2397 3028 2403 3032
rect 2333 2977 2355 2983
rect 2285 2968 2291 2972
rect 2189 2928 2195 2932
rect 2269 2928 2275 2952
rect 2317 2928 2323 2952
rect 2333 2928 2339 2977
rect 2365 2948 2371 3012
rect 2477 2968 2483 3172
rect 2493 3148 2499 3232
rect 2509 3228 2515 3232
rect 2509 3108 2515 3212
rect 2589 3108 2595 3332
rect 2621 3328 2627 3537
rect 2653 3508 2659 3552
rect 2701 3508 2707 3672
rect 2685 3348 2691 3392
rect 2701 3368 2707 3392
rect 2717 3328 2723 3672
rect 2733 3548 2739 3712
rect 2749 3708 2755 3712
rect 2749 3588 2755 3592
rect 2781 3508 2787 3552
rect 2733 3408 2739 3432
rect 2749 3348 2755 3492
rect 2781 3363 2787 3372
rect 2776 3357 2787 3363
rect 2813 3344 2819 3432
rect 2829 3428 2835 3712
rect 2845 3688 2851 3712
rect 2893 3688 2899 3712
rect 2845 3508 2851 3592
rect 2861 3588 2867 3632
rect 2877 3508 2883 3532
rect 2893 3508 2899 3572
rect 2957 3488 2963 3632
rect 2973 3488 2979 3492
rect 2829 3348 2835 3352
rect 2621 3308 2627 3312
rect 2717 3188 2723 3232
rect 2477 2948 2483 2952
rect 2493 2948 2499 2952
rect 1821 2908 1827 2912
rect 1768 2657 1779 2663
rect 1773 2648 1779 2657
rect 1725 2548 1731 2612
rect 1741 2548 1747 2552
rect 1789 2548 1795 2832
rect 1805 2768 1811 2892
rect 1805 2708 1811 2752
rect 1821 2708 1827 2812
rect 1869 2688 1875 2892
rect 1917 2828 1923 2832
rect 2029 2808 2035 2832
rect 2029 2708 2035 2752
rect 1917 2688 1923 2692
rect 2077 2688 2083 2712
rect 2093 2708 2099 2832
rect 2157 2808 2163 2832
rect 2125 2668 2131 2752
rect 2189 2708 2195 2792
rect 2141 2688 2147 2692
rect 2189 2677 2200 2683
rect 1837 2583 1843 2632
rect 1821 2577 1843 2583
rect 1757 2448 1763 2452
rect 1757 2343 1763 2432
rect 1757 2337 1779 2343
rect 1704 2257 1715 2263
rect 1645 2148 1651 2232
rect 1709 2168 1715 2257
rect 1725 2188 1731 2292
rect 1773 2288 1779 2337
rect 1773 2168 1779 2252
rect 1597 2128 1603 2132
rect 1709 2128 1715 2152
rect 1821 2148 1827 2577
rect 1885 2568 1891 2652
rect 1901 2648 1907 2652
rect 2061 2648 2067 2652
rect 2109 2628 2115 2632
rect 2125 2568 2131 2632
rect 2173 2628 2179 2632
rect 1837 2528 1843 2552
rect 2189 2548 2195 2677
rect 2221 2688 2227 2832
rect 2253 2668 2259 2812
rect 2285 2708 2291 2772
rect 2317 2768 2323 2912
rect 2397 2828 2403 2832
rect 2349 2708 2355 2812
rect 2477 2788 2483 2912
rect 2237 2568 2243 2632
rect 1885 2148 1891 2312
rect 1917 2188 1923 2472
rect 1933 2328 1939 2432
rect 2045 2388 2051 2532
rect 2269 2528 2275 2632
rect 2301 2563 2307 2632
rect 2365 2588 2371 2692
rect 2477 2668 2483 2772
rect 2525 2688 2531 2992
rect 2557 2968 2563 3092
rect 2573 2948 2579 3032
rect 2637 2963 2643 3032
rect 2653 2988 2659 3032
rect 2685 2968 2691 3092
rect 2749 3088 2755 3232
rect 2845 3208 2851 3312
rect 2845 3148 2851 3192
rect 2861 3088 2867 3272
rect 2909 3148 2915 3212
rect 2941 3088 2947 3412
rect 2973 3408 2979 3432
rect 2989 3368 2995 3452
rect 3021 3348 3027 3632
rect 3037 3508 3043 3812
rect 3085 3748 3091 3792
rect 3117 3763 3123 3772
rect 3112 3757 3123 3763
rect 3133 3663 3139 4063
rect 3197 3948 3203 4063
rect 3309 4028 3315 4063
rect 3405 3968 3411 4063
rect 3149 3808 3155 3832
rect 3165 3763 3171 3892
rect 3181 3828 3187 3892
rect 3245 3888 3251 3932
rect 3272 3857 3283 3863
rect 3277 3848 3283 3857
rect 3213 3808 3219 3832
rect 3149 3757 3171 3763
rect 3149 3728 3155 3757
rect 3176 3737 3224 3743
rect 3133 3657 3155 3663
rect 3069 3508 3075 3612
rect 3085 3508 3091 3512
rect 3037 3448 3043 3492
rect 3149 3368 3155 3657
rect 3165 3488 3171 3672
rect 3213 3568 3219 3712
rect 3229 3508 3235 3552
rect 3181 3468 3187 3492
rect 3037 3328 3043 3332
rect 3149 3328 3155 3352
rect 3165 3348 3171 3432
rect 3197 3428 3203 3432
rect 3277 3383 3283 3592
rect 3293 3528 3299 3892
rect 3325 3868 3331 3872
rect 3373 3828 3379 3876
rect 3309 3728 3315 3732
rect 3325 3728 3331 3752
rect 3293 3508 3299 3512
rect 3309 3488 3315 3692
rect 3341 3503 3347 3812
rect 3405 3728 3411 3952
rect 3485 3908 3491 4063
rect 3533 3908 3539 4063
rect 3581 4028 3587 4063
rect 3613 4008 3619 4063
rect 3581 3908 3587 3992
rect 3421 3748 3427 3752
rect 3421 3728 3427 3732
rect 3357 3648 3363 3712
rect 3357 3588 3363 3632
rect 3341 3497 3352 3503
rect 3325 3488 3331 3492
rect 3261 3377 3283 3383
rect 3213 3368 3219 3372
rect 3261 3348 3267 3377
rect 3341 3368 3347 3497
rect 3373 3488 3379 3572
rect 3373 3383 3379 3472
rect 3357 3377 3379 3383
rect 3357 3348 3363 3377
rect 3373 3348 3379 3352
rect 3021 3188 3027 3212
rect 2989 3108 2995 3152
rect 2701 3068 2707 3072
rect 2749 3068 2755 3072
rect 2717 3008 2723 3032
rect 2765 2968 2771 3052
rect 2781 2988 2787 3052
rect 2637 2957 2648 2963
rect 2797 2943 2803 3012
rect 2792 2937 2803 2943
rect 2717 2928 2723 2932
rect 2669 2908 2675 2912
rect 2557 2748 2563 2832
rect 2685 2768 2691 2912
rect 2749 2788 2755 2792
rect 2557 2708 2563 2732
rect 2573 2708 2579 2752
rect 2781 2708 2787 2832
rect 2653 2697 2680 2703
rect 2541 2668 2547 2692
rect 2653 2683 2659 2697
rect 2648 2677 2659 2683
rect 2605 2657 2616 2663
rect 2605 2648 2611 2657
rect 2285 2557 2307 2563
rect 2013 2303 2019 2312
rect 2013 2297 2024 2303
rect 1933 2248 1939 2276
rect 1901 2128 1907 2152
rect 1325 2028 1331 2032
rect 1389 1908 1395 2012
rect 1357 1888 1363 1892
rect 1325 1788 1331 1876
rect 1453 1883 1459 2032
rect 1485 1903 1491 1912
rect 1549 1908 1555 2072
rect 1565 1908 1571 2052
rect 1629 2048 1635 2112
rect 1581 2028 1587 2032
rect 1480 1897 1491 1903
rect 1453 1877 1480 1883
rect 1373 1863 1379 1872
rect 1357 1857 1379 1863
rect 1357 1788 1363 1857
rect 1421 1848 1427 1852
rect 1373 1788 1379 1812
rect 1240 1777 1251 1783
rect 1533 1768 1539 1876
rect 1549 1768 1555 1772
rect 1597 1748 1603 1832
rect 1613 1808 1619 1832
rect 1661 1743 1667 1892
rect 1656 1737 1667 1743
rect 1197 1708 1203 1712
rect 1229 1548 1235 1592
rect 1245 1588 1251 1732
rect 1165 1528 1171 1532
rect 1133 1488 1139 1512
rect 877 1457 888 1463
rect 877 1448 883 1457
rect 1021 1428 1027 1432
rect 1037 1428 1043 1452
rect 1101 1428 1107 1452
rect 797 1328 803 1332
rect 781 1228 787 1232
rect 797 1148 803 1292
rect 813 1123 819 1232
rect 861 1128 867 1332
rect 973 1308 979 1332
rect 1053 1328 1059 1372
rect 1117 1363 1123 1432
rect 1197 1388 1203 1472
rect 1117 1357 1128 1363
rect 1069 1348 1075 1352
rect 1229 1348 1235 1432
rect 1144 1337 1155 1343
rect 1149 1328 1155 1337
rect 1245 1343 1251 1492
rect 1261 1408 1267 1512
rect 1277 1488 1283 1552
rect 1293 1528 1299 1692
rect 1309 1608 1315 1712
rect 1421 1708 1427 1712
rect 1325 1528 1331 1672
rect 1293 1488 1299 1492
rect 1245 1337 1267 1343
rect 1197 1328 1203 1332
rect 1229 1328 1235 1332
rect 1053 1303 1059 1312
rect 1053 1297 1064 1303
rect 973 1168 979 1292
rect 925 1128 931 1152
rect 797 1117 819 1123
rect 733 1088 739 1092
rect 797 1068 803 1117
rect 669 1028 675 1032
rect 669 968 675 992
rect 13 728 19 732
rect 93 708 99 732
rect 653 728 659 932
rect 669 928 675 952
rect 701 868 707 1052
rect 733 944 739 1012
rect 797 944 803 1052
rect 813 1028 819 1032
rect 717 908 723 932
rect 845 928 851 1052
rect 861 1028 867 1072
rect 56 697 67 703
rect 61 688 67 697
rect 93 637 104 643
rect 13 528 19 532
rect 61 523 67 532
rect 93 528 99 637
rect 269 548 275 672
rect 317 668 323 712
rect 669 708 675 852
rect 717 703 723 712
rect 717 697 728 703
rect 221 528 227 532
rect 56 517 67 523
rect 269 488 275 532
rect 317 528 323 552
rect 429 508 435 512
rect 93 437 104 443
rect 13 328 19 332
rect 93 308 99 437
rect 221 308 227 432
rect 56 297 67 303
rect 61 288 67 297
rect 269 288 275 472
rect 333 308 339 432
rect 445 288 451 672
rect 573 668 579 692
rect 589 668 595 672
rect 605 588 611 692
rect 813 688 819 832
rect 829 728 835 832
rect 845 708 851 832
rect 717 648 723 672
rect 541 568 547 572
rect 605 548 611 552
rect 621 548 627 552
rect 637 548 643 592
rect 749 548 755 652
rect 493 488 499 532
rect 765 528 771 632
rect 829 588 835 652
rect 845 608 851 632
rect 861 563 867 1012
rect 877 948 883 972
rect 909 948 915 1032
rect 925 948 931 1112
rect 941 1088 947 1092
rect 989 1088 995 1232
rect 1005 1108 1011 1152
rect 1021 1108 1027 1252
rect 1213 1188 1219 1292
rect 1229 1163 1235 1232
rect 1261 1228 1267 1337
rect 1357 1328 1363 1692
rect 1469 1668 1475 1712
rect 1389 1488 1395 1512
rect 1469 1508 1475 1632
rect 1517 1508 1523 1612
rect 1549 1508 1555 1532
rect 1213 1157 1235 1163
rect 1037 1068 1043 1092
rect 989 968 995 1032
rect 1069 983 1075 1092
rect 1085 1088 1091 1112
rect 1133 1088 1139 1092
rect 1213 1088 1219 1157
rect 1293 1148 1299 1232
rect 1261 1128 1267 1132
rect 1325 1108 1331 1132
rect 1341 1088 1347 1272
rect 1357 1108 1363 1312
rect 1373 1308 1379 1392
rect 1437 1388 1443 1472
rect 1485 1408 1491 1432
rect 1453 1348 1459 1352
rect 1389 1288 1395 1312
rect 1405 1148 1411 1312
rect 1469 1288 1475 1332
rect 1533 1308 1539 1492
rect 1565 1448 1571 1492
rect 1597 1488 1603 1572
rect 1629 1528 1635 1692
rect 1661 1563 1667 1712
rect 1677 1588 1683 1732
rect 1693 1728 1699 2112
rect 1757 1968 1763 2112
rect 1917 2088 1923 2152
rect 1709 1948 1715 1952
rect 1725 1948 1731 1952
rect 1736 1897 1747 1903
rect 1661 1557 1683 1563
rect 1661 1508 1667 1532
rect 1613 1488 1619 1492
rect 1549 1328 1555 1332
rect 1565 1308 1571 1392
rect 1629 1388 1635 1432
rect 1645 1328 1651 1392
rect 1677 1388 1683 1557
rect 1741 1508 1747 1897
rect 1773 1868 1779 1876
rect 1757 1648 1763 1732
rect 1773 1728 1779 1732
rect 1757 1568 1763 1632
rect 1789 1588 1795 2032
rect 1837 1988 1843 2052
rect 1869 1988 1875 1992
rect 1821 1888 1827 1932
rect 1805 1763 1811 1832
rect 1805 1757 1827 1763
rect 1805 1608 1811 1692
rect 1821 1588 1827 1757
rect 1837 1708 1843 1912
rect 1853 1788 1859 1912
rect 1901 1908 1907 1932
rect 1997 1888 2003 2032
rect 2013 1928 2019 2112
rect 2029 2108 2035 2112
rect 2045 2108 2051 2372
rect 2077 2288 2083 2312
rect 2157 2288 2163 2392
rect 2109 2183 2115 2272
rect 2125 2208 2131 2232
rect 2109 2177 2120 2183
rect 2141 2168 2147 2172
rect 2077 2117 2088 2123
rect 2077 2108 2083 2117
rect 2045 1968 2051 2092
rect 1917 1868 1923 1872
rect 2013 1868 2019 1912
rect 1885 1788 1891 1852
rect 2061 1828 2067 1872
rect 2013 1748 2019 1792
rect 2077 1788 2083 1852
rect 2029 1768 2035 1772
rect 2077 1768 2083 1772
rect 2093 1768 2099 1952
rect 1837 1688 1843 1692
rect 1709 1388 1715 1492
rect 1741 1488 1747 1492
rect 1853 1488 1859 1712
rect 1880 1697 1891 1703
rect 1869 1588 1875 1672
rect 1885 1548 1891 1697
rect 2045 1688 2051 1752
rect 2109 1748 2115 2152
rect 2173 2088 2179 2492
rect 2285 2448 2291 2557
rect 2317 2523 2323 2552
rect 2333 2528 2339 2572
rect 2413 2548 2419 2552
rect 2301 2517 2323 2523
rect 2253 2368 2259 2432
rect 2269 2423 2275 2432
rect 2269 2417 2291 2423
rect 2221 2288 2227 2332
rect 2285 2308 2291 2417
rect 2205 2148 2211 2212
rect 2269 2168 2275 2252
rect 2253 2128 2259 2132
rect 2141 1908 2147 2012
rect 2157 1868 2163 2072
rect 2221 2068 2227 2112
rect 2173 1888 2179 2032
rect 2189 2028 2195 2032
rect 2173 1768 2179 1772
rect 2157 1737 2168 1743
rect 2045 1528 2051 1632
rect 2077 1568 2083 1732
rect 2157 1728 2163 1737
rect 1725 1468 1731 1472
rect 1821 1468 1827 1472
rect 1773 1448 1779 1452
rect 1901 1448 1907 1492
rect 1933 1443 1939 1476
rect 1917 1437 1939 1443
rect 1725 1388 1731 1412
rect 1837 1368 1843 1432
rect 1549 1108 1555 1252
rect 1565 1088 1571 1172
rect 1661 1108 1667 1112
rect 1677 1083 1683 1332
rect 1693 1328 1699 1352
rect 1672 1077 1683 1083
rect 1165 1048 1171 1052
rect 1101 1008 1107 1032
rect 1064 977 1075 983
rect 1101 948 1107 972
rect 877 688 883 772
rect 1005 768 1011 932
rect 1181 908 1187 1072
rect 1213 948 1219 1052
rect 1229 1028 1235 1072
rect 1501 1068 1507 1072
rect 1405 1048 1411 1052
rect 1213 928 1219 932
rect 1229 908 1235 1012
rect 1277 968 1283 1032
rect 1261 944 1267 952
rect 1309 928 1315 952
rect 893 648 899 652
rect 909 648 915 652
rect 861 557 883 563
rect 877 548 883 557
rect 461 308 467 432
rect 573 348 579 472
rect 797 388 803 432
rect 333 237 344 243
rect 88 157 99 163
rect 13 128 19 132
rect 61 123 67 132
rect 93 128 99 157
rect 109 128 115 232
rect 301 163 307 232
rect 285 157 307 163
rect 56 117 67 123
rect 141 123 147 132
rect 285 128 291 157
rect 301 128 307 132
rect 333 128 339 237
rect 509 188 515 272
rect 605 148 611 272
rect 701 248 707 272
rect 749 268 755 312
rect 813 306 819 512
rect 861 468 867 532
rect 909 508 915 572
rect 957 568 963 752
rect 1053 688 1059 812
rect 1069 688 1075 892
rect 1117 888 1123 892
rect 1149 888 1155 892
rect 1005 628 1011 652
rect 1085 588 1091 872
rect 1133 828 1139 832
rect 1101 728 1107 732
rect 1181 688 1187 812
rect 1197 748 1203 832
rect 1261 708 1267 852
rect 1261 688 1267 692
rect 1277 688 1283 892
rect 1293 888 1299 892
rect 1309 868 1315 912
rect 1309 828 1315 832
rect 1325 748 1331 872
rect 1357 688 1363 812
rect 1373 748 1379 932
rect 1421 783 1427 912
rect 1416 777 1427 783
rect 1421 728 1427 732
rect 1437 708 1443 712
rect 1197 568 1203 632
rect 1293 568 1299 632
rect 1357 588 1363 672
rect 1453 668 1459 1032
rect 1469 988 1475 1012
rect 1501 668 1507 1052
rect 1581 988 1587 992
rect 1565 948 1571 972
rect 1549 748 1555 912
rect 1453 568 1459 652
rect 1565 628 1571 672
rect 1517 568 1523 612
rect 1565 588 1571 612
rect 957 508 963 552
rect 1277 548 1283 552
rect 1517 548 1523 552
rect 973 528 979 532
rect 1021 528 1027 532
rect 1133 528 1139 532
rect 1053 448 1059 472
rect 1053 288 1059 312
rect 1069 308 1075 372
rect 141 117 152 123
rect 397 123 403 132
rect 392 117 403 123
rect 637 128 643 232
rect 749 188 755 232
rect 813 188 819 252
rect 845 188 851 272
rect 877 168 883 192
rect 669 123 675 132
rect 1005 128 1011 232
rect 669 117 680 123
rect 1069 123 1075 132
rect 1064 117 1075 123
rect 781 108 787 112
rect 845 108 851 112
rect 189 -43 195 32
rect 205 28 211 32
rect 237 -43 243 12
rect 253 -37 259 32
rect 253 -43 275 -37
rect 349 -43 355 32
rect 717 -43 723 32
rect 893 -43 899 32
rect 1021 28 1027 32
rect 989 -43 995 12
rect 1149 -37 1155 532
rect 1229 508 1235 512
rect 1245 508 1251 532
rect 1325 528 1331 532
rect 1325 488 1331 512
rect 1197 303 1203 432
rect 1309 408 1315 432
rect 1389 428 1395 432
rect 1197 297 1208 303
rect 1181 288 1187 292
rect 1229 288 1235 332
rect 1309 328 1315 392
rect 1437 388 1443 492
rect 1501 468 1507 532
rect 1549 508 1555 552
rect 1581 528 1587 532
rect 1597 488 1603 492
rect 1533 308 1539 412
rect 1277 148 1283 172
rect 1309 128 1315 232
rect 1405 148 1411 272
rect 1533 208 1539 292
rect 1549 268 1555 272
rect 1581 268 1587 352
rect 1597 288 1603 292
rect 1341 123 1347 132
rect 1565 128 1571 232
rect 1341 117 1352 123
rect 1485 108 1491 112
rect 1133 -43 1155 -37
rect 1181 -43 1187 12
rect 1229 -43 1235 12
rect 1389 -43 1395 32
rect 1613 -43 1619 912
rect 1629 868 1635 1070
rect 1693 1048 1699 1076
rect 1645 948 1651 952
rect 1677 928 1683 932
rect 1709 908 1715 1332
rect 1773 1328 1779 1332
rect 1757 1268 1763 1312
rect 1885 1303 1891 1332
rect 1869 1297 1891 1303
rect 1757 1068 1763 1092
rect 1725 988 1731 1032
rect 1773 968 1779 972
rect 1789 948 1795 1032
rect 1821 1028 1827 1092
rect 1853 1008 1859 1092
rect 1869 1088 1875 1297
rect 1901 1288 1907 1312
rect 1917 1108 1923 1437
rect 1997 1388 2003 1512
rect 2013 1388 2019 1492
rect 1949 1308 1955 1332
rect 2029 1328 2035 1432
rect 2045 1348 2051 1372
rect 2061 1168 2067 1492
rect 2093 1348 2099 1572
rect 2109 1508 2115 1692
rect 2125 1628 2131 1712
rect 2125 1488 2131 1512
rect 2189 1508 2195 1992
rect 2221 1908 2227 1972
rect 2301 1928 2307 2517
rect 2365 2428 2371 2432
rect 2349 2308 2355 2392
rect 2429 2283 2435 2632
rect 2477 2548 2483 2592
rect 2621 2528 2627 2612
rect 2669 2548 2675 2632
rect 2669 2528 2675 2532
rect 2509 2348 2515 2432
rect 2525 2308 2531 2512
rect 2589 2468 2595 2492
rect 2605 2348 2611 2492
rect 2685 2488 2691 2612
rect 2669 2308 2675 2432
rect 2717 2388 2723 2432
rect 2781 2408 2787 2432
rect 2717 2308 2723 2352
rect 2813 2323 2819 3032
rect 2861 3008 2867 3052
rect 2925 3048 2931 3052
rect 2861 2963 2867 2972
rect 2856 2957 2867 2963
rect 2893 2944 2899 2952
rect 2909 2948 2915 3012
rect 2941 3008 2947 3072
rect 3021 2968 3027 3032
rect 2925 2948 2931 2952
rect 3021 2788 3027 2832
rect 2829 2568 2835 2752
rect 2893 2708 2899 2712
rect 2797 2317 2819 2323
rect 2733 2308 2739 2312
rect 2424 2277 2435 2283
rect 2237 1768 2243 1852
rect 2237 1688 2243 1752
rect 2285 1588 2291 1752
rect 2317 1748 2323 2232
rect 2381 2188 2387 2212
rect 2360 2117 2371 2123
rect 2349 1988 2355 2012
rect 2349 1908 2355 1972
rect 2365 1883 2371 2117
rect 2461 2088 2467 2092
rect 2413 1988 2419 2072
rect 2445 2028 2451 2032
rect 2429 1888 2435 1932
rect 2445 1908 2451 1952
rect 2461 1888 2467 1892
rect 2349 1877 2371 1883
rect 2349 1788 2355 1877
rect 2413 1768 2419 1832
rect 2429 1788 2435 1872
rect 2461 1788 2467 1852
rect 2477 1748 2483 2292
rect 2525 2168 2531 2252
rect 2541 2188 2547 2272
rect 2605 2183 2611 2292
rect 2637 2188 2643 2272
rect 2653 2228 2659 2272
rect 2701 2188 2707 2232
rect 2605 2177 2627 2183
rect 2605 2148 2611 2152
rect 2509 2108 2515 2132
rect 2541 1908 2547 2132
rect 2557 2128 2563 2132
rect 2621 2128 2627 2177
rect 2749 2168 2755 2252
rect 2765 2188 2771 2232
rect 2573 2028 2579 2032
rect 2621 1968 2627 2112
rect 2637 2088 2643 2092
rect 2669 1988 2675 2072
rect 2696 2037 2707 2043
rect 2509 1888 2515 1892
rect 2685 1888 2691 1912
rect 2701 1908 2707 2037
rect 2765 1928 2771 2152
rect 2797 2128 2803 2317
rect 2829 2308 2835 2312
rect 2877 2288 2883 2352
rect 2829 2063 2835 2152
rect 2861 2148 2867 2272
rect 2893 2268 2899 2552
rect 2909 2548 2915 2772
rect 3021 2708 3027 2712
rect 2925 2668 2931 2692
rect 2973 2608 2979 2676
rect 2909 2288 2915 2532
rect 2925 2528 2931 2592
rect 2941 2288 2947 2332
rect 2957 2268 2963 2592
rect 3021 2548 3027 2632
rect 3037 2628 3043 3312
rect 3165 3248 3171 3332
rect 3101 3108 3107 3232
rect 3181 3228 3187 3312
rect 3053 3088 3059 3092
rect 3133 3068 3139 3192
rect 3181 3148 3187 3172
rect 3181 3108 3187 3132
rect 3053 2948 3059 3032
rect 3085 2963 3091 2972
rect 3080 2957 3091 2963
rect 3117 2928 3123 2952
rect 3133 2948 3139 3052
rect 3053 2548 3059 2772
rect 3133 2768 3139 2872
rect 3085 2728 3091 2732
rect 3085 2688 3091 2712
rect 3149 2688 3155 3032
rect 3197 2948 3203 3232
rect 3213 3108 3219 3112
rect 3229 3048 3235 3232
rect 3245 3108 3251 3112
rect 3277 3028 3283 3332
rect 3389 3208 3395 3432
rect 3405 3208 3411 3712
rect 3469 3628 3475 3632
rect 3485 3603 3491 3892
rect 3501 3728 3507 3892
rect 3533 3828 3539 3892
rect 3549 3888 3555 3892
rect 3549 3748 3555 3872
rect 3533 3708 3539 3712
rect 3597 3688 3603 3712
rect 3597 3648 3603 3652
rect 3469 3597 3491 3603
rect 3469 3468 3475 3597
rect 3565 3548 3571 3612
rect 3485 3508 3491 3512
rect 3597 3488 3603 3632
rect 3597 3468 3603 3472
rect 3448 3457 3459 3463
rect 3421 3328 3427 3452
rect 3453 3448 3459 3457
rect 3533 3428 3539 3432
rect 3565 3428 3571 3432
rect 3437 3328 3443 3412
rect 3485 3368 3491 3412
rect 3453 3328 3459 3332
rect 3421 3183 3427 3312
rect 3453 3228 3459 3252
rect 3421 3177 3443 3183
rect 3421 3088 3427 3112
rect 3437 3088 3443 3177
rect 3453 3108 3459 3112
rect 3485 3108 3491 3152
rect 3501 3108 3507 3272
rect 3213 2968 3219 2972
rect 3293 2943 3299 3032
rect 3309 2963 3315 3032
rect 3309 2957 3320 2963
rect 3373 2963 3379 3032
rect 3373 2957 3384 2963
rect 3293 2937 3304 2943
rect 3181 2808 3187 2912
rect 3197 2748 3203 2912
rect 3165 2708 3171 2712
rect 3245 2708 3251 2912
rect 3373 2888 3379 2932
rect 3405 2928 3411 2932
rect 3261 2728 3267 2872
rect 3341 2748 3347 2832
rect 3261 2688 3267 2712
rect 3245 2668 3251 2672
rect 3101 2568 3107 2632
rect 3197 2628 3203 2632
rect 3117 2548 3123 2552
rect 3053 2428 3059 2432
rect 3069 2308 3075 2432
rect 3133 2428 3139 2492
rect 3149 2468 3155 2512
rect 3165 2488 3171 2532
rect 3117 2288 3123 2292
rect 2877 2168 2883 2232
rect 2909 2228 2915 2232
rect 2925 2228 2931 2252
rect 2957 2248 2963 2252
rect 3133 2248 3139 2272
rect 2893 2188 2899 2192
rect 2813 2057 2835 2063
rect 2493 1788 2499 1832
rect 2557 1808 2563 1872
rect 2621 1788 2627 1832
rect 2637 1748 2643 1792
rect 2157 1328 2163 1432
rect 2173 1428 2179 1476
rect 2221 1468 2227 1492
rect 2237 1388 2243 1412
rect 2221 1328 2227 1372
rect 2285 1368 2291 1572
rect 2317 1528 2323 1712
rect 2397 1588 2403 1732
rect 2605 1728 2611 1732
rect 2653 1728 2659 1792
rect 2669 1728 2675 1732
rect 2589 1708 2595 1712
rect 2685 1708 2691 1712
rect 2445 1608 2451 1632
rect 2525 1628 2531 1652
rect 2557 1648 2563 1692
rect 2365 1528 2371 1552
rect 2413 1528 2419 1532
rect 2445 1528 2451 1592
rect 2509 1588 2515 1612
rect 2493 1528 2499 1552
rect 2525 1548 2531 1612
rect 2557 1588 2563 1592
rect 2573 1548 2579 1552
rect 2333 1488 2339 1492
rect 2301 1428 2307 1472
rect 2381 1468 2387 1512
rect 2397 1508 2403 1512
rect 2589 1508 2595 1672
rect 2621 1648 2627 1692
rect 2717 1608 2723 1892
rect 2797 1888 2803 1932
rect 2813 1868 2819 2057
rect 2829 2008 2835 2032
rect 2829 1888 2835 1892
rect 2845 1888 2851 1932
rect 2845 1868 2851 1872
rect 2877 1868 2883 2132
rect 2925 2128 2931 2172
rect 2989 2148 2995 2232
rect 3085 2168 3091 2172
rect 3053 2128 3059 2152
rect 3101 2148 3107 2172
rect 2893 2088 2899 2092
rect 2941 1888 2947 1892
rect 2893 1877 2904 1883
rect 2893 1848 2899 1877
rect 2909 1848 2915 1852
rect 2749 1748 2755 1832
rect 2797 1788 2803 1832
rect 2861 1763 2867 1832
rect 2973 1788 2979 1792
rect 2845 1757 2867 1763
rect 2845 1728 2851 1757
rect 2909 1744 2915 1772
rect 2669 1528 2675 1572
rect 2733 1528 2739 1632
rect 2765 1588 2771 1712
rect 2813 1648 2819 1692
rect 2317 1408 2323 1452
rect 2349 1428 2355 1432
rect 2397 1408 2403 1492
rect 2509 1488 2515 1492
rect 2429 1388 2435 1392
rect 2333 1328 2339 1332
rect 2397 1328 2403 1332
rect 2429 1328 2435 1372
rect 2013 1108 2019 1152
rect 1837 968 1843 972
rect 1837 948 1843 952
rect 1917 948 1923 952
rect 1661 888 1667 892
rect 1853 888 1859 932
rect 1933 928 1939 972
rect 1629 688 1635 832
rect 1709 708 1715 792
rect 1741 728 1747 832
rect 1645 628 1651 632
rect 1677 548 1683 572
rect 1725 568 1731 652
rect 1773 543 1779 852
rect 1821 808 1827 832
rect 1885 728 1891 812
rect 1821 688 1827 712
rect 1869 708 1875 712
rect 1949 688 1955 892
rect 1853 668 1859 672
rect 1949 668 1955 672
rect 1901 628 1907 652
rect 1917 637 1928 643
rect 1917 568 1923 637
rect 1773 537 1795 543
rect 1645 308 1651 392
rect 1661 388 1667 532
rect 1709 508 1715 532
rect 1677 388 1683 392
rect 1741 348 1747 492
rect 1757 468 1763 532
rect 1773 508 1779 512
rect 1789 508 1795 537
rect 1805 508 1811 512
rect 1885 508 1891 532
rect 1821 468 1827 472
rect 1853 468 1859 472
rect 1709 308 1715 312
rect 1629 248 1635 292
rect 1741 288 1747 332
rect 1757 308 1763 372
rect 1773 328 1779 392
rect 1725 123 1731 132
rect 1725 117 1736 123
rect 1693 -43 1699 32
rect 1757 28 1763 292
rect 1789 268 1795 372
rect 1864 317 1875 323
rect 1869 308 1875 317
rect 1837 128 1843 132
rect 1741 -43 1747 12
rect 1773 -43 1779 32
rect 1821 -43 1827 12
rect 1853 -43 1859 272
rect 1885 268 1891 492
rect 1901 388 1907 532
rect 1949 348 1955 452
rect 1981 408 1987 892
rect 2029 708 2035 1152
rect 2125 1143 2131 1232
rect 2125 1137 2147 1143
rect 2125 1128 2131 1137
rect 2141 1128 2147 1137
rect 2173 1128 2179 1152
rect 2189 1143 2195 1232
rect 2269 1188 2275 1312
rect 2189 1137 2211 1143
rect 2141 1048 2147 1072
rect 2045 988 2051 1012
rect 2173 988 2179 1032
rect 2189 1008 2195 1092
rect 2205 1088 2211 1137
rect 2285 1108 2291 1272
rect 2429 1188 2435 1292
rect 2461 1248 2467 1312
rect 2477 1308 2483 1472
rect 2621 1468 2627 1472
rect 2525 1368 2531 1372
rect 2605 1344 2611 1352
rect 2317 1128 2323 1172
rect 2365 1128 2371 1132
rect 2237 1048 2243 1072
rect 2301 1028 2307 1092
rect 2237 988 2243 992
rect 2381 988 2387 1092
rect 2429 1028 2435 1092
rect 2445 1068 2451 1132
rect 2461 1128 2467 1232
rect 2509 1168 2515 1332
rect 2509 1088 2515 1092
rect 2525 1068 2531 1332
rect 2621 1303 2627 1452
rect 2669 1428 2675 1512
rect 2733 1448 2739 1492
rect 2813 1488 2819 1632
rect 2845 1508 2851 1612
rect 2861 1608 2867 1732
rect 2941 1728 2947 1752
rect 2893 1548 2899 1552
rect 2925 1508 2931 1712
rect 2957 1648 2963 1732
rect 3005 1728 3011 1912
rect 3021 1768 3027 1792
rect 3037 1788 3043 2032
rect 3069 1948 3075 2012
rect 3069 1868 3075 1932
rect 3133 1928 3139 2112
rect 3149 2108 3155 2132
rect 3165 2128 3171 2412
rect 3181 2297 3192 2303
rect 3181 2263 3187 2297
rect 3181 2257 3203 2263
rect 3197 2188 3203 2257
rect 3213 2168 3219 2652
rect 3277 2628 3283 2692
rect 3389 2683 3395 2892
rect 3384 2677 3395 2683
rect 3277 2608 3283 2612
rect 3277 2388 3283 2592
rect 3309 2583 3315 2632
rect 3293 2577 3315 2583
rect 3293 2548 3299 2577
rect 3325 2563 3331 2592
rect 3320 2557 3331 2563
rect 3389 2528 3395 2532
rect 3405 2528 3411 2912
rect 3453 2768 3459 3092
rect 3469 2928 3475 2932
rect 3485 2928 3491 3072
rect 3501 2968 3507 3092
rect 3517 3008 3523 3312
rect 3565 3108 3571 3192
rect 3597 3108 3603 3352
rect 3613 3328 3619 3972
rect 3661 3908 3667 4063
rect 3677 3908 3683 3972
rect 3645 3888 3651 3892
rect 3677 3888 3683 3892
rect 3645 3868 3651 3872
rect 3693 3788 3699 3832
rect 3661 3748 3667 3772
rect 3693 3768 3699 3772
rect 3661 3508 3667 3732
rect 3677 3728 3683 3732
rect 3709 3728 3715 4063
rect 3757 3988 3763 4063
rect 3885 3988 3891 4063
rect 3997 4028 4003 4063
rect 4045 4028 4051 4063
rect 4173 4028 4179 4063
rect 3757 3908 3763 3972
rect 3725 3888 3731 3892
rect 3773 3728 3779 3872
rect 3805 3788 3811 3952
rect 3965 3908 3971 3972
rect 3997 3908 4003 4012
rect 4077 3908 4083 4012
rect 4125 3908 4131 4012
rect 4173 3908 4179 4012
rect 4221 3908 4227 4012
rect 4365 4008 4371 4063
rect 4269 3908 4275 3932
rect 4317 3908 4323 3972
rect 4365 3908 4371 3992
rect 4861 3928 4867 4063
rect 5853 3988 5859 4063
rect 3821 3748 3827 3892
rect 3885 3888 3891 3892
rect 3853 3848 3859 3852
rect 3821 3723 3827 3732
rect 3853 3728 3859 3832
rect 3869 3728 3875 3792
rect 3949 3768 3955 3872
rect 3949 3728 3955 3752
rect 3965 3728 3971 3892
rect 4013 3868 4019 3892
rect 3821 3717 3832 3723
rect 3693 3708 3699 3712
rect 3677 3548 3683 3692
rect 3709 3688 3715 3712
rect 3757 3708 3763 3712
rect 3917 3708 3923 3712
rect 3965 3708 3971 3712
rect 4029 3668 4035 3892
rect 4077 3868 4083 3872
rect 4045 3728 4051 3852
rect 4093 3728 4099 3892
rect 4109 3768 4115 3892
rect 4445 3888 4451 3892
rect 4653 3883 4659 3892
rect 4648 3877 4659 3883
rect 4429 3848 4435 3872
rect 4509 3868 4515 3872
rect 4573 3868 4579 3872
rect 4701 3868 4707 3872
rect 4509 3848 4515 3852
rect 4157 3828 4163 3832
rect 4189 3788 4195 3832
rect 4189 3768 4195 3772
rect 4285 3763 4291 3772
rect 4280 3757 4291 3763
rect 4093 3703 4099 3712
rect 4077 3697 4099 3703
rect 3741 3628 3747 3632
rect 3741 3588 3747 3592
rect 3629 3428 3635 3432
rect 3629 3368 3635 3412
rect 3677 3328 3683 3532
rect 3709 3448 3715 3452
rect 3709 3343 3715 3432
rect 3693 3337 3715 3343
rect 3693 3328 3699 3337
rect 3725 3323 3731 3512
rect 3757 3328 3763 3652
rect 3789 3508 3795 3592
rect 3773 3388 3779 3476
rect 3805 3408 3811 3632
rect 3997 3588 4003 3632
rect 4013 3508 4019 3512
rect 4077 3508 4083 3697
rect 4093 3588 4099 3672
rect 4141 3643 4147 3712
rect 4136 3637 4147 3643
rect 4125 3508 4131 3632
rect 4205 3568 4211 3732
rect 4317 3728 4323 3832
rect 4333 3748 4339 3792
rect 4381 3748 4387 3812
rect 4397 3768 4403 3832
rect 4461 3828 4467 3832
rect 4525 3808 4531 3832
rect 4589 3828 4595 3832
rect 4637 3828 4643 3852
rect 4717 3828 4723 3832
rect 4477 3763 4483 3772
rect 4472 3757 4483 3763
rect 4541 3748 4547 3772
rect 4717 3768 4723 3792
rect 4765 3788 4771 3872
rect 4829 3868 4835 3872
rect 4781 3768 4787 3832
rect 4845 3828 4851 3832
rect 4205 3528 4211 3552
rect 3773 3368 3779 3372
rect 3720 3317 3731 3323
rect 3613 3128 3619 3312
rect 3661 3308 3667 3312
rect 3661 3108 3667 3132
rect 3565 3068 3571 3092
rect 3501 2928 3507 2932
rect 3517 2928 3523 2992
rect 3565 2948 3571 2952
rect 3581 2928 3587 2932
rect 3485 2828 3491 2912
rect 3581 2848 3587 2912
rect 3421 2523 3427 2552
rect 3437 2548 3443 2632
rect 3453 2588 3459 2692
rect 3485 2628 3491 2672
rect 3421 2517 3443 2523
rect 3229 2288 3235 2292
rect 3181 2008 3187 2132
rect 3229 1988 3235 2112
rect 3245 1968 3251 2312
rect 3277 2288 3283 2352
rect 3272 2257 3283 2263
rect 3261 2228 3267 2232
rect 3261 2188 3267 2212
rect 3277 2028 3283 2257
rect 3309 2088 3315 2372
rect 3341 2268 3347 2292
rect 3373 2288 3379 2292
rect 3421 2288 3427 2492
rect 3437 2268 3443 2517
rect 3453 2308 3459 2572
rect 3517 2548 3523 2632
rect 3533 2568 3539 2772
rect 3597 2768 3603 2832
rect 3613 2828 3619 3092
rect 3645 3028 3651 3032
rect 3645 2908 3651 2952
rect 3661 2903 3667 3092
rect 3693 3063 3699 3312
rect 3741 3208 3747 3232
rect 3725 3108 3731 3112
rect 3677 3057 3699 3063
rect 3677 2928 3683 3057
rect 3693 2948 3699 3032
rect 3725 3003 3731 3092
rect 3725 2997 3747 3003
rect 3725 2963 3731 2972
rect 3720 2957 3731 2963
rect 3661 2897 3683 2903
rect 3645 2808 3651 2892
rect 3565 2708 3571 2732
rect 3565 2688 3571 2692
rect 3581 2688 3587 2692
rect 3549 2488 3555 2672
rect 3597 2568 3603 2752
rect 3629 2628 3635 2652
rect 3581 2548 3587 2552
rect 3597 2548 3603 2552
rect 3560 2437 3571 2443
rect 3469 2308 3475 2432
rect 3437 2248 3443 2252
rect 3485 2228 3491 2432
rect 3565 2348 3571 2437
rect 3565 2308 3571 2332
rect 3597 2308 3603 2472
rect 3501 2228 3507 2232
rect 3341 2008 3347 2092
rect 3293 1988 3299 1992
rect 3197 1928 3203 1952
rect 3213 1908 3219 1932
rect 3261 1908 3267 1972
rect 3309 1908 3315 1972
rect 3165 1863 3171 1892
rect 3229 1868 3235 1872
rect 3149 1857 3171 1863
rect 3085 1808 3091 1832
rect 3149 1788 3155 1857
rect 3053 1728 3059 1752
rect 3117 1728 3123 1732
rect 3005 1708 3011 1712
rect 2797 1457 2808 1463
rect 2637 1388 2643 1412
rect 2733 1388 2739 1432
rect 2781 1388 2787 1432
rect 2797 1388 2803 1457
rect 2605 1297 2627 1303
rect 2557 1148 2563 1272
rect 1997 588 2003 612
rect 2061 568 2067 792
rect 2077 748 2083 912
rect 2093 897 2104 903
rect 2093 788 2099 897
rect 2093 708 2099 712
rect 2109 548 2115 632
rect 2141 608 2147 912
rect 2173 728 2179 892
rect 2189 788 2195 912
rect 2205 728 2211 812
rect 2285 748 2291 932
rect 2349 688 2355 752
rect 2397 708 2403 952
rect 2429 868 2435 912
rect 2477 888 2483 932
rect 2493 928 2499 952
rect 2413 788 2419 792
rect 2445 708 2451 712
rect 2397 688 2403 692
rect 2253 668 2259 672
rect 2285 668 2291 672
rect 2205 568 2211 652
rect 2253 628 2259 652
rect 2029 388 2035 512
rect 2045 388 2051 512
rect 2077 428 2083 432
rect 1949 288 1955 332
rect 1901 128 1907 172
rect 1885 -37 1891 32
rect 1885 -43 1907 -37
rect 1933 -43 1939 12
rect 1981 -43 1987 32
rect 2029 -37 2035 332
rect 2045 308 2051 332
rect 2061 328 2067 392
rect 2125 306 2131 412
rect 2045 268 2051 292
rect 2125 223 2131 252
rect 2141 228 2147 432
rect 2109 217 2131 223
rect 2077 148 2083 172
rect 2109 148 2115 217
rect 2125 208 2131 217
rect 2141 148 2147 212
rect 2157 168 2163 432
rect 2221 408 2227 492
rect 2253 448 2259 472
rect 2269 268 2275 632
rect 2333 528 2339 532
rect 2429 528 2435 592
rect 2461 528 2467 532
rect 2317 448 2323 512
rect 2349 508 2355 512
rect 2397 508 2403 512
rect 2477 508 2483 812
rect 2493 528 2499 912
rect 2509 908 2515 1012
rect 2525 1008 2531 1052
rect 2509 688 2515 692
rect 2525 668 2531 712
rect 2541 688 2547 692
rect 2557 563 2563 1132
rect 2573 1108 2579 1152
rect 2589 1128 2595 1292
rect 2573 1028 2579 1092
rect 2573 948 2579 992
rect 2573 728 2579 932
rect 2589 748 2595 1112
rect 2605 1108 2611 1297
rect 2621 1108 2627 1172
rect 2637 948 2643 1192
rect 2669 1148 2675 1372
rect 2813 1368 2819 1412
rect 2701 1348 2707 1352
rect 2685 1188 2691 1312
rect 2717 1288 2723 1332
rect 2749 1308 2755 1332
rect 2765 1308 2771 1312
rect 2669 1128 2675 1132
rect 2781 1108 2787 1192
rect 2653 948 2659 1032
rect 2701 988 2707 1092
rect 2733 948 2739 1032
rect 2797 1003 2803 1032
rect 2781 997 2803 1003
rect 2749 937 2760 943
rect 2621 928 2627 932
rect 2669 923 2675 932
rect 2664 917 2675 923
rect 2605 748 2611 872
rect 2589 588 2595 592
rect 2552 557 2563 563
rect 2509 488 2515 492
rect 2333 288 2339 292
rect 2157 128 2163 152
rect 2237 128 2243 212
rect 2253 128 2259 232
rect 2349 168 2355 232
rect 2397 228 2403 232
rect 2397 148 2403 192
rect 2285 123 2291 132
rect 2445 128 2451 132
rect 2285 117 2296 123
rect 2541 68 2547 552
rect 2605 508 2611 732
rect 2621 668 2627 912
rect 2637 688 2643 912
rect 2685 828 2691 832
rect 2733 808 2739 912
rect 2749 768 2755 937
rect 2765 788 2771 912
rect 2781 903 2787 997
rect 2813 988 2819 1252
rect 2829 1108 2835 1212
rect 2845 1188 2851 1492
rect 2877 1488 2883 1492
rect 2893 1388 2899 1392
rect 2941 1388 2947 1592
rect 3069 1588 3075 1672
rect 2957 1528 2963 1532
rect 3133 1508 3139 1532
rect 3181 1528 3187 1832
rect 3229 1768 3235 1852
rect 3277 1848 3283 1852
rect 3213 1748 3219 1752
rect 3197 1588 3203 1732
rect 3277 1708 3283 1732
rect 3293 1708 3299 1712
rect 3229 1528 3235 1592
rect 3277 1528 3283 1612
rect 3325 1528 3331 1992
rect 3373 1948 3379 2112
rect 3341 1768 3347 1832
rect 3341 1548 3347 1632
rect 3048 1497 3096 1503
rect 3133 1488 3139 1492
rect 3261 1488 3267 1512
rect 3373 1508 3379 1792
rect 3389 1748 3395 2052
rect 3405 1888 3411 2072
rect 3437 1888 3443 2212
rect 3453 2088 3459 2132
rect 3469 2028 3475 2152
rect 3485 2128 3491 2132
rect 3501 2128 3507 2192
rect 3581 2128 3587 2232
rect 3613 2208 3619 2552
rect 3629 2548 3635 2572
rect 3661 2508 3667 2832
rect 3677 2768 3683 2897
rect 3741 2708 3747 2997
rect 3757 2988 3763 3072
rect 3773 2948 3779 3132
rect 3757 2908 3763 2912
rect 3789 2908 3795 3212
rect 3821 2988 3827 3492
rect 3853 3363 3859 3432
rect 3848 3357 3859 3363
rect 3848 3337 3859 3343
rect 3853 3328 3859 3337
rect 3869 3328 3875 3432
rect 3901 3368 3907 3492
rect 3917 3488 3923 3492
rect 3933 3428 3939 3492
rect 4141 3488 4147 3492
rect 4221 3483 4227 3632
rect 4333 3548 4339 3732
rect 4381 3508 4387 3512
rect 4397 3508 4403 3732
rect 4509 3528 4515 3712
rect 4525 3708 4531 3732
rect 4525 3568 4531 3692
rect 4493 3508 4499 3512
rect 4557 3508 4563 3512
rect 4573 3508 4579 3712
rect 4589 3668 4595 3732
rect 4717 3728 4723 3752
rect 4797 3743 4803 3812
rect 4829 3748 4835 3752
rect 4845 3748 4851 3752
rect 4792 3737 4803 3743
rect 4861 3723 4867 3912
rect 4957 3908 4963 3912
rect 5005 3908 5011 3912
rect 4893 3828 4899 3872
rect 4973 3808 4979 3892
rect 4845 3717 4867 3723
rect 4589 3628 4595 3652
rect 4653 3648 4659 3712
rect 4685 3648 4691 3692
rect 4621 3528 4627 3632
rect 4205 3477 4227 3483
rect 3997 3468 4003 3472
rect 3885 3328 3891 3352
rect 3869 3108 3875 3172
rect 3901 3148 3907 3272
rect 3917 3108 3923 3172
rect 3837 3088 3843 3092
rect 3757 2708 3763 2892
rect 3773 2748 3779 2852
rect 3805 2848 3811 2912
rect 3837 2863 3843 3032
rect 3853 2948 3859 2992
rect 3901 2928 3907 2932
rect 3821 2857 3843 2863
rect 3821 2708 3827 2857
rect 3837 2828 3843 2832
rect 3837 2708 3843 2812
rect 3869 2708 3875 2912
rect 3917 2708 3923 2832
rect 3933 2768 3939 3412
rect 4056 3377 4072 3383
rect 3949 3348 3955 3372
rect 4109 3368 4115 3412
rect 4109 3344 4115 3352
rect 4157 3343 4163 3432
rect 4189 3428 4195 3476
rect 4205 3448 4211 3477
rect 4413 3488 4419 3492
rect 4637 3488 4643 3512
rect 4685 3508 4691 3632
rect 4221 3368 4227 3432
rect 4253 3408 4259 3476
rect 4344 3457 4355 3463
rect 4349 3448 4355 3457
rect 4269 3363 4275 3372
rect 4264 3357 4275 3363
rect 4237 3348 4243 3352
rect 4157 3337 4168 3343
rect 4061 3328 4067 3332
rect 4125 3328 4131 3332
rect 4301 3328 4307 3392
rect 4365 3328 4371 3412
rect 4397 3388 4403 3472
rect 4477 3468 4483 3472
rect 4525 3363 4531 3432
rect 4520 3357 4531 3363
rect 4520 3337 4531 3343
rect 4445 3328 4451 3332
rect 4525 3328 4531 3337
rect 4045 3308 4051 3312
rect 3981 3108 3987 3172
rect 4029 2988 4035 3292
rect 4189 3268 4195 3292
rect 4301 3268 4307 3312
rect 4317 3308 4323 3312
rect 4429 3303 4435 3312
rect 4429 3297 4451 3303
rect 4445 3268 4451 3297
rect 4541 3288 4547 3472
rect 4664 3457 4675 3463
rect 4669 3448 4675 3457
rect 4573 3348 4579 3372
rect 4589 3368 4595 3432
rect 4557 3283 4563 3312
rect 4557 3277 4579 3283
rect 4029 2708 4035 2872
rect 4045 2848 4051 3076
rect 4061 2928 4067 3152
rect 4125 3108 4131 3112
rect 4141 3108 4147 3112
rect 4189 3108 4195 3252
rect 4205 3148 4211 3232
rect 4205 3088 4211 3092
rect 4253 3088 4259 3092
rect 4077 2948 4083 3032
rect 4093 2968 4099 3032
rect 4157 2968 4163 3032
rect 4173 3008 4179 3072
rect 4317 3068 4323 3092
rect 4381 3088 4387 3212
rect 4397 3108 4403 3232
rect 4445 3108 4451 3252
rect 4280 3057 4291 3063
rect 4285 3048 4291 3057
rect 4408 3057 4419 3063
rect 4136 2937 4147 2943
rect 4141 2928 4147 2937
rect 4173 2928 4179 2992
rect 4189 2948 4195 3012
rect 4317 3008 4323 3052
rect 4413 3048 4419 3057
rect 4445 3008 4451 3092
rect 4477 2968 4483 3232
rect 4525 3068 4531 3152
rect 4541 3148 4547 3272
rect 4541 3088 4547 3092
rect 4557 3028 4563 3192
rect 4573 3108 4579 3277
rect 4621 3108 4627 3412
rect 4648 3337 4659 3343
rect 4653 3328 4659 3337
rect 4685 3328 4691 3492
rect 4701 3408 4707 3492
rect 4717 3488 4723 3672
rect 4845 3648 4851 3717
rect 4893 3708 4899 3712
rect 4733 3568 4739 3632
rect 4797 3608 4803 3632
rect 4813 3508 4819 3512
rect 4845 3508 4851 3632
rect 4781 3468 4787 3472
rect 4813 3428 4819 3492
rect 4909 3488 4915 3732
rect 4925 3728 4931 3792
rect 4989 3728 4995 3752
rect 5005 3543 5011 3892
rect 5053 3768 5059 3952
rect 5069 3908 5075 3912
rect 5805 3897 5816 3903
rect 5101 3848 5107 3892
rect 5053 3688 5059 3752
rect 5005 3537 5027 3543
rect 5021 3508 5027 3537
rect 4984 3457 4995 3463
rect 4989 3448 4995 3457
rect 4925 3428 4931 3432
rect 4781 3363 4787 3372
rect 4776 3357 4787 3363
rect 4701 3348 4707 3352
rect 4749 3348 4755 3352
rect 4701 3168 4707 3332
rect 4813 3328 4819 3392
rect 4845 3368 4851 3372
rect 5021 3348 5027 3492
rect 5053 3488 5059 3492
rect 5069 3488 5075 3772
rect 5101 3663 5107 3832
rect 5149 3748 5155 3872
rect 5181 3848 5187 3872
rect 5165 3768 5171 3772
rect 5197 3743 5203 3832
rect 5229 3788 5235 3876
rect 5293 3868 5299 3892
rect 5405 3888 5411 3892
rect 5437 3888 5443 3892
rect 5309 3868 5315 3872
rect 5373 3868 5379 3872
rect 5261 3768 5267 3832
rect 5325 3768 5331 3832
rect 5197 3737 5208 3743
rect 5304 3737 5315 3743
rect 5309 3728 5315 3737
rect 5341 3668 5347 3712
rect 5085 3657 5107 3663
rect 5085 3408 5091 3657
rect 5117 3623 5123 3632
rect 5101 3617 5123 3623
rect 4717 3208 4723 3232
rect 4637 3108 4643 3132
rect 4765 3108 4771 3112
rect 4781 3108 4787 3252
rect 4813 3108 4819 3312
rect 4893 3303 4899 3332
rect 4877 3297 4899 3303
rect 4829 3088 4835 3112
rect 4205 2948 4211 2952
rect 4317 2948 4323 2952
rect 4477 2948 4483 2952
rect 4269 2928 4275 2932
rect 4493 2928 4499 2992
rect 4509 2928 4515 2992
rect 4557 2928 4563 3012
rect 4061 2788 4067 2912
rect 4045 2708 4051 2752
rect 4061 2708 4067 2752
rect 4077 2748 4083 2832
rect 4093 2788 4099 2892
rect 4301 2848 4307 2912
rect 4109 2708 4115 2712
rect 4189 2708 4195 2772
rect 3677 2628 3683 2672
rect 3693 2648 3699 2652
rect 3741 2648 3747 2692
rect 3805 2688 3811 2692
rect 3885 2668 3891 2692
rect 3677 2528 3683 2612
rect 3709 2608 3715 2632
rect 3741 2548 3747 2552
rect 3757 2528 3763 2532
rect 3709 2488 3715 2512
rect 3773 2508 3779 2632
rect 3869 2608 3875 2632
rect 3869 2563 3875 2572
rect 3864 2557 3875 2563
rect 3917 2548 3923 2572
rect 3789 2528 3795 2532
rect 3901 2488 3907 2512
rect 3709 2428 3715 2432
rect 3677 2288 3683 2332
rect 3725 2308 3731 2312
rect 3629 2248 3635 2252
rect 3597 2148 3603 2172
rect 3613 2168 3619 2192
rect 3629 2128 3635 2132
rect 3421 1868 3427 1872
rect 3421 1808 3427 1852
rect 3405 1648 3411 1752
rect 3437 1743 3443 1752
rect 3453 1743 3459 1892
rect 3469 1788 3475 2012
rect 3533 1928 3539 2032
rect 3512 1917 3523 1923
rect 3517 1908 3523 1917
rect 3581 1848 3587 2112
rect 3645 2048 3651 2232
rect 3677 2128 3683 2232
rect 3672 2037 3683 2043
rect 3613 1908 3619 1972
rect 3629 1928 3635 1992
rect 3661 1948 3667 1952
rect 3677 1948 3683 2037
rect 3597 1868 3603 1892
rect 3437 1737 3459 1743
rect 3389 1628 3395 1632
rect 3421 1628 3427 1632
rect 3389 1528 3395 1612
rect 3453 1528 3459 1737
rect 3501 1608 3507 1632
rect 3533 1528 3539 1832
rect 3549 1768 3555 1832
rect 3565 1828 3571 1832
rect 3565 1803 3571 1812
rect 3565 1797 3587 1803
rect 3565 1768 3571 1772
rect 3581 1748 3587 1797
rect 3549 1728 3555 1732
rect 3661 1688 3667 1932
rect 3693 1908 3699 2232
rect 3709 2128 3715 2292
rect 3741 2148 3747 2312
rect 3757 2168 3763 2192
rect 3757 1908 3763 2152
rect 3789 2128 3795 2392
rect 3805 2328 3811 2432
rect 3789 2048 3795 2112
rect 3805 2028 3811 2252
rect 3821 2068 3827 2272
rect 3837 2108 3843 2472
rect 3933 2308 3939 2652
rect 3981 2648 3987 2692
rect 3949 2528 3955 2552
rect 3997 2528 4003 2572
rect 3949 2508 3955 2512
rect 3981 2328 3987 2432
rect 4029 2308 4035 2632
rect 3853 2128 3859 2132
rect 3885 2128 3891 2252
rect 3917 2088 3923 2232
rect 3933 2128 3939 2272
rect 3965 2248 3971 2252
rect 3949 2128 3955 2192
rect 3917 2028 3923 2032
rect 3789 1908 3795 1912
rect 3693 1768 3699 1792
rect 3725 1708 3731 1732
rect 3741 1668 3747 1832
rect 3757 1688 3763 1832
rect 3821 1768 3827 1772
rect 3837 1648 3843 1712
rect 3741 1637 3752 1643
rect 3629 1628 3635 1632
rect 3037 1468 3043 1472
rect 3101 1468 3107 1472
rect 3325 1468 3331 1472
rect 3053 1448 3059 1452
rect 3053 1428 3059 1432
rect 3069 1383 3075 1432
rect 3053 1377 3075 1383
rect 3053 1368 3059 1377
rect 2877 1308 2883 1332
rect 2861 1208 2867 1232
rect 2845 1128 2851 1172
rect 2829 1088 2835 1092
rect 2877 1068 2883 1092
rect 2893 1088 2899 1112
rect 2909 928 2915 932
rect 2781 897 2792 903
rect 2845 848 2851 912
rect 2861 788 2867 912
rect 2925 908 2931 1252
rect 2941 1128 2947 1232
rect 2957 1108 2963 1292
rect 3053 1128 3059 1132
rect 2941 1008 2947 1092
rect 2989 1088 2995 1112
rect 3069 1108 3075 1112
rect 3021 988 3027 1092
rect 3053 1028 3059 1032
rect 3085 968 3091 1392
rect 3101 1188 3107 1412
rect 3117 1368 3123 1372
rect 3128 1337 3139 1343
rect 3133 1328 3139 1337
rect 3197 1328 3203 1452
rect 3213 1437 3224 1443
rect 3213 1348 3219 1437
rect 3245 1368 3251 1412
rect 3165 1188 3171 1192
rect 3149 1148 3155 1172
rect 3181 1128 3187 1212
rect 3181 1083 3187 1112
rect 3165 1077 3187 1083
rect 3165 968 3171 1077
rect 2941 948 2947 952
rect 3085 948 3091 952
rect 3181 948 3187 1052
rect 3197 988 3203 1092
rect 3213 1088 3219 1192
rect 3245 1088 3251 1352
rect 3341 1348 3347 1432
rect 3389 1428 3395 1472
rect 3437 1468 3443 1472
rect 3373 1328 3379 1372
rect 3421 1348 3427 1452
rect 3437 1437 3448 1443
rect 3437 1328 3443 1437
rect 3485 1388 3491 1492
rect 3501 1488 3507 1492
rect 3581 1488 3587 1572
rect 3661 1508 3667 1612
rect 3613 1488 3619 1492
rect 3677 1488 3683 1512
rect 3533 1468 3539 1472
rect 3581 1468 3587 1472
rect 3517 1448 3523 1452
rect 3277 1108 3283 1272
rect 3325 1128 3331 1312
rect 3437 1088 3443 1292
rect 3453 1268 3459 1312
rect 3469 1128 3475 1332
rect 3485 1248 3491 1352
rect 3501 1308 3507 1352
rect 3533 1348 3539 1352
rect 3549 1328 3555 1432
rect 3565 1348 3571 1432
rect 3613 1308 3619 1312
rect 3245 1068 3251 1072
rect 3261 1043 3267 1072
rect 3325 1068 3331 1072
rect 3373 1068 3379 1072
rect 3261 1037 3283 1043
rect 3277 968 3283 1037
rect 3309 988 3315 1032
rect 3325 963 3331 1032
rect 3320 957 3331 963
rect 2685 688 2691 752
rect 2733 708 2739 712
rect 2861 648 2867 732
rect 2637 637 2648 643
rect 2621 568 2627 572
rect 2621 528 2627 532
rect 2637 528 2643 637
rect 2685 568 2691 612
rect 2765 608 2771 632
rect 2717 548 2723 592
rect 2813 568 2819 572
rect 2877 548 2883 812
rect 2893 788 2899 792
rect 2925 728 2931 892
rect 3069 888 3075 932
rect 3181 868 3187 932
rect 3053 788 3059 832
rect 2925 648 2931 672
rect 2973 668 2979 692
rect 3085 688 3091 732
rect 3117 708 3123 772
rect 3197 728 3203 952
rect 3261 948 3267 952
rect 3341 948 3347 972
rect 3229 928 3235 932
rect 3117 688 3123 692
rect 2824 537 2835 543
rect 2829 528 2835 537
rect 2925 508 2931 632
rect 2957 528 2963 532
rect 2973 528 2979 652
rect 3197 588 3203 712
rect 3037 508 3043 572
rect 3053 508 3059 552
rect 3133 548 3139 552
rect 3133 528 3139 532
rect 3213 528 3219 692
rect 3261 688 3267 852
rect 3261 548 3267 672
rect 3277 648 3283 672
rect 3325 668 3331 852
rect 3357 788 3363 892
rect 3373 868 3379 1052
rect 3389 968 3395 1032
rect 3405 948 3411 952
rect 3437 948 3443 1072
rect 3485 1068 3491 1232
rect 3533 1088 3539 1232
rect 3581 1128 3587 1192
rect 3597 1108 3603 1232
rect 3629 1108 3635 1432
rect 3645 1108 3651 1312
rect 3661 1108 3667 1432
rect 3693 1368 3699 1552
rect 3725 1508 3731 1512
rect 3741 1508 3747 1637
rect 3789 1488 3795 1512
rect 3805 1468 3811 1632
rect 3837 1528 3843 1632
rect 3837 1488 3843 1492
rect 3693 1348 3699 1352
rect 3773 1328 3779 1332
rect 3853 1328 3859 1752
rect 3869 1748 3875 1832
rect 3917 1568 3923 1872
rect 3933 1868 3939 1872
rect 3933 1744 3939 1832
rect 3965 1788 3971 2232
rect 4045 2128 4051 2692
rect 4061 2563 4067 2692
rect 4109 2608 4115 2692
rect 4061 2557 4083 2563
rect 4061 2428 4067 2432
rect 4061 2308 4067 2332
rect 4061 2128 4067 2272
rect 4077 2228 4083 2557
rect 4237 2548 4243 2632
rect 4120 2537 4131 2543
rect 4125 2528 4131 2537
rect 4157 2488 4163 2512
rect 4189 2488 4195 2512
rect 4093 2308 4099 2412
rect 4109 2308 4115 2312
rect 4157 2308 4163 2312
rect 4093 2128 4099 2132
rect 4109 2128 4115 2172
rect 4029 1808 4035 2032
rect 4045 1988 4051 2092
rect 4125 2068 4131 2232
rect 4157 2128 4163 2212
rect 4141 1928 4147 2032
rect 4173 1968 4179 2292
rect 4189 2268 4195 2332
rect 4221 2328 4227 2432
rect 4253 2328 4259 2832
rect 4269 2568 4275 2632
rect 4301 2548 4307 2692
rect 4317 2688 4323 2852
rect 4349 2748 4355 2912
rect 4365 2708 4371 2812
rect 4317 2588 4323 2672
rect 4397 2668 4403 2912
rect 4205 2288 4211 2292
rect 4061 1848 4067 1872
rect 3965 1728 3971 1752
rect 3997 1728 4003 1772
rect 4029 1768 4035 1772
rect 4061 1648 4067 1832
rect 3917 1508 3923 1512
rect 3933 1488 3939 1592
rect 4077 1588 4083 1872
rect 4136 1837 4147 1843
rect 4093 1768 4099 1772
rect 4093 1728 4099 1752
rect 4125 1748 4131 1812
rect 4141 1788 4147 1837
rect 4205 1788 4211 1992
rect 4221 1888 4227 2232
rect 4237 2228 4243 2232
rect 4253 2143 4259 2312
rect 4269 2308 4275 2512
rect 4301 2408 4307 2432
rect 4248 2137 4259 2143
rect 4269 2088 4275 2232
rect 4285 2168 4291 2272
rect 4317 2128 4323 2192
rect 4285 2108 4291 2112
rect 4285 2008 4291 2092
rect 4253 1928 4259 1992
rect 4237 1868 4243 1872
rect 4141 1548 4147 1712
rect 4189 1648 4195 1732
rect 4237 1728 4243 1792
rect 4317 1768 4323 1972
rect 4333 1788 4339 2632
rect 4365 2548 4371 2592
rect 4397 2563 4403 2632
rect 4392 2557 4403 2563
rect 4397 2428 4403 2432
rect 4349 2308 4355 2392
rect 4413 2343 4419 2912
rect 4589 2908 4595 3072
rect 4653 2963 4659 2972
rect 4701 2968 4707 2992
rect 4717 2988 4723 3072
rect 4856 3057 4867 3063
rect 4861 3048 4867 3057
rect 4648 2957 4659 2963
rect 4621 2948 4627 2952
rect 4701 2948 4707 2952
rect 4429 2748 4435 2832
rect 4525 2808 4531 2832
rect 4429 2708 4435 2712
rect 4397 2337 4419 2343
rect 4365 2308 4371 2312
rect 4397 2148 4403 2337
rect 4429 2323 4435 2692
rect 4445 2688 4451 2772
rect 4493 2708 4499 2732
rect 4509 2688 4515 2752
rect 4541 2708 4547 2732
rect 4589 2688 4595 2752
rect 4605 2708 4611 2712
rect 4461 2608 4467 2632
rect 4445 2568 4451 2572
rect 4509 2548 4515 2552
rect 4456 2537 4467 2543
rect 4461 2528 4467 2537
rect 4493 2488 4499 2512
rect 4525 2488 4531 2672
rect 4637 2648 4643 2652
rect 4573 2583 4579 2632
rect 4557 2577 4579 2583
rect 4557 2548 4563 2577
rect 4589 2563 4595 2572
rect 4584 2557 4595 2563
rect 4637 2548 4643 2612
rect 4653 2568 4659 2632
rect 4653 2548 4659 2552
rect 4669 2548 4675 2912
rect 4717 2683 4723 2692
rect 4712 2677 4723 2683
rect 4733 2543 4739 3032
rect 4749 2928 4755 3012
rect 4797 2968 4803 3032
rect 4877 2988 4883 3297
rect 4909 3188 4915 3332
rect 4957 3328 4963 3332
rect 5069 3308 5075 3332
rect 4989 3188 4995 3212
rect 4845 2963 4851 2972
rect 4909 2968 4915 2972
rect 4840 2957 4851 2963
rect 4813 2948 4819 2952
rect 4941 2928 4947 3092
rect 4957 3068 4963 3092
rect 4973 3048 4979 3072
rect 4973 3008 4979 3032
rect 4893 2908 4899 2912
rect 4749 2708 4755 2732
rect 4845 2708 4851 2872
rect 4861 2688 4867 2692
rect 4765 2628 4771 2672
rect 4829 2668 4835 2672
rect 4893 2608 4899 2632
rect 4909 2628 4915 2632
rect 4829 2568 4835 2572
rect 4765 2548 4771 2552
rect 4733 2537 4744 2543
rect 4493 2328 4499 2472
rect 4429 2317 4440 2323
rect 4413 2308 4419 2312
rect 4445 2288 4451 2292
rect 4525 2288 4531 2432
rect 4557 2328 4563 2352
rect 4557 2308 4563 2312
rect 4605 2308 4611 2532
rect 4397 2128 4403 2132
rect 4413 2123 4419 2272
rect 4429 2188 4435 2232
rect 4509 2188 4515 2232
rect 4525 2148 4531 2232
rect 4557 2148 4563 2212
rect 4573 2168 4579 2172
rect 4477 2128 4483 2132
rect 4413 2117 4424 2123
rect 4365 1908 4371 1972
rect 4461 1908 4467 2032
rect 4477 1908 4483 1952
rect 4493 1908 4499 2012
rect 4509 2008 4515 2032
rect 4605 1968 4611 2232
rect 4621 2088 4627 2512
rect 4637 2448 4643 2532
rect 4797 2528 4803 2532
rect 4877 2508 4883 2532
rect 4701 2328 4707 2432
rect 4717 2428 4723 2432
rect 4845 2428 4851 2432
rect 4909 2408 4915 2432
rect 4717 2283 4723 2292
rect 4712 2277 4723 2283
rect 4637 2248 4643 2252
rect 4653 2208 4659 2232
rect 4701 2148 4707 2152
rect 4733 2148 4739 2332
rect 4749 2308 4755 2352
rect 4797 2288 4803 2292
rect 4829 2283 4835 2312
rect 4925 2303 4931 2912
rect 4941 2628 4947 2912
rect 4973 2908 4979 2912
rect 4957 2688 4963 2692
rect 4968 2657 4979 2663
rect 4973 2648 4979 2657
rect 4989 2628 4995 2932
rect 5005 2708 5011 3272
rect 5021 3028 5027 3092
rect 5037 2928 5043 2932
rect 5053 2908 5059 2912
rect 5069 2788 5075 3292
rect 5101 3268 5107 3617
rect 5133 3508 5139 3632
rect 5197 3568 5203 3652
rect 5117 3488 5123 3492
rect 5197 3488 5203 3552
rect 5245 3528 5251 3632
rect 5245 3488 5251 3492
rect 5149 3368 5155 3432
rect 5181 3408 5187 3476
rect 5261 3468 5267 3572
rect 5325 3488 5331 3512
rect 5357 3468 5363 3492
rect 5197 3437 5208 3443
rect 5117 3328 5123 3332
rect 5197 3288 5203 3437
rect 5213 3328 5219 3332
rect 5261 3328 5267 3452
rect 5277 3368 5283 3432
rect 5341 3368 5347 3372
rect 5309 3328 5315 3332
rect 5373 3328 5379 3852
rect 5389 3788 5395 3872
rect 5512 3857 5523 3863
rect 5517 3848 5523 3857
rect 5437 3768 5443 3772
rect 5453 3708 5459 3832
rect 5549 3828 5555 3876
rect 5805 3888 5811 3897
rect 5565 3868 5571 3872
rect 5549 3783 5555 3812
rect 5533 3777 5555 3783
rect 5517 3748 5523 3772
rect 5469 3728 5475 3732
rect 5389 3508 5395 3632
rect 5469 3508 5475 3712
rect 5501 3488 5507 3672
rect 5533 3528 5539 3777
rect 5581 3743 5587 3832
rect 5645 3788 5651 3832
rect 5661 3788 5667 3872
rect 5677 3868 5683 3876
rect 5741 3868 5747 3876
rect 5677 3848 5683 3852
rect 5709 3768 5715 3832
rect 5741 3768 5747 3772
rect 5757 3748 5763 3872
rect 5805 3763 5811 3772
rect 5805 3757 5816 3763
rect 5837 3748 5843 3752
rect 5917 3748 5923 3832
rect 5581 3737 5592 3743
rect 5549 3508 5555 3512
rect 5389 3348 5395 3432
rect 5229 3228 5235 3232
rect 5261 3108 5267 3272
rect 5325 3188 5331 3212
rect 5149 3083 5155 3092
rect 5213 3088 5219 3092
rect 5144 3077 5155 3083
rect 5144 3057 5155 3063
rect 5149 2988 5155 3057
rect 5197 3008 5203 3072
rect 5245 2968 5251 3092
rect 5288 3057 5299 3063
rect 5293 2988 5299 3057
rect 5165 2908 5171 2932
rect 5181 2928 5187 2932
rect 4973 2568 4979 2592
rect 5005 2568 5011 2692
rect 5053 2648 5059 2672
rect 5053 2548 5059 2632
rect 4989 2528 4995 2532
rect 4925 2297 4936 2303
rect 4829 2277 4851 2283
rect 4829 2248 4835 2252
rect 4733 2128 4739 2132
rect 4605 1908 4611 1952
rect 4653 1908 4659 1952
rect 4701 1908 4707 2052
rect 4717 2008 4723 2032
rect 4509 1888 4515 1892
rect 4349 1783 4355 1876
rect 4541 1868 4547 1892
rect 4429 1848 4435 1852
rect 4349 1777 4360 1783
rect 4445 1763 4451 1832
rect 4477 1768 4483 1852
rect 4557 1768 4563 1832
rect 4573 1768 4579 1832
rect 4440 1757 4451 1763
rect 4285 1728 4291 1732
rect 4173 1543 4179 1632
rect 4157 1537 4179 1543
rect 4013 1468 4019 1472
rect 3869 1388 3875 1432
rect 3885 1428 3891 1432
rect 3901 1348 3907 1392
rect 4029 1388 4035 1472
rect 4093 1468 4099 1532
rect 4141 1488 4147 1492
rect 4157 1468 4163 1537
rect 4173 1508 4179 1512
rect 4189 1488 4195 1632
rect 4045 1348 4051 1372
rect 4205 1368 4211 1452
rect 4221 1428 4227 1712
rect 4237 1548 4243 1552
rect 4253 1508 4259 1532
rect 4269 1528 4275 1572
rect 4317 1568 4323 1752
rect 4440 1737 4451 1743
rect 4333 1688 4339 1732
rect 4445 1728 4451 1737
rect 4477 1728 4483 1752
rect 4621 1748 4627 1752
rect 4568 1737 4579 1743
rect 4573 1728 4579 1737
rect 4653 1728 4659 1752
rect 4349 1528 4355 1552
rect 4301 1508 4307 1512
rect 4381 1488 4387 1532
rect 4477 1528 4483 1712
rect 4605 1568 4611 1712
rect 4493 1488 4499 1532
rect 4605 1508 4611 1552
rect 4621 1508 4627 1512
rect 4669 1508 4675 1672
rect 4685 1668 4691 1832
rect 4701 1788 4707 1892
rect 4733 1888 4739 1932
rect 4749 1908 4755 2192
rect 4797 2028 4803 2032
rect 4813 1988 4819 2232
rect 4829 2148 4835 2172
rect 4845 2168 4851 2277
rect 4909 2283 4915 2292
rect 4904 2277 4915 2283
rect 4904 2257 4915 2263
rect 4909 2188 4915 2257
rect 4925 2208 4931 2297
rect 4829 2088 4835 2112
rect 4829 1908 4835 2072
rect 4861 1948 4867 2132
rect 4941 2128 4947 2212
rect 4973 2108 4979 2232
rect 4989 2128 4995 2472
rect 5021 2103 5027 2272
rect 5053 2128 5059 2132
rect 5037 2108 5043 2112
rect 5053 2108 5059 2112
rect 5005 2097 5027 2103
rect 4781 1783 4787 1832
rect 4765 1777 4787 1783
rect 4701 1768 4707 1772
rect 4765 1748 4771 1777
rect 4797 1763 4803 1832
rect 4813 1768 4819 1792
rect 4792 1757 4803 1763
rect 4701 1728 4707 1732
rect 4813 1728 4819 1752
rect 4829 1728 4835 1892
rect 4845 1888 4851 1912
rect 4893 1908 4899 1992
rect 4861 1728 4867 1812
rect 4925 1748 4931 2052
rect 5005 2048 5011 2097
rect 5069 2088 5075 2112
rect 4941 1768 4947 1972
rect 4984 1877 4995 1883
rect 4989 1848 4995 1877
rect 5005 1828 5011 2032
rect 5085 1908 5091 2892
rect 5277 2828 5283 2832
rect 5309 2828 5315 2952
rect 5325 2928 5331 2932
rect 5325 2908 5331 2912
rect 5341 2848 5347 2912
rect 5197 2708 5203 2792
rect 5341 2708 5347 2812
rect 5101 2668 5107 2672
rect 5117 2648 5123 2652
rect 5165 2528 5171 2692
rect 5213 2688 5219 2692
rect 5213 2588 5219 2672
rect 5293 2648 5299 2692
rect 5309 2668 5315 2672
rect 5245 2608 5251 2632
rect 5261 2563 5267 2632
rect 5293 2583 5299 2632
rect 5288 2577 5299 2583
rect 5256 2557 5267 2563
rect 5229 2548 5235 2552
rect 5181 2528 5187 2532
rect 5165 2328 5171 2512
rect 5197 2428 5203 2432
rect 5229 2308 5235 2312
rect 5245 2308 5251 2532
rect 5309 2508 5315 2512
rect 5325 2463 5331 2672
rect 5357 2668 5363 3232
rect 5421 3208 5427 3232
rect 5421 3108 5427 3152
rect 5373 2948 5379 3032
rect 5389 2928 5395 2992
rect 5421 2968 5427 3012
rect 5437 2988 5443 3470
rect 5453 3428 5459 3432
rect 5485 3363 5491 3372
rect 5480 3357 5491 3363
rect 5517 3348 5523 3432
rect 5533 3348 5539 3412
rect 5565 3408 5571 3632
rect 5629 3528 5635 3712
rect 5661 3488 5667 3632
rect 5693 3488 5699 3732
rect 5885 3608 5891 3712
rect 5917 3628 5923 3632
rect 5837 3508 5843 3512
rect 5869 3508 5875 3512
rect 5677 3468 5683 3476
rect 5565 3348 5571 3372
rect 5629 3348 5635 3432
rect 5645 3368 5651 3432
rect 5693 3428 5699 3472
rect 5725 3468 5731 3492
rect 5757 3343 5763 3432
rect 5773 3363 5779 3432
rect 5773 3357 5784 3363
rect 5805 3348 5811 3492
rect 5837 3388 5843 3472
rect 5757 3337 5768 3343
rect 5517 3308 5523 3312
rect 5517 3103 5523 3292
rect 5512 3097 5523 3103
rect 5453 2988 5459 3032
rect 5469 2948 5475 3032
rect 5373 2808 5379 2832
rect 5469 2828 5475 2832
rect 5485 2828 5491 2832
rect 5437 2708 5443 2812
rect 5501 2708 5507 3092
rect 5533 2983 5539 3032
rect 5549 3028 5555 3232
rect 5565 3108 5571 3332
rect 5597 3328 5603 3332
rect 5693 3328 5699 3332
rect 5869 3328 5875 3472
rect 5581 3308 5587 3312
rect 5725 3308 5731 3312
rect 5805 3308 5811 3312
rect 5661 3208 5667 3232
rect 5725 3228 5731 3292
rect 5613 3108 5619 3132
rect 5613 3028 5619 3092
rect 5517 2977 5539 2983
rect 5517 2948 5523 2977
rect 5549 2963 5555 2972
rect 5544 2957 5555 2963
rect 5581 2944 5587 3012
rect 5613 2968 5619 2972
rect 5645 2943 5651 3032
rect 5640 2937 5651 2943
rect 5677 2928 5683 2932
rect 5693 2928 5699 3172
rect 5741 3108 5747 3212
rect 5789 3068 5795 3072
rect 5389 2608 5395 2632
rect 5357 2548 5363 2592
rect 5389 2563 5395 2572
rect 5384 2557 5395 2563
rect 5421 2544 5427 2572
rect 5453 2568 5459 2632
rect 5453 2528 5459 2532
rect 5469 2528 5475 2612
rect 5309 2457 5331 2463
rect 5309 2388 5315 2457
rect 5325 2428 5331 2432
rect 5437 2308 5443 2452
rect 5453 2308 5459 2332
rect 5128 2257 5139 2263
rect 5133 2248 5139 2257
rect 5149 2188 5155 2272
rect 5101 2128 5107 2152
rect 5117 2128 5123 2152
rect 5165 2128 5171 2292
rect 5181 2288 5187 2292
rect 5181 2228 5187 2272
rect 5277 2248 5283 2272
rect 5181 2148 5187 2192
rect 5149 1908 5155 1952
rect 4941 1708 4947 1752
rect 4973 1728 4979 1772
rect 5037 1768 5043 1872
rect 5021 1728 5027 1732
rect 5085 1728 5091 1892
rect 5101 1788 5107 1892
rect 5133 1788 5139 1832
rect 5197 1808 5203 2232
rect 5325 2168 5331 2272
rect 5421 2268 5427 2272
rect 5421 2168 5427 2252
rect 5229 2148 5235 2152
rect 5405 2148 5411 2152
rect 5437 2148 5443 2292
rect 5469 2188 5475 2232
rect 5485 2168 5491 2432
rect 5517 2328 5523 2632
rect 5533 2528 5539 2792
rect 5597 2708 5603 2712
rect 5645 2708 5651 2852
rect 5661 2828 5667 2832
rect 5677 2688 5683 2912
rect 5693 2868 5699 2912
rect 5693 2708 5699 2832
rect 5549 2588 5555 2676
rect 5549 2528 5555 2532
rect 5613 2528 5619 2632
rect 5693 2508 5699 2512
rect 5597 2428 5603 2432
rect 5501 2308 5507 2312
rect 5533 2308 5539 2352
rect 5517 2288 5523 2292
rect 5597 2288 5603 2372
rect 5613 2308 5619 2332
rect 5693 2328 5699 2432
rect 5709 2428 5715 3032
rect 5773 2983 5779 3032
rect 5805 3008 5811 3092
rect 5853 3068 5859 3072
rect 5757 2977 5779 2983
rect 5725 2963 5731 2972
rect 5725 2957 5736 2963
rect 5757 2948 5763 2977
rect 5757 2708 5763 2712
rect 5773 2703 5779 2952
rect 5805 2928 5811 2952
rect 5837 2943 5843 3032
rect 5869 2968 5875 3076
rect 5885 3048 5891 3312
rect 5901 3268 5907 3432
rect 5933 3328 5939 3492
rect 5901 3128 5907 3232
rect 5928 3057 5939 3063
rect 5832 2937 5843 2943
rect 5768 2697 5779 2703
rect 5821 2688 5827 2712
rect 5741 2583 5747 2672
rect 5869 2668 5875 2692
rect 5805 2648 5811 2652
rect 5736 2577 5747 2583
rect 5789 2568 5795 2632
rect 5853 2628 5859 2632
rect 5693 2308 5699 2312
rect 5741 2308 5747 2412
rect 5757 2368 5763 2512
rect 5725 2288 5731 2292
rect 5565 2163 5571 2172
rect 5597 2168 5603 2272
rect 5560 2157 5571 2163
rect 5645 2143 5651 2232
rect 5661 2163 5667 2232
rect 5661 2157 5672 2163
rect 5645 2137 5656 2143
rect 5453 2128 5459 2132
rect 5485 2128 5491 2132
rect 5613 2128 5619 2132
rect 5709 2128 5715 2172
rect 5741 2148 5747 2292
rect 5757 2128 5763 2232
rect 5773 2228 5779 2512
rect 5789 2308 5795 2312
rect 5821 2308 5827 2352
rect 5789 2148 5795 2192
rect 5261 2117 5272 2123
rect 5229 2048 5235 2112
rect 5229 1928 5235 2032
rect 5261 1948 5267 2117
rect 5341 2108 5347 2112
rect 5357 2108 5363 2112
rect 5693 2108 5699 2112
rect 5261 1928 5267 1932
rect 5261 1908 5267 1912
rect 5133 1748 5139 1752
rect 5101 1728 5107 1732
rect 5149 1728 5155 1752
rect 5181 1728 5187 1752
rect 4685 1568 4691 1632
rect 4717 1508 4723 1652
rect 4781 1508 4787 1512
rect 4813 1508 4819 1692
rect 4829 1508 4835 1552
rect 4845 1508 4851 1632
rect 4589 1483 4595 1492
rect 4781 1488 4787 1492
rect 4584 1477 4595 1483
rect 4093 1348 4099 1352
rect 4253 1348 4259 1432
rect 4333 1408 4339 1432
rect 3725 1208 3731 1232
rect 3869 1208 3875 1312
rect 3885 1108 3891 1152
rect 3901 1108 3907 1272
rect 3965 1108 3971 1112
rect 3549 1068 3555 1072
rect 3485 1048 3491 1052
rect 3629 1043 3635 1072
rect 3645 1068 3651 1072
rect 3677 1063 3683 1092
rect 3661 1057 3683 1063
rect 3629 1037 3651 1043
rect 3501 1008 3507 1032
rect 3453 968 3459 972
rect 3485 943 3491 992
rect 3485 937 3496 943
rect 3437 908 3443 932
rect 3485 908 3491 912
rect 3549 908 3555 952
rect 3565 948 3571 952
rect 3581 948 3587 952
rect 3629 928 3635 932
rect 3645 868 3651 1037
rect 3661 1028 3667 1057
rect 3677 968 3683 1032
rect 3709 923 3715 1032
rect 3709 917 3720 923
rect 3421 837 3432 843
rect 3309 563 3315 632
rect 3373 608 3379 832
rect 3309 557 3320 563
rect 3336 537 3347 543
rect 3341 528 3347 537
rect 2557 308 2563 432
rect 2029 -43 2051 -37
rect 2093 -43 2099 12
rect 2205 -43 2211 32
rect 2253 -43 2259 12
rect 2333 -43 2339 32
rect 2381 -43 2387 12
rect 2429 -43 2435 12
rect 2477 -43 2483 52
rect 2573 -43 2579 492
rect 2685 288 2691 372
rect 2733 292 2739 352
rect 2749 308 2755 432
rect 2605 268 2611 272
rect 2605 188 2611 252
rect 2669 188 2675 276
rect 2701 143 2707 232
rect 2733 168 2739 276
rect 2781 148 2787 192
rect 2845 148 2851 252
rect 2701 137 2712 143
rect 2605 123 2611 132
rect 2605 117 2616 123
rect 2653 -43 2659 32
rect 2957 -37 2963 492
rect 3005 488 3011 492
rect 3053 308 3059 312
rect 3069 288 3075 312
rect 3149 308 3155 492
rect 3213 488 3219 512
rect 3277 368 3283 432
rect 3389 408 3395 512
rect 3357 308 3363 332
rect 3085 128 3091 232
rect 3117 168 3123 292
rect 3405 288 3411 292
rect 3421 288 3427 837
rect 3437 788 3443 792
rect 3437 588 3443 752
rect 3501 688 3507 732
rect 3565 688 3571 752
rect 3629 708 3635 712
rect 3517 648 3523 652
rect 3581 648 3587 652
rect 3597 628 3603 632
rect 3501 548 3507 592
rect 3629 544 3635 552
rect 3645 548 3651 832
rect 3677 668 3683 832
rect 3741 703 3747 1092
rect 3821 1088 3827 1092
rect 3773 828 3779 1052
rect 3837 988 3843 1052
rect 3885 1048 3891 1092
rect 3949 1048 3955 1092
rect 3805 968 3811 972
rect 3853 948 3859 1032
rect 3917 963 3923 1032
rect 3917 957 3928 963
rect 3869 888 3875 952
rect 3917 928 3923 932
rect 3773 708 3779 712
rect 3821 708 3827 832
rect 3885 748 3891 832
rect 3741 697 3752 703
rect 3693 688 3699 692
rect 3853 688 3859 692
rect 3949 688 3955 792
rect 3981 788 3987 932
rect 3709 648 3715 652
rect 3709 568 3715 632
rect 3725 608 3731 632
rect 3853 568 3859 572
rect 3869 548 3875 572
rect 3592 537 3603 543
rect 3597 528 3603 537
rect 3693 368 3699 532
rect 3917 528 3923 652
rect 3965 648 3971 652
rect 3965 548 3971 632
rect 4029 523 4035 1232
rect 4045 1088 4051 1252
rect 4045 1068 4051 1072
rect 4061 1068 4067 1092
rect 4077 1063 4083 1312
rect 4125 1088 4131 1232
rect 4157 1228 4163 1232
rect 4141 1188 4147 1192
rect 4205 1188 4211 1332
rect 4317 1288 4323 1332
rect 4333 1268 4339 1352
rect 4349 1308 4355 1432
rect 4381 1348 4387 1372
rect 4173 1088 4179 1152
rect 4136 1077 4147 1083
rect 4077 1057 4099 1063
rect 4077 968 4083 1032
rect 4072 937 4083 943
rect 4077 788 4083 937
rect 4045 688 4051 732
rect 4061 668 4067 672
rect 4061 568 4067 652
rect 4093 583 4099 1057
rect 4125 928 4131 1052
rect 4141 1008 4147 1077
rect 4157 988 4163 1052
rect 4221 988 4227 1232
rect 4429 1188 4435 1332
rect 4541 1328 4547 1392
rect 4589 1368 4595 1432
rect 4573 1337 4584 1343
rect 4573 1328 4579 1337
rect 4717 1328 4723 1472
rect 4797 1468 4803 1472
rect 4733 1348 4739 1412
rect 4845 1363 4851 1372
rect 4840 1357 4851 1363
rect 4877 1328 4883 1352
rect 4237 1117 4248 1123
rect 4237 1108 4243 1117
rect 4333 1088 4339 1132
rect 4269 1028 4275 1032
rect 4237 963 4243 972
rect 4232 957 4243 963
rect 4205 948 4211 952
rect 4269 944 4275 1012
rect 4301 948 4307 1072
rect 4333 948 4339 972
rect 4381 968 4387 1032
rect 4413 968 4419 1052
rect 4429 1048 4435 1072
rect 4445 1068 4451 1232
rect 4493 1088 4499 1132
rect 4525 1088 4531 1312
rect 4573 1088 4579 1292
rect 4637 1208 4643 1232
rect 4701 1228 4707 1312
rect 4520 1057 4531 1063
rect 4445 1028 4451 1052
rect 4525 1048 4531 1057
rect 4477 968 4483 992
rect 4541 968 4547 992
rect 4525 948 4531 952
rect 4109 688 4115 732
rect 4125 688 4131 912
rect 4173 688 4179 832
rect 4253 708 4259 832
rect 4301 688 4307 932
rect 4317 688 4323 812
rect 4365 708 4371 832
rect 4429 708 4435 832
rect 4557 788 4563 832
rect 4477 688 4483 712
rect 4557 688 4563 752
rect 4573 688 4579 1072
rect 4637 1068 4643 1072
rect 4701 1068 4707 1072
rect 4589 963 4595 1032
rect 4653 1008 4659 1032
rect 4589 957 4600 963
rect 4669 948 4675 992
rect 4685 928 4691 932
rect 4717 928 4723 1072
rect 4733 928 4739 1252
rect 4797 1108 4803 1112
rect 4829 1108 4835 1152
rect 4765 1068 4771 1072
rect 4589 788 4595 792
rect 4637 708 4643 712
rect 4621 688 4627 692
rect 4125 648 4131 652
rect 4189 648 4195 652
rect 4088 577 4099 583
rect 4125 568 4131 612
rect 4189 568 4195 612
rect 4029 517 4040 523
rect 4109 508 4115 532
rect 3789 306 3795 312
rect 3901 288 3907 432
rect 3965 308 3971 312
rect 4061 308 4067 332
rect 4125 317 4136 323
rect 4125 308 4131 317
rect 3272 277 3283 283
rect 3197 188 3203 252
rect 3277 248 3283 277
rect 3421 268 3427 272
rect 3517 268 3523 272
rect 3565 248 3571 272
rect 3757 248 3763 272
rect 3736 237 3747 243
rect 3277 188 3283 232
rect 3469 208 3475 232
rect 3117 123 3123 132
rect 3117 117 3128 123
rect 3565 123 3571 132
rect 3629 128 3635 192
rect 3741 148 3747 237
rect 3757 168 3763 232
rect 3917 203 3923 232
rect 3917 197 3939 203
rect 4077 208 4083 272
rect 3869 148 3875 172
rect 3725 128 3731 132
rect 3933 128 3939 197
rect 4125 163 4131 292
rect 4141 188 4147 272
rect 4173 248 4179 532
rect 4205 528 4211 652
rect 4269 568 4275 632
rect 4301 588 4307 672
rect 4317 668 4323 672
rect 4381 668 4387 672
rect 4461 648 4467 652
rect 4317 588 4323 612
rect 4381 568 4387 632
rect 4573 588 4579 652
rect 4589 588 4595 652
rect 4461 563 4467 572
rect 4637 568 4643 592
rect 4685 588 4691 672
rect 4701 668 4707 852
rect 4733 688 4739 912
rect 4781 788 4787 912
rect 4813 692 4819 772
rect 4829 703 4835 1092
rect 4845 1028 4851 1032
rect 4861 948 4867 1172
rect 4877 1108 4883 1312
rect 4893 1308 4899 1632
rect 5005 1528 5011 1632
rect 5101 1508 5107 1632
rect 5197 1508 5203 1732
rect 5229 1723 5235 1812
rect 5245 1743 5251 1892
rect 5245 1737 5267 1743
rect 5261 1728 5267 1737
rect 5229 1717 5240 1723
rect 5245 1508 5251 1512
rect 5277 1508 5283 2072
rect 5373 2068 5379 2072
rect 5485 1908 5491 2032
rect 5533 1908 5539 1912
rect 5293 1728 5299 1832
rect 5309 1828 5315 1892
rect 5325 1888 5331 1892
rect 5373 1888 5379 1892
rect 5421 1888 5427 1892
rect 5341 1728 5347 1732
rect 5373 1728 5379 1872
rect 5389 1808 5395 1872
rect 5389 1728 5395 1732
rect 5357 1708 5363 1712
rect 5373 1508 5379 1712
rect 5405 1668 5411 1872
rect 5485 1868 5491 1892
rect 5581 1888 5587 2092
rect 5741 1948 5747 2032
rect 5805 1988 5811 2272
rect 5645 1908 5651 1912
rect 5437 1728 5443 1772
rect 5453 1748 5459 1832
rect 5517 1768 5523 1772
rect 5517 1723 5523 1732
rect 5501 1717 5523 1723
rect 5453 1708 5459 1712
rect 5405 1508 5411 1612
rect 4909 1348 4915 1392
rect 5005 1348 5011 1472
rect 5261 1468 5267 1492
rect 5293 1468 5299 1492
rect 5421 1468 5427 1492
rect 5453 1457 5464 1463
rect 5453 1448 5459 1457
rect 5021 1248 5027 1432
rect 5085 1348 5091 1392
rect 5117 1343 5123 1432
rect 5325 1363 5331 1432
rect 5341 1388 5347 1432
rect 5501 1428 5507 1717
rect 5533 1508 5539 1792
rect 5549 1728 5555 1872
rect 5565 1488 5571 1832
rect 5597 1728 5603 1792
rect 5613 1788 5619 1872
rect 5677 1768 5683 1832
rect 5693 1783 5699 1832
rect 5725 1828 5731 1892
rect 5725 1788 5731 1812
rect 5693 1777 5715 1783
rect 5645 1728 5651 1752
rect 5693 1743 5699 1752
rect 5709 1748 5715 1777
rect 5821 1783 5827 1832
rect 5837 1808 5843 2532
rect 5869 2308 5875 2632
rect 5885 2468 5891 2912
rect 5901 2728 5907 3032
rect 5917 2588 5923 2832
rect 5933 2623 5939 3057
rect 5949 2928 5955 3312
rect 5965 3028 5971 3032
rect 5933 2617 5955 2623
rect 5928 2537 5939 2543
rect 5933 2388 5939 2537
rect 5901 2308 5907 2312
rect 5869 2188 5875 2292
rect 5885 2188 5891 2212
rect 5885 1908 5891 2112
rect 5853 1868 5859 1892
rect 5869 1888 5875 1892
rect 5901 1808 5907 1892
rect 5821 1777 5843 1783
rect 5837 1748 5843 1777
rect 5677 1737 5699 1743
rect 5677 1728 5683 1737
rect 5773 1728 5779 1732
rect 5901 1728 5907 1772
rect 5645 1508 5651 1512
rect 5709 1508 5715 1512
rect 5549 1468 5555 1476
rect 5357 1368 5363 1372
rect 5325 1357 5336 1363
rect 5277 1348 5283 1352
rect 5117 1337 5128 1343
rect 5165 1328 5171 1332
rect 5213 1328 5219 1332
rect 5261 1328 5267 1332
rect 5181 1308 5187 1312
rect 5373 1308 5379 1332
rect 5405 1328 5411 1412
rect 4877 1088 4883 1092
rect 4877 948 4883 1072
rect 4909 1008 4915 1032
rect 4925 928 4931 1092
rect 4941 1088 4947 1232
rect 4957 1108 4963 1232
rect 5101 1188 5107 1232
rect 5101 1088 5107 1132
rect 5165 1108 5171 1292
rect 5229 1108 5235 1152
rect 5293 1108 5299 1192
rect 5373 1108 5379 1292
rect 4968 1057 4979 1063
rect 4973 1048 4979 1057
rect 5053 1048 5059 1072
rect 5128 1057 5139 1063
rect 5133 1048 5139 1057
rect 5053 988 5059 1032
rect 4845 788 4851 912
rect 4957 708 4963 712
rect 4829 697 4840 703
rect 4717 608 4723 632
rect 4749 608 4755 676
rect 4456 557 4467 563
rect 4717 563 4723 572
rect 4712 557 4723 563
rect 4285 488 4291 532
rect 4285 388 4291 392
rect 4221 283 4227 292
rect 4317 288 4323 312
rect 4381 308 4387 552
rect 4429 548 4435 552
rect 4557 528 4563 552
rect 4685 548 4691 552
rect 4493 488 4499 512
rect 4525 508 4531 512
rect 4541 408 4547 512
rect 4621 488 4627 532
rect 4749 528 4755 592
rect 4765 548 4771 652
rect 4813 528 4819 676
rect 4877 608 4883 632
rect 4941 628 4947 692
rect 4989 668 4995 952
rect 5085 948 5091 972
rect 5133 948 5139 1012
rect 5229 1008 5235 1092
rect 5405 1088 5411 1312
rect 5517 1308 5523 1432
rect 5533 1388 5539 1392
rect 5549 1388 5555 1452
rect 5549 1363 5555 1372
rect 5581 1368 5587 1432
rect 5533 1357 5555 1363
rect 5421 1108 5427 1132
rect 5181 988 5187 992
rect 5277 968 5283 972
rect 5325 968 5331 1052
rect 5261 928 5267 932
rect 5005 688 5011 732
rect 4216 277 4227 283
rect 4333 268 4339 292
rect 4445 288 4451 372
rect 4381 208 4387 272
rect 4461 268 4467 292
rect 4477 268 4483 332
rect 4701 308 4707 452
rect 4717 308 4723 392
rect 4813 283 4819 512
rect 4861 388 4867 392
rect 4829 308 4835 312
rect 4877 308 4883 572
rect 4893 568 4899 572
rect 4909 528 4915 612
rect 4925 328 4931 332
rect 4957 328 4963 512
rect 4973 388 4979 612
rect 4989 588 4995 652
rect 5069 628 5075 912
rect 5101 748 5107 832
rect 5101 608 5107 692
rect 5117 688 5123 712
rect 5181 708 5187 832
rect 5181 588 5187 672
rect 5213 648 5219 912
rect 5293 728 5299 832
rect 5261 683 5267 692
rect 5357 688 5363 832
rect 5373 788 5379 1072
rect 5389 968 5395 1032
rect 5405 948 5411 1052
rect 5421 1028 5427 1052
rect 5453 948 5459 1032
rect 5469 948 5475 1292
rect 5485 1108 5491 1112
rect 5517 1108 5523 1212
rect 5533 1148 5539 1357
rect 5709 1348 5715 1472
rect 5741 1468 5747 1632
rect 5805 1528 5811 1712
rect 5736 1437 5747 1443
rect 5672 1337 5683 1343
rect 5549 1308 5555 1332
rect 5677 1328 5683 1337
rect 5565 1168 5571 1312
rect 5533 1108 5539 1132
rect 5613 1108 5619 1152
rect 5677 1108 5683 1112
rect 5693 1103 5699 1332
rect 5725 1328 5731 1412
rect 5688 1097 5699 1103
rect 5581 1048 5587 1052
rect 5565 968 5571 1032
rect 5581 944 5587 1012
rect 5645 948 5651 1032
rect 5389 768 5395 912
rect 5453 708 5459 892
rect 5469 743 5475 872
rect 5485 788 5491 912
rect 5469 737 5491 743
rect 5437 688 5443 692
rect 5256 677 5267 683
rect 5384 657 5395 663
rect 5005 528 5011 532
rect 5213 528 5219 592
rect 5165 428 5171 512
rect 4973 348 4979 372
rect 5005 308 5011 312
rect 4813 277 4835 283
rect 4221 168 4227 192
rect 4525 168 4531 272
rect 4749 248 4755 252
rect 4685 228 4691 232
rect 4120 157 4131 163
rect 4269 148 4275 152
rect 4077 128 4083 132
rect 3565 117 3576 123
rect 4157 123 4163 132
rect 4157 117 4168 123
rect 4477 123 4483 132
rect 4477 117 4488 123
rect 4589 123 4595 132
rect 4621 128 4627 212
rect 4637 168 4643 172
rect 4829 168 4835 277
rect 4685 148 4691 152
rect 4925 148 4931 232
rect 4957 168 4963 212
rect 5021 188 5027 352
rect 5149 328 5155 332
rect 5245 328 5251 592
rect 5277 548 5283 572
rect 5293 568 5299 652
rect 5389 648 5395 657
rect 5309 528 5315 632
rect 5341 588 5347 592
rect 5437 563 5443 572
rect 5432 557 5443 563
rect 5405 548 5411 552
rect 5245 308 5251 312
rect 5309 303 5315 512
rect 5325 328 5331 512
rect 5325 308 5331 312
rect 5421 308 5427 532
rect 5469 528 5475 672
rect 5485 528 5491 737
rect 5549 708 5555 752
rect 5565 708 5571 912
rect 5645 768 5651 912
rect 5645 708 5651 732
rect 5677 708 5683 1092
rect 5725 988 5731 1312
rect 5741 948 5747 1437
rect 5821 1343 5827 1372
rect 5837 1363 5843 1432
rect 5853 1388 5859 1432
rect 5837 1357 5848 1363
rect 5821 1337 5832 1343
rect 5869 1268 5875 1632
rect 5901 1508 5907 1692
rect 5885 1448 5891 1492
rect 5917 1488 5923 1492
rect 5917 1448 5923 1452
rect 5757 1088 5763 1112
rect 5805 1108 5811 1232
rect 5768 1057 5779 1063
rect 5773 1048 5779 1057
rect 5517 568 5523 632
rect 5533 588 5539 592
rect 5549 588 5555 692
rect 5533 528 5539 572
rect 5581 543 5587 632
rect 5613 628 5619 692
rect 5661 688 5667 692
rect 5725 668 5731 932
rect 5757 688 5763 972
rect 5773 948 5779 972
rect 5805 968 5811 1092
rect 5789 943 5795 952
rect 5789 937 5811 943
rect 5805 928 5811 937
rect 5821 728 5827 1072
rect 5837 1028 5843 1032
rect 5837 928 5843 952
rect 5853 928 5859 1252
rect 5869 1128 5875 1232
rect 5869 1088 5875 1092
rect 5885 1088 5891 1432
rect 5901 1108 5907 1292
rect 5885 1068 5891 1072
rect 5869 988 5875 1032
rect 5693 563 5699 632
rect 5709 568 5715 632
rect 5725 568 5731 612
rect 5688 557 5699 563
rect 5581 537 5592 543
rect 5688 537 5699 543
rect 5693 528 5699 537
rect 5725 528 5731 552
rect 5757 548 5763 652
rect 5773 603 5779 632
rect 5773 597 5795 603
rect 5773 528 5779 572
rect 5437 308 5443 312
rect 5304 297 5315 303
rect 5117 268 5123 272
rect 5069 188 5075 232
rect 5117 188 5123 192
rect 5133 188 5139 292
rect 5469 288 5475 512
rect 5485 288 5491 512
rect 5597 288 5603 392
rect 5613 288 5619 412
rect 5629 408 5635 432
rect 5741 308 5747 432
rect 5693 288 5699 292
rect 5229 228 5235 272
rect 5597 268 5603 272
rect 5677 268 5683 272
rect 5245 188 5251 232
rect 5277 223 5283 232
rect 5277 217 5299 223
rect 5181 163 5187 172
rect 5176 157 5187 163
rect 4584 117 4595 123
rect 4893 123 4899 132
rect 5213 128 5219 172
rect 5277 148 5283 192
rect 5293 168 5299 217
rect 5357 208 5363 232
rect 5341 148 5347 172
rect 5469 168 5475 232
rect 5485 188 5491 252
rect 5533 168 5539 232
rect 5549 208 5555 232
rect 5389 144 5395 152
rect 5357 128 5363 132
rect 5517 144 5523 152
rect 5581 148 5587 192
rect 5597 168 5603 172
rect 5661 163 5667 232
rect 5661 157 5672 163
rect 5709 163 5715 212
rect 5725 188 5731 232
rect 5709 157 5720 163
rect 5613 148 5619 152
rect 5773 148 5779 332
rect 5789 283 5795 597
rect 5805 588 5811 692
rect 5837 688 5843 912
rect 5853 688 5859 912
rect 5885 863 5891 1052
rect 5933 968 5939 1832
rect 5949 1788 5955 2617
rect 5965 2128 5971 2432
rect 5981 1988 5987 3872
rect 5997 2708 6003 2772
rect 5965 1328 5971 1452
rect 5949 988 5955 1032
rect 5869 857 5891 863
rect 5821 668 5827 672
rect 5837 668 5843 672
rect 5869 568 5875 857
rect 5917 708 5923 712
rect 5965 708 5971 1312
rect 5885 588 5891 592
rect 5805 348 5811 432
rect 5821 308 5827 432
rect 5917 388 5923 672
rect 5933 568 5939 572
rect 5981 388 5987 532
rect 5869 308 5875 372
rect 5933 288 5939 312
rect 5789 277 5800 283
rect 5789 208 5795 232
rect 5789 168 5795 172
rect 5837 148 5843 192
rect 5853 168 5859 232
rect 5901 188 5907 232
rect 5981 188 5987 352
rect 5453 128 5459 132
rect 5949 144 5955 152
rect 4893 117 4904 123
rect 3245 108 3251 112
rect 5533 108 5539 112
rect 2957 -43 2979 -37
rect 3069 -43 3075 32
rect 3117 -43 3123 12
rect 3165 -43 3171 32
rect 3213 -43 3219 12
rect 3245 -37 3251 92
rect 3245 -43 3267 -37
rect 3613 -43 3619 32
rect 3661 28 3667 32
rect 3677 -37 3683 32
rect 3709 28 3715 32
rect 3661 -43 3683 -37
rect 3693 -37 3699 12
rect 3693 -43 3715 -37
rect 3741 -43 3747 12
rect 3789 -43 3795 12
rect 3965 -43 3971 32
rect 4205 -43 4211 32
rect 4525 -43 4531 32
rect 4541 28 4547 32
rect 4573 -43 4579 12
rect 4941 -43 4947 32
<< m3contact >>
rect 392 4012 408 4028
rect 344 3912 360 3928
rect 472 4012 504 4028
rect 24 3792 40 3808
rect 8 3772 24 3788
rect 72 3852 88 3868
rect 40 3752 56 3768
rect 8 3732 24 3748
rect 200 3832 216 3848
rect 136 3792 152 3808
rect 168 3792 184 3808
rect 168 3752 184 3768
rect 216 3752 232 3768
rect 328 3872 344 3888
rect 440 3872 456 3888
rect 360 3852 376 3868
rect 408 3852 424 3868
rect 456 3832 472 3848
rect 376 3812 392 3828
rect 296 3792 312 3808
rect 360 3792 376 3808
rect 312 3772 328 3788
rect 392 3772 408 3788
rect 424 3752 440 3768
rect 925 4002 961 4018
rect 888 3972 904 3988
rect 536 3912 552 3928
rect 1144 3952 1160 3968
rect 1192 3952 1208 3968
rect 1048 3912 1064 3928
rect 488 3892 504 3908
rect 584 3892 600 3908
rect 520 3852 552 3868
rect 504 3732 520 3748
rect 680 3832 696 3848
rect 744 3832 760 3848
rect 552 3812 568 3828
rect 632 3812 648 3828
rect 632 3752 648 3768
rect 680 3752 696 3768
rect 552 3732 568 3748
rect 600 3732 616 3748
rect 184 3712 200 3728
rect 88 3692 104 3708
rect 40 3512 56 3528
rect 168 3512 184 3528
rect 248 3652 264 3668
rect 56 3492 72 3508
rect 184 3492 200 3508
rect 56 3472 72 3488
rect 456 3532 472 3548
rect 424 3512 440 3528
rect 568 3692 584 3708
rect 520 3612 536 3628
rect 568 3572 584 3588
rect 632 3732 648 3748
rect 808 3832 824 3848
rect 936 3872 952 3888
rect 2104 3992 2120 4008
rect 1176 3892 1192 3908
rect 1320 3892 1336 3908
rect 1416 3892 1432 3908
rect 952 3852 968 3868
rect 904 3832 920 3848
rect 824 3812 840 3828
rect 776 3792 792 3808
rect 744 3752 760 3768
rect 776 3752 792 3768
rect 824 3752 840 3768
rect 856 3772 872 3788
rect 792 3732 808 3748
rect 872 3732 888 3748
rect 1032 3792 1048 3808
rect 968 3772 984 3788
rect 1176 3872 1192 3888
rect 1224 3872 1240 3888
rect 1128 3852 1144 3868
rect 1208 3852 1224 3868
rect 1096 3812 1112 3828
rect 968 3752 984 3768
rect 1064 3752 1080 3768
rect 872 3712 888 3728
rect 936 3712 952 3728
rect 888 3692 904 3708
rect 728 3672 744 3688
rect 824 3672 840 3688
rect 632 3552 648 3568
rect 472 3512 488 3528
rect 616 3512 632 3528
rect 328 3492 344 3508
rect 424 3492 440 3508
rect 552 3492 568 3508
rect 616 3492 632 3508
rect 88 3452 120 3468
rect 24 3332 40 3348
rect 72 3332 88 3348
rect 248 3472 264 3488
rect 808 3632 824 3648
rect 664 3492 680 3508
rect 344 3452 360 3468
rect 568 3472 584 3488
rect 648 3472 664 3488
rect 840 3632 856 3648
rect 925 3602 961 3618
rect 840 3552 856 3568
rect 856 3492 872 3508
rect 792 3452 808 3468
rect 232 3432 248 3448
rect 280 3432 296 3448
rect 472 3432 488 3448
rect 664 3432 680 3448
rect 120 3372 136 3388
rect 248 3392 264 3408
rect 392 3392 408 3408
rect 392 3372 408 3388
rect 440 3372 456 3388
rect 376 3352 392 3368
rect 616 3412 632 3428
rect 552 3392 568 3408
rect 584 3392 600 3408
rect 568 3352 584 3368
rect 664 3392 680 3408
rect 632 3372 648 3388
rect 200 3332 216 3348
rect 232 3332 248 3348
rect 376 3332 392 3348
rect 360 3272 376 3288
rect 56 3212 72 3228
rect 200 3232 216 3248
rect 360 3112 376 3128
rect 280 3092 296 3108
rect 328 3092 344 3108
rect 392 3272 424 3288
rect 88 3052 104 3068
rect 24 3012 56 3028
rect 8 2972 24 2988
rect 8 2932 24 2948
rect 88 2972 104 2988
rect 120 2972 136 2988
rect 56 2952 72 2968
rect 56 2692 72 2708
rect 216 3072 232 3088
rect 264 3072 280 3088
rect 440 3232 456 3248
rect 568 3212 600 3228
rect 440 3092 456 3108
rect 552 3092 568 3108
rect 488 3072 504 3088
rect 488 3052 504 3068
rect 168 3012 184 3028
rect 184 2992 200 3008
rect 120 2952 136 2968
rect 136 2952 152 2968
rect 168 2952 184 2968
rect 104 2912 120 2928
rect 376 3032 392 3048
rect 376 3012 392 3028
rect 328 2992 344 3008
rect 376 2992 392 3008
rect 232 2972 248 2988
rect 312 2972 328 2988
rect 312 2952 328 2968
rect 408 2972 424 2988
rect 248 2932 264 2948
rect 392 2932 408 2948
rect 456 2932 472 2948
rect 264 2912 280 2928
rect 200 2872 216 2888
rect 232 2872 248 2888
rect 296 2872 312 2888
rect 104 2712 120 2728
rect 24 2552 40 2568
rect 40 2552 56 2568
rect 8 2512 24 2528
rect 40 2352 56 2368
rect 88 2652 104 2668
rect 72 2592 88 2608
rect 72 2512 88 2528
rect 104 2352 120 2368
rect 136 2432 152 2448
rect 296 2732 312 2748
rect 232 2712 248 2728
rect 504 2992 520 3008
rect 632 3152 648 3168
rect 648 3092 664 3108
rect 712 3392 728 3408
rect 776 3352 792 3368
rect 824 3452 840 3468
rect 1016 3712 1032 3728
rect 1048 3712 1064 3728
rect 1080 3712 1096 3728
rect 1192 3812 1208 3828
rect 1144 3752 1160 3768
rect 1128 3712 1144 3728
rect 1272 3872 1288 3888
rect 1336 3872 1352 3888
rect 1384 3872 1400 3888
rect 1448 3876 1480 3888
rect 1448 3872 1464 3876
rect 1464 3872 1480 3876
rect 1400 3832 1416 3848
rect 1288 3812 1304 3828
rect 1240 3792 1256 3808
rect 1352 3792 1368 3808
rect 1400 3792 1416 3808
rect 1208 3772 1224 3788
rect 1240 3772 1256 3788
rect 1096 3692 1112 3708
rect 1144 3692 1160 3708
rect 1064 3672 1080 3688
rect 1112 3672 1128 3688
rect 1160 3652 1176 3668
rect 1016 3612 1032 3628
rect 1032 3552 1048 3568
rect 1032 3512 1048 3528
rect 984 3492 1000 3508
rect 1096 3492 1112 3508
rect 936 3472 952 3488
rect 1096 3472 1112 3488
rect 920 3392 936 3408
rect 968 3392 984 3408
rect 856 3372 872 3388
rect 808 3332 824 3348
rect 1096 3452 1112 3468
rect 1064 3392 1080 3408
rect 1032 3332 1048 3348
rect 1048 3332 1064 3348
rect 824 3312 840 3328
rect 872 3312 904 3328
rect 808 3292 824 3308
rect 744 3272 760 3288
rect 776 3272 792 3288
rect 760 3172 776 3188
rect 616 3076 632 3088
rect 616 3072 632 3076
rect 616 3052 632 3068
rect 1064 3312 1080 3328
rect 1048 3272 1064 3288
rect 824 3252 840 3268
rect 1160 3512 1176 3528
rect 1144 3492 1160 3508
rect 1320 3732 1336 3748
rect 1272 3712 1288 3728
rect 1480 3792 1496 3808
rect 1448 3744 1464 3748
rect 1448 3732 1464 3744
rect 1464 3692 1480 3708
rect 1336 3672 1352 3688
rect 1256 3552 1272 3568
rect 1480 3632 1496 3648
rect 1592 3932 1608 3948
rect 1912 3932 1928 3948
rect 2008 3932 2024 3948
rect 1592 3892 1608 3908
rect 1656 3892 1672 3908
rect 1528 3872 1544 3888
rect 1512 3812 1528 3828
rect 1512 3792 1528 3808
rect 1448 3552 1464 3568
rect 1352 3532 1368 3548
rect 1400 3532 1416 3548
rect 1240 3492 1256 3508
rect 1336 3492 1352 3508
rect 1416 3492 1432 3508
rect 1336 3472 1352 3488
rect 1352 3472 1368 3488
rect 1400 3472 1416 3488
rect 1288 3452 1304 3468
rect 1176 3432 1192 3448
rect 1224 3432 1240 3448
rect 1304 3432 1320 3448
rect 1192 3412 1208 3428
rect 1272 3392 1288 3408
rect 1336 3392 1352 3408
rect 1096 3344 1112 3348
rect 1112 3344 1128 3348
rect 1096 3332 1128 3344
rect 1160 3332 1176 3348
rect 840 3232 856 3248
rect 904 3212 920 3228
rect 925 3202 961 3218
rect 888 3112 904 3128
rect 1080 3232 1096 3248
rect 1176 3312 1192 3328
rect 1224 3312 1240 3328
rect 1320 3292 1336 3308
rect 1320 3232 1336 3248
rect 1160 3172 1176 3188
rect 1144 3112 1160 3128
rect 872 3052 888 3068
rect 600 3032 632 3048
rect 648 3032 664 3048
rect 744 3032 760 3048
rect 824 3032 840 3048
rect 584 2972 600 2988
rect 520 2932 536 2948
rect 360 2852 376 2868
rect 344 2692 360 2708
rect 248 2672 264 2688
rect 328 2672 344 2688
rect 168 2652 184 2668
rect 200 2652 216 2668
rect 184 2572 200 2588
rect 216 2572 232 2588
rect 248 2572 264 2588
rect 200 2532 216 2548
rect 168 2432 184 2448
rect 152 2352 168 2368
rect 184 2292 200 2308
rect 232 2552 248 2568
rect 344 2572 360 2588
rect 328 2552 344 2568
rect 440 2832 456 2848
rect 456 2812 472 2828
rect 424 2712 440 2728
rect 584 2892 600 2908
rect 520 2832 536 2848
rect 488 2712 504 2728
rect 472 2692 488 2708
rect 472 2652 488 2668
rect 360 2552 376 2568
rect 264 2532 280 2548
rect 600 2732 616 2748
rect 536 2692 552 2708
rect 696 3012 712 3028
rect 664 2952 680 2968
rect 776 2952 792 2968
rect 840 2992 856 3008
rect 1288 3112 1304 3128
rect 1096 3092 1128 3108
rect 1176 3092 1192 3108
rect 1288 3092 1304 3108
rect 1096 3072 1112 3088
rect 968 3052 984 3068
rect 1080 3052 1096 3068
rect 872 3012 888 3028
rect 904 3012 920 3028
rect 712 2912 728 2928
rect 808 2912 824 2928
rect 696 2892 712 2908
rect 632 2772 648 2788
rect 616 2712 632 2728
rect 808 2852 824 2868
rect 776 2832 792 2848
rect 728 2752 744 2768
rect 856 2912 872 2928
rect 600 2672 616 2688
rect 808 2672 824 2688
rect 840 2652 856 2668
rect 680 2632 696 2648
rect 568 2612 584 2628
rect 504 2552 520 2568
rect 584 2552 600 2568
rect 584 2532 600 2548
rect 696 2532 712 2548
rect 744 2512 760 2528
rect 568 2492 584 2508
rect 664 2492 680 2508
rect 648 2472 664 2488
rect 392 2432 408 2448
rect 312 2412 328 2428
rect 376 2412 392 2428
rect 360 2372 376 2388
rect 424 2372 440 2388
rect 376 2332 392 2348
rect 392 2312 408 2328
rect 472 2352 488 2368
rect 520 2292 536 2308
rect 648 2372 664 2388
rect 584 2292 600 2308
rect 616 2292 632 2308
rect 392 2272 408 2288
rect 728 2472 744 2488
rect 952 2952 968 2968
rect 952 2932 968 2948
rect 936 2832 952 2848
rect 872 2672 888 2688
rect 856 2552 872 2568
rect 872 2532 888 2548
rect 888 2512 904 2528
rect 808 2492 824 2508
rect 760 2432 776 2448
rect 200 2252 216 2268
rect 264 2252 280 2268
rect 552 2252 568 2268
rect 72 2212 88 2228
rect 8 2192 24 2208
rect 136 2172 152 2188
rect 8 2152 24 2168
rect 72 2152 88 2168
rect 136 2152 152 2168
rect 200 2132 216 2148
rect 232 2132 248 2148
rect 184 2112 200 2128
rect 152 2092 168 2108
rect 56 2072 72 2088
rect 40 1912 56 1928
rect 40 1872 56 1888
rect 72 2032 88 2048
rect 72 1912 88 1928
rect 8 1852 24 1868
rect 56 1852 72 1868
rect 8 1792 24 1808
rect 280 2132 296 2148
rect 424 2212 440 2228
rect 408 2152 424 2168
rect 632 2212 648 2228
rect 536 2192 552 2208
rect 568 2192 584 2208
rect 504 2172 520 2188
rect 376 2132 392 2148
rect 552 2132 568 2148
rect 600 2132 616 2148
rect 632 2132 648 2148
rect 664 2132 680 2148
rect 312 2112 328 2128
rect 472 2112 488 2128
rect 648 2112 664 2128
rect 232 2092 264 2108
rect 504 2092 520 2108
rect 120 2072 136 2088
rect 184 2072 200 2088
rect 264 2072 280 2088
rect 360 2072 376 2088
rect 104 2032 120 2048
rect 136 2032 152 2048
rect 216 2032 232 2048
rect 328 2032 344 2048
rect 200 2012 216 2028
rect 168 1912 184 1928
rect 200 1892 216 1908
rect 344 2012 360 2028
rect 248 1912 264 1928
rect 280 1912 296 1928
rect 328 1892 344 1908
rect 152 1872 168 1888
rect 264 1852 280 1868
rect 136 1812 152 1828
rect 248 1792 264 1808
rect 88 1772 104 1788
rect 152 1772 168 1788
rect 104 1752 120 1768
rect 120 1732 136 1748
rect 216 1752 232 1768
rect 24 1712 40 1728
rect 184 1712 200 1728
rect 40 1692 56 1708
rect 56 1592 72 1608
rect 8 1552 24 1568
rect 168 1552 184 1568
rect 248 1712 264 1728
rect 280 1712 296 1728
rect 216 1612 232 1628
rect 312 1692 328 1708
rect 376 1852 392 1868
rect 360 1832 376 1848
rect 408 2032 424 2048
rect 712 2292 728 2308
rect 712 2232 728 2248
rect 792 2212 808 2228
rect 728 2152 744 2168
rect 776 2152 792 2168
rect 888 2352 904 2368
rect 925 2802 961 2818
rect 1176 3072 1192 3088
rect 1208 3072 1224 3088
rect 1256 3072 1272 3088
rect 1272 3072 1288 3088
rect 1192 3052 1208 3068
rect 1176 2992 1192 3008
rect 1000 2952 1016 2968
rect 1048 2952 1064 2968
rect 1112 2932 1128 2948
rect 1160 2932 1176 2948
rect 1208 2972 1224 2988
rect 1224 2932 1240 2948
rect 1416 3372 1432 3388
rect 1400 3332 1416 3348
rect 1448 3272 1464 3288
rect 1496 3332 1512 3348
rect 1480 3312 1496 3328
rect 1464 3232 1480 3248
rect 1496 3272 1512 3288
rect 1368 3152 1384 3168
rect 1480 3152 1496 3168
rect 1368 3132 1384 3148
rect 1448 3112 1464 3128
rect 1480 3112 1496 3128
rect 1384 3092 1400 3108
rect 1496 3092 1512 3108
rect 1768 3872 1784 3888
rect 1832 3876 1864 3888
rect 1832 3872 1848 3876
rect 1848 3872 1864 3876
rect 1736 3832 1752 3848
rect 1640 3812 1672 3828
rect 1576 3732 1592 3748
rect 1576 3712 1592 3728
rect 1800 3812 1816 3828
rect 1688 3752 1704 3768
rect 1768 3752 1784 3768
rect 2088 3912 2104 3928
rect 2216 4012 2232 4028
rect 2248 4012 2264 4028
rect 2200 3972 2216 3988
rect 2152 3912 2168 3928
rect 2120 3892 2136 3908
rect 2168 3892 2184 3908
rect 1864 3792 1880 3808
rect 1933 3802 1969 3818
rect 2008 3872 2024 3888
rect 1864 3752 1880 3768
rect 1896 3752 1912 3768
rect 1992 3752 2008 3768
rect 1832 3732 1848 3748
rect 1944 3732 1960 3748
rect 2120 3792 2136 3808
rect 2120 3772 2136 3788
rect 2072 3732 2088 3748
rect 1640 3712 1656 3728
rect 1704 3712 1736 3728
rect 1848 3712 1864 3728
rect 1912 3712 1928 3728
rect 1992 3712 2008 3728
rect 2088 3712 2104 3728
rect 1592 3692 1608 3708
rect 1544 3632 1560 3648
rect 1528 3552 1544 3568
rect 1560 3612 1576 3628
rect 1608 3532 1624 3548
rect 1560 3512 1576 3528
rect 1736 3632 1752 3648
rect 1800 3512 1816 3528
rect 1656 3492 1672 3508
rect 1704 3492 1720 3508
rect 1784 3492 1800 3508
rect 1864 3552 1880 3568
rect 1864 3512 1880 3528
rect 2120 3692 2136 3708
rect 2056 3652 2072 3668
rect 2104 3652 2120 3668
rect 2040 3532 2056 3548
rect 2200 3872 2216 3888
rect 2248 3992 2264 4008
rect 2504 3952 2520 3968
rect 2568 3952 2584 3968
rect 2440 3932 2456 3948
rect 2296 3912 2312 3928
rect 2344 3912 2360 3928
rect 2392 3912 2408 3928
rect 2232 3892 2248 3908
rect 2264 3892 2280 3908
rect 2376 3892 2392 3908
rect 2456 3892 2472 3908
rect 2248 3872 2264 3888
rect 2280 3872 2296 3888
rect 2312 3732 2328 3748
rect 2184 3712 2200 3728
rect 2216 3712 2232 3728
rect 2168 3692 2184 3708
rect 2264 3692 2280 3708
rect 2328 3692 2344 3708
rect 2152 3632 2168 3648
rect 2120 3592 2136 3608
rect 2376 3872 2392 3888
rect 2424 3812 2440 3828
rect 2360 3772 2376 3788
rect 2360 3732 2376 3748
rect 2488 3792 2504 3808
rect 2440 3732 2456 3748
rect 2520 3912 2536 3928
rect 2536 3892 2552 3908
rect 2552 3752 2568 3768
rect 2472 3712 2488 3728
rect 2584 3912 2600 3928
rect 2744 4012 2760 4028
rect 2648 3972 2664 3988
rect 2632 3892 2648 3908
rect 2616 3812 2632 3828
rect 2744 3892 2760 3908
rect 2920 4012 2936 4028
rect 2872 3972 2888 3988
rect 2840 3892 2856 3908
rect 2680 3872 2696 3888
rect 2712 3872 2744 3888
rect 2776 3872 2808 3888
rect 2664 3832 2680 3848
rect 2696 3772 2712 3788
rect 2760 3772 2776 3788
rect 2680 3752 2696 3768
rect 2920 3892 2936 3908
rect 2973 4002 3009 4018
rect 2840 3872 2856 3888
rect 2872 3872 2888 3888
rect 2904 3872 2920 3888
rect 2952 3872 2984 3888
rect 2872 3852 2888 3868
rect 3000 3832 3016 3848
rect 2968 3772 2984 3788
rect 2904 3752 2920 3768
rect 3000 3752 3016 3768
rect 3080 3912 3096 3928
rect 3048 3892 3064 3908
rect 3032 3812 3048 3828
rect 3112 3812 3128 3828
rect 2616 3712 2632 3728
rect 2728 3712 2744 3728
rect 2952 3712 2968 3728
rect 2984 3712 3000 3728
rect 3016 3712 3032 3728
rect 2328 3652 2360 3668
rect 2184 3612 2200 3628
rect 2312 3592 2328 3608
rect 2216 3572 2232 3588
rect 2280 3572 2296 3588
rect 2184 3512 2200 3528
rect 1896 3492 1912 3508
rect 1912 3492 1928 3508
rect 1992 3492 2008 3508
rect 1576 3472 1592 3488
rect 1720 3476 1736 3488
rect 1720 3472 1736 3476
rect 1832 3476 1848 3488
rect 1848 3476 1864 3488
rect 1832 3472 1864 3476
rect 1672 3452 1688 3468
rect 1736 3452 1752 3468
rect 1928 3452 1944 3468
rect 1736 3432 1752 3448
rect 1576 3392 1592 3408
rect 1544 3332 1560 3348
rect 1624 3412 1640 3428
rect 1656 3412 1672 3428
rect 1672 3352 1688 3368
rect 1608 3332 1624 3348
rect 1640 3332 1656 3348
rect 1720 3412 1736 3428
rect 1752 3412 1768 3428
rect 1752 3392 1768 3408
rect 1933 3402 1969 3418
rect 2424 3692 2440 3708
rect 2408 3592 2424 3608
rect 2376 3532 2392 3548
rect 2360 3512 2376 3528
rect 2504 3632 2520 3648
rect 2472 3592 2504 3608
rect 2536 3572 2552 3588
rect 2264 3492 2280 3508
rect 2328 3492 2344 3508
rect 2376 3492 2392 3508
rect 2424 3492 2440 3508
rect 2216 3432 2232 3448
rect 1992 3412 2008 3428
rect 2024 3412 2040 3428
rect 1976 3372 1992 3388
rect 1848 3352 1864 3368
rect 1880 3352 1896 3368
rect 1528 3312 1544 3328
rect 1784 3312 1800 3328
rect 1960 3312 1976 3328
rect 1592 3292 1608 3308
rect 1592 3232 1608 3248
rect 1800 3232 1816 3248
rect 1528 3132 1544 3148
rect 1656 3132 1672 3148
rect 1608 3112 1624 3128
rect 1544 3092 1560 3108
rect 1608 3092 1624 3108
rect 1640 3092 1656 3108
rect 1960 3212 1976 3228
rect 1880 3112 1912 3128
rect 1736 3092 1752 3108
rect 1512 3072 1544 3088
rect 1656 3072 1672 3088
rect 1528 3052 1544 3068
rect 1352 3032 1368 3048
rect 1416 2992 1432 3008
rect 1336 2972 1352 2988
rect 1352 2952 1368 2968
rect 1368 2952 1384 2968
rect 1256 2912 1272 2928
rect 1304 2912 1336 2928
rect 984 2852 1000 2868
rect 1016 2832 1032 2848
rect 920 2732 936 2748
rect 1000 2672 1016 2688
rect 936 2652 952 2668
rect 936 2612 952 2628
rect 1128 2772 1144 2788
rect 1224 2772 1240 2788
rect 1176 2712 1192 2728
rect 1080 2692 1096 2708
rect 1128 2672 1144 2688
rect 1080 2632 1096 2648
rect 1064 2572 1080 2588
rect 1416 2912 1432 2928
rect 1448 2912 1464 2928
rect 1480 2912 1496 2928
rect 1656 3012 1672 3028
rect 1640 2992 1656 3008
rect 1640 2972 1656 2988
rect 2104 3372 2120 3388
rect 2184 3372 2200 3388
rect 2056 3352 2072 3368
rect 2136 3352 2152 3368
rect 2168 3352 2184 3368
rect 2088 3332 2104 3348
rect 2008 3312 2024 3328
rect 2216 3292 2232 3308
rect 2120 3272 2136 3288
rect 2280 3412 2296 3428
rect 2360 3472 2376 3488
rect 2440 3472 2456 3488
rect 2296 3372 2312 3388
rect 2328 3372 2344 3388
rect 2568 3552 2584 3568
rect 2552 3532 2584 3548
rect 2648 3692 2664 3708
rect 2696 3692 2712 3708
rect 2696 3672 2728 3688
rect 2632 3552 2664 3568
rect 2488 3492 2504 3508
rect 2536 3472 2552 3488
rect 2520 3452 2536 3468
rect 2552 3432 2568 3448
rect 2600 3492 2616 3508
rect 2584 3472 2616 3488
rect 2568 3412 2584 3428
rect 2536 3392 2552 3408
rect 2536 3332 2552 3348
rect 2264 3312 2280 3328
rect 2584 3332 2600 3348
rect 2568 3292 2584 3308
rect 2088 3252 2104 3268
rect 1992 3192 2024 3208
rect 2024 3112 2040 3128
rect 1864 3072 1880 3088
rect 1944 3072 1960 3088
rect 1800 3052 1816 3068
rect 1752 3032 1768 3048
rect 1832 3032 1848 3048
rect 1672 2992 1688 3008
rect 1720 2992 1736 3008
rect 1672 2952 1688 2968
rect 1512 2892 1524 2908
rect 1524 2892 1528 2908
rect 1576 2892 1608 2908
rect 1400 2832 1416 2848
rect 1432 2832 1448 2848
rect 1368 2792 1384 2808
rect 1336 2772 1352 2788
rect 1288 2752 1304 2768
rect 1336 2752 1368 2768
rect 1368 2712 1384 2728
rect 1560 2832 1576 2848
rect 1528 2752 1544 2768
rect 1272 2692 1288 2708
rect 1416 2692 1432 2708
rect 1448 2692 1464 2708
rect 1544 2732 1560 2748
rect 1240 2672 1256 2688
rect 1192 2652 1208 2668
rect 1160 2612 1176 2628
rect 936 2552 952 2568
rect 1032 2552 1048 2568
rect 1128 2552 1144 2568
rect 920 2532 936 2548
rect 1000 2532 1016 2548
rect 1048 2532 1064 2548
rect 1112 2532 1128 2548
rect 1176 2532 1192 2548
rect 1224 2532 1240 2548
rect 1256 2532 1272 2548
rect 984 2492 1000 2508
rect 1080 2472 1096 2488
rect 1016 2452 1032 2468
rect 925 2402 961 2418
rect 968 2392 984 2408
rect 936 2352 952 2368
rect 872 2252 888 2268
rect 696 2144 712 2148
rect 696 2132 712 2144
rect 760 2144 776 2148
rect 760 2132 776 2144
rect 792 2132 808 2148
rect 840 2212 856 2228
rect 840 2192 856 2208
rect 856 2152 872 2168
rect 1000 2292 1016 2308
rect 984 2192 1000 2208
rect 952 2152 968 2168
rect 1400 2632 1416 2648
rect 1304 2572 1320 2588
rect 1368 2512 1384 2528
rect 1160 2372 1176 2388
rect 1272 2372 1288 2388
rect 1352 2352 1368 2368
rect 1288 2332 1320 2348
rect 1080 2312 1096 2328
rect 1112 2312 1128 2328
rect 1192 2312 1208 2328
rect 1032 2212 1048 2228
rect 1096 2232 1112 2248
rect 1064 2152 1080 2168
rect 1080 2152 1096 2168
rect 1112 2152 1128 2168
rect 1032 2144 1048 2148
rect 1032 2132 1048 2144
rect 1096 2112 1112 2128
rect 824 2072 840 2088
rect 680 2052 696 2068
rect 520 2032 536 2048
rect 488 1932 504 1948
rect 472 1912 488 1928
rect 424 1832 440 1848
rect 440 1832 456 1848
rect 376 1772 408 1788
rect 344 1752 360 1768
rect 360 1732 376 1748
rect 344 1712 360 1728
rect 584 2012 600 2028
rect 824 2012 840 2028
rect 712 1932 728 1948
rect 760 1912 776 1928
rect 696 1892 712 1908
rect 504 1872 520 1888
rect 472 1792 488 1808
rect 456 1772 472 1788
rect 584 1872 600 1888
rect 600 1872 616 1888
rect 648 1872 664 1888
rect 744 1892 760 1908
rect 792 1892 808 1908
rect 632 1852 648 1868
rect 520 1752 552 1768
rect 392 1732 408 1748
rect 408 1712 424 1728
rect 440 1692 456 1708
rect 536 1692 552 1708
rect 344 1672 360 1688
rect 328 1652 344 1668
rect 456 1652 472 1668
rect 264 1572 280 1588
rect 184 1532 200 1548
rect 424 1532 440 1548
rect 88 1492 104 1508
rect 152 1492 168 1508
rect 328 1506 344 1508
rect 328 1492 344 1506
rect 392 1492 408 1508
rect 440 1492 456 1508
rect 40 1472 56 1488
rect 104 1472 120 1488
rect 536 1552 552 1568
rect 504 1532 520 1548
rect 520 1492 536 1508
rect 136 1372 152 1388
rect 296 1372 312 1388
rect 8 1312 24 1328
rect 408 1372 424 1388
rect 232 1314 248 1328
rect 232 1312 248 1314
rect 104 1152 120 1168
rect 88 1132 104 1148
rect 8 1112 24 1128
rect 328 1106 344 1108
rect 328 1092 344 1106
rect 424 1152 440 1168
rect 424 1132 440 1148
rect 392 1092 408 1108
rect 136 972 152 988
rect 56 952 72 968
rect 8 912 24 928
rect 40 912 56 928
rect 408 1052 424 1068
rect 424 972 440 988
rect 408 952 424 968
rect 360 932 376 948
rect 152 912 168 928
rect 328 914 344 928
rect 328 912 344 914
rect 392 912 408 928
rect 488 1452 504 1468
rect 568 1812 584 1828
rect 616 1732 632 1748
rect 680 1732 696 1748
rect 600 1712 616 1728
rect 728 1752 744 1768
rect 925 2002 961 2018
rect 1016 1992 1032 2008
rect 1000 1972 1016 1988
rect 1000 1952 1016 1968
rect 904 1932 920 1948
rect 840 1912 856 1928
rect 888 1912 904 1928
rect 968 1912 984 1928
rect 920 1892 936 1908
rect 952 1832 968 1848
rect 808 1812 824 1828
rect 1192 2192 1208 2208
rect 1272 2212 1288 2228
rect 1416 2612 1432 2628
rect 1720 2852 1736 2868
rect 1672 2752 1688 2768
rect 1704 2752 1720 2768
rect 1640 2692 1656 2708
rect 1480 2632 1496 2648
rect 1624 2632 1640 2648
rect 1448 2592 1464 2608
rect 1656 2632 1672 2648
rect 1576 2572 1592 2588
rect 1608 2572 1624 2588
rect 1640 2572 1656 2588
rect 1480 2552 1496 2568
rect 1512 2552 1544 2568
rect 1400 2544 1416 2548
rect 1400 2532 1416 2544
rect 1464 2512 1480 2528
rect 1624 2552 1640 2568
rect 1496 2492 1512 2508
rect 1384 2312 1400 2328
rect 1384 2292 1400 2308
rect 1336 2252 1352 2268
rect 1416 2252 1432 2268
rect 1304 2192 1320 2208
rect 1304 2152 1320 2168
rect 1368 2152 1384 2168
rect 1144 2132 1160 2148
rect 1192 2132 1208 2148
rect 1128 2092 1144 2108
rect 1128 2032 1144 2048
rect 1128 1932 1144 1948
rect 1208 1892 1224 1908
rect 1064 1872 1080 1888
rect 1080 1872 1096 1888
rect 1000 1792 1016 1808
rect 824 1772 840 1788
rect 872 1772 888 1788
rect 1112 1812 1128 1828
rect 776 1732 792 1748
rect 808 1732 824 1748
rect 856 1744 872 1748
rect 856 1732 872 1744
rect 904 1732 920 1748
rect 952 1732 968 1748
rect 1048 1732 1064 1748
rect 568 1652 584 1668
rect 632 1652 648 1668
rect 744 1652 760 1668
rect 728 1632 744 1648
rect 600 1612 632 1628
rect 584 1572 600 1588
rect 616 1592 632 1608
rect 504 1392 520 1408
rect 552 1392 568 1408
rect 552 1352 568 1368
rect 584 1332 600 1348
rect 664 1572 680 1588
rect 872 1692 888 1708
rect 808 1672 824 1688
rect 936 1672 952 1688
rect 968 1632 984 1648
rect 925 1602 961 1618
rect 760 1552 776 1568
rect 888 1552 904 1568
rect 744 1512 760 1528
rect 616 1412 632 1428
rect 680 1492 696 1508
rect 744 1492 760 1508
rect 776 1492 792 1508
rect 808 1492 824 1508
rect 904 1492 920 1508
rect 648 1472 664 1488
rect 712 1472 728 1488
rect 824 1472 840 1488
rect 776 1452 792 1468
rect 808 1452 824 1468
rect 696 1432 712 1448
rect 744 1432 760 1448
rect 728 1412 744 1428
rect 632 1392 648 1408
rect 664 1332 680 1348
rect 696 1332 712 1348
rect 616 1312 632 1328
rect 600 1292 616 1308
rect 536 1232 552 1248
rect 552 1212 568 1228
rect 520 1152 536 1168
rect 456 892 472 908
rect 600 1152 616 1168
rect 648 1232 664 1248
rect 616 1072 632 1088
rect 616 952 632 968
rect 632 952 648 968
rect 680 1072 696 1088
rect 760 1412 776 1428
rect 792 1352 808 1368
rect 1032 1612 1048 1628
rect 1080 1592 1096 1608
rect 1048 1532 1064 1548
rect 1128 1744 1144 1748
rect 1128 1732 1144 1744
rect 1256 2092 1272 2108
rect 1288 2072 1304 2088
rect 1272 1932 1288 1948
rect 1400 2192 1416 2208
rect 1528 2432 1544 2448
rect 1464 2352 1480 2368
rect 1496 2352 1512 2368
rect 1608 2412 1624 2428
rect 1672 2452 1688 2468
rect 1528 2332 1544 2348
rect 1608 2332 1624 2348
rect 1656 2332 1672 2348
rect 1512 2292 1528 2308
rect 1560 2292 1576 2308
rect 1544 2272 1560 2288
rect 1448 2212 1480 2228
rect 1512 2212 1544 2228
rect 1512 2152 1528 2168
rect 1432 2132 1448 2148
rect 1480 2132 1496 2148
rect 1736 2832 1752 2848
rect 1976 3052 1992 3068
rect 2024 3052 2040 3068
rect 1880 3012 1896 3028
rect 1864 2972 1880 2988
rect 1784 2952 1800 2968
rect 1848 2952 1864 2968
rect 1933 3002 1969 3018
rect 1928 2972 1944 2988
rect 2056 2992 2072 3008
rect 2136 3232 2152 3248
rect 2120 3112 2136 3128
rect 2104 3072 2120 3088
rect 2168 3076 2200 3088
rect 2168 3072 2184 3076
rect 2184 3072 2200 3076
rect 2136 2992 2152 3008
rect 2200 2992 2216 3008
rect 2360 3272 2376 3288
rect 2392 3272 2408 3288
rect 2296 3252 2312 3268
rect 2360 3252 2376 3268
rect 2248 3112 2264 3128
rect 2232 3092 2248 3108
rect 2296 3092 2312 3108
rect 2328 3092 2344 3108
rect 2312 3072 2328 3088
rect 2504 3232 2520 3248
rect 2424 3172 2440 3188
rect 2472 3172 2488 3188
rect 2424 3112 2440 3128
rect 2376 3072 2392 3088
rect 2216 2972 2232 2988
rect 2200 2952 2216 2968
rect 2360 3012 2376 3028
rect 2392 3012 2408 3028
rect 2280 2952 2296 2968
rect 2312 2952 2328 2968
rect 2344 2952 2360 2968
rect 2504 3212 2520 3228
rect 2488 3132 2504 3148
rect 2520 3112 2536 3128
rect 2696 3492 2712 3508
rect 2664 3472 2680 3488
rect 2680 3392 2712 3408
rect 2744 3692 2760 3708
rect 2744 3592 2760 3608
rect 2776 3552 2792 3568
rect 2728 3532 2744 3548
rect 2792 3512 2808 3528
rect 2744 3492 2760 3508
rect 2728 3392 2744 3408
rect 2792 3472 2808 3488
rect 2808 3432 2824 3448
rect 2840 3672 2856 3688
rect 2888 3672 2904 3688
rect 2840 3592 2856 3608
rect 2856 3572 2872 3588
rect 2888 3572 2904 3588
rect 2872 3532 2888 3548
rect 2973 3602 3009 3618
rect 2856 3472 2872 3488
rect 2952 3472 2984 3488
rect 2920 3452 2936 3468
rect 2984 3452 3000 3468
rect 2824 3412 2840 3428
rect 2936 3412 2952 3428
rect 2872 3372 2888 3388
rect 2824 3352 2840 3368
rect 2712 3312 2728 3328
rect 2616 3292 2632 3308
rect 2648 3232 2664 3248
rect 2744 3232 2760 3248
rect 2712 3172 2728 3188
rect 2488 3092 2504 3108
rect 2600 3092 2616 3108
rect 2520 2992 2536 3008
rect 2504 2972 2520 2988
rect 2488 2952 2504 2968
rect 2472 2932 2488 2948
rect 1768 2912 1784 2928
rect 1832 2912 1848 2928
rect 1912 2912 1928 2928
rect 2008 2912 2024 2928
rect 2184 2912 2200 2928
rect 2264 2912 2280 2928
rect 2328 2912 2344 2928
rect 2472 2912 2488 2928
rect 1816 2892 1832 2908
rect 1864 2892 1880 2908
rect 1784 2832 1800 2848
rect 1720 2612 1736 2628
rect 1736 2552 1752 2568
rect 1816 2812 1832 2828
rect 1800 2752 1816 2768
rect 1912 2812 1928 2828
rect 2024 2792 2040 2808
rect 2024 2752 2040 2768
rect 2072 2712 2088 2728
rect 1912 2692 1928 2708
rect 1960 2692 1976 2708
rect 2040 2692 2056 2708
rect 2152 2792 2168 2808
rect 2184 2792 2200 2808
rect 2120 2752 2136 2768
rect 2088 2692 2104 2708
rect 2136 2692 2152 2708
rect 1800 2552 1816 2568
rect 1736 2532 1752 2548
rect 1752 2452 1768 2468
rect 1704 2392 1720 2408
rect 1688 2332 1704 2348
rect 1704 2292 1720 2308
rect 1752 2292 1768 2308
rect 1656 2272 1672 2288
rect 1768 2152 1784 2168
rect 1592 2132 1608 2148
rect 1688 2132 1704 2148
rect 1896 2632 1912 2648
rect 1976 2632 1992 2648
rect 2056 2632 2072 2648
rect 2120 2632 2136 2648
rect 1933 2602 1969 2618
rect 2104 2612 2120 2628
rect 2168 2612 2184 2628
rect 1832 2552 1848 2568
rect 1880 2552 1896 2568
rect 1976 2552 1992 2568
rect 2136 2552 2152 2568
rect 2248 2812 2264 2828
rect 2216 2672 2232 2688
rect 2280 2772 2296 2788
rect 2344 2812 2360 2828
rect 2392 2812 2408 2828
rect 2312 2752 2328 2768
rect 2392 2772 2408 2788
rect 2472 2772 2488 2788
rect 2328 2692 2344 2708
rect 2200 2552 2216 2568
rect 2232 2552 2248 2568
rect 1912 2532 1928 2548
rect 1976 2532 1992 2548
rect 2040 2532 2056 2548
rect 2184 2532 2200 2548
rect 2200 2532 2216 2548
rect 1864 2512 1880 2528
rect 1912 2472 1928 2488
rect 2024 2472 2040 2488
rect 1848 2372 1864 2388
rect 1880 2312 1896 2328
rect 1832 2292 1848 2308
rect 1832 2272 1848 2288
rect 1832 2152 1848 2168
rect 1896 2292 1912 2308
rect 2456 2672 2472 2688
rect 2488 2692 2504 2708
rect 2568 3032 2584 3048
rect 2552 2952 2568 2968
rect 2584 2952 2600 2968
rect 2648 2972 2664 2988
rect 2856 3272 2872 3288
rect 2840 3192 2856 3208
rect 2840 3132 2856 3148
rect 2808 3112 2824 3128
rect 2904 3232 2920 3248
rect 2904 3212 2920 3228
rect 2968 3392 2984 3408
rect 3080 3792 3096 3808
rect 3304 4012 3320 4028
rect 3400 3952 3416 3968
rect 3192 3932 3208 3948
rect 3240 3932 3256 3948
rect 3320 3932 3336 3948
rect 3384 3932 3400 3948
rect 3160 3892 3176 3908
rect 3144 3792 3160 3808
rect 3288 3892 3304 3908
rect 3304 3892 3320 3908
rect 3192 3872 3208 3888
rect 3176 3812 3192 3828
rect 3208 3792 3224 3808
rect 3272 3712 3288 3728
rect 3064 3612 3080 3628
rect 3080 3512 3096 3528
rect 3112 3492 3128 3508
rect 3032 3432 3048 3448
rect 3112 3432 3128 3448
rect 3272 3592 3288 3608
rect 3208 3552 3240 3568
rect 3176 3492 3192 3508
rect 3256 3492 3272 3508
rect 3240 3472 3256 3488
rect 3160 3432 3176 3448
rect 3112 3352 3128 3368
rect 3016 3332 3048 3348
rect 3192 3412 3208 3428
rect 3320 3872 3336 3888
rect 3320 3852 3336 3868
rect 3384 3872 3400 3888
rect 3336 3812 3352 3828
rect 3368 3812 3384 3828
rect 3320 3752 3336 3768
rect 3304 3732 3320 3748
rect 3304 3692 3320 3708
rect 3288 3512 3304 3528
rect 3576 4012 3592 4028
rect 3576 3992 3592 4008
rect 3608 3992 3624 4008
rect 3608 3972 3624 3988
rect 3432 3892 3448 3908
rect 3496 3892 3512 3908
rect 3576 3892 3592 3908
rect 3448 3872 3464 3888
rect 3416 3752 3432 3768
rect 3416 3732 3432 3748
rect 3432 3712 3448 3728
rect 3368 3692 3384 3708
rect 3352 3632 3368 3648
rect 3352 3572 3384 3588
rect 3304 3472 3320 3488
rect 3320 3472 3336 3488
rect 3208 3352 3224 3368
rect 3272 3352 3288 3368
rect 3368 3352 3384 3368
rect 3144 3312 3160 3328
rect 2973 3202 3009 3218
rect 3016 3212 3032 3228
rect 2984 3152 3000 3168
rect 2696 3052 2712 3068
rect 2744 3052 2760 3068
rect 2712 2992 2728 3008
rect 2792 3012 2808 3028
rect 2776 2972 2792 2988
rect 2680 2952 2696 2968
rect 2760 2952 2776 2968
rect 2776 2952 2792 2968
rect 2648 2932 2664 2948
rect 2712 2932 2728 2948
rect 2664 2892 2680 2908
rect 2600 2852 2616 2868
rect 2536 2832 2552 2848
rect 2552 2832 2568 2848
rect 2792 2892 2808 2908
rect 2728 2832 2744 2848
rect 2776 2832 2792 2848
rect 2744 2792 2760 2808
rect 2568 2752 2584 2768
rect 2680 2752 2696 2768
rect 2552 2732 2568 2748
rect 2536 2692 2552 2708
rect 2520 2672 2536 2688
rect 2712 2692 2728 2708
rect 2664 2672 2680 2688
rect 2728 2672 2744 2688
rect 2424 2632 2440 2648
rect 2664 2632 2680 2648
rect 2328 2572 2344 2588
rect 2360 2572 2376 2588
rect 2056 2512 2072 2528
rect 2088 2512 2104 2528
rect 2168 2512 2184 2528
rect 2264 2512 2280 2528
rect 2072 2492 2084 2508
rect 2084 2492 2088 2508
rect 2088 2492 2104 2508
rect 2136 2492 2152 2508
rect 2168 2492 2184 2508
rect 2152 2392 2168 2408
rect 2040 2372 2056 2388
rect 1928 2312 1944 2328
rect 2008 2272 2024 2288
rect 1928 2232 1944 2248
rect 1933 2202 1969 2218
rect 1912 2172 1928 2188
rect 1912 2152 1928 2168
rect 1816 2132 1832 2148
rect 1576 2112 1592 2128
rect 1688 2112 1720 2128
rect 1896 2112 1912 2128
rect 1544 2072 1560 2088
rect 1320 2012 1336 2028
rect 1384 2012 1400 2028
rect 1432 1892 1448 1908
rect 1352 1872 1368 1888
rect 1560 2052 1576 2068
rect 1640 2092 1656 2108
rect 1624 2032 1640 2048
rect 1576 2012 1592 2028
rect 1576 1892 1592 1908
rect 1624 1892 1640 1908
rect 1672 1892 1688 1908
rect 1416 1852 1432 1868
rect 1368 1812 1384 1828
rect 1288 1772 1304 1788
rect 1320 1772 1336 1788
rect 1592 1832 1608 1848
rect 1544 1772 1560 1788
rect 1176 1752 1192 1768
rect 1528 1752 1544 1768
rect 1608 1792 1624 1808
rect 1608 1752 1624 1768
rect 1176 1732 1192 1748
rect 1240 1732 1256 1748
rect 1320 1744 1336 1748
rect 1320 1732 1336 1744
rect 1528 1732 1544 1748
rect 1592 1732 1608 1748
rect 1176 1712 1192 1728
rect 1192 1692 1208 1708
rect 1224 1692 1240 1708
rect 1160 1632 1176 1648
rect 1224 1592 1240 1608
rect 1112 1572 1128 1588
rect 1208 1572 1224 1588
rect 1256 1712 1272 1728
rect 1400 1712 1416 1728
rect 1432 1712 1448 1728
rect 1480 1712 1496 1728
rect 1560 1712 1576 1728
rect 1288 1692 1304 1708
rect 1240 1572 1256 1588
rect 1272 1552 1288 1568
rect 1160 1532 1176 1548
rect 1128 1512 1144 1528
rect 984 1492 1000 1508
rect 1064 1492 1080 1508
rect 1096 1492 1112 1508
rect 1240 1492 1256 1508
rect 1080 1472 1096 1488
rect 1192 1472 1208 1488
rect 936 1452 952 1468
rect 1016 1412 1048 1428
rect 1096 1412 1112 1428
rect 840 1392 856 1408
rect 1048 1372 1064 1388
rect 792 1332 808 1348
rect 824 1332 840 1348
rect 872 1332 888 1348
rect 840 1312 856 1328
rect 792 1292 808 1308
rect 776 1212 792 1228
rect 808 1232 824 1248
rect 792 1132 808 1148
rect 760 1112 776 1128
rect 904 1312 920 1328
rect 1064 1352 1080 1368
rect 1224 1432 1240 1448
rect 1192 1372 1208 1388
rect 1176 1344 1192 1348
rect 1176 1332 1192 1344
rect 1224 1332 1240 1348
rect 1352 1692 1368 1708
rect 1416 1692 1432 1708
rect 1320 1672 1336 1688
rect 1304 1592 1320 1608
rect 1336 1532 1352 1548
rect 1288 1512 1304 1528
rect 1304 1492 1320 1508
rect 1288 1472 1304 1488
rect 1256 1392 1272 1408
rect 1192 1312 1208 1328
rect 968 1292 984 1308
rect 1208 1292 1224 1308
rect 925 1202 961 1218
rect 1016 1252 1032 1268
rect 920 1152 936 1168
rect 968 1152 984 1168
rect 888 1132 904 1148
rect 728 1092 744 1108
rect 712 1072 728 1088
rect 824 1112 840 1128
rect 856 1112 872 1128
rect 904 1092 920 1108
rect 696 1052 712 1068
rect 728 1052 744 1068
rect 664 1012 680 1028
rect 664 992 680 1008
rect 664 952 680 968
rect 584 932 600 948
rect 552 914 568 928
rect 552 912 568 914
rect 616 912 632 928
rect 88 732 104 748
rect 328 732 344 748
rect 8 712 24 728
rect 728 1012 744 1028
rect 808 1012 824 1028
rect 856 1012 872 1028
rect 840 912 856 928
rect 664 852 680 868
rect 696 852 712 868
rect 312 712 328 728
rect 648 712 664 728
rect 232 706 248 708
rect 232 692 248 706
rect 296 692 312 708
rect 8 512 24 528
rect 808 832 824 848
rect 456 706 472 708
rect 456 692 472 706
rect 552 692 568 708
rect 568 692 584 708
rect 648 692 664 708
rect 216 532 232 548
rect 312 512 328 528
rect 424 492 440 508
rect 264 472 280 488
rect 8 312 24 328
rect 216 432 232 448
rect 296 432 312 448
rect 584 672 600 688
rect 536 652 552 668
rect 584 652 600 668
rect 824 712 840 728
rect 840 692 856 708
rect 776 672 792 688
rect 744 652 760 668
rect 632 632 648 648
rect 712 632 728 648
rect 632 592 648 608
rect 536 572 552 588
rect 600 572 616 588
rect 568 552 584 568
rect 616 552 632 568
rect 584 532 600 548
rect 600 532 616 548
rect 632 544 648 548
rect 632 532 648 544
rect 840 592 856 608
rect 808 552 824 568
rect 872 972 888 988
rect 888 952 904 968
rect 1000 1152 1016 1168
rect 1240 1272 1256 1288
rect 1208 1172 1224 1188
rect 1304 1332 1320 1348
rect 1464 1652 1480 1668
rect 1464 1632 1480 1648
rect 1496 1632 1512 1648
rect 1512 1612 1528 1628
rect 1592 1572 1608 1588
rect 1544 1532 1560 1548
rect 1528 1512 1544 1528
rect 1432 1492 1448 1508
rect 1368 1476 1384 1488
rect 1368 1472 1384 1476
rect 1432 1472 1448 1488
rect 1368 1392 1384 1408
rect 1272 1272 1288 1288
rect 1256 1212 1272 1228
rect 1080 1112 1096 1128
rect 936 1072 952 1088
rect 984 1072 1000 1088
rect 1032 1052 1048 1068
rect 984 1032 1000 1048
rect 1128 1092 1144 1108
rect 1256 1132 1272 1148
rect 1288 1132 1304 1148
rect 1320 1132 1336 1148
rect 1304 1092 1320 1108
rect 1480 1392 1496 1408
rect 1448 1332 1464 1348
rect 1480 1312 1496 1328
rect 1512 1312 1528 1328
rect 2008 2112 2024 2128
rect 1848 2072 1864 2088
rect 1912 2072 1928 2088
rect 1832 2052 1848 2068
rect 1784 2032 1800 2048
rect 1704 1952 1720 1968
rect 1752 1952 1768 1968
rect 1720 1932 1736 1948
rect 1736 1912 1752 1928
rect 1720 1652 1736 1668
rect 1672 1572 1688 1588
rect 1656 1532 1672 1548
rect 1624 1512 1640 1528
rect 1640 1512 1656 1528
rect 1608 1472 1624 1488
rect 1560 1432 1576 1448
rect 1624 1432 1640 1448
rect 1560 1392 1576 1408
rect 1544 1332 1560 1348
rect 1640 1392 1656 1408
rect 1752 1892 1768 1908
rect 1768 1852 1784 1868
rect 1768 1732 1784 1748
rect 1752 1632 1768 1648
rect 1992 2032 2008 2048
rect 1864 1992 1880 2008
rect 1816 1932 1832 1948
rect 1896 1932 1912 1948
rect 1832 1912 1848 1928
rect 1800 1732 1816 1748
rect 1800 1592 1816 1608
rect 2088 2292 2104 2308
rect 2104 2272 2120 2288
rect 2136 2252 2152 2268
rect 2120 2192 2136 2208
rect 2136 2172 2152 2188
rect 2104 2152 2120 2168
rect 2072 2132 2088 2148
rect 2024 2092 2056 2108
rect 2040 1952 2056 1968
rect 2088 1952 2104 1968
rect 2040 1932 2056 1948
rect 2008 1912 2024 1928
rect 1880 1852 1896 1868
rect 1912 1852 1928 1868
rect 1944 1852 1960 1868
rect 1933 1802 1969 1818
rect 2056 1812 2072 1828
rect 2008 1792 2024 1808
rect 2024 1772 2040 1788
rect 2072 1772 2088 1788
rect 2040 1752 2056 1768
rect 2072 1752 2088 1768
rect 1912 1744 1928 1748
rect 1912 1732 1928 1744
rect 1832 1672 1848 1688
rect 1816 1572 1832 1588
rect 1752 1552 1768 1568
rect 2136 2132 2152 2148
rect 2312 2552 2328 2568
rect 2296 2532 2312 2548
rect 2392 2552 2408 2568
rect 2408 2552 2424 2568
rect 2280 2432 2296 2448
rect 2248 2352 2264 2368
rect 2216 2332 2232 2348
rect 2248 2292 2264 2308
rect 2264 2272 2280 2288
rect 2200 2252 2216 2268
rect 2264 2252 2280 2268
rect 2200 2232 2216 2248
rect 2200 2212 2216 2228
rect 2248 2132 2264 2148
rect 2152 2072 2184 2088
rect 2136 2012 2152 2028
rect 2216 2052 2232 2068
rect 2168 2032 2184 2048
rect 2184 2012 2200 2028
rect 2184 1992 2200 2008
rect 2152 1852 2168 1868
rect 2168 1772 2184 1788
rect 2040 1672 2056 1688
rect 2040 1632 2056 1648
rect 1880 1532 1896 1548
rect 2104 1692 2120 1708
rect 2088 1572 2104 1588
rect 2072 1552 2088 1568
rect 1992 1512 2008 1528
rect 2040 1512 2056 1528
rect 1912 1492 1928 1508
rect 1976 1492 1992 1508
rect 1736 1472 1752 1488
rect 1848 1472 1864 1488
rect 1720 1452 1736 1468
rect 1768 1452 1784 1468
rect 1816 1452 1832 1468
rect 1832 1452 1848 1468
rect 1832 1432 1848 1448
rect 1896 1432 1912 1448
rect 1720 1412 1736 1428
rect 1704 1372 1720 1388
rect 1656 1332 1672 1348
rect 1672 1332 1688 1348
rect 1576 1312 1592 1328
rect 1608 1312 1624 1328
rect 1528 1292 1544 1308
rect 1464 1272 1480 1288
rect 1528 1272 1544 1288
rect 1544 1252 1560 1268
rect 1416 1112 1432 1128
rect 1560 1172 1576 1188
rect 1352 1092 1368 1108
rect 1480 1092 1496 1108
rect 1544 1092 1560 1108
rect 1656 1112 1672 1128
rect 1176 1072 1192 1088
rect 1336 1072 1352 1088
rect 1352 1072 1368 1088
rect 1768 1332 1784 1348
rect 1848 1332 1864 1348
rect 1688 1312 1704 1328
rect 1160 1032 1176 1048
rect 1096 992 1112 1008
rect 1096 972 1112 988
rect 968 952 984 968
rect 920 932 936 948
rect 1000 932 1016 948
rect 904 912 920 928
rect 925 802 961 818
rect 872 772 888 788
rect 1128 912 1144 928
rect 1208 1052 1224 1068
rect 1352 1052 1368 1068
rect 1400 1052 1416 1068
rect 1496 1052 1512 1068
rect 1400 1032 1416 1048
rect 1224 1012 1240 1028
rect 1208 912 1224 928
rect 1256 952 1288 968
rect 1304 952 1320 968
rect 1352 952 1368 968
rect 1272 932 1288 948
rect 1064 892 1080 908
rect 1144 892 1160 908
rect 1176 892 1192 908
rect 1224 892 1240 908
rect 1272 892 1288 908
rect 1048 812 1064 828
rect 952 752 968 768
rect 1000 752 1016 768
rect 904 652 920 668
rect 888 632 904 648
rect 904 572 920 588
rect 696 512 712 528
rect 808 512 824 528
rect 552 492 568 508
rect 744 492 760 508
rect 488 472 504 488
rect 568 472 584 488
rect 456 432 472 448
rect 520 432 536 448
rect 792 372 808 388
rect 744 312 760 328
rect 664 306 680 308
rect 664 292 680 306
rect 728 292 744 308
rect 8 112 24 128
rect 536 232 552 248
rect 504 172 520 188
rect 968 692 984 708
rect 1080 872 1096 888
rect 1112 872 1128 888
rect 1000 672 1016 688
rect 1064 672 1080 688
rect 1000 652 1016 668
rect 1016 632 1032 648
rect 1000 612 1016 628
rect 1256 852 1272 868
rect 1224 832 1240 848
rect 1128 812 1144 828
rect 1176 812 1192 828
rect 1096 732 1112 748
rect 1144 712 1160 728
rect 1192 732 1208 748
rect 1224 732 1240 748
rect 1240 712 1256 728
rect 1256 692 1272 708
rect 1288 872 1304 888
rect 1304 852 1320 868
rect 1304 812 1320 828
rect 1352 812 1368 828
rect 1320 732 1336 748
rect 1336 712 1352 728
rect 1400 912 1416 928
rect 1432 912 1448 928
rect 1368 732 1384 748
rect 1384 732 1400 748
rect 1416 732 1432 748
rect 1432 712 1448 728
rect 1400 692 1416 708
rect 1432 692 1448 708
rect 1112 672 1128 688
rect 1208 652 1224 668
rect 1032 572 1048 588
rect 1464 1012 1480 1028
rect 1480 972 1496 988
rect 1480 692 1496 708
rect 1480 672 1496 688
rect 1608 1032 1624 1048
rect 1576 992 1592 1008
rect 1560 972 1576 988
rect 1544 932 1560 948
rect 1512 912 1528 928
rect 1608 912 1624 928
rect 1528 752 1544 768
rect 1544 732 1560 748
rect 1592 712 1608 728
rect 1448 652 1464 668
rect 1496 652 1512 668
rect 1512 612 1528 628
rect 1560 612 1576 628
rect 1560 572 1576 588
rect 952 552 968 568
rect 1160 552 1176 568
rect 1192 552 1208 568
rect 1256 552 1272 568
rect 1272 552 1304 568
rect 1512 552 1528 568
rect 1544 552 1560 568
rect 968 532 984 548
rect 1016 532 1032 548
rect 1128 532 1160 548
rect 1320 532 1336 548
rect 1432 532 1448 548
rect 1016 512 1032 528
rect 984 472 1000 488
rect 1048 472 1064 488
rect 856 452 872 468
rect 968 452 984 468
rect 1048 432 1064 448
rect 925 402 961 418
rect 1064 372 1080 388
rect 984 292 1000 308
rect 1096 292 1112 308
rect 1128 292 1144 308
rect 1000 272 1016 288
rect 1112 272 1128 288
rect 808 252 824 268
rect 632 232 648 248
rect 696 232 712 248
rect 744 232 760 248
rect 232 112 248 128
rect 296 112 312 128
rect 936 232 952 248
rect 1000 232 1016 248
rect 872 192 888 208
rect 840 172 856 188
rect 568 114 584 128
rect 568 112 584 114
rect 856 112 872 128
rect 776 92 792 108
rect 840 92 856 108
rect 200 12 216 28
rect 232 12 248 28
rect 925 2 961 18
rect 984 12 1000 28
rect 1016 12 1032 28
rect 1224 492 1256 508
rect 1432 492 1448 508
rect 1320 472 1336 488
rect 1160 292 1176 308
rect 1384 412 1400 428
rect 1304 392 1320 408
rect 1224 332 1240 348
rect 1576 532 1592 548
rect 1576 492 1608 508
rect 1496 452 1512 468
rect 1576 452 1592 468
rect 1528 412 1544 428
rect 1304 312 1320 328
rect 1576 352 1592 368
rect 1352 292 1368 308
rect 1464 292 1480 308
rect 1496 292 1512 308
rect 1176 272 1192 288
rect 1480 272 1496 288
rect 1240 232 1256 248
rect 1304 232 1320 248
rect 1272 172 1288 188
rect 1592 272 1608 288
rect 1544 252 1560 268
rect 1576 252 1592 268
rect 1528 192 1544 208
rect 1416 152 1432 168
rect 1400 132 1416 148
rect 1448 132 1464 148
rect 1512 132 1528 148
rect 1240 114 1256 128
rect 1240 112 1256 114
rect 1400 112 1416 128
rect 1480 92 1496 108
rect 1176 12 1192 28
rect 1224 12 1240 28
rect 1688 1032 1704 1048
rect 1640 932 1656 948
rect 1672 932 1688 948
rect 1800 1312 1816 1328
rect 1864 1312 1880 1328
rect 1752 1252 1768 1268
rect 1832 1112 1844 1128
rect 1844 1112 1848 1128
rect 1848 1112 1864 1128
rect 1720 1072 1736 1088
rect 1800 1072 1816 1088
rect 1752 1052 1768 1068
rect 1720 972 1736 988
rect 1768 972 1784 988
rect 1816 1012 1832 1028
rect 1896 1272 1912 1288
rect 1933 1402 1969 1418
rect 2024 1432 2040 1448
rect 2008 1372 2024 1388
rect 1928 1332 1944 1348
rect 2040 1332 2056 1348
rect 2120 1612 2136 1628
rect 2216 1972 2232 1988
rect 2360 2412 2376 2428
rect 2344 2392 2360 2408
rect 2312 2272 2328 2288
rect 2616 2612 2632 2628
rect 2472 2592 2488 2608
rect 2440 2552 2456 2568
rect 2504 2552 2520 2568
rect 2456 2532 2472 2548
rect 2536 2532 2552 2548
rect 2680 2612 2696 2628
rect 2632 2532 2648 2548
rect 2664 2532 2680 2548
rect 2520 2512 2536 2528
rect 2504 2332 2520 2348
rect 2648 2492 2664 2508
rect 2584 2452 2600 2468
rect 2568 2432 2584 2448
rect 2760 2552 2776 2568
rect 2760 2532 2776 2548
rect 2664 2452 2680 2468
rect 2664 2432 2680 2448
rect 2776 2392 2792 2408
rect 2712 2372 2728 2388
rect 2712 2352 2728 2368
rect 2728 2312 2744 2328
rect 2776 2312 2792 2328
rect 2888 3032 2904 3048
rect 2920 3032 2936 3048
rect 2904 3012 2920 3028
rect 2856 2992 2872 3008
rect 2888 2952 2904 2968
rect 2840 2932 2856 2948
rect 2936 2992 2952 3008
rect 3016 2952 3032 2968
rect 2920 2932 2936 2948
rect 2936 2932 2952 2948
rect 2968 2852 2984 2868
rect 2973 2802 3009 2818
rect 2904 2772 2920 2788
rect 3016 2772 3032 2788
rect 2824 2752 2840 2768
rect 2888 2692 2904 2708
rect 2840 2672 2856 2688
rect 2888 2552 2904 2568
rect 2872 2532 2888 2548
rect 2872 2352 2888 2368
rect 2456 2292 2472 2308
rect 2504 2292 2520 2308
rect 2392 2252 2408 2268
rect 2392 2232 2408 2248
rect 2456 2232 2472 2248
rect 2296 1912 2312 1928
rect 2248 1892 2264 1908
rect 2264 1892 2280 1908
rect 2296 1892 2312 1908
rect 2200 1872 2216 1888
rect 2280 1872 2296 1888
rect 2232 1852 2248 1868
rect 2280 1752 2296 1768
rect 2200 1712 2216 1728
rect 2264 1732 2280 1748
rect 2232 1672 2248 1688
rect 2376 2212 2392 2228
rect 2376 2152 2392 2168
rect 2408 2132 2424 2148
rect 2456 2132 2472 2148
rect 2344 2012 2360 2028
rect 2344 1972 2360 1988
rect 2328 1892 2344 1908
rect 2408 2072 2424 2088
rect 2456 2072 2472 2088
rect 2440 2012 2456 2028
rect 2440 1952 2456 1968
rect 2424 1932 2440 1948
rect 2376 1912 2392 1928
rect 2456 1872 2472 1888
rect 2456 1852 2472 1868
rect 2424 1772 2440 1788
rect 2568 2272 2584 2288
rect 2520 2252 2536 2268
rect 2744 2252 2760 2268
rect 2648 2212 2664 2228
rect 2600 2152 2616 2168
rect 2536 2132 2552 2148
rect 2488 2112 2504 2128
rect 2504 2092 2520 2108
rect 2632 2172 2648 2188
rect 2696 2172 2712 2188
rect 2760 2172 2776 2188
rect 2696 2132 2712 2148
rect 2728 2132 2744 2148
rect 2552 2112 2568 2128
rect 2648 2112 2664 2128
rect 2568 2012 2584 2028
rect 2632 2072 2648 2088
rect 2616 1952 2632 1968
rect 2648 1932 2664 1948
rect 2584 1892 2600 1908
rect 2648 1892 2664 1908
rect 2824 2312 2840 2328
rect 2808 2276 2824 2288
rect 2808 2272 2824 2276
rect 2840 2272 2856 2288
rect 2856 2272 2872 2288
rect 2824 2152 2840 2168
rect 2792 2112 2808 2128
rect 2808 2112 2824 2128
rect 2936 2712 2952 2728
rect 3016 2712 3032 2728
rect 2920 2652 2936 2668
rect 2920 2592 2936 2608
rect 2952 2592 2984 2608
rect 2936 2332 2952 2348
rect 2904 2272 2920 2288
rect 3128 3272 3144 3288
rect 3096 3232 3112 3248
rect 3160 3232 3176 3248
rect 3192 3232 3208 3248
rect 3176 3212 3192 3228
rect 3128 3192 3144 3208
rect 3080 3092 3096 3108
rect 3048 3072 3064 3088
rect 3176 3172 3192 3188
rect 3176 3132 3192 3148
rect 3144 3092 3160 3108
rect 3160 3072 3176 3088
rect 3128 3052 3144 3068
rect 3048 3032 3064 3048
rect 3112 3032 3128 3048
rect 3112 2952 3128 2968
rect 3144 3032 3160 3048
rect 3048 2772 3064 2788
rect 3032 2612 3048 2628
rect 3128 2752 3144 2768
rect 3080 2732 3096 2748
rect 3080 2712 3096 2728
rect 3064 2692 3080 2708
rect 3128 2692 3144 2708
rect 3208 3092 3224 3108
rect 3240 3112 3256 3128
rect 3256 3092 3272 3108
rect 3224 3032 3240 3048
rect 3368 3312 3384 3328
rect 3464 3612 3480 3628
rect 3544 3872 3560 3888
rect 3528 3812 3544 3828
rect 3592 3852 3608 3868
rect 3544 3732 3560 3748
rect 3496 3712 3528 3728
rect 3528 3692 3544 3708
rect 3592 3672 3608 3688
rect 3592 3652 3608 3668
rect 3576 3632 3608 3648
rect 3560 3612 3576 3628
rect 3416 3472 3432 3488
rect 3480 3512 3496 3528
rect 3496 3472 3512 3488
rect 3416 3452 3432 3468
rect 3464 3452 3480 3468
rect 3512 3452 3528 3468
rect 3592 3452 3608 3468
rect 3432 3412 3448 3428
rect 3480 3412 3496 3428
rect 3528 3412 3544 3428
rect 3560 3412 3576 3428
rect 3592 3352 3608 3368
rect 3448 3332 3464 3348
rect 3560 3312 3592 3328
rect 3384 3192 3416 3208
rect 3496 3272 3512 3288
rect 3448 3252 3464 3268
rect 3448 3212 3464 3228
rect 3416 3112 3432 3128
rect 3336 3092 3352 3108
rect 3400 3092 3416 3108
rect 3480 3152 3496 3168
rect 3448 3092 3464 3108
rect 3352 3072 3368 3088
rect 3432 3072 3448 3088
rect 3272 3012 3288 3028
rect 3208 2952 3224 2968
rect 3192 2932 3208 2948
rect 3256 2932 3272 2948
rect 3400 2932 3416 2948
rect 3176 2912 3192 2928
rect 3192 2912 3208 2928
rect 3176 2792 3192 2808
rect 3160 2712 3176 2728
rect 3416 2912 3432 2928
rect 3384 2892 3400 2908
rect 3368 2872 3384 2888
rect 3320 2772 3336 2788
rect 3336 2732 3352 2748
rect 3256 2712 3272 2728
rect 3240 2692 3256 2708
rect 3352 2692 3368 2708
rect 3144 2672 3160 2688
rect 3160 2672 3176 2688
rect 3240 2672 3256 2688
rect 3192 2612 3208 2628
rect 3096 2552 3128 2568
rect 3160 2552 3176 2568
rect 3048 2532 3064 2548
rect 3160 2532 3176 2548
rect 3096 2512 3112 2528
rect 3128 2492 3144 2508
rect 2973 2402 3009 2418
rect 3048 2412 3064 2428
rect 3192 2512 3208 2528
rect 3144 2452 3160 2468
rect 3128 2412 3144 2428
rect 3160 2412 3176 2428
rect 3112 2312 3128 2328
rect 3032 2292 3064 2308
rect 3112 2292 3128 2308
rect 3144 2292 3160 2308
rect 3064 2272 3080 2288
rect 2888 2252 2904 2268
rect 2920 2252 2936 2268
rect 2872 2232 2888 2248
rect 2952 2232 2968 2248
rect 3128 2232 3144 2248
rect 2904 2212 2936 2228
rect 2888 2192 2904 2208
rect 2920 2172 2936 2188
rect 2872 2132 2888 2148
rect 2792 1932 2808 1948
rect 2760 1912 2776 1928
rect 2504 1872 2520 1888
rect 2568 1872 2584 1888
rect 2680 1872 2696 1888
rect 2552 1792 2568 1808
rect 2632 1792 2664 1808
rect 2488 1772 2504 1788
rect 2616 1772 2632 1788
rect 2520 1752 2536 1768
rect 2312 1732 2328 1748
rect 2472 1732 2488 1748
rect 2552 1732 2568 1748
rect 2264 1572 2280 1588
rect 2280 1572 2296 1588
rect 2232 1532 2248 1548
rect 2200 1512 2216 1528
rect 2152 1432 2168 1448
rect 2216 1452 2232 1468
rect 2232 1452 2248 1468
rect 2168 1412 2184 1428
rect 2232 1412 2248 1428
rect 2216 1372 2232 1388
rect 2376 1632 2392 1648
rect 2664 1732 2680 1748
rect 2424 1712 2440 1728
rect 2488 1712 2504 1728
rect 2600 1712 2616 1728
rect 2664 1712 2680 1728
rect 2696 1712 2712 1728
rect 2584 1692 2600 1708
rect 2680 1692 2696 1708
rect 2520 1652 2536 1668
rect 2440 1632 2456 1648
rect 2584 1672 2600 1688
rect 2552 1632 2568 1648
rect 2504 1612 2536 1628
rect 2440 1592 2456 1608
rect 2360 1552 2376 1568
rect 2488 1552 2504 1568
rect 2552 1592 2568 1608
rect 2568 1552 2584 1568
rect 2312 1512 2328 1528
rect 2392 1512 2424 1528
rect 2456 1512 2472 1528
rect 2328 1492 2344 1508
rect 2616 1632 2632 1648
rect 2824 1992 2840 2008
rect 2840 1932 2856 1948
rect 2824 1872 2840 1888
rect 3064 2172 3080 2188
rect 3080 2172 3096 2188
rect 3048 2152 3064 2168
rect 2936 2132 2952 2148
rect 3096 2132 3112 2148
rect 3000 2112 3016 2128
rect 3128 2112 3144 2128
rect 2888 2072 2904 2088
rect 2973 2002 3009 2018
rect 2888 1932 2904 1948
rect 3000 1912 3016 1928
rect 2984 1892 3000 1908
rect 2840 1852 2856 1868
rect 2936 1872 2952 1888
rect 2760 1832 2776 1848
rect 2792 1832 2808 1848
rect 2888 1832 2920 1848
rect 2968 1792 2984 1808
rect 2904 1772 2920 1788
rect 2856 1732 2872 1748
rect 2936 1752 2952 1768
rect 2712 1592 2728 1608
rect 2664 1572 2680 1588
rect 2696 1572 2712 1588
rect 2824 1692 2828 1708
rect 2828 1692 2840 1708
rect 2808 1632 2824 1648
rect 2760 1572 2776 1588
rect 2600 1512 2616 1528
rect 2648 1512 2660 1528
rect 2660 1512 2664 1528
rect 2728 1512 2744 1528
rect 2584 1492 2600 1508
rect 2632 1492 2648 1508
rect 2376 1452 2392 1468
rect 2296 1412 2312 1428
rect 2344 1412 2360 1428
rect 2472 1472 2488 1488
rect 2504 1472 2520 1488
rect 2312 1392 2328 1408
rect 2392 1392 2408 1408
rect 2424 1392 2440 1408
rect 2424 1372 2440 1388
rect 2280 1352 2296 1368
rect 2344 1352 2360 1368
rect 2408 1352 2424 1368
rect 2280 1332 2296 1348
rect 2360 1332 2376 1348
rect 2392 1332 2408 1348
rect 2072 1312 2088 1328
rect 2328 1312 2344 1328
rect 2392 1312 2408 1328
rect 2456 1312 2472 1328
rect 2008 1152 2040 1168
rect 2056 1152 2072 1168
rect 1960 1112 1976 1128
rect 1976 1092 1992 1108
rect 1864 1072 1880 1088
rect 2008 1072 2024 1088
rect 1912 1032 1928 1048
rect 1848 992 1864 1008
rect 1933 1002 1969 1018
rect 1832 972 1848 988
rect 1928 972 1944 988
rect 1752 932 1768 948
rect 1832 932 1848 948
rect 1896 932 1928 948
rect 1704 892 1720 908
rect 1960 932 1976 948
rect 2008 944 2024 948
rect 2008 932 2024 944
rect 1944 892 1960 908
rect 1656 872 1672 888
rect 1688 872 1704 888
rect 1720 872 1736 888
rect 1848 872 1864 888
rect 1912 872 1928 888
rect 1624 852 1640 868
rect 1768 852 1784 868
rect 1624 832 1640 848
rect 1672 832 1688 848
rect 1704 792 1720 808
rect 1736 712 1752 728
rect 1720 692 1736 708
rect 1752 692 1768 708
rect 1736 672 1752 688
rect 1656 652 1672 668
rect 1720 652 1736 668
rect 1672 632 1688 648
rect 1640 612 1656 628
rect 1672 572 1688 588
rect 1624 552 1640 568
rect 1736 572 1752 588
rect 1656 532 1672 548
rect 1704 532 1720 548
rect 1880 812 1896 828
rect 1816 792 1832 808
rect 1784 732 1800 748
rect 1848 732 1864 748
rect 1816 712 1832 728
rect 1864 712 1880 728
rect 1896 692 1912 708
rect 1848 672 1864 688
rect 1896 672 1912 688
rect 1944 672 1960 688
rect 1896 652 1912 668
rect 1896 612 1912 628
rect 1933 602 1969 618
rect 1896 552 1912 568
rect 1912 552 1928 568
rect 1944 552 1960 568
rect 1624 492 1640 508
rect 1640 392 1656 408
rect 1736 492 1752 508
rect 1688 452 1704 468
rect 1672 392 1688 408
rect 1656 372 1672 388
rect 1848 532 1864 548
rect 1896 532 1912 548
rect 1928 532 1944 548
rect 1768 492 1784 508
rect 1800 492 1816 508
rect 1880 492 1896 508
rect 1752 452 1768 468
rect 1800 452 1816 468
rect 1816 452 1832 468
rect 1848 452 1864 468
rect 1768 392 1784 408
rect 1752 372 1768 388
rect 1704 312 1720 328
rect 1720 292 1736 308
rect 1784 372 1800 388
rect 1736 272 1752 288
rect 1624 232 1640 248
rect 1688 32 1704 48
rect 1848 292 1864 308
rect 1800 272 1816 288
rect 1848 272 1864 288
rect 1784 112 1800 128
rect 1832 112 1848 128
rect 1816 32 1832 48
rect 1736 12 1768 28
rect 1816 12 1832 28
rect 1944 452 1960 468
rect 1912 372 1928 388
rect 2168 1152 2184 1168
rect 2424 1292 2440 1308
rect 2120 1112 2136 1128
rect 2056 1092 2072 1108
rect 2120 1092 2136 1108
rect 2136 1032 2152 1048
rect 2168 1032 2184 1048
rect 2040 1012 2056 1028
rect 2616 1452 2632 1468
rect 2520 1372 2536 1388
rect 2600 1352 2616 1368
rect 2488 1332 2504 1348
rect 2472 1292 2488 1308
rect 2312 1172 2328 1188
rect 2360 1132 2376 1148
rect 2440 1132 2456 1148
rect 2328 1112 2344 1128
rect 2408 1112 2424 1128
rect 2280 1092 2296 1108
rect 2200 1072 2216 1088
rect 2280 1072 2296 1088
rect 2216 1052 2232 1068
rect 2232 1032 2248 1048
rect 2296 1012 2312 1028
rect 2184 992 2200 1008
rect 2232 992 2248 1008
rect 2472 1152 2488 1168
rect 2504 1152 2520 1168
rect 2456 1112 2472 1128
rect 2504 1092 2520 1108
rect 2584 1292 2600 1308
rect 2680 1492 2696 1508
rect 2728 1492 2744 1508
rect 2840 1612 2856 1628
rect 2872 1712 2888 1728
rect 2936 1712 2952 1728
rect 2856 1592 2872 1608
rect 2872 1572 2888 1588
rect 2888 1552 2904 1568
rect 3016 1872 3032 1888
rect 3016 1792 3032 1808
rect 3064 2012 3080 2028
rect 3064 1932 3080 1948
rect 3048 1872 3064 1888
rect 3192 2272 3208 2288
rect 3176 2232 3192 2248
rect 3384 2632 3400 2648
rect 3272 2612 3288 2628
rect 3272 2592 3288 2608
rect 3256 2552 3272 2568
rect 3240 2532 3256 2548
rect 3256 2512 3272 2528
rect 3320 2592 3336 2608
rect 3384 2532 3400 2548
rect 3480 3072 3496 3088
rect 3528 3272 3544 3288
rect 3560 3192 3576 3208
rect 3672 3972 3688 3988
rect 3624 3892 3640 3908
rect 3656 3892 3672 3908
rect 3640 3872 3656 3888
rect 3672 3872 3688 3888
rect 3640 3852 3656 3868
rect 3656 3772 3672 3788
rect 3688 3772 3704 3788
rect 3688 3752 3704 3768
rect 3656 3732 3688 3748
rect 3640 3692 3656 3708
rect 3992 4012 4008 4028
rect 4040 4012 4056 4028
rect 4072 4012 4088 4028
rect 4120 4012 4136 4028
rect 4168 4012 4184 4028
rect 4216 4012 4232 4028
rect 3752 3972 3768 3988
rect 3880 3972 3896 3988
rect 3960 3972 3976 3988
rect 3800 3952 3816 3968
rect 3752 3892 3768 3908
rect 3720 3872 3736 3888
rect 3768 3872 3784 3888
rect 4360 3992 4376 4008
rect 4312 3972 4328 3988
rect 4264 3932 4280 3948
rect 5021 4002 5057 4018
rect 5048 3952 5064 3968
rect 4856 3912 4872 3928
rect 4952 3912 4968 3928
rect 3896 3892 3912 3908
rect 3992 3892 4008 3908
rect 4088 3892 4104 3908
rect 4104 3892 4120 3908
rect 4200 3892 4216 3908
rect 4296 3892 4312 3908
rect 4440 3892 4456 3908
rect 4488 3892 4504 3908
rect 4552 3892 4568 3908
rect 4680 3892 4696 3908
rect 3880 3872 3896 3888
rect 3944 3872 3960 3888
rect 3848 3852 3864 3868
rect 3816 3732 3832 3748
rect 3768 3712 3784 3728
rect 3864 3792 3880 3808
rect 3944 3752 3960 3768
rect 3976 3872 3992 3888
rect 4008 3852 4024 3868
rect 3981 3802 4017 3818
rect 3848 3712 3864 3728
rect 3928 3712 3944 3728
rect 4008 3712 4024 3728
rect 3672 3692 3704 3708
rect 3752 3692 3768 3708
rect 3912 3692 3928 3708
rect 3960 3692 3976 3708
rect 3704 3672 3720 3688
rect 3880 3672 3896 3688
rect 4040 3852 4056 3868
rect 4072 3852 4088 3868
rect 4264 3872 4280 3888
rect 4360 3872 4376 3888
rect 4424 3876 4440 3888
rect 4424 3872 4440 3876
rect 4744 3876 4760 3888
rect 4744 3872 4760 3876
rect 4808 3876 4824 3888
rect 4808 3872 4824 3876
rect 4504 3852 4520 3868
rect 4568 3852 4584 3868
rect 4696 3852 4712 3868
rect 4184 3832 4200 3848
rect 4312 3832 4328 3848
rect 4424 3832 4440 3848
rect 4504 3832 4520 3848
rect 4152 3812 4168 3828
rect 4104 3752 4120 3768
rect 4184 3752 4200 3768
rect 4248 3732 4264 3748
rect 3752 3652 3768 3668
rect 4024 3652 4040 3668
rect 3736 3612 3752 3628
rect 3736 3592 3752 3608
rect 3672 3532 3688 3548
rect 3624 3412 3640 3428
rect 3624 3352 3640 3368
rect 3720 3512 3736 3528
rect 3704 3452 3720 3468
rect 3672 3312 3688 3328
rect 3784 3592 3800 3608
rect 3992 3572 4008 3588
rect 4008 3512 4024 3528
rect 4088 3672 4104 3688
rect 4104 3652 4120 3668
rect 4120 3632 4136 3648
rect 4376 3812 4392 3828
rect 4328 3792 4344 3808
rect 4456 3812 4472 3828
rect 4584 3812 4600 3828
rect 4632 3812 4648 3828
rect 4712 3812 4728 3828
rect 4520 3792 4536 3808
rect 4712 3792 4728 3808
rect 4824 3852 4840 3868
rect 4760 3772 4776 3788
rect 4792 3812 4808 3828
rect 4840 3812 4856 3828
rect 4712 3752 4728 3768
rect 4440 3732 4456 3748
rect 4536 3732 4552 3748
rect 4200 3552 4216 3568
rect 4200 3512 4216 3528
rect 3944 3492 3960 3508
rect 3992 3492 4008 3508
rect 4072 3492 4088 3508
rect 4200 3492 4216 3508
rect 3800 3392 3816 3408
rect 3768 3372 3784 3388
rect 3768 3352 3784 3368
rect 3656 3292 3672 3308
rect 3624 3252 3640 3268
rect 3656 3132 3672 3148
rect 3608 3112 3624 3128
rect 3608 3092 3624 3108
rect 3560 3052 3576 3068
rect 3544 3032 3560 3048
rect 3512 2992 3528 3008
rect 3496 2952 3512 2968
rect 3496 2932 3512 2948
rect 3560 2952 3576 2968
rect 3576 2932 3592 2948
rect 3464 2912 3480 2928
rect 3496 2912 3512 2928
rect 3592 2852 3608 2868
rect 3576 2832 3608 2848
rect 3480 2812 3496 2828
rect 3528 2772 3544 2788
rect 3448 2752 3464 2768
rect 3416 2692 3448 2708
rect 3432 2632 3448 2648
rect 3336 2512 3352 2528
rect 3480 2672 3496 2688
rect 3480 2612 3496 2628
rect 3448 2572 3464 2588
rect 3416 2492 3432 2508
rect 3352 2432 3368 2448
rect 3272 2372 3288 2388
rect 3304 2372 3320 2388
rect 3272 2352 3288 2368
rect 3240 2312 3256 2328
rect 3224 2272 3240 2288
rect 3160 2112 3176 2128
rect 3144 2092 3160 2108
rect 3176 1992 3192 2008
rect 3224 1972 3240 1988
rect 3256 2232 3272 2248
rect 3256 2212 3272 2228
rect 3384 2292 3400 2308
rect 3368 2272 3384 2288
rect 3640 3012 3656 3028
rect 3624 2932 3640 2948
rect 3640 2892 3656 2908
rect 3784 3232 3800 3248
rect 3784 3212 3800 3228
rect 3736 3192 3752 3208
rect 3768 3172 3784 3188
rect 3768 3132 3784 3148
rect 3720 3112 3736 3128
rect 3736 3072 3752 3088
rect 3672 2912 3688 2928
rect 3608 2812 3624 2828
rect 3640 2792 3656 2808
rect 3592 2752 3608 2768
rect 3560 2732 3576 2748
rect 3560 2692 3592 2708
rect 3544 2676 3560 2688
rect 3544 2672 3560 2676
rect 3624 2692 3640 2708
rect 3624 2672 3640 2688
rect 3624 2612 3640 2628
rect 3624 2572 3640 2588
rect 3576 2552 3592 2568
rect 3592 2532 3608 2548
rect 3544 2472 3560 2488
rect 3592 2472 3608 2488
rect 3448 2292 3464 2308
rect 3448 2272 3464 2288
rect 3336 2252 3352 2268
rect 3432 2232 3448 2248
rect 3560 2332 3576 2348
rect 3512 2292 3528 2308
rect 3544 2232 3560 2248
rect 3576 2232 3592 2248
rect 3432 2212 3448 2228
rect 3480 2212 3512 2228
rect 3352 2132 3368 2148
rect 3416 2132 3432 2148
rect 3320 2112 3336 2128
rect 3400 2112 3416 2128
rect 3288 2052 3304 2068
rect 3272 2012 3288 2028
rect 3288 1992 3304 2008
rect 3320 1992 3352 2008
rect 3256 1972 3272 1988
rect 3304 1972 3320 1988
rect 3192 1952 3208 1968
rect 3240 1952 3256 1968
rect 3208 1932 3224 1948
rect 3128 1912 3144 1928
rect 3112 1872 3128 1888
rect 3128 1872 3144 1888
rect 3128 1852 3144 1868
rect 3224 1872 3240 1888
rect 3080 1792 3096 1808
rect 3224 1852 3240 1868
rect 3176 1832 3192 1848
rect 3032 1772 3048 1788
rect 3048 1752 3064 1768
rect 3112 1732 3128 1748
rect 3160 1732 3176 1748
rect 3000 1712 3016 1728
rect 2952 1632 2968 1648
rect 2936 1592 2952 1608
rect 2973 1602 3009 1618
rect 2920 1492 2936 1508
rect 2728 1432 2744 1448
rect 2632 1412 2648 1428
rect 2664 1412 2680 1428
rect 2808 1412 2824 1428
rect 2648 1372 2664 1388
rect 2664 1372 2680 1388
rect 2776 1372 2792 1388
rect 2552 1272 2568 1288
rect 2568 1172 2584 1188
rect 2568 1152 2584 1168
rect 2552 1132 2568 1148
rect 2440 1052 2456 1068
rect 2424 1012 2440 1028
rect 2504 1012 2520 1028
rect 2296 952 2312 968
rect 2392 952 2408 968
rect 2056 932 2072 948
rect 2200 912 2216 928
rect 2248 912 2264 928
rect 2056 792 2072 808
rect 2040 692 2056 708
rect 1992 632 2008 648
rect 1992 612 2008 628
rect 2072 732 2088 748
rect 2088 712 2104 728
rect 2104 712 2120 728
rect 2104 632 2120 648
rect 2088 552 2104 568
rect 2168 892 2184 908
rect 2152 772 2168 788
rect 2200 812 2216 828
rect 2184 772 2200 788
rect 2360 912 2376 928
rect 2328 892 2344 908
rect 2344 752 2360 768
rect 2216 732 2232 748
rect 2280 732 2296 748
rect 2168 712 2184 728
rect 2312 712 2328 728
rect 2152 692 2168 708
rect 2200 692 2216 708
rect 2360 732 2376 748
rect 2376 712 2392 728
rect 2408 944 2424 948
rect 2408 932 2424 944
rect 2440 932 2456 948
rect 2488 912 2504 928
rect 2472 872 2488 888
rect 2424 852 2440 868
rect 2472 812 2488 828
rect 2408 792 2424 808
rect 2440 712 2456 728
rect 2392 692 2408 708
rect 2248 672 2264 688
rect 2200 652 2216 668
rect 2216 652 2232 668
rect 2280 652 2296 668
rect 2136 592 2152 608
rect 2248 612 2264 628
rect 2184 532 2200 548
rect 2232 512 2248 528
rect 1976 392 1992 408
rect 2072 412 2088 428
rect 2120 412 2136 428
rect 2056 392 2072 408
rect 2024 372 2040 388
rect 1944 332 1960 348
rect 2024 332 2040 348
rect 2040 332 2056 348
rect 1880 252 1896 268
rect 1960 252 1976 268
rect 1933 202 1969 218
rect 1880 32 1896 48
rect 1976 32 1992 48
rect 1928 12 1944 28
rect 2040 252 2056 268
rect 2072 172 2088 188
rect 2136 212 2152 228
rect 2120 192 2136 208
rect 2120 152 2136 168
rect 2248 432 2264 448
rect 2216 392 2232 408
rect 2424 592 2440 608
rect 2296 532 2312 548
rect 2408 532 2424 548
rect 2456 532 2472 548
rect 2328 512 2344 528
rect 2376 512 2392 528
rect 2520 992 2536 1008
rect 2520 912 2536 928
rect 2504 892 2520 908
rect 2536 872 2552 888
rect 2520 852 2536 868
rect 2520 712 2536 728
rect 2504 692 2520 708
rect 2536 672 2552 688
rect 2520 652 2536 668
rect 2568 1012 2584 1028
rect 2568 992 2584 1008
rect 2632 1192 2648 1208
rect 2616 1172 2632 1188
rect 2696 1352 2712 1368
rect 2776 1352 2792 1368
rect 2744 1332 2760 1348
rect 2824 1332 2840 1348
rect 2760 1292 2776 1308
rect 2712 1272 2728 1288
rect 2776 1272 2792 1288
rect 2808 1252 2824 1268
rect 2776 1192 2792 1208
rect 2680 1172 2696 1188
rect 2664 1132 2680 1148
rect 2792 1112 2808 1128
rect 2680 1092 2696 1108
rect 2760 1092 2776 1108
rect 2712 1072 2728 1088
rect 2616 932 2632 948
rect 2648 932 2680 948
rect 2728 932 2744 948
rect 2632 912 2648 928
rect 2600 872 2616 888
rect 2584 732 2600 748
rect 2568 712 2584 728
rect 2584 672 2600 688
rect 2584 652 2600 668
rect 2584 592 2600 608
rect 2520 512 2536 528
rect 2344 492 2360 508
rect 2392 492 2408 508
rect 2504 492 2520 508
rect 2312 432 2328 448
rect 2360 292 2376 308
rect 2280 272 2296 288
rect 2328 272 2344 288
rect 2376 272 2392 288
rect 2312 232 2328 248
rect 2344 232 2360 248
rect 2232 212 2248 228
rect 2152 152 2168 168
rect 2104 132 2120 148
rect 2392 212 2408 228
rect 2392 192 2408 208
rect 2360 132 2376 148
rect 2440 132 2456 148
rect 2040 114 2056 128
rect 2040 112 2056 114
rect 2104 112 2120 128
rect 2184 112 2200 128
rect 2552 532 2568 548
rect 2680 812 2696 828
rect 2728 792 2744 808
rect 2696 772 2712 788
rect 2824 1212 2840 1228
rect 2872 1472 2888 1488
rect 2920 1472 2936 1488
rect 2888 1392 2904 1408
rect 3064 1572 3080 1588
rect 2952 1532 2968 1548
rect 3112 1532 3128 1548
rect 3128 1532 3144 1548
rect 3112 1512 3128 1528
rect 3272 1832 3288 1848
rect 3224 1752 3240 1768
rect 3272 1752 3288 1768
rect 3208 1732 3224 1748
rect 3240 1732 3256 1748
rect 3272 1732 3288 1748
rect 3304 1744 3320 1748
rect 3304 1732 3320 1744
rect 3272 1692 3304 1708
rect 3224 1652 3240 1668
rect 3272 1612 3288 1628
rect 3224 1592 3240 1608
rect 3192 1572 3208 1588
rect 3400 2072 3416 2088
rect 3384 2052 3400 2068
rect 3368 1932 3384 1948
rect 3368 1852 3384 1868
rect 3368 1792 3384 1808
rect 3336 1752 3352 1768
rect 3352 1692 3368 1708
rect 3336 1532 3352 1548
rect 3256 1512 3272 1528
rect 3320 1512 3336 1528
rect 3496 2192 3512 2208
rect 3448 2072 3464 2088
rect 3672 2752 3688 2768
rect 3752 2972 3768 2988
rect 3768 2932 3784 2948
rect 3800 3032 3816 3048
rect 3912 3472 3928 3488
rect 4136 3472 4152 3488
rect 4360 3632 4376 3648
rect 4328 3532 4344 3548
rect 4376 3512 4392 3528
rect 4520 3692 4536 3708
rect 4520 3552 4536 3568
rect 4488 3512 4520 3528
rect 4552 3512 4568 3528
rect 4824 3752 4840 3768
rect 4840 3732 4856 3748
rect 4872 3892 4888 3908
rect 5000 3892 5016 3908
rect 4920 3872 4936 3888
rect 4888 3812 4904 3828
rect 4920 3792 4936 3808
rect 4968 3792 4984 3808
rect 4904 3732 4920 3748
rect 4584 3652 4600 3668
rect 4680 3692 4696 3708
rect 4712 3672 4728 3688
rect 4648 3632 4664 3648
rect 4584 3612 4600 3628
rect 4616 3512 4648 3528
rect 4392 3492 4408 3508
rect 4440 3492 4456 3508
rect 4568 3492 4584 3508
rect 3992 3452 4008 3468
rect 3928 3412 3944 3428
rect 3880 3352 3912 3368
rect 3864 3312 3880 3328
rect 3896 3312 3912 3328
rect 3864 3172 3880 3188
rect 3912 3172 3928 3188
rect 3896 3132 3912 3148
rect 3832 3092 3848 3108
rect 3864 3052 3880 3068
rect 3832 3032 3848 3048
rect 3912 3032 3928 3048
rect 3816 2972 3832 2988
rect 3752 2892 3768 2908
rect 3768 2852 3784 2868
rect 3816 2872 3832 2888
rect 3848 2992 3864 3008
rect 3896 2932 3912 2948
rect 3800 2832 3816 2848
rect 3832 2812 3848 2828
rect 3981 3402 4017 3418
rect 4104 3412 4120 3428
rect 3944 3372 3960 3388
rect 4040 3372 4056 3388
rect 4104 3352 4120 3368
rect 4680 3492 4696 3508
rect 4200 3432 4216 3448
rect 4184 3412 4200 3428
rect 4264 3472 4280 3488
rect 4312 3472 4328 3488
rect 4408 3472 4424 3488
rect 4456 3472 4472 3488
rect 4536 3472 4552 3488
rect 4360 3412 4376 3428
rect 4248 3392 4264 3408
rect 4296 3392 4312 3408
rect 4184 3352 4200 3368
rect 4216 3352 4248 3368
rect 4472 3452 4488 3468
rect 4392 3372 4408 3388
rect 4456 3352 4472 3368
rect 4056 3312 4072 3328
rect 4120 3312 4136 3328
rect 4312 3312 4328 3328
rect 4344 3312 4360 3328
rect 4376 3312 4392 3328
rect 4440 3312 4456 3328
rect 4024 3292 4056 3308
rect 4184 3292 4200 3308
rect 3976 3172 3992 3188
rect 3976 3092 3992 3108
rect 3960 3072 3976 3088
rect 3981 3002 4017 3018
rect 4312 3292 4328 3308
rect 4600 3432 4616 3448
rect 4568 3372 4584 3388
rect 4616 3412 4632 3428
rect 4584 3352 4600 3368
rect 4552 3312 4568 3328
rect 4536 3272 4552 3288
rect 4584 3292 4600 3308
rect 4184 3252 4200 3268
rect 4296 3252 4312 3268
rect 4440 3252 4456 3268
rect 4120 3232 4136 3248
rect 4056 3152 4072 3168
rect 4024 2972 4040 2988
rect 3960 2952 3976 2968
rect 3944 2932 3960 2948
rect 4024 2872 4040 2888
rect 3944 2772 3960 2788
rect 3928 2752 3944 2768
rect 4120 3112 4152 3128
rect 4376 3212 4392 3228
rect 4200 3132 4216 3148
rect 4344 3112 4360 3128
rect 4200 3092 4216 3108
rect 4248 3092 4264 3108
rect 4168 3072 4184 3088
rect 4472 3232 4488 3248
rect 4392 3092 4408 3108
rect 4328 3072 4344 3088
rect 4216 3052 4232 3068
rect 4312 3052 4328 3068
rect 4184 3012 4200 3028
rect 4168 2992 4184 3008
rect 4088 2952 4104 2968
rect 4120 2952 4136 2968
rect 4152 2952 4168 2968
rect 4072 2932 4088 2948
rect 4456 3072 4472 3088
rect 4312 2992 4328 3008
rect 4440 2992 4456 3008
rect 4520 3152 4536 3168
rect 4504 3072 4520 3088
rect 4552 3192 4568 3208
rect 4536 3132 4552 3148
rect 4536 3072 4552 3088
rect 4600 3112 4616 3128
rect 4632 3352 4648 3368
rect 4888 3692 4904 3708
rect 4856 3672 4872 3688
rect 4840 3632 4856 3648
rect 4792 3592 4808 3608
rect 4728 3552 4744 3568
rect 4728 3512 4744 3528
rect 4760 3492 4776 3508
rect 4808 3492 4824 3508
rect 4712 3472 4728 3488
rect 4776 3452 4792 3468
rect 4984 3712 5000 3728
rect 4952 3632 4968 3648
rect 5128 3932 5144 3948
rect 5064 3912 5080 3928
rect 5096 3892 5112 3908
rect 5160 3892 5176 3908
rect 5288 3892 5304 3908
rect 5336 3892 5352 3908
rect 5608 3892 5624 3908
rect 5144 3872 5160 3888
rect 5064 3772 5080 3788
rect 5048 3672 5064 3688
rect 5021 3602 5057 3618
rect 4904 3472 4920 3488
rect 4952 3472 4968 3488
rect 4888 3432 4904 3448
rect 4808 3412 4824 3428
rect 4920 3412 4936 3428
rect 4696 3392 4712 3408
rect 4808 3392 4824 3408
rect 4696 3352 4712 3368
rect 4744 3352 4760 3368
rect 4680 3312 4696 3328
rect 4840 3352 4856 3368
rect 5176 3832 5192 3848
rect 5160 3772 5176 3788
rect 5240 3872 5256 3888
rect 5384 3872 5400 3888
rect 5400 3872 5416 3888
rect 5432 3872 5448 3888
rect 5480 3872 5496 3888
rect 5288 3852 5320 3868
rect 5368 3852 5384 3868
rect 5224 3772 5240 3788
rect 5224 3752 5240 3768
rect 5256 3752 5272 3768
rect 5288 3752 5304 3768
rect 5320 3752 5336 3768
rect 5048 3472 5064 3488
rect 5192 3652 5208 3668
rect 5336 3652 5352 3668
rect 5096 3632 5112 3648
rect 5128 3632 5144 3648
rect 5160 3632 5176 3648
rect 5080 3392 5096 3408
rect 5032 3352 5048 3368
rect 4824 3332 4840 3348
rect 4904 3332 4920 3348
rect 4952 3332 4968 3348
rect 5000 3332 5016 3348
rect 5016 3332 5032 3348
rect 5080 3344 5096 3348
rect 5080 3332 5096 3344
rect 4872 3312 4888 3328
rect 4776 3252 4792 3268
rect 4712 3192 4728 3208
rect 4664 3152 4680 3168
rect 4696 3152 4712 3168
rect 4648 3112 4664 3128
rect 4760 3112 4776 3128
rect 4824 3112 4840 3128
rect 4616 3092 4632 3108
rect 4632 3092 4648 3108
rect 4696 3092 4712 3108
rect 4808 3092 4824 3108
rect 4584 3072 4600 3088
rect 4552 3012 4568 3028
rect 4488 2992 4520 3008
rect 4312 2952 4328 2968
rect 4472 2952 4488 2968
rect 4200 2932 4216 2948
rect 4216 2932 4232 2948
rect 4264 2932 4280 2948
rect 4344 2932 4360 2948
rect 4408 2912 4424 2928
rect 4456 2912 4472 2928
rect 4040 2832 4056 2848
rect 4088 2892 4104 2908
rect 4056 2772 4072 2788
rect 4040 2752 4072 2768
rect 4312 2852 4328 2868
rect 4296 2832 4312 2848
rect 4184 2772 4200 2788
rect 4072 2732 4088 2748
rect 4104 2712 4120 2728
rect 3752 2692 3768 2708
rect 3800 2692 3816 2708
rect 3864 2692 3880 2708
rect 3912 2692 3928 2708
rect 3880 2652 3896 2668
rect 3928 2652 3944 2668
rect 3688 2632 3704 2648
rect 3736 2632 3752 2648
rect 3912 2632 3928 2648
rect 3672 2612 3688 2628
rect 3704 2592 3720 2608
rect 3736 2552 3752 2568
rect 3752 2532 3768 2548
rect 3672 2512 3688 2528
rect 3656 2492 3672 2508
rect 3864 2592 3880 2608
rect 3912 2572 3928 2588
rect 3784 2532 3800 2548
rect 3832 2532 3848 2548
rect 3720 2492 3736 2508
rect 3768 2492 3784 2508
rect 3656 2472 3672 2488
rect 3688 2472 3704 2488
rect 3704 2472 3720 2488
rect 3832 2472 3848 2488
rect 3896 2472 3912 2488
rect 3704 2412 3720 2428
rect 3784 2392 3800 2408
rect 3752 2372 3768 2388
rect 3672 2332 3688 2348
rect 3720 2312 3752 2328
rect 3624 2252 3640 2268
rect 3688 2252 3704 2268
rect 3672 2232 3704 2248
rect 3608 2192 3624 2208
rect 3592 2172 3608 2188
rect 3608 2152 3624 2168
rect 3624 2132 3640 2148
rect 3480 2112 3496 2128
rect 3608 2112 3624 2128
rect 3544 2092 3560 2108
rect 3464 2012 3480 2028
rect 3448 1892 3464 1908
rect 3416 1872 3432 1888
rect 3416 1792 3432 1808
rect 3400 1752 3416 1768
rect 3528 1912 3544 1928
rect 3496 1872 3512 1888
rect 3640 2032 3656 2048
rect 3624 1992 3640 2008
rect 3608 1972 3624 1988
rect 3656 1952 3672 1968
rect 3672 1932 3688 1948
rect 3640 1892 3656 1908
rect 3592 1852 3608 1868
rect 3640 1852 3656 1868
rect 3528 1832 3544 1848
rect 3576 1832 3592 1848
rect 3464 1772 3480 1788
rect 3432 1712 3448 1728
rect 3384 1632 3416 1648
rect 3384 1612 3400 1628
rect 3416 1612 3432 1628
rect 3464 1712 3480 1728
rect 3512 1712 3528 1728
rect 3496 1592 3512 1608
rect 3560 1812 3576 1828
rect 3560 1772 3576 1788
rect 3544 1752 3560 1768
rect 3544 1712 3560 1728
rect 3624 1692 3640 1708
rect 3768 2292 3784 2308
rect 3752 2192 3768 2208
rect 3752 2152 3768 2168
rect 3704 2112 3720 2128
rect 3704 2072 3720 2088
rect 3800 2312 3816 2328
rect 3768 2112 3784 2128
rect 3784 2032 3800 2048
rect 3976 2632 3992 2648
rect 4024 2632 4040 2648
rect 3981 2602 4017 2618
rect 3992 2572 4008 2588
rect 3944 2552 3960 2568
rect 4008 2512 4024 2528
rect 3944 2492 3960 2508
rect 3992 2332 4008 2348
rect 3976 2312 3992 2328
rect 4024 2292 4040 2308
rect 3880 2276 3896 2288
rect 3880 2272 3896 2276
rect 3928 2272 3944 2288
rect 3880 2252 3896 2268
rect 3848 2132 3864 2148
rect 3864 2112 3880 2128
rect 3832 2092 3848 2108
rect 3960 2252 3976 2268
rect 3944 2192 3960 2208
rect 3912 2072 3928 2088
rect 3816 2052 3832 2068
rect 3816 2032 3832 2048
rect 3800 2012 3816 2028
rect 3912 2012 3928 2028
rect 3864 1952 3880 1968
rect 3928 1952 3944 1968
rect 3784 1912 3800 1928
rect 3752 1892 3768 1908
rect 3832 1892 3848 1908
rect 3688 1872 3704 1888
rect 3800 1872 3832 1888
rect 3928 1872 3944 1888
rect 3688 1792 3704 1808
rect 3672 1732 3688 1748
rect 3720 1692 3736 1708
rect 3656 1672 3672 1688
rect 3816 1772 3832 1788
rect 3848 1752 3864 1768
rect 3768 1732 3784 1748
rect 3816 1732 3832 1748
rect 3832 1712 3848 1728
rect 3752 1672 3768 1688
rect 3736 1652 3752 1668
rect 3624 1612 3640 1628
rect 3656 1612 3672 1628
rect 3576 1572 3592 1588
rect 3496 1512 3512 1528
rect 3288 1492 3320 1508
rect 3480 1492 3512 1508
rect 3128 1472 3144 1488
rect 3224 1472 3240 1488
rect 3256 1472 3272 1488
rect 3032 1452 3048 1468
rect 3096 1452 3112 1468
rect 3128 1452 3144 1468
rect 3320 1452 3336 1468
rect 3048 1432 3064 1448
rect 3048 1412 3064 1428
rect 3096 1412 3112 1428
rect 3080 1392 3096 1408
rect 3064 1352 3080 1368
rect 3048 1332 3064 1348
rect 2872 1292 2888 1308
rect 2952 1292 2968 1308
rect 2920 1252 2936 1268
rect 2856 1192 2872 1208
rect 2840 1172 2856 1188
rect 2840 1112 2856 1128
rect 2824 1092 2840 1108
rect 2872 1052 2888 1068
rect 2840 1032 2856 1048
rect 2792 972 2808 988
rect 2888 952 2904 968
rect 2904 932 2920 948
rect 2840 832 2856 848
rect 2936 1112 2952 1128
rect 3000 1232 3016 1248
rect 2973 1202 3009 1218
rect 3048 1132 3064 1148
rect 2984 1112 3000 1128
rect 3064 1112 3080 1128
rect 2984 1072 3000 1088
rect 2936 992 2952 1008
rect 3048 1012 3064 1028
rect 3112 1372 3128 1388
rect 3176 1332 3192 1348
rect 3240 1412 3256 1428
rect 3224 1352 3240 1368
rect 3304 1352 3320 1368
rect 3160 1312 3176 1328
rect 3176 1212 3192 1228
rect 3160 1192 3176 1208
rect 3144 1172 3160 1188
rect 3208 1192 3224 1208
rect 3144 1092 3160 1108
rect 3176 1052 3192 1068
rect 2936 952 2952 968
rect 3160 952 3176 968
rect 3432 1452 3448 1468
rect 3384 1412 3400 1428
rect 3368 1372 3384 1388
rect 3288 1332 3304 1348
rect 3336 1332 3352 1348
rect 3592 1552 3608 1568
rect 3688 1552 3704 1568
rect 3608 1492 3624 1508
rect 3528 1452 3544 1468
rect 3576 1452 3592 1468
rect 3512 1432 3528 1448
rect 3560 1432 3576 1448
rect 3656 1432 3672 1448
rect 3480 1352 3496 1368
rect 3464 1332 3480 1348
rect 3272 1272 3288 1288
rect 3256 1232 3272 1248
rect 3432 1292 3448 1308
rect 3352 1232 3368 1248
rect 3320 1112 3336 1128
rect 3352 1112 3368 1128
rect 3336 1092 3352 1108
rect 3416 1092 3432 1108
rect 3448 1252 3464 1268
rect 3512 1332 3528 1348
rect 3528 1332 3544 1348
rect 3592 1352 3624 1368
rect 3496 1292 3512 1308
rect 3608 1292 3624 1308
rect 3480 1232 3496 1248
rect 3528 1232 3544 1248
rect 3240 1072 3256 1088
rect 3368 1072 3384 1088
rect 3416 1072 3432 1088
rect 3448 1072 3464 1088
rect 3224 1032 3240 1048
rect 3320 1052 3336 1068
rect 3192 972 3208 988
rect 3320 1032 3336 1048
rect 3304 972 3320 988
rect 3192 952 3208 968
rect 3208 952 3224 968
rect 3256 952 3288 968
rect 3336 972 3352 988
rect 3080 932 3096 948
rect 2952 912 2968 928
rect 3032 912 3048 928
rect 2888 872 2904 888
rect 2872 812 2888 828
rect 2760 772 2776 788
rect 2840 772 2856 788
rect 2856 772 2872 788
rect 2680 752 2696 768
rect 2744 752 2760 768
rect 2728 712 2744 728
rect 2824 712 2840 728
rect 2792 692 2824 708
rect 2840 692 2856 708
rect 2744 672 2760 688
rect 2616 652 2632 668
rect 2616 572 2632 588
rect 2856 632 2872 648
rect 2680 612 2696 628
rect 2712 592 2728 608
rect 2760 592 2776 608
rect 2680 552 2696 568
rect 2760 572 2776 588
rect 2808 572 2824 588
rect 2888 792 2904 808
rect 3160 912 3176 928
rect 3064 872 3080 888
rect 3128 872 3144 888
rect 3176 852 3192 868
rect 3048 832 3064 848
rect 2973 802 3009 818
rect 3000 772 3016 788
rect 3112 772 3128 788
rect 3016 732 3032 748
rect 3080 732 3096 748
rect 2920 712 2936 728
rect 2984 712 3000 728
rect 2968 692 2984 708
rect 3000 692 3016 708
rect 3144 732 3160 748
rect 3176 732 3192 748
rect 3224 932 3240 948
rect 3256 912 3272 928
rect 3240 892 3256 908
rect 3352 892 3368 908
rect 3208 872 3224 888
rect 3256 852 3272 868
rect 3320 852 3336 868
rect 3128 712 3144 728
rect 3224 712 3240 728
rect 3112 692 3128 708
rect 3176 692 3192 708
rect 2920 632 2936 648
rect 2904 572 2920 588
rect 2888 552 2904 568
rect 2616 512 2632 528
rect 2856 512 2872 528
rect 2952 532 2968 548
rect 3176 632 3192 648
rect 3208 692 3224 708
rect 3032 572 3048 588
rect 3192 572 3208 588
rect 2968 512 2984 528
rect 3016 512 3032 528
rect 3048 552 3064 568
rect 3096 552 3112 568
rect 3128 552 3144 568
rect 3064 532 3096 548
rect 3144 532 3160 548
rect 3240 572 3256 588
rect 3400 952 3416 968
rect 3576 1192 3592 1208
rect 3720 1512 3736 1528
rect 3800 1632 3816 1648
rect 3784 1512 3800 1528
rect 3832 1512 3848 1528
rect 3816 1492 3832 1508
rect 3832 1472 3848 1488
rect 3752 1432 3768 1448
rect 3688 1352 3704 1368
rect 3672 1332 3688 1348
rect 3736 1332 3752 1348
rect 3768 1332 3784 1348
rect 3896 1772 3912 1788
rect 3880 1752 3896 1768
rect 3928 1832 3944 1848
rect 3981 2202 4017 2218
rect 4168 2632 4184 2648
rect 4104 2592 4120 2608
rect 4056 2412 4072 2428
rect 4056 2332 4072 2348
rect 4056 2292 4072 2308
rect 4056 2272 4072 2288
rect 4104 2552 4120 2568
rect 4232 2532 4248 2548
rect 4168 2512 4184 2528
rect 4200 2512 4216 2528
rect 4152 2472 4168 2488
rect 4184 2472 4200 2488
rect 4088 2412 4104 2428
rect 4184 2332 4200 2348
rect 4104 2312 4120 2328
rect 4152 2312 4168 2328
rect 4088 2292 4104 2308
rect 4072 2212 4088 2228
rect 4104 2172 4120 2188
rect 4088 2132 4104 2148
rect 4040 2112 4056 2128
rect 4072 2112 4088 2128
rect 4040 2092 4056 2108
rect 3976 1872 3992 1888
rect 4008 1852 4024 1868
rect 3981 1802 4017 1818
rect 4152 2212 4168 2228
rect 4120 2052 4136 2068
rect 4264 2552 4280 2568
rect 4360 2812 4376 2828
rect 4344 2732 4360 2748
rect 4376 2692 4392 2708
rect 4392 2652 4408 2668
rect 4312 2572 4328 2588
rect 4280 2532 4296 2548
rect 4296 2532 4312 2548
rect 4312 2512 4328 2528
rect 4216 2312 4232 2328
rect 4200 2292 4216 2308
rect 4216 2232 4232 2248
rect 4184 2052 4200 2068
rect 4200 1992 4216 2008
rect 4168 1952 4184 1968
rect 4136 1912 4152 1928
rect 4184 1892 4200 1908
rect 4184 1872 4200 1888
rect 4056 1832 4072 1848
rect 4024 1792 4040 1808
rect 3960 1772 3976 1788
rect 3992 1772 4008 1788
rect 3960 1752 3976 1768
rect 3944 1732 3960 1748
rect 4024 1752 4040 1768
rect 4008 1732 4024 1748
rect 3928 1712 3944 1728
rect 4056 1632 4072 1648
rect 3928 1592 3944 1608
rect 3912 1552 3928 1568
rect 3912 1512 3928 1528
rect 4120 1812 4136 1828
rect 4088 1772 4104 1788
rect 4088 1752 4104 1768
rect 4232 2212 4248 2228
rect 4232 2152 4248 2168
rect 4296 2392 4312 2408
rect 4264 2292 4280 2308
rect 4296 2252 4312 2268
rect 4312 2232 4328 2248
rect 4312 2192 4328 2208
rect 4280 2152 4296 2168
rect 4280 2092 4296 2108
rect 4296 2092 4312 2108
rect 4232 2052 4248 2068
rect 4248 1992 4264 2008
rect 4280 1992 4296 2008
rect 4312 1972 4328 1988
rect 4248 1892 4264 1908
rect 4296 1892 4312 1908
rect 4232 1872 4248 1888
rect 4232 1792 4248 1808
rect 4136 1772 4152 1788
rect 4136 1712 4152 1728
rect 4072 1572 4088 1588
rect 4360 2592 4376 2608
rect 4392 2412 4408 2428
rect 4344 2392 4360 2408
rect 4696 2992 4712 3008
rect 4616 2952 4632 2968
rect 4712 2972 4728 2988
rect 4696 2952 4712 2968
rect 4664 2912 4680 2928
rect 4680 2912 4696 2928
rect 4712 2912 4728 2928
rect 4584 2892 4600 2908
rect 4584 2872 4600 2888
rect 4520 2792 4536 2808
rect 4440 2772 4456 2788
rect 4424 2732 4440 2748
rect 4424 2712 4440 2728
rect 4360 2292 4376 2308
rect 4408 2312 4424 2328
rect 4504 2752 4520 2768
rect 4584 2752 4600 2768
rect 4488 2732 4504 2748
rect 4536 2732 4552 2748
rect 4600 2712 4616 2728
rect 4520 2672 4536 2688
rect 4456 2592 4472 2608
rect 4440 2572 4456 2588
rect 4504 2552 4520 2568
rect 4632 2652 4648 2668
rect 4632 2612 4648 2628
rect 4648 2552 4664 2568
rect 4696 2652 4712 2668
rect 4600 2532 4616 2548
rect 4664 2544 4680 2548
rect 4664 2532 4680 2544
rect 4744 3012 4760 3028
rect 4920 3312 4936 3328
rect 4968 3312 4984 3328
rect 5064 3292 5080 3308
rect 5000 3272 5016 3288
rect 4984 3212 5000 3228
rect 4904 3172 4920 3188
rect 4904 3112 4920 3128
rect 4888 3092 4904 3108
rect 4936 3092 4952 3108
rect 4920 3072 4936 3088
rect 4872 2972 4888 2988
rect 4792 2952 4824 2968
rect 4904 2952 4920 2968
rect 4952 3052 4968 3068
rect 4968 3032 4984 3048
rect 4968 2992 4984 3008
rect 4952 2932 4968 2948
rect 4872 2912 4888 2928
rect 4920 2912 4936 2928
rect 4888 2892 4904 2908
rect 4840 2872 4856 2888
rect 4744 2732 4760 2748
rect 4776 2692 4792 2708
rect 4824 2672 4840 2688
rect 4856 2672 4872 2688
rect 4760 2612 4776 2628
rect 4904 2612 4920 2628
rect 4888 2592 4904 2608
rect 4824 2552 4840 2568
rect 4888 2552 4904 2568
rect 4760 2532 4776 2548
rect 4792 2532 4808 2548
rect 4488 2472 4504 2488
rect 4520 2472 4536 2488
rect 4488 2312 4504 2328
rect 4440 2292 4456 2308
rect 4472 2292 4488 2308
rect 4552 2352 4568 2368
rect 4552 2312 4568 2328
rect 4600 2292 4616 2308
rect 4424 2272 4456 2288
rect 4520 2272 4536 2288
rect 4584 2272 4600 2288
rect 4392 2132 4408 2148
rect 4376 2112 4392 2128
rect 4600 2232 4616 2248
rect 4424 2172 4440 2188
rect 4504 2172 4520 2188
rect 4552 2212 4568 2228
rect 4568 2172 4584 2188
rect 4472 2132 4488 2148
rect 4520 2132 4536 2148
rect 4584 2132 4600 2148
rect 4536 2112 4552 2128
rect 4360 2052 4376 2068
rect 4360 1972 4376 1988
rect 4488 2012 4504 2028
rect 4472 1952 4488 1968
rect 4504 1992 4520 2008
rect 4872 2492 4888 2508
rect 4632 2432 4648 2448
rect 4712 2412 4728 2428
rect 4840 2412 4856 2428
rect 4904 2392 4920 2408
rect 4744 2352 4760 2368
rect 4728 2332 4744 2348
rect 4696 2312 4712 2328
rect 4632 2252 4648 2268
rect 4696 2252 4712 2268
rect 4648 2192 4664 2208
rect 4632 2152 4648 2168
rect 4824 2312 4840 2328
rect 4776 2292 4792 2308
rect 4792 2292 4808 2308
rect 4840 2292 4856 2308
rect 4968 2892 4984 2908
rect 4952 2692 4968 2708
rect 5021 3202 5057 3218
rect 5016 3012 5032 3028
rect 5032 2932 5048 2948
rect 5048 2892 5064 2908
rect 5021 2802 5057 2818
rect 5192 3552 5208 3568
rect 5112 3492 5128 3508
rect 5256 3572 5272 3588
rect 5240 3512 5256 3528
rect 5240 3492 5256 3508
rect 5112 3472 5128 3488
rect 5320 3512 5336 3528
rect 5336 3492 5352 3508
rect 5304 3476 5320 3488
rect 5304 3472 5320 3476
rect 5256 3452 5272 3468
rect 5352 3452 5368 3468
rect 5176 3392 5192 3408
rect 5144 3352 5160 3368
rect 5176 3352 5192 3368
rect 5112 3332 5128 3348
rect 5160 3332 5176 3348
rect 5208 3332 5224 3348
rect 5272 3352 5288 3368
rect 5336 3352 5352 3368
rect 5304 3332 5320 3348
rect 5432 3752 5448 3768
rect 5416 3712 5432 3728
rect 5624 3872 5640 3888
rect 5656 3872 5672 3888
rect 5560 3852 5576 3868
rect 5544 3812 5560 3828
rect 5512 3772 5528 3788
rect 5496 3752 5512 3768
rect 5464 3732 5480 3748
rect 5496 3732 5512 3748
rect 5448 3692 5464 3708
rect 5496 3672 5512 3688
rect 5384 3492 5400 3508
rect 5464 3492 5480 3508
rect 5688 3872 5704 3888
rect 5864 3872 5880 3888
rect 5672 3852 5688 3868
rect 5736 3852 5752 3868
rect 5672 3832 5688 3848
rect 5640 3772 5656 3788
rect 5608 3752 5624 3768
rect 5704 3752 5720 3768
rect 5736 3752 5752 3768
rect 5832 3752 5848 3768
rect 5688 3732 5704 3748
rect 5752 3732 5768 3748
rect 5912 3732 5928 3748
rect 5624 3712 5640 3728
rect 5544 3632 5560 3648
rect 5528 3512 5560 3528
rect 5400 3472 5416 3488
rect 5400 3352 5416 3368
rect 5288 3312 5304 3328
rect 5368 3312 5384 3328
rect 5192 3272 5208 3288
rect 5256 3272 5272 3288
rect 5096 3252 5112 3268
rect 5128 3232 5144 3248
rect 5224 3212 5240 3228
rect 5320 3212 5336 3228
rect 5176 3092 5192 3108
rect 5208 3072 5224 3088
rect 5192 2992 5208 3008
rect 5272 3072 5288 3088
rect 5336 3032 5352 3048
rect 5240 2952 5256 2968
rect 5096 2932 5112 2948
rect 5176 2932 5192 2948
rect 5256 2932 5272 2948
rect 5112 2912 5128 2928
rect 5208 2912 5224 2928
rect 5080 2892 5096 2908
rect 5160 2892 5176 2908
rect 5064 2772 5080 2788
rect 4936 2612 4952 2628
rect 4984 2612 5000 2628
rect 4968 2592 4984 2608
rect 5032 2632 5048 2648
rect 5048 2632 5064 2648
rect 4952 2552 4968 2568
rect 5000 2552 5016 2568
rect 4936 2532 4952 2548
rect 5048 2532 5064 2548
rect 4984 2512 5000 2528
rect 5032 2512 5048 2528
rect 4984 2472 5000 2488
rect 4824 2232 4840 2248
rect 4744 2192 4760 2208
rect 4648 2132 4664 2148
rect 4696 2132 4712 2148
rect 4680 2112 4696 2128
rect 4616 2072 4632 2088
rect 4696 2052 4712 2068
rect 4600 1952 4616 1968
rect 4648 1952 4664 1968
rect 4712 1992 4728 2008
rect 4728 1932 4744 1948
rect 4456 1892 4472 1908
rect 4648 1892 4664 1908
rect 4712 1892 4728 1908
rect 4328 1772 4344 1788
rect 4376 1872 4392 1888
rect 4408 1872 4424 1888
rect 4504 1872 4520 1888
rect 4552 1872 4568 1888
rect 4616 1872 4632 1888
rect 4472 1852 4488 1868
rect 4536 1852 4552 1868
rect 4424 1832 4440 1848
rect 4552 1832 4568 1848
rect 4472 1752 4488 1768
rect 4568 1752 4584 1768
rect 4616 1752 4632 1768
rect 4648 1752 4664 1768
rect 4280 1732 4296 1748
rect 4296 1712 4312 1728
rect 4184 1632 4200 1648
rect 4088 1532 4104 1548
rect 4136 1532 4152 1548
rect 4008 1492 4024 1508
rect 4024 1472 4040 1488
rect 4072 1472 4088 1488
rect 3928 1452 3944 1468
rect 3992 1452 4008 1468
rect 4008 1452 4024 1468
rect 3880 1412 3896 1428
rect 3896 1392 3912 1408
rect 3981 1402 4017 1418
rect 3864 1372 3880 1388
rect 3880 1352 3896 1368
rect 4104 1512 4120 1528
rect 4136 1492 4152 1508
rect 4168 1512 4184 1528
rect 4184 1472 4200 1488
rect 4184 1432 4200 1448
rect 4040 1372 4056 1388
rect 4264 1672 4280 1688
rect 4264 1572 4280 1588
rect 4232 1552 4248 1568
rect 4248 1532 4264 1548
rect 4632 1712 4648 1728
rect 4376 1692 4392 1708
rect 4328 1672 4344 1688
rect 4312 1552 4328 1568
rect 4344 1552 4360 1568
rect 4376 1532 4392 1548
rect 4296 1512 4312 1528
rect 4664 1672 4680 1688
rect 4600 1552 4616 1568
rect 4488 1532 4504 1548
rect 4392 1512 4408 1528
rect 4472 1512 4488 1528
rect 4456 1492 4472 1508
rect 4616 1512 4632 1528
rect 4760 2092 4776 2108
rect 4792 2012 4808 2028
rect 4824 2172 4840 2188
rect 4952 2272 4968 2288
rect 4936 2212 4952 2228
rect 4920 2192 4936 2208
rect 4824 2112 4840 2128
rect 4824 2072 4840 2088
rect 4808 1972 4824 1988
rect 4872 2112 4888 2128
rect 4920 2112 4936 2128
rect 5016 2452 5032 2468
rect 5021 2402 5057 2418
rect 5000 2292 5016 2308
rect 5016 2272 5032 2288
rect 5032 2272 5048 2288
rect 4968 2092 4984 2108
rect 5048 2132 5064 2148
rect 4968 2072 4984 2088
rect 4920 2052 4936 2068
rect 4888 1992 4904 2008
rect 4856 1932 4872 1948
rect 4840 1912 4856 1928
rect 4744 1892 4760 1908
rect 4696 1772 4712 1788
rect 4696 1752 4728 1768
rect 4808 1792 4824 1808
rect 4808 1752 4824 1768
rect 4696 1732 4712 1748
rect 4856 1832 4872 1848
rect 4856 1812 4872 1828
rect 5032 2092 5064 2108
rect 5064 2072 5080 2088
rect 5000 2032 5016 2048
rect 4936 1972 4952 1988
rect 4952 1852 4968 1868
rect 5021 2002 5057 2018
rect 5320 2932 5336 2948
rect 5320 2892 5336 2908
rect 5336 2832 5352 2848
rect 5272 2812 5288 2828
rect 5304 2812 5320 2828
rect 5336 2812 5352 2828
rect 5192 2792 5208 2808
rect 5128 2692 5144 2708
rect 5160 2692 5176 2708
rect 5096 2652 5112 2668
rect 5112 2632 5128 2648
rect 5128 2532 5144 2548
rect 5208 2672 5224 2688
rect 5304 2652 5320 2668
rect 5288 2632 5304 2648
rect 5240 2592 5256 2608
rect 5208 2572 5224 2588
rect 5224 2552 5240 2568
rect 5240 2532 5256 2548
rect 5096 2512 5112 2528
rect 5160 2512 5176 2528
rect 5176 2512 5192 2528
rect 5112 2492 5128 2508
rect 5192 2412 5208 2428
rect 5160 2312 5176 2328
rect 5224 2312 5240 2328
rect 5304 2492 5320 2508
rect 5416 3192 5432 3208
rect 5416 3152 5432 3168
rect 5416 3012 5432 3028
rect 5384 2992 5400 3008
rect 5368 2932 5384 2948
rect 5448 3412 5464 3428
rect 5528 3412 5544 3428
rect 5624 3512 5640 3528
rect 5592 3492 5608 3508
rect 5576 3472 5592 3488
rect 5656 3472 5672 3488
rect 5704 3712 5720 3728
rect 5768 3712 5784 3728
rect 5864 3632 5880 3648
rect 5912 3612 5928 3628
rect 5880 3592 5896 3608
rect 5832 3512 5848 3528
rect 5704 3492 5720 3508
rect 5864 3492 5880 3508
rect 5688 3472 5704 3488
rect 5672 3452 5688 3468
rect 5560 3392 5576 3408
rect 5560 3372 5576 3388
rect 5608 3352 5624 3368
rect 5720 3452 5736 3468
rect 5688 3412 5704 3428
rect 5640 3352 5656 3368
rect 5448 3332 5464 3348
rect 5512 3332 5528 3348
rect 5560 3332 5576 3348
rect 5816 3472 5832 3488
rect 5832 3472 5848 3488
rect 5864 3472 5880 3488
rect 5800 3332 5816 3348
rect 5512 3292 5528 3308
rect 5432 2972 5464 2988
rect 5432 2932 5448 2948
rect 5464 2932 5480 2948
rect 5432 2812 5448 2828
rect 5464 2812 5496 2828
rect 5368 2792 5384 2808
rect 5368 2772 5384 2788
rect 5528 3072 5544 3088
rect 5592 3312 5608 3328
rect 5688 3312 5704 3328
rect 5864 3312 5880 3328
rect 5576 3292 5592 3308
rect 5720 3292 5736 3308
rect 5800 3292 5816 3308
rect 5752 3232 5768 3248
rect 5720 3212 5752 3228
rect 5656 3192 5672 3208
rect 5688 3172 5704 3188
rect 5608 3132 5624 3148
rect 5592 3072 5608 3088
rect 5672 3072 5688 3088
rect 5544 3012 5560 3028
rect 5576 3012 5592 3028
rect 5608 3012 5624 3028
rect 5608 2972 5624 2988
rect 5592 2932 5608 2948
rect 5672 2932 5688 2948
rect 5720 3092 5736 3108
rect 5720 3072 5736 3088
rect 5784 3072 5800 3088
rect 5784 3052 5800 3068
rect 5704 3032 5720 3048
rect 5640 2852 5656 2868
rect 5528 2792 5544 2808
rect 5416 2692 5432 2708
rect 5480 2692 5496 2708
rect 5496 2692 5512 2708
rect 5496 2672 5512 2688
rect 5352 2652 5368 2668
rect 5352 2592 5368 2608
rect 5384 2592 5400 2608
rect 5416 2572 5432 2588
rect 5464 2612 5480 2628
rect 5448 2552 5464 2568
rect 5448 2532 5464 2548
rect 5432 2512 5448 2528
rect 5432 2452 5448 2468
rect 5320 2412 5336 2428
rect 5448 2332 5464 2348
rect 5176 2292 5192 2308
rect 5432 2292 5448 2308
rect 5096 2272 5112 2288
rect 5144 2272 5160 2288
rect 5096 2152 5128 2168
rect 5320 2272 5336 2288
rect 5256 2252 5272 2268
rect 5272 2232 5288 2248
rect 5176 2212 5192 2228
rect 5176 2192 5192 2208
rect 5176 2144 5192 2148
rect 5176 2132 5192 2144
rect 5160 2112 5176 2128
rect 5144 1952 5160 1968
rect 5016 1892 5032 1908
rect 5000 1812 5016 1828
rect 4968 1772 4984 1788
rect 4792 1712 4808 1728
rect 4824 1712 4840 1728
rect 5032 1752 5048 1768
rect 5016 1732 5032 1748
rect 5176 1832 5192 1848
rect 5304 2172 5320 2188
rect 5416 2252 5432 2268
rect 5368 2232 5384 2248
rect 5224 2152 5240 2168
rect 5320 2152 5336 2168
rect 5400 2152 5416 2168
rect 5464 2172 5480 2188
rect 5592 2712 5608 2728
rect 5656 2812 5672 2828
rect 5640 2692 5656 2708
rect 5688 2852 5704 2868
rect 5688 2832 5704 2848
rect 5560 2672 5576 2688
rect 5672 2672 5688 2688
rect 5544 2572 5560 2588
rect 5544 2532 5560 2548
rect 5656 2572 5672 2588
rect 5528 2512 5544 2528
rect 5560 2512 5576 2528
rect 5688 2512 5704 2528
rect 5688 2492 5704 2508
rect 5688 2432 5704 2448
rect 5592 2412 5608 2428
rect 5592 2372 5608 2388
rect 5528 2352 5544 2368
rect 5496 2312 5528 2328
rect 5608 2332 5624 2348
rect 5848 3052 5864 3068
rect 5800 2992 5816 3008
rect 5768 2952 5784 2968
rect 5752 2712 5768 2728
rect 5944 3472 5960 3488
rect 5896 3252 5912 3268
rect 5896 3112 5912 3128
rect 5928 3072 5944 3088
rect 5880 3032 5896 3048
rect 5864 2952 5880 2968
rect 5848 2932 5864 2948
rect 5800 2912 5816 2928
rect 5880 2912 5896 2928
rect 5784 2832 5800 2848
rect 5864 2832 5880 2848
rect 5816 2712 5832 2728
rect 5736 2672 5752 2688
rect 5720 2632 5736 2648
rect 5864 2652 5880 2668
rect 5800 2632 5816 2648
rect 5864 2632 5880 2648
rect 5848 2612 5864 2628
rect 5784 2552 5800 2568
rect 5832 2552 5848 2568
rect 5832 2532 5864 2548
rect 5768 2512 5784 2528
rect 5704 2412 5720 2428
rect 5736 2412 5752 2428
rect 5688 2312 5704 2328
rect 5752 2352 5768 2368
rect 5720 2292 5736 2308
rect 5512 2272 5528 2288
rect 5560 2272 5576 2288
rect 5720 2272 5736 2288
rect 5480 2152 5496 2168
rect 5592 2152 5608 2168
rect 5448 2132 5464 2148
rect 5480 2132 5496 2148
rect 5528 2132 5544 2148
rect 5704 2172 5720 2188
rect 5736 2132 5752 2148
rect 5816 2352 5832 2368
rect 5784 2312 5800 2328
rect 5800 2292 5816 2308
rect 5800 2272 5816 2288
rect 5768 2212 5784 2228
rect 5784 2192 5800 2208
rect 5224 2032 5240 2048
rect 5288 2112 5304 2128
rect 5592 2112 5608 2128
rect 5608 2112 5624 2128
rect 5336 2092 5368 2108
rect 5496 2092 5512 2108
rect 5576 2092 5592 2108
rect 5688 2092 5704 2108
rect 5272 2072 5288 2088
rect 5368 2072 5384 2088
rect 5256 1932 5272 1948
rect 5224 1912 5240 1928
rect 5256 1912 5272 1928
rect 5240 1892 5256 1908
rect 5208 1872 5224 1888
rect 5224 1852 5240 1868
rect 5224 1812 5240 1828
rect 5192 1792 5208 1808
rect 5096 1772 5112 1788
rect 5128 1772 5144 1788
rect 5144 1752 5160 1768
rect 5176 1752 5192 1768
rect 5096 1732 5112 1748
rect 5128 1732 5144 1748
rect 5160 1712 5176 1728
rect 4808 1692 4824 1708
rect 4936 1692 4952 1708
rect 4680 1652 4696 1668
rect 4712 1652 4728 1668
rect 4680 1552 4696 1568
rect 4744 1532 4760 1548
rect 4776 1512 4792 1528
rect 4888 1632 4904 1648
rect 5096 1632 5112 1648
rect 4824 1552 4840 1568
rect 4600 1492 4616 1508
rect 4728 1492 4744 1508
rect 4808 1492 4824 1508
rect 4840 1492 4856 1508
rect 4872 1492 4888 1508
rect 4280 1472 4296 1488
rect 4424 1472 4440 1488
rect 4504 1472 4520 1488
rect 4712 1472 4728 1488
rect 4776 1472 4792 1488
rect 4424 1452 4440 1468
rect 4504 1452 4520 1468
rect 4584 1452 4600 1468
rect 4584 1432 4600 1448
rect 4216 1412 4232 1428
rect 4088 1352 4104 1368
rect 4200 1352 4216 1368
rect 4328 1392 4344 1408
rect 4328 1352 4344 1368
rect 3944 1332 3960 1348
rect 4040 1332 4056 1348
rect 4104 1332 4120 1348
rect 3816 1312 3832 1328
rect 3928 1312 3944 1328
rect 3960 1312 3976 1328
rect 3752 1292 3768 1308
rect 3704 1272 3720 1288
rect 3784 1272 3800 1288
rect 3768 1232 3784 1248
rect 3896 1272 3912 1288
rect 3720 1192 3736 1208
rect 3864 1192 3880 1208
rect 3880 1152 3896 1168
rect 3704 1112 3720 1128
rect 4040 1252 4056 1268
rect 3960 1112 3976 1128
rect 3592 1092 3608 1108
rect 3624 1092 3656 1108
rect 3736 1092 3752 1108
rect 3816 1092 3832 1108
rect 3960 1092 3976 1108
rect 3576 1072 3592 1088
rect 3640 1072 3656 1088
rect 3544 1052 3560 1068
rect 3480 1032 3496 1048
rect 3480 992 3512 1008
rect 3448 952 3464 968
rect 3432 932 3448 948
rect 3544 952 3560 968
rect 3576 952 3592 968
rect 3512 932 3528 948
rect 3528 912 3544 928
rect 3560 932 3576 948
rect 3624 912 3640 928
rect 3432 892 3448 908
rect 3480 892 3496 908
rect 3672 1032 3688 1048
rect 3656 1012 3672 1028
rect 3688 972 3704 988
rect 3368 852 3384 868
rect 3640 852 3656 868
rect 3272 632 3288 648
rect 3384 692 3400 708
rect 3368 592 3384 608
rect 3256 532 3272 548
rect 3352 532 3368 548
rect 3128 512 3144 528
rect 3192 512 3208 528
rect 3400 512 3416 528
rect 2568 492 2584 508
rect 2600 492 2616 508
rect 2920 492 2936 508
rect 2952 492 2968 508
rect 3000 492 3016 508
rect 3080 492 3096 508
rect 3144 492 3160 508
rect 2552 432 2568 448
rect 2472 52 2488 68
rect 2536 52 2552 68
rect 2088 12 2104 28
rect 2248 12 2264 28
rect 2376 12 2392 28
rect 2424 12 2440 28
rect 2600 432 2616 448
rect 2680 372 2696 388
rect 2632 312 2648 328
rect 2728 352 2744 368
rect 2776 292 2792 308
rect 2840 306 2856 308
rect 2840 292 2856 306
rect 2600 252 2616 268
rect 2600 172 2616 188
rect 2776 192 2792 208
rect 2840 132 2856 148
rect 2696 112 2712 128
rect 2744 112 2760 128
rect 2808 114 2824 128
rect 2808 112 2824 114
rect 2973 402 3009 418
rect 3048 312 3064 328
rect 2984 292 3000 308
rect 3208 472 3224 488
rect 3384 392 3400 408
rect 3272 352 3288 368
rect 3368 312 3384 328
rect 3160 292 3176 308
rect 3224 306 3240 308
rect 3224 292 3240 306
rect 3352 292 3368 308
rect 2984 232 3000 248
rect 3080 232 3096 248
rect 3640 832 3656 848
rect 3432 792 3448 808
rect 3432 752 3448 768
rect 3560 752 3576 768
rect 3496 732 3512 748
rect 3448 692 3464 708
rect 3624 712 3640 728
rect 3528 672 3544 688
rect 3512 632 3528 648
rect 3576 632 3592 648
rect 3592 612 3608 628
rect 3496 592 3512 608
rect 3528 552 3544 568
rect 3576 552 3592 568
rect 3624 552 3640 568
rect 3688 692 3704 708
rect 3752 1072 3768 1088
rect 3800 1052 3816 1068
rect 3832 1052 3848 1068
rect 3976 1072 3992 1088
rect 3880 1032 3896 1048
rect 3944 1032 3960 1048
rect 3800 972 3816 988
rect 3832 972 3848 988
rect 3981 1002 4017 1018
rect 3784 932 3800 948
rect 3912 912 3928 928
rect 3944 892 3960 908
rect 3864 872 3880 888
rect 3768 812 3784 828
rect 3768 712 3784 728
rect 3944 792 3960 808
rect 3880 732 3896 748
rect 3912 712 3928 728
rect 3816 692 3832 708
rect 3864 692 3880 708
rect 3896 692 3912 708
rect 3800 672 3816 688
rect 3848 672 3864 688
rect 3672 652 3688 668
rect 3784 652 3800 668
rect 3912 652 3928 668
rect 3704 632 3720 648
rect 3848 632 3864 648
rect 3720 592 3736 608
rect 3848 572 3880 588
rect 3832 552 3848 568
rect 3768 532 3784 548
rect 3816 532 3832 548
rect 3640 492 3656 508
rect 3464 432 3480 448
rect 3512 432 3528 448
rect 3960 632 3976 648
rect 3981 602 4017 618
rect 3976 572 3992 588
rect 3768 512 3784 528
rect 3912 512 3928 528
rect 4056 1092 4072 1108
rect 4040 1052 4056 1068
rect 4120 1232 4136 1248
rect 4104 1092 4120 1108
rect 4152 1212 4168 1228
rect 4136 1192 4152 1208
rect 4264 1312 4280 1328
rect 4264 1292 4280 1308
rect 4312 1272 4328 1288
rect 4536 1392 4552 1408
rect 4376 1372 4392 1388
rect 4440 1352 4456 1368
rect 4504 1352 4520 1368
rect 4440 1332 4456 1348
rect 4504 1332 4520 1348
rect 4360 1312 4376 1328
rect 4376 1292 4392 1308
rect 4328 1252 4344 1268
rect 4200 1172 4216 1188
rect 4168 1152 4184 1168
rect 4200 1132 4216 1148
rect 4040 952 4056 968
rect 4072 952 4088 968
rect 4040 732 4056 748
rect 4056 672 4072 688
rect 4120 1052 4136 1068
rect 4152 1052 4168 1068
rect 4184 1052 4200 1068
rect 4136 992 4152 1008
rect 4792 1452 4808 1468
rect 4856 1452 4872 1468
rect 4728 1412 4744 1428
rect 4760 1352 4776 1368
rect 4872 1352 4888 1368
rect 4760 1332 4776 1348
rect 4808 1332 4824 1348
rect 4696 1312 4712 1328
rect 4440 1232 4456 1248
rect 4424 1172 4440 1188
rect 4328 1132 4344 1148
rect 4344 1092 4360 1108
rect 4248 1072 4264 1088
rect 4392 1072 4408 1088
rect 4264 1032 4280 1048
rect 4264 1012 4280 1028
rect 4216 972 4232 988
rect 4200 952 4216 968
rect 4408 1052 4424 1068
rect 4328 972 4344 988
rect 4488 1132 4504 1148
rect 4456 1112 4472 1128
rect 4568 1292 4584 1308
rect 4552 1092 4568 1108
rect 4664 1232 4680 1248
rect 4776 1272 4792 1288
rect 4728 1252 4744 1268
rect 4696 1212 4712 1228
rect 4632 1192 4648 1208
rect 4696 1132 4712 1148
rect 4616 1092 4632 1108
rect 4680 1092 4696 1108
rect 4520 1072 4536 1088
rect 4712 1072 4728 1088
rect 4424 1032 4440 1048
rect 4440 1012 4456 1028
rect 4472 992 4488 1008
rect 4536 992 4552 1008
rect 4344 952 4360 968
rect 4376 952 4392 968
rect 4520 952 4536 968
rect 4280 932 4296 948
rect 4296 932 4312 948
rect 4392 932 4408 948
rect 4456 932 4472 948
rect 4104 732 4120 748
rect 4248 832 4264 848
rect 4136 692 4152 708
rect 4200 712 4216 728
rect 4232 692 4248 708
rect 4264 692 4280 708
rect 4488 832 4504 848
rect 4312 812 4328 828
rect 4392 752 4408 768
rect 4520 772 4536 788
rect 4552 772 4568 788
rect 4552 752 4568 768
rect 4472 712 4488 728
rect 4520 712 4536 728
rect 4328 692 4344 708
rect 4440 692 4456 708
rect 4632 1052 4648 1068
rect 4696 1052 4712 1068
rect 4648 992 4680 1008
rect 4584 932 4600 948
rect 4680 932 4696 948
rect 4856 1172 4872 1188
rect 4824 1152 4840 1168
rect 4792 1092 4808 1108
rect 4744 1076 4760 1088
rect 4744 1072 4760 1076
rect 4760 1052 4776 1068
rect 4808 972 4824 988
rect 4792 932 4808 948
rect 4616 912 4632 928
rect 4648 912 4664 928
rect 4776 912 4792 928
rect 4696 852 4712 868
rect 4584 792 4600 808
rect 4632 712 4648 728
rect 4120 672 4136 688
rect 4312 672 4328 688
rect 4568 672 4584 688
rect 4616 672 4632 688
rect 4648 672 4664 688
rect 4200 652 4216 668
rect 4120 632 4136 648
rect 4184 632 4200 648
rect 4120 612 4136 628
rect 4184 612 4200 628
rect 4056 552 4072 568
rect 4120 552 4136 568
rect 4152 552 4168 568
rect 4056 512 4072 528
rect 4104 492 4120 508
rect 3688 352 3704 368
rect 3528 312 3544 328
rect 3784 312 3800 328
rect 3432 292 3448 308
rect 3496 292 3512 308
rect 3592 306 3608 308
rect 3592 292 3608 306
rect 3928 372 3944 388
rect 4056 332 4072 348
rect 3960 312 3976 328
rect 4072 312 4088 328
rect 3192 252 3208 268
rect 3400 272 3416 288
rect 3512 272 3528 288
rect 3896 272 3912 288
rect 4072 272 4088 288
rect 3416 252 3432 268
rect 3480 252 3496 268
rect 3272 232 3288 248
rect 3560 232 3576 248
rect 3464 192 3480 208
rect 3624 192 3640 208
rect 3192 172 3208 188
rect 3112 152 3128 168
rect 3304 152 3320 168
rect 3352 132 3368 148
rect 3320 112 3336 128
rect 3384 114 3400 128
rect 3752 232 3768 248
rect 3981 202 4017 218
rect 3864 172 3880 188
rect 3752 152 3768 168
rect 3736 132 3752 148
rect 4072 192 4088 208
rect 4088 172 4104 188
rect 4264 632 4280 648
rect 4376 652 4392 668
rect 4584 652 4600 668
rect 4376 632 4392 648
rect 4456 632 4472 648
rect 4312 612 4328 628
rect 4296 572 4312 588
rect 4632 592 4648 608
rect 4232 552 4248 568
rect 4376 552 4392 568
rect 4424 552 4440 568
rect 4744 872 4760 888
rect 4776 772 4792 788
rect 4808 772 4824 788
rect 4776 752 4792 768
rect 4840 1012 4856 1028
rect 5021 1602 5057 1618
rect 5000 1512 5016 1528
rect 5256 1712 5272 1728
rect 5240 1512 5256 1528
rect 5368 2052 5384 2068
rect 5480 2032 5496 2048
rect 5528 1912 5544 1928
rect 5464 1892 5480 1908
rect 5320 1872 5336 1888
rect 5368 1872 5384 1888
rect 5416 1872 5432 1888
rect 5304 1812 5320 1828
rect 5336 1732 5352 1748
rect 5384 1792 5400 1808
rect 5384 1732 5400 1748
rect 5368 1712 5384 1728
rect 5352 1692 5368 1708
rect 5304 1632 5320 1648
rect 5624 2032 5640 2048
rect 5816 2132 5832 2148
rect 5816 2112 5832 2128
rect 5816 2072 5832 2088
rect 5736 1932 5752 1948
rect 5640 1912 5656 1928
rect 5640 1892 5656 1908
rect 5768 1892 5784 1908
rect 5576 1876 5592 1888
rect 5592 1876 5608 1888
rect 5576 1872 5608 1876
rect 5624 1872 5640 1888
rect 5480 1852 5496 1868
rect 5432 1772 5448 1788
rect 5528 1792 5544 1808
rect 5512 1772 5528 1788
rect 5448 1732 5464 1748
rect 5496 1732 5512 1748
rect 5448 1692 5464 1708
rect 5400 1652 5416 1668
rect 5400 1632 5416 1648
rect 5448 1632 5464 1648
rect 5400 1612 5416 1628
rect 5080 1492 5096 1508
rect 5144 1492 5160 1508
rect 4904 1472 4920 1488
rect 4952 1432 4968 1448
rect 4904 1392 4920 1408
rect 5480 1472 5496 1488
rect 5256 1452 5272 1468
rect 5288 1452 5304 1468
rect 5416 1452 5432 1468
rect 4904 1312 4920 1328
rect 4888 1292 4904 1308
rect 5080 1392 5096 1408
rect 5144 1352 5160 1368
rect 5592 1792 5608 1808
rect 5608 1772 5624 1788
rect 5752 1872 5768 1888
rect 5720 1812 5736 1828
rect 5640 1752 5656 1768
rect 5672 1752 5688 1768
rect 5608 1732 5624 1748
rect 5720 1772 5736 1788
rect 5896 2712 5912 2728
rect 5896 2692 5912 2708
rect 5960 3012 5976 3028
rect 5944 2912 5960 2928
rect 5944 2632 5960 2648
rect 5912 2572 5928 2588
rect 5896 2552 5912 2568
rect 5880 2452 5896 2468
rect 5880 2432 5896 2448
rect 5896 2312 5912 2328
rect 5848 2232 5864 2248
rect 5880 2212 5896 2228
rect 5864 2172 5880 2188
rect 5928 2132 5944 2148
rect 5880 2112 5896 2128
rect 5864 1892 5880 1908
rect 5848 1852 5864 1868
rect 5832 1792 5848 1808
rect 5896 1792 5912 1808
rect 5816 1752 5832 1768
rect 5896 1772 5912 1788
rect 5880 1732 5896 1748
rect 5608 1712 5624 1728
rect 5768 1712 5784 1728
rect 5640 1512 5656 1528
rect 5704 1512 5720 1528
rect 5560 1472 5576 1488
rect 5608 1472 5624 1488
rect 5704 1472 5720 1488
rect 5544 1452 5560 1468
rect 5400 1412 5416 1428
rect 5496 1412 5512 1428
rect 5336 1372 5352 1388
rect 5352 1352 5368 1368
rect 5208 1332 5224 1348
rect 5272 1332 5288 1348
rect 5320 1332 5336 1348
rect 5368 1344 5400 1348
rect 5368 1332 5384 1344
rect 5384 1332 5400 1344
rect 5160 1312 5176 1328
rect 5224 1312 5240 1328
rect 5256 1312 5272 1328
rect 5448 1332 5464 1348
rect 5480 1332 5496 1348
rect 5432 1312 5448 1328
rect 5048 1292 5064 1308
rect 5160 1292 5192 1308
rect 5368 1292 5384 1308
rect 4936 1232 4952 1248
rect 5016 1232 5032 1248
rect 4920 1092 4936 1108
rect 4872 1072 4888 1088
rect 4888 1072 4904 1088
rect 4904 992 4920 1008
rect 5021 1202 5057 1218
rect 5096 1172 5112 1188
rect 5096 1132 5112 1148
rect 4952 1092 4968 1108
rect 5000 1092 5016 1108
rect 5288 1232 5304 1248
rect 5288 1192 5304 1208
rect 5224 1152 5240 1168
rect 5176 1132 5192 1148
rect 5240 1112 5256 1128
rect 5160 1092 5176 1108
rect 5176 1072 5192 1088
rect 5032 1032 5048 1048
rect 5048 1032 5064 1048
rect 5128 1012 5144 1028
rect 5048 972 5064 988
rect 5080 972 5096 988
rect 4936 952 4952 968
rect 4984 952 5000 968
rect 4920 912 4936 928
rect 4840 772 4856 788
rect 4904 732 4920 748
rect 4952 712 4968 728
rect 4968 692 4984 708
rect 4728 672 4744 688
rect 4696 652 4712 668
rect 4760 672 4776 688
rect 4760 652 4776 668
rect 4712 592 4728 608
rect 4744 592 4760 608
rect 4680 572 4696 588
rect 4552 552 4568 568
rect 4680 552 4696 568
rect 4328 512 4344 528
rect 4280 472 4296 488
rect 4280 392 4296 408
rect 4312 312 4328 328
rect 4248 292 4264 308
rect 4504 532 4520 548
rect 4488 512 4504 528
rect 4536 512 4552 528
rect 4552 512 4568 528
rect 4520 492 4536 508
rect 4488 472 4504 488
rect 4824 672 4840 688
rect 5528 1392 5544 1408
rect 5672 1432 5688 1448
rect 5544 1372 5560 1388
rect 5464 1292 5480 1308
rect 5512 1292 5528 1308
rect 5416 1132 5432 1148
rect 5240 1072 5256 1088
rect 5400 1072 5416 1088
rect 5448 1072 5464 1088
rect 5176 992 5192 1008
rect 5224 992 5240 1008
rect 5272 972 5288 988
rect 5144 952 5160 968
rect 5320 952 5336 968
rect 5336 952 5352 968
rect 5224 932 5240 948
rect 5320 932 5336 948
rect 5208 912 5224 928
rect 5256 912 5272 928
rect 5021 802 5057 818
rect 5000 732 5016 748
rect 4984 652 5000 668
rect 4904 612 4920 628
rect 4936 612 4952 628
rect 4968 612 4984 628
rect 4872 592 4888 608
rect 4872 572 4904 588
rect 4840 532 4856 548
rect 4776 512 4792 528
rect 4824 512 4840 528
rect 4648 492 4664 508
rect 4616 472 4632 488
rect 4696 452 4712 468
rect 4536 392 4552 408
rect 4440 372 4456 388
rect 4328 292 4344 308
rect 4376 292 4392 308
rect 4264 272 4280 288
rect 4472 332 4488 348
rect 4456 292 4472 308
rect 4344 272 4360 288
rect 4392 272 4408 288
rect 4200 252 4216 268
rect 4328 252 4344 268
rect 4168 232 4184 248
rect 4712 392 4728 408
rect 4760 312 4776 328
rect 4488 292 4504 308
rect 4552 306 4568 308
rect 4552 292 4568 306
rect 4792 272 4808 288
rect 4856 392 4872 408
rect 4824 312 4840 328
rect 4936 552 4952 568
rect 4920 332 4936 348
rect 5128 752 5144 768
rect 5096 732 5112 748
rect 5112 712 5128 728
rect 5064 612 5080 628
rect 5176 692 5192 708
rect 5096 592 5112 608
rect 5288 712 5304 728
rect 5288 692 5320 708
rect 5400 1052 5432 1068
rect 5384 952 5400 968
rect 5416 1012 5432 1028
rect 5512 1212 5528 1228
rect 5480 1112 5496 1128
rect 5576 1352 5592 1368
rect 5656 1352 5672 1368
rect 5896 1692 5912 1708
rect 5800 1512 5816 1528
rect 5800 1492 5816 1508
rect 5752 1476 5768 1488
rect 5752 1472 5768 1476
rect 5784 1472 5800 1488
rect 5736 1452 5752 1468
rect 5720 1412 5736 1428
rect 5688 1344 5720 1348
rect 5688 1332 5704 1344
rect 5704 1332 5720 1344
rect 5592 1312 5608 1328
rect 5544 1292 5560 1308
rect 5608 1232 5624 1248
rect 5560 1152 5576 1168
rect 5608 1152 5624 1168
rect 5528 1132 5544 1148
rect 5672 1112 5688 1128
rect 5624 1092 5640 1108
rect 5704 1092 5720 1108
rect 5576 1052 5592 1068
rect 5544 972 5560 988
rect 5576 1012 5592 1028
rect 5528 952 5544 968
rect 5560 952 5576 968
rect 5448 932 5464 948
rect 5512 932 5528 948
rect 5640 932 5656 948
rect 5416 912 5432 928
rect 5448 912 5464 928
rect 5480 912 5496 928
rect 5560 912 5576 928
rect 5368 772 5384 788
rect 5448 892 5464 908
rect 5384 752 5400 768
rect 5544 752 5560 768
rect 5432 692 5448 708
rect 5320 672 5336 688
rect 5416 676 5432 688
rect 5416 672 5432 676
rect 5464 672 5480 688
rect 5240 652 5256 668
rect 5288 652 5304 668
rect 5208 632 5224 648
rect 5208 592 5224 608
rect 5240 592 5256 608
rect 5112 572 5128 588
rect 5000 532 5016 548
rect 5096 532 5112 548
rect 5224 532 5240 548
rect 5080 512 5096 528
rect 5144 512 5160 528
rect 5224 472 5240 488
rect 5021 402 5057 418
rect 5160 412 5176 428
rect 5160 372 5176 388
rect 5016 352 5032 368
rect 4968 332 4984 348
rect 4952 312 4968 328
rect 5000 312 5016 328
rect 4936 292 4952 308
rect 4392 252 4408 268
rect 4216 192 4232 208
rect 4376 192 4392 208
rect 4136 172 4152 188
rect 4744 252 4760 268
rect 4808 252 4824 268
rect 4616 212 4632 228
rect 4680 212 4696 228
rect 4264 152 4280 168
rect 4520 152 4536 168
rect 4072 132 4088 148
rect 3384 112 3400 114
rect 3672 112 3688 128
rect 3720 112 3736 128
rect 3896 114 3912 128
rect 3896 112 3912 114
rect 3928 112 3944 128
rect 4104 112 4120 128
rect 4232 112 4248 128
rect 4296 114 4312 128
rect 4296 112 4312 114
rect 4632 172 4648 188
rect 4680 152 4696 168
rect 4824 152 4840 168
rect 4952 212 4968 228
rect 5112 332 5128 348
rect 5144 332 5160 348
rect 5272 572 5288 588
rect 5304 632 5320 648
rect 5336 592 5352 608
rect 5400 552 5416 568
rect 5416 532 5432 548
rect 5320 512 5336 528
rect 5352 512 5368 528
rect 5240 312 5256 328
rect 5288 292 5304 308
rect 5640 752 5656 768
rect 5640 732 5656 748
rect 5688 1072 5704 1088
rect 5720 972 5736 988
rect 5720 952 5736 968
rect 5752 1372 5768 1388
rect 5816 1372 5832 1388
rect 5848 1372 5864 1388
rect 5784 1312 5800 1328
rect 5912 1492 5928 1508
rect 5880 1432 5896 1448
rect 5912 1432 5928 1448
rect 5800 1252 5816 1268
rect 5848 1252 5880 1268
rect 5800 1232 5816 1248
rect 5752 1112 5768 1128
rect 5752 972 5784 988
rect 5704 932 5720 948
rect 5736 932 5752 948
rect 5672 692 5688 708
rect 5496 672 5512 688
rect 5496 572 5512 588
rect 5528 592 5544 608
rect 5528 572 5560 588
rect 5512 552 5528 568
rect 5656 672 5672 688
rect 5816 1072 5832 1088
rect 5800 952 5816 968
rect 5832 1012 5848 1028
rect 5832 952 5848 968
rect 5864 1112 5880 1128
rect 5864 1092 5880 1108
rect 5896 1344 5912 1348
rect 5896 1332 5912 1344
rect 5896 1292 5912 1308
rect 5880 1072 5896 1088
rect 5912 1076 5928 1088
rect 5912 1072 5928 1076
rect 5864 1032 5880 1048
rect 5816 712 5832 728
rect 5736 676 5752 688
rect 5736 672 5752 676
rect 5720 652 5736 668
rect 5752 652 5768 668
rect 5608 612 5624 628
rect 5608 552 5624 568
rect 5720 612 5736 628
rect 5704 552 5736 568
rect 5768 572 5784 588
rect 5736 532 5752 548
rect 5432 312 5448 328
rect 5320 292 5336 308
rect 5384 292 5400 308
rect 5112 272 5128 288
rect 5112 192 5128 208
rect 5560 432 5576 448
rect 5736 432 5752 448
rect 5608 412 5624 428
rect 5592 392 5608 408
rect 5496 292 5512 308
rect 5576 292 5592 308
rect 5624 392 5640 408
rect 5768 332 5784 348
rect 5192 276 5224 288
rect 5192 272 5208 276
rect 5208 272 5224 276
rect 5464 272 5480 288
rect 5624 276 5640 288
rect 5624 272 5640 276
rect 5688 272 5704 288
rect 5752 276 5768 288
rect 5752 272 5768 276
rect 5480 252 5496 268
rect 5592 252 5608 268
rect 5672 252 5688 268
rect 5240 232 5256 248
rect 5224 212 5240 228
rect 5272 192 5288 208
rect 5064 172 5080 188
rect 5128 172 5144 188
rect 5208 172 5224 188
rect 4920 132 4936 148
rect 4968 132 4984 148
rect 5144 132 5160 148
rect 4648 112 4664 128
rect 4712 114 4728 128
rect 5352 192 5368 208
rect 5336 172 5352 188
rect 5320 152 5336 168
rect 5544 192 5560 208
rect 5576 192 5592 208
rect 5384 152 5400 168
rect 5512 152 5544 168
rect 5352 132 5368 148
rect 5400 132 5416 148
rect 5592 172 5608 188
rect 5608 152 5624 168
rect 5704 212 5720 228
rect 5720 172 5736 188
rect 5960 2112 5976 2128
rect 5992 2772 6008 2788
rect 5976 1972 5992 1988
rect 5960 1472 5976 1488
rect 5960 1452 5976 1468
rect 5944 972 5960 988
rect 5896 932 5912 948
rect 5832 672 5848 688
rect 5816 652 5832 668
rect 5800 572 5816 588
rect 5944 772 5960 788
rect 5912 712 5928 728
rect 5896 692 5912 708
rect 5912 672 5928 688
rect 5880 652 5896 668
rect 5880 592 5896 608
rect 5864 552 5880 568
rect 5848 532 5864 548
rect 5800 332 5816 348
rect 5928 572 5944 588
rect 5864 372 5880 388
rect 5976 352 5992 368
rect 5928 312 5944 328
rect 5880 292 5896 308
rect 5944 292 5960 308
rect 5896 232 5912 248
rect 5784 192 5800 208
rect 5832 192 5848 208
rect 5784 172 5800 188
rect 5944 152 5960 168
rect 5736 132 5752 148
rect 5928 132 5944 148
rect 4712 112 4728 114
rect 5000 112 5016 128
rect 5080 112 5112 128
rect 5416 112 5432 128
rect 5448 112 5464 128
rect 5544 112 5560 128
rect 5864 112 5880 128
rect 3240 92 3256 108
rect 5528 92 5544 108
rect 5800 92 5816 108
rect 2973 2 3009 18
rect 3112 12 3128 28
rect 3208 12 3224 28
rect 3672 32 3688 48
rect 3656 12 3672 28
rect 3688 12 3720 28
rect 3736 12 3752 28
rect 3784 12 3800 28
rect 4536 12 4552 28
rect 4568 12 4584 28
rect 5021 2 5057 18
<< metal3 >>
rect 408 4017 472 4023
rect 504 4017 792 4023
rect 2232 4017 2248 4023
rect 2120 3997 2248 4003
rect 3656 4017 3992 4023
rect 4056 4017 4072 4023
rect 4088 4017 4120 4023
rect 4184 4017 4216 4023
rect 3592 3997 3608 4003
rect 3736 3997 4360 4003
rect 728 3977 888 3983
rect 904 3977 2024 3983
rect 2216 3977 2648 3983
rect 2888 3977 3608 3983
rect 3688 3977 3752 3983
rect 3896 3977 3960 3983
rect 4280 3977 4312 3983
rect 1160 3957 1192 3963
rect 1208 3957 1352 3963
rect 1368 3957 2504 3963
rect 2584 3957 3400 3963
rect 3816 3957 5048 3963
rect 1224 3937 1592 3943
rect 1928 3937 2008 3943
rect 2040 3937 2440 3943
rect 3256 3937 3320 3943
rect 3352 3937 3384 3943
rect 4840 3937 5128 3943
rect 216 3917 344 3923
rect 360 3917 536 3923
rect 552 3917 968 3923
rect 1064 3917 2088 3923
rect 2104 3917 2136 3923
rect 2168 3917 2296 3923
rect 2312 3917 2328 3923
rect 2360 3917 2392 3923
rect 2536 3917 2584 3923
rect 2600 3917 3080 3923
rect 3096 3917 4856 3923
rect 4872 3917 4952 3923
rect 4968 3917 5064 3923
rect 504 3897 584 3903
rect 600 3897 648 3903
rect 1192 3897 1203 3903
rect 1336 3897 1416 3903
rect 1608 3897 1656 3903
rect 1672 3897 2120 3903
rect 2184 3897 2232 3903
rect 2248 3897 2264 3903
rect 2280 3897 2376 3903
rect 2392 3897 2456 3903
rect 2472 3897 2536 3903
rect 2552 3897 2632 3903
rect 2648 3897 2744 3903
rect 2760 3897 2840 3903
rect 2856 3897 2920 3903
rect 3064 3897 3160 3903
rect 3176 3897 3288 3903
rect 3320 3897 3432 3903
rect 3512 3897 3576 3903
rect 3640 3897 3656 3903
rect 3768 3897 3896 3903
rect 4008 3897 4088 3903
rect 4120 3897 4200 3903
rect 4216 3897 4296 3903
rect 4317 3897 4440 3903
rect 941 3888 947 3892
rect 3725 3888 3731 3892
rect 317 3877 328 3883
rect 408 3877 440 3883
rect 456 3877 936 3883
rect 1192 3877 1224 3883
rect 1288 3877 1336 3883
rect 1400 3877 1448 3883
rect 1480 3877 1528 3883
rect 1544 3877 1624 3883
rect 1784 3877 1832 3883
rect 1864 3877 2008 3883
rect 2024 3877 2200 3883
rect 2568 3877 2680 3883
rect 2744 3877 2776 3883
rect 2856 3877 2872 3883
rect 2920 3877 2952 3883
rect 3208 3877 3320 3883
rect 3400 3877 3448 3883
rect 3560 3877 3640 3883
rect 3784 3877 3880 3883
rect 3896 3877 3944 3883
rect 3992 3877 4248 3883
rect 4317 3883 4323 3897
rect 4504 3897 4552 3903
rect 4568 3897 4680 3903
rect 4696 3897 4872 3903
rect 4888 3897 5000 3903
rect 5112 3897 5160 3903
rect 5304 3897 5320 3903
rect 5352 3897 5608 3903
rect 4280 3877 4323 3883
rect 4440 3877 4600 3883
rect 4616 3877 4744 3883
rect 4760 3877 4808 3883
rect 4824 3877 4920 3883
rect 5160 3877 5240 3883
rect 5256 3877 5384 3883
rect 5448 3877 5480 3883
rect 5640 3877 5656 3883
rect 5672 3877 5688 3883
rect 88 3857 360 3863
rect 424 3857 520 3863
rect 552 3857 952 3863
rect 968 3857 1128 3863
rect 1144 3857 1208 3863
rect 1224 3857 2872 3863
rect 3336 3857 3592 3863
rect 3656 3857 3848 3863
rect 3864 3857 4008 3863
rect 4024 3857 4040 3863
rect 4088 3857 4504 3863
rect 4536 3857 4568 3863
rect 4600 3857 4696 3863
rect 4712 3857 4824 3863
rect 4840 3857 5288 3863
rect 5320 3857 5368 3863
rect 5384 3857 5560 3863
rect 5688 3857 5736 3863
rect 216 3837 456 3843
rect 696 3837 744 3843
rect 824 3837 904 3843
rect 936 3837 1400 3843
rect 1416 3837 1720 3843
rect 1752 3837 2664 3843
rect 2680 3837 3000 3843
rect 3016 3837 4184 3843
rect 4328 3837 4424 3843
rect 4520 3837 5176 3843
rect 5192 3837 5672 3843
rect 392 3817 552 3823
rect 648 3817 824 3823
rect 840 3817 1096 3823
rect 1208 3817 1267 3823
rect 40 3797 136 3803
rect 184 3797 296 3803
rect 312 3797 360 3803
rect 376 3797 776 3803
rect 792 3797 1032 3803
rect 1048 3797 1240 3803
rect 1261 3803 1267 3817
rect 1528 3817 1640 3823
rect 1672 3817 1800 3823
rect 1261 3797 1352 3803
rect 1416 3797 1480 3803
rect 1528 3797 1864 3803
rect 2440 3817 2616 3823
rect 3048 3817 3112 3823
rect 3128 3817 3176 3823
rect 3192 3817 3336 3823
rect 3352 3817 3368 3823
rect 3464 3817 3528 3823
rect 2136 3797 2488 3803
rect 3096 3797 3144 3803
rect 3320 3797 3720 3803
rect 3736 3797 3864 3803
rect 4392 3817 4456 3823
rect 4648 3817 4712 3823
rect 4808 3817 4840 3823
rect 4872 3817 4888 3823
rect 4904 3817 5544 3823
rect 4029 3797 4328 3803
rect 328 3777 392 3783
rect 872 3777 968 3783
rect 1256 3777 2120 3783
rect 2376 3777 2696 3783
rect 2984 3777 3656 3783
rect 4029 3783 4035 3797
rect 4360 3797 4520 3803
rect 4728 3797 4920 3803
rect 4936 3797 4968 3803
rect 3704 3777 4035 3783
rect 4264 3777 4760 3783
rect 4776 3777 5064 3783
rect 5080 3777 5160 3783
rect 5176 3777 5224 3783
rect 5528 3777 5640 3783
rect 56 3757 168 3763
rect 184 3757 216 3763
rect 232 3757 424 3763
rect 440 3757 632 3763
rect 696 3757 744 3763
rect 792 3757 824 3763
rect 984 3757 1064 3763
rect 1160 3757 1688 3763
rect 1784 3757 1864 3763
rect 1912 3757 1992 3763
rect 2008 3757 2552 3763
rect 2920 3757 3000 3763
rect 3016 3757 3320 3763
rect 3336 3757 3416 3763
rect 3544 3757 3688 3763
rect 3960 3757 4104 3763
rect 4200 3757 4712 3763
rect 5240 3757 5256 3763
rect 5304 3757 5320 3763
rect 5448 3757 5496 3763
rect 5624 3757 5704 3763
rect 5752 3757 5832 3763
rect 4829 3748 4835 3752
rect 4845 3748 4851 3752
rect 520 3737 552 3743
rect 616 3737 632 3743
rect 808 3737 856 3743
rect 888 3737 1320 3743
rect 1464 3737 1576 3743
rect 1592 3737 1832 3743
rect 1960 3737 1971 3743
rect 1981 3737 2072 3743
rect 200 3717 872 3723
rect 952 3717 1016 3723
rect 1037 3717 1048 3723
rect 1096 3717 1128 3723
rect 1288 3717 1560 3723
rect 1592 3717 1640 3723
rect 1656 3717 1704 3723
rect 1736 3717 1848 3723
rect 1864 3717 1896 3723
rect 1981 3723 1987 3737
rect 2088 3737 2312 3743
rect 2328 3737 2360 3743
rect 3432 3737 3544 3743
rect 3688 3737 3816 3743
rect 4264 3737 4344 3743
rect 4456 3737 4536 3743
rect 4920 3737 5464 3743
rect 5512 3737 5688 3743
rect 5704 3737 5752 3743
rect 5800 3737 5912 3743
rect 3309 3728 3315 3732
rect 1928 3717 1987 3723
rect 2008 3717 2088 3723
rect 2232 3717 2296 3723
rect 2312 3717 2472 3723
rect 2632 3717 2728 3723
rect 3000 3717 3016 3723
rect 3032 3717 3256 3723
rect 3480 3717 3496 3723
rect 3528 3717 3768 3723
rect 3864 3717 3928 3723
rect 3960 3717 4008 3723
rect 4024 3717 4648 3723
rect 4664 3717 4984 3723
rect 5432 3717 5624 3723
rect 104 3697 568 3703
rect 904 3697 1080 3703
rect 1112 3697 1144 3703
rect 1480 3697 1592 3703
rect 1608 3697 1928 3703
rect 2136 3697 2168 3703
rect 2344 3697 2424 3703
rect 2712 3697 2744 3703
rect 2760 3697 2931 3703
rect 744 3677 824 3683
rect 1080 3677 1112 3683
rect 1352 3677 2696 3683
rect 2728 3677 2840 3683
rect 2925 3683 2931 3697
rect 3320 3697 3368 3703
rect 3416 3697 3528 3703
rect 3656 3697 3672 3703
rect 3768 3697 3784 3703
rect 3981 3697 4520 3703
rect 2925 3677 3592 3683
rect 3688 3677 3704 3683
rect 3981 3683 3987 3697
rect 4696 3697 4888 3703
rect 5416 3697 5448 3703
rect 3896 3677 3987 3683
rect 4104 3677 4712 3683
rect 5064 3677 5496 3683
rect 264 3657 1160 3663
rect 2072 3657 2104 3663
rect 2120 3657 2328 3663
rect 2360 3657 3592 3663
rect 3640 3657 3752 3663
rect 3768 3657 4024 3663
rect 4600 3657 5192 3663
rect 744 3637 808 3643
rect 856 3637 1480 3643
rect 1560 3637 1736 3643
rect 1864 3637 2152 3643
rect 2520 3637 3128 3643
rect 3368 3637 3416 3643
rect 3608 3637 4120 3643
rect 4664 3637 4840 3643
rect 5112 3637 5128 3643
rect 5848 3637 5864 3643
rect 536 3617 872 3623
rect 1032 3617 1304 3623
rect 1576 3617 2184 3623
rect 2136 3597 2312 3603
rect 2328 3597 2408 3603
rect 2424 3597 2472 3603
rect 2504 3597 2744 3603
rect 2856 3597 2872 3603
rect 3080 3617 3464 3623
rect 3752 3617 4584 3623
rect 3288 3597 3736 3603
rect 3800 3597 4792 3603
rect 5816 3617 5912 3623
rect 5736 3597 5880 3603
rect 584 3577 2200 3583
rect 2232 3577 2280 3583
rect 2552 3577 2856 3583
rect 2904 3577 3352 3583
rect 3384 3577 3992 3583
rect 4008 3577 5256 3583
rect 648 3557 840 3563
rect 1048 3557 1256 3563
rect 1272 3557 1448 3563
rect 1464 3557 1528 3563
rect 1880 3557 2568 3563
rect 2664 3557 2776 3563
rect 2792 3557 3208 3563
rect 3240 3557 4200 3563
rect 4536 3557 4664 3563
rect 5208 3557 5752 3563
rect 472 3537 1352 3543
rect 1416 3537 1608 3543
rect 2056 3537 2376 3543
rect 2488 3537 2552 3543
rect 2584 3537 2728 3543
rect 2744 3537 2872 3543
rect 2888 3537 3672 3543
rect 4344 3537 5336 3543
rect 56 3517 168 3523
rect 184 3517 424 3523
rect 632 3517 1032 3523
rect 1176 3517 1560 3523
rect 1816 3517 1864 3523
rect 2200 3517 2360 3523
rect 2536 3517 2792 3523
rect 2888 3517 3080 3523
rect 3096 3517 3288 3523
rect 3304 3517 3480 3523
rect 3512 3517 3720 3523
rect 3736 3517 4008 3523
rect 4216 3517 4376 3523
rect 4392 3517 4488 3523
rect 4520 3517 4552 3523
rect 4568 3517 4616 3523
rect 4648 3517 4728 3523
rect 5224 3517 5240 3523
rect 5336 3517 5528 3523
rect 5640 3517 5704 3523
rect 5720 3517 5832 3523
rect 200 3497 328 3503
rect 440 3497 552 3503
rect 568 3497 616 3503
rect 680 3497 856 3503
rect 1000 3497 1096 3503
rect 1160 3497 1240 3503
rect 1352 3497 1416 3503
rect 1672 3497 1704 3503
rect 1720 3497 1784 3503
rect 1800 3497 1896 3503
rect 2008 3497 2232 3503
rect 2280 3497 2328 3503
rect 2392 3497 2424 3503
rect 2440 3497 2488 3503
rect 2504 3497 2600 3503
rect 2760 3497 3112 3503
rect 3192 3497 3256 3503
rect 3448 3497 3944 3503
rect 4008 3497 4072 3503
rect 4216 3497 4392 3503
rect 4456 3497 4568 3503
rect 4584 3497 4680 3503
rect 4696 3497 4760 3503
rect 4824 3497 5112 3503
rect 5256 3497 5336 3503
rect 5352 3497 5384 3503
rect 5480 3497 5592 3503
rect 5720 3497 5864 3503
rect 72 3477 248 3483
rect 584 3477 648 3483
rect 664 3477 936 3483
rect 1112 3477 1336 3483
rect 1368 3477 1400 3483
rect 1592 3477 1720 3483
rect 1736 3477 1832 3483
rect 2376 3477 2440 3483
rect 2456 3477 2536 3483
rect 2616 3477 2664 3483
rect 2808 3477 2856 3483
rect 2872 3477 2952 3483
rect 3256 3477 3304 3483
rect 3336 3477 3416 3483
rect 3512 3477 3528 3483
rect 3981 3477 4136 3483
rect 120 3457 344 3463
rect 360 3457 792 3463
rect 808 3457 824 3463
rect 840 3457 1096 3463
rect 1304 3457 1656 3463
rect 1688 3457 1736 3463
rect 1944 3457 2520 3463
rect 2536 3457 2920 3463
rect 3000 3457 3336 3463
rect 3432 3457 3464 3463
rect 3528 3457 3592 3463
rect 3981 3463 3987 3477
rect 4168 3477 4264 3483
rect 4328 3477 4408 3483
rect 4472 3477 4536 3483
rect 4728 3477 4904 3483
rect 4968 3477 5048 3483
rect 5128 3477 5240 3483
rect 5256 3477 5304 3483
rect 5320 3477 5400 3483
rect 5592 3477 5656 3483
rect 5704 3477 5816 3483
rect 5880 3477 5944 3483
rect 3720 3457 3987 3463
rect 4008 3457 4472 3463
rect 4488 3457 4776 3463
rect 5272 3457 5352 3463
rect 5384 3457 5672 3463
rect 5688 3457 5720 3463
rect 248 3437 280 3443
rect 296 3437 472 3443
rect 488 3437 664 3443
rect 1144 3437 1176 3443
rect 1240 3437 1304 3443
rect 1752 3437 2216 3443
rect 2248 3437 2552 3443
rect 2584 3437 2808 3443
rect 2824 3437 3032 3443
rect 3128 3437 3139 3443
rect 3176 3437 4200 3443
rect 5453 3428 5459 3432
rect 632 3417 1192 3423
rect 1640 3417 1656 3423
rect 1736 3417 1752 3423
rect 264 3397 392 3403
rect 568 3397 584 3403
rect 680 3397 712 3403
rect 936 3397 968 3403
rect 1080 3397 1272 3403
rect 1352 3397 1576 3403
rect 1592 3397 1752 3403
rect 2008 3417 2024 3423
rect 2296 3417 2568 3423
rect 2840 3417 2936 3423
rect 2968 3417 3192 3423
rect 3448 3417 3480 3423
rect 3496 3417 3512 3423
rect 3640 3417 3928 3423
rect 2712 3397 2728 3403
rect 2760 3397 2968 3403
rect 3192 3397 3800 3403
rect 4120 3417 4184 3423
rect 4200 3417 4360 3423
rect 4632 3417 4808 3423
rect 4872 3417 4920 3423
rect 5544 3417 5688 3423
rect 4264 3397 4296 3403
rect 4712 3397 4808 3403
rect 4824 3397 5080 3403
rect 5096 3397 5176 3403
rect 72 3377 120 3383
rect 136 3377 392 3383
rect 456 3377 632 3383
rect 872 3377 1416 3383
rect 1432 3377 1976 3383
rect 2120 3377 2131 3383
rect 2312 3377 2328 3383
rect 2344 3377 2872 3383
rect 2888 3377 3768 3383
rect 3960 3377 4040 3383
rect 4072 3377 4392 3383
rect 4408 3377 4568 3383
rect 4584 3377 5560 3383
rect 392 3357 568 3363
rect 792 3357 1672 3363
rect 1864 3357 1880 3363
rect 2072 3357 2136 3363
rect 2184 3357 2824 3363
rect 2840 3357 3096 3363
rect 3128 3357 3176 3363
rect 3224 3357 3272 3363
rect 3608 3357 3624 3363
rect 3784 3357 3880 3363
rect 3912 3357 4104 3363
rect 4200 3357 4216 3363
rect 4280 3357 4456 3363
rect 4600 3357 4632 3363
rect 4680 3357 4696 3363
rect 4760 3357 4840 3363
rect 5048 3357 5144 3363
rect 5192 3357 5272 3363
rect 5352 3357 5400 3363
rect 5624 3357 5640 3363
rect 40 3337 72 3343
rect 216 3337 232 3343
rect 392 3337 728 3343
rect 824 3337 1032 3343
rect 1064 3337 1096 3343
rect 1128 3337 1160 3343
rect 1389 3337 1400 3343
rect 1528 3337 1544 3343
rect 1624 3337 1640 3343
rect 2104 3337 2344 3343
rect 2600 3337 3016 3343
rect 3048 3337 3448 3343
rect 3464 3337 4600 3343
rect 4632 3337 4824 3343
rect 4840 3337 4904 3343
rect 4968 3337 5000 3343
rect 5032 3337 5064 3343
rect 5128 3337 5160 3343
rect 5224 3337 5304 3343
rect 5320 3337 5336 3343
rect 5464 3337 5512 3343
rect 5576 3337 5800 3343
rect 840 3317 872 3323
rect 904 3317 1064 3323
rect 1192 3317 1224 3323
rect 1496 3317 1528 3323
rect 1800 3317 1960 3323
rect 1976 3317 2008 3323
rect 2280 3317 2712 3323
rect 3032 3317 3144 3323
rect 3160 3317 3368 3323
rect 3592 3317 3672 3323
rect 3704 3317 3864 3323
rect 3912 3317 4056 3323
rect 4072 3317 4104 3323
rect 4136 3317 4312 3323
rect 4392 3317 4440 3323
rect 4456 3317 4536 3323
rect 4568 3317 4680 3323
rect 4696 3317 4872 3323
rect 4888 3317 4920 3323
rect 5304 3317 5368 3323
rect 5384 3317 5592 3323
rect 5608 3317 5688 3323
rect 5784 3317 5864 3323
rect 824 3297 1320 3303
rect 1336 3297 1592 3303
rect 1704 3297 2216 3303
rect 2232 3297 2568 3303
rect 2632 3297 3155 3303
rect 376 3277 392 3283
rect 424 3277 744 3283
rect 760 3277 776 3283
rect 792 3277 1048 3283
rect 1064 3277 1448 3283
rect 1464 3277 1496 3283
rect 2136 3277 2360 3283
rect 2408 3277 2616 3283
rect 2872 3277 3128 3283
rect 3149 3283 3155 3297
rect 3224 3297 3656 3303
rect 3672 3297 3816 3303
rect 4056 3297 4184 3303
rect 4328 3297 4584 3303
rect 5080 3297 5512 3303
rect 5736 3297 5800 3303
rect 3149 3277 3496 3283
rect 3544 3277 4536 3283
rect 5016 3277 5192 3283
rect 5272 3277 5448 3283
rect 2104 3257 2296 3263
rect 2376 3257 3448 3263
rect 3640 3257 3736 3263
rect 4200 3257 4296 3263
rect 4312 3257 4440 3263
rect 4792 3257 5096 3263
rect 856 3237 1080 3243
rect 1336 3237 1464 3243
rect 1480 3237 1592 3243
rect 1608 3237 1800 3243
rect 1928 3237 2136 3243
rect 2520 3237 2648 3243
rect 2760 3237 2904 3243
rect 3112 3237 3160 3243
rect 3208 3237 3784 3243
rect 4488 3237 5128 3243
rect 5229 3228 5235 3232
rect 72 3217 568 3223
rect 600 3217 904 3223
rect 1976 3217 2504 3223
rect 973 3197 1992 3203
rect 973 3183 979 3197
rect 2024 3197 2840 3203
rect 3032 3217 3176 3223
rect 3464 3217 3784 3223
rect 4392 3217 4984 3223
rect 3144 3197 3384 3203
rect 3416 3197 3560 3203
rect 3752 3197 4216 3203
rect 4568 3197 4712 3203
rect 5336 3217 5720 3223
rect 5128 3197 5416 3203
rect 5448 3197 5656 3203
rect 776 3177 979 3183
rect 1176 3177 2424 3183
rect 2488 3177 2712 3183
rect 3192 3177 3768 3183
rect 3784 3177 3864 3183
rect 3880 3177 3912 3183
rect 3992 3177 4568 3183
rect 4920 3177 5688 3183
rect 648 3157 1368 3163
rect 1496 3157 2984 3163
rect 3000 3157 3480 3163
rect 3496 3157 4056 3163
rect 4536 3157 4664 3163
rect 4712 3157 5416 3163
rect 5432 3157 5688 3163
rect 1384 3137 1528 3143
rect 1672 3137 2488 3143
rect 2856 3137 3176 3143
rect 3272 3137 3656 3143
rect 3784 3137 3896 3143
rect 3976 3137 4200 3143
rect 4552 3137 5608 3143
rect 376 3117 888 3123
rect 904 3117 1128 3123
rect 1160 3117 1288 3123
rect 1464 3117 1480 3123
rect 1624 3117 1880 3123
rect 1912 3117 2024 3123
rect 2136 3117 2248 3123
rect 2264 3117 2392 3123
rect 2440 3117 2520 3123
rect 2824 3117 3080 3123
rect 3256 3117 3416 3123
rect 3432 3117 3480 3123
rect 3736 3117 4120 3123
rect 4152 3117 4344 3123
rect 4472 3117 4600 3123
rect 4664 3117 4760 3123
rect 4840 3117 4904 3123
rect 5656 3117 5896 3123
rect 296 3097 328 3103
rect 456 3097 552 3103
rect 1128 3097 1176 3103
rect 1304 3097 1384 3103
rect 1400 3097 1496 3103
rect 1512 3097 1544 3103
rect 1560 3097 1608 3103
rect 1656 3097 1736 3103
rect 2248 3097 2296 3103
rect 2312 3097 2328 3103
rect 2344 3097 2488 3103
rect 2504 3097 2600 3103
rect 2616 3097 3080 3103
rect 3096 3097 3144 3103
rect 3160 3097 3208 3103
rect 3224 3097 3256 3103
rect 3352 3097 3400 3103
rect 3416 3097 3448 3103
rect 3848 3097 3976 3103
rect 4264 3097 4392 3103
rect 4440 3097 4616 3103
rect 4712 3097 4808 3103
rect 4824 3097 4888 3103
rect 4904 3097 4936 3103
rect 4952 3097 5176 3103
rect 4205 3088 4211 3092
rect 232 3077 264 3083
rect 504 3077 616 3083
rect 1112 3077 1160 3083
rect 1192 3077 1208 3083
rect 1240 3077 1256 3083
rect 1288 3077 1512 3083
rect 1544 3077 1656 3083
rect 1880 3077 1944 3083
rect 1960 3077 2104 3083
rect 2120 3077 2168 3083
rect 2200 3077 2312 3083
rect 2328 3077 2360 3083
rect 2392 3077 3016 3083
rect 3176 3077 3352 3083
rect 3368 3077 3384 3083
rect 3448 3077 3480 3083
rect 3752 3077 3955 3083
rect 104 3057 488 3063
rect 632 3057 872 3063
rect 888 3057 968 3063
rect 984 3057 1080 3063
rect 1096 3057 1192 3063
rect 1544 3057 1800 3063
rect 1816 3057 1976 3063
rect 1992 3057 2024 3063
rect 2712 3057 2744 3063
rect 2765 3057 3128 3063
rect 392 3037 600 3043
rect 632 3037 648 3043
rect 664 3037 744 3043
rect 840 3037 1352 3043
rect 1768 3037 1832 3043
rect 2765 3043 2771 3057
rect 3576 3057 3832 3063
rect 3949 3063 3955 3077
rect 3976 3077 4168 3083
rect 4344 3077 4456 3083
rect 4520 3077 4536 3083
rect 4600 3077 4904 3083
rect 5224 3077 5272 3083
rect 5517 3077 5528 3083
rect 5608 3077 5672 3083
rect 5688 3077 5720 3083
rect 5736 3077 5784 3083
rect 5832 3077 5928 3083
rect 3949 3057 4216 3063
rect 4328 3057 4568 3063
rect 5800 3057 5848 3063
rect 2584 3037 2771 3043
rect 3064 3037 3112 3043
rect 3160 3037 3224 3043
rect 3533 3037 3544 3043
rect 3816 3037 3832 3043
rect 3933 3037 4968 3043
rect 56 3017 168 3023
rect 184 3017 376 3023
rect 888 3017 904 3023
rect 1672 3017 1880 3023
rect 1896 3017 1912 3023
rect 200 2997 328 3003
rect 392 2997 435 3003
rect 24 2977 88 2983
rect 136 2977 232 2983
rect 328 2977 408 2983
rect 429 2983 435 2997
rect 520 2997 840 3003
rect 1192 2997 1416 3003
rect 1432 2997 1640 3003
rect 1656 2997 1672 3003
rect 1736 2997 1891 3003
rect 2376 3017 2392 3023
rect 2808 3017 2904 3023
rect 2920 3017 3272 3023
rect 3933 3023 3939 3037
rect 5720 3037 5880 3043
rect 5965 3028 5971 3032
rect 3656 3017 3939 3023
rect 429 2977 584 2983
rect 1224 2977 1336 2983
rect 1656 2977 1864 2983
rect 1885 2983 1891 2997
rect 2152 2997 2200 3003
rect 2536 2997 2712 3003
rect 2872 2997 2936 3003
rect 2952 2997 3512 3003
rect 3544 2997 3848 3003
rect 3864 2997 3960 3003
rect 4200 3017 4552 3023
rect 4584 3017 4744 3023
rect 4760 3017 5000 3023
rect 5432 3017 5544 3023
rect 5592 3017 5608 3023
rect 4184 2997 4312 3003
rect 4456 2997 4488 3003
rect 4520 2997 4696 3003
rect 4984 2997 5192 3003
rect 5208 2997 5384 3003
rect 5400 2997 5800 3003
rect 1885 2977 1928 2983
rect 1944 2977 2216 2983
rect 2680 2977 2776 2983
rect 2792 2977 3176 2983
rect 3768 2977 3816 2983
rect 3832 2977 4024 2983
rect 4056 2977 4712 2983
rect 4728 2977 4872 2983
rect 4888 2977 5347 2983
rect 72 2957 120 2963
rect 152 2957 168 2963
rect 328 2957 632 2963
rect 680 2957 776 2963
rect 968 2957 1000 2963
rect 1064 2957 1352 2963
rect 1384 2957 1672 2963
rect 1800 2957 1848 2963
rect 2216 2957 2280 2963
rect 2328 2957 2344 2963
rect 2504 2957 2552 2963
rect 2568 2957 2584 2963
rect 2600 2957 2680 2963
rect 2696 2957 2760 2963
rect 2792 2957 2888 2963
rect 2904 2957 3016 2963
rect 3032 2957 3112 2963
rect 3133 2957 3208 2963
rect 24 2937 184 2943
rect 264 2937 392 2943
rect 408 2937 456 2943
rect 472 2937 520 2943
rect 536 2937 952 2943
rect 1176 2937 1224 2943
rect 1240 2937 2472 2943
rect 2728 2937 2808 2943
rect 3133 2943 3139 2957
rect 3512 2957 3544 2963
rect 3576 2957 3912 2963
rect 3976 2957 4088 2963
rect 4136 2957 4152 2963
rect 4328 2957 4472 2963
rect 4632 2957 4680 2963
rect 4712 2957 4792 2963
rect 4824 2957 4904 2963
rect 5256 2957 5288 2963
rect 5341 2963 5347 2977
rect 5464 2977 5608 2983
rect 5341 2957 5768 2963
rect 5784 2957 5864 2963
rect 2952 2937 3139 2943
rect 3208 2937 3256 2943
rect 3416 2937 3496 2943
rect 3640 2937 3768 2943
rect 3912 2937 3944 2943
rect 4088 2937 4200 2943
rect 4232 2937 4264 2943
rect 4360 2937 4952 2943
rect 4968 2937 5032 2943
rect 5048 2937 5096 2943
rect 5112 2937 5176 2943
rect 5272 2937 5304 2943
rect 5336 2937 5368 2943
rect 5448 2937 5464 2943
rect 5608 2937 5672 2943
rect 120 2917 264 2923
rect 824 2917 856 2923
rect 1272 2917 1304 2923
rect 1336 2917 1416 2923
rect 1464 2917 1480 2923
rect 1784 2917 1832 2923
rect 1848 2917 1912 2923
rect 2024 2917 2184 2923
rect 2280 2917 2328 2923
rect 2488 2917 3176 2923
rect 3384 2917 3416 2923
rect 3512 2917 3672 2923
rect 3688 2917 4408 2923
rect 4472 2917 4664 2923
rect 4888 2917 4920 2923
rect 4936 2917 4952 2923
rect 4968 2917 5112 2923
rect 5224 2917 5800 2923
rect 5896 2917 5944 2923
rect 600 2897 696 2903
rect 1528 2897 1576 2903
rect 1608 2897 1816 2903
rect 1880 2897 2664 2903
rect 2680 2897 2792 2903
rect 3400 2897 3528 2903
rect 3656 2897 3752 2903
rect 4104 2897 4584 2903
rect 4680 2897 4888 2903
rect 4904 2897 4968 2903
rect 5064 2897 5080 2903
rect 5096 2897 5160 2903
rect 5176 2897 5320 2903
rect 216 2877 232 2883
rect 248 2877 296 2883
rect 3384 2877 3688 2883
rect 3832 2877 3944 2883
rect 4040 2877 4584 2883
rect 4856 2877 5176 2883
rect 376 2857 808 2863
rect 1736 2857 2600 2863
rect 3229 2857 3592 2863
rect 456 2837 520 2843
rect 952 2837 1016 2843
rect 1416 2837 1432 2843
rect 1576 2837 1736 2843
rect 1800 2837 2536 2843
rect 2568 2837 2728 2843
rect 3229 2843 3235 2857
rect 3784 2857 4136 2863
rect 4328 2857 4728 2863
rect 5656 2857 5688 2863
rect 2792 2837 3235 2843
rect 3256 2837 3576 2843
rect 3608 2837 3800 2843
rect 3816 2837 3848 2843
rect 3864 2837 4040 2843
rect 4920 2837 5336 2843
rect 5352 2837 5688 2843
rect 5768 2837 5784 2843
rect 5853 2837 5864 2843
rect 472 2817 840 2823
rect 1832 2817 1912 2823
rect 1928 2817 2248 2823
rect 2360 2817 2392 2823
rect 1384 2797 2024 2803
rect 2168 2797 2184 2803
rect 2328 2797 2744 2803
rect 3048 2817 3480 2823
rect 3496 2817 3528 2823
rect 3624 2817 3667 2823
rect 3192 2797 3640 2803
rect 3661 2803 3667 2817
rect 3848 2817 4360 2823
rect 3661 2797 4024 2803
rect 4056 2797 4520 2803
rect 5288 2817 5304 2823
rect 5320 2817 5336 2823
rect 5448 2817 5464 2823
rect 5496 2817 5512 2823
rect 5384 2797 5528 2803
rect 648 2777 1128 2783
rect 1240 2777 1336 2783
rect 2296 2777 2392 2783
rect 2408 2777 2472 2783
rect 2920 2777 3016 2783
rect 3064 2777 3320 2783
rect 3544 2777 3944 2783
rect 4072 2777 4184 2783
rect 4232 2777 4440 2783
rect 4456 2777 5064 2783
rect 5384 2777 5704 2783
rect 5720 2777 5992 2783
rect 744 2757 1288 2763
rect 1368 2757 1528 2763
rect 1688 2757 1704 2763
rect 1720 2757 1800 2763
rect 1816 2757 2024 2763
rect 2040 2757 2120 2763
rect 2136 2757 2312 2763
rect 2328 2757 2568 2763
rect 2584 2757 2680 2763
rect 2840 2757 3128 2763
rect 3240 2757 3448 2763
rect 3464 2757 3592 2763
rect 3688 2757 3848 2763
rect 3944 2757 4040 2763
rect 4136 2757 4504 2763
rect 4520 2757 4584 2763
rect 4600 2757 5576 2763
rect 312 2737 600 2743
rect 936 2737 1544 2743
rect 1912 2737 2552 2743
rect 3096 2737 3336 2743
rect 3576 2737 4072 2743
rect 4504 2737 4536 2743
rect 4552 2737 4744 2743
rect 4760 2737 5064 2743
rect 120 2717 232 2723
rect 248 2717 424 2723
rect 440 2717 488 2723
rect 504 2717 616 2723
rect 1192 2717 1368 2723
rect 2536 2717 2936 2723
rect 3032 2717 3080 2723
rect 3176 2717 3256 2723
rect 3368 2717 3416 2723
rect 3432 2717 4104 2723
rect 5608 2717 5752 2723
rect 5832 2717 5896 2723
rect 360 2697 472 2703
rect 552 2697 1064 2703
rect 1096 2697 1272 2703
rect 1464 2697 1640 2703
rect 1928 2697 1960 2703
rect 2056 2697 2088 2703
rect 2104 2697 2136 2703
rect 2344 2697 2488 2703
rect 2552 2697 2712 2703
rect 2728 2697 2888 2703
rect 2904 2697 3064 2703
rect 3080 2697 3128 2703
rect 3144 2697 3240 2703
rect 3256 2697 3352 2703
rect 3368 2697 3416 2703
rect 3448 2697 3560 2703
rect 3640 2697 3656 2703
rect 3768 2697 3800 2703
rect 3816 2697 3864 2703
rect 3885 2697 3912 2703
rect 264 2677 328 2683
rect 344 2677 456 2683
rect 616 2677 808 2683
rect 824 2677 872 2683
rect 1016 2677 1128 2683
rect 1256 2677 2216 2683
rect 2472 2677 2520 2683
rect 2680 2677 2712 2683
rect 2744 2677 2840 2683
rect 2856 2677 3144 2683
rect 3176 2677 3240 2683
rect 3496 2677 3544 2683
rect 3581 2683 3587 2692
rect 3576 2677 3587 2683
rect 3608 2677 3624 2683
rect 3885 2683 3891 2697
rect 4392 2697 4776 2703
rect 4968 2697 5128 2703
rect 5176 2697 5416 2703
rect 5432 2697 5480 2703
rect 5656 2697 5896 2703
rect 3656 2677 3891 2683
rect 3928 2677 4520 2683
rect 4840 2677 4856 2683
rect 4872 2677 5208 2683
rect 5512 2677 5544 2683
rect 5688 2677 5736 2683
rect 184 2657 200 2663
rect 488 2657 840 2663
rect 856 2657 936 2663
rect 952 2657 1192 2663
rect 1208 2657 2920 2663
rect 2936 2657 3880 2663
rect 3896 2657 3928 2663
rect 4408 2657 4472 2663
rect 4648 2657 4696 2663
rect 5112 2657 5304 2663
rect 5320 2657 5352 2663
rect 696 2637 808 2643
rect 824 2637 1080 2643
rect 1416 2637 1480 2643
rect 1640 2637 1656 2643
rect 1672 2637 1896 2643
rect 1992 2637 2056 2643
rect 2136 2637 2424 2643
rect 2680 2637 3032 2643
rect 3064 2637 3384 2643
rect 3448 2637 3640 2643
rect 3752 2637 3912 2643
rect 3928 2637 3976 2643
rect 3992 2637 4024 2643
rect 4200 2637 5032 2643
rect 5064 2637 5112 2643
rect 5128 2637 5288 2643
rect 5736 2637 5800 2643
rect 5880 2637 5944 2643
rect 2109 2628 2115 2632
rect 5853 2628 5859 2632
rect 952 2617 1160 2623
rect 1432 2617 1720 2623
rect 88 2597 1448 2603
rect 2632 2617 2680 2623
rect 2696 2617 3032 2623
rect 3288 2617 3480 2623
rect 3640 2617 3672 2623
rect 2488 2597 2904 2603
rect 2936 2597 2952 2603
rect 2984 2597 3272 2603
rect 3336 2597 3704 2603
rect 4648 2617 4760 2623
rect 4952 2617 4968 2623
rect 5000 2617 5464 2623
rect 4376 2597 4456 2603
rect 4904 2597 4968 2603
rect 5368 2597 5384 2603
rect 200 2577 216 2583
rect 264 2577 344 2583
rect 360 2577 1064 2583
rect 1320 2577 1560 2583
rect 1592 2577 1608 2583
rect 1656 2577 2328 2583
rect 2344 2577 2360 2583
rect 2376 2577 3448 2583
rect 3928 2577 3992 2583
rect 4008 2577 4312 2583
rect 5224 2577 5416 2583
rect 5432 2577 5544 2583
rect 5560 2577 5656 2583
rect 4445 2568 4451 2572
rect 56 2557 232 2563
rect 248 2557 328 2563
rect 344 2557 360 2563
rect 520 2557 584 2563
rect 872 2557 936 2563
rect 1048 2557 1128 2563
rect 1496 2557 1512 2563
rect 1544 2557 1624 2563
rect 1752 2557 1800 2563
rect 1816 2557 1832 2563
rect 1848 2557 1880 2563
rect 1992 2557 2136 2563
rect 2216 2557 2232 2563
rect 2328 2557 2392 2563
rect 2456 2557 2467 2563
rect 2776 2557 2888 2563
rect 2920 2557 3096 2563
rect 3128 2557 3160 2563
rect 3592 2557 3736 2563
rect 3752 2557 3944 2563
rect 4120 2557 4264 2563
rect 4520 2557 4648 2563
rect 4840 2557 4888 2563
rect 4968 2557 5000 2563
rect 5240 2557 5448 2563
rect 5800 2557 5832 2563
rect 216 2537 264 2543
rect 600 2537 696 2543
rect 888 2537 920 2543
rect 1016 2537 1048 2543
rect 1128 2537 1176 2543
rect 1240 2537 1256 2543
rect 1272 2537 1400 2543
rect 1416 2537 1736 2543
rect 1992 2537 2003 2543
rect 2056 2537 2184 2543
rect 2216 2537 2227 2543
rect 2413 2543 2419 2552
rect 2413 2537 2424 2543
rect 2472 2537 2536 2543
rect 2648 2537 2664 2543
rect 2888 2537 3048 2543
rect 3176 2537 3224 2543
rect 3608 2537 3752 2543
rect 3800 2537 3832 2543
rect 4248 2537 4280 2543
rect 4312 2537 4600 2543
rect 4616 2537 4664 2543
rect 4776 2537 4792 2543
rect 4808 2537 4936 2543
rect 4952 2537 5048 2543
rect 5464 2537 5544 2543
rect 5560 2537 5832 2543
rect -51 2517 8 2523
rect 24 2517 72 2523
rect 760 2517 888 2523
rect 1384 2517 1464 2523
rect 1880 2517 2040 2523
rect 2072 2517 2088 2523
rect 2184 2517 2264 2523
rect 2280 2517 2520 2523
rect 3112 2517 3192 2523
rect 3240 2517 3256 2523
rect 3352 2517 3432 2523
rect 3688 2517 3960 2523
rect 4024 2517 4152 2523
rect 4184 2517 4200 2523
rect 4216 2517 4312 2523
rect 5000 2517 5032 2523
rect 5112 2517 5160 2523
rect 5192 2517 5400 2523
rect 5416 2517 5432 2523
rect 5544 2517 5560 2523
rect 5704 2517 5720 2523
rect 5736 2517 5768 2523
rect 584 2497 664 2503
rect 680 2497 808 2503
rect 824 2497 984 2503
rect 1000 2497 1496 2503
rect 2104 2497 2136 2503
rect 2152 2497 2168 2503
rect 2664 2497 3128 2503
rect 3432 2497 3656 2503
rect 3736 2497 3768 2503
rect 3960 2497 4856 2503
rect 4888 2497 5112 2503
rect 5320 2497 5688 2503
rect 664 2477 728 2483
rect 744 2477 1080 2483
rect 1096 2477 1912 2483
rect 2040 2477 3112 2483
rect 3560 2477 3592 2483
rect 3672 2477 3688 2483
rect 3720 2477 3832 2483
rect 3912 2477 4152 2483
rect 4168 2477 4184 2483
rect 4200 2477 4296 2483
rect 4312 2477 4488 2483
rect 4536 2477 4984 2483
rect 776 2457 1016 2463
rect 1688 2457 1752 2463
rect 2600 2457 2664 2463
rect 3160 2457 3240 2463
rect 3256 2457 3448 2463
rect 3464 2457 4472 2463
rect 5000 2457 5016 2463
rect 5448 2457 5880 2463
rect 152 2437 168 2443
rect 776 2437 792 2443
rect 1544 2437 2280 2443
rect 2584 2437 2664 2443
rect 3368 2437 4632 2443
rect 4648 2437 5688 2443
rect 3053 2428 3059 2432
rect 328 2417 376 2423
rect 1624 2417 2136 2423
rect 2376 2417 2808 2423
rect 984 2397 1704 2403
rect 1720 2397 2152 2403
rect 2360 2397 2776 2403
rect 3144 2417 3160 2423
rect 4072 2417 4088 2423
rect 4136 2417 4392 2423
rect 3560 2397 3784 2403
rect 4312 2397 4344 2403
rect 4440 2397 4904 2403
rect 5224 2417 5320 2423
rect 5720 2417 5736 2423
rect 376 2377 424 2383
rect 440 2377 648 2383
rect 1176 2377 1240 2383
rect 1288 2377 1848 2383
rect 1864 2377 2040 2383
rect 2088 2377 2712 2383
rect 3288 2377 3304 2383
rect 3768 2377 4568 2383
rect 5544 2377 5592 2383
rect 56 2357 104 2363
rect 120 2357 152 2363
rect 168 2357 472 2363
rect 488 2357 808 2363
rect 904 2357 936 2363
rect 1368 2357 1464 2363
rect 1512 2357 2088 2363
rect 2264 2357 2712 2363
rect 2888 2357 2952 2363
rect 2968 2357 3272 2363
rect 4568 2357 4744 2363
rect 5336 2357 5528 2363
rect 5544 2357 5752 2363
rect 5768 2357 5816 2363
rect 392 2337 1288 2343
rect 1320 2337 1528 2343
rect 1624 2337 1656 2343
rect 1704 2337 2216 2343
rect 2520 2337 2776 2343
rect 2952 2337 3560 2343
rect 3688 2337 3992 2343
rect 4072 2337 4184 2343
rect 4200 2337 4728 2343
rect 5464 2337 5576 2343
rect 5592 2337 5608 2343
rect -51 2317 392 2323
rect 1096 2317 1112 2323
rect 1208 2317 1384 2323
rect 1896 2317 1928 2323
rect 2744 2317 2776 2323
rect 2840 2317 3096 2323
rect 3128 2317 3240 2323
rect 3752 2317 3800 2323
rect 3992 2317 4104 2323
rect 4168 2317 4216 2323
rect 4424 2317 4488 2323
rect 4504 2317 4552 2323
rect 4712 2317 4824 2323
rect 5176 2317 5224 2323
rect 5240 2317 5320 2323
rect 5704 2317 5784 2323
rect 5800 2317 5896 2323
rect 3725 2308 3731 2312
rect 5501 2308 5507 2312
rect 200 2297 520 2303
rect 605 2297 616 2303
rect 728 2297 984 2303
rect 1016 2297 1384 2303
rect 1501 2297 1512 2303
rect 1576 2297 1704 2303
rect 1768 2297 1816 2303
rect 1848 2297 1896 2303
rect 1928 2297 2088 2303
rect 2264 2297 2456 2303
rect 2520 2297 3032 2303
rect 3064 2297 3096 2303
rect 3128 2297 3144 2303
rect 3352 2297 3384 2303
rect 3464 2297 3512 2303
rect 3752 2297 3768 2303
rect 4040 2297 4056 2303
rect 4104 2297 4200 2303
rect 4280 2297 4360 2303
rect 4376 2297 4440 2303
rect 4488 2297 4600 2303
rect 4616 2297 4776 2303
rect 4808 2297 4840 2303
rect 4984 2297 5000 2303
rect 5192 2297 5432 2303
rect 5736 2297 5752 2303
rect 5784 2297 5800 2303
rect 3229 2288 3235 2292
rect 408 2277 696 2283
rect 808 2277 1544 2283
rect 1672 2277 1832 2283
rect 2024 2277 2072 2283
rect 2120 2277 2264 2283
rect 2328 2277 2339 2283
rect 2557 2277 2568 2283
rect 2824 2277 2840 2283
rect 2872 2277 2904 2283
rect 3080 2277 3144 2283
rect 3160 2277 3192 2283
rect 3384 2277 3448 2283
rect 3496 2277 3880 2283
rect 4072 2277 4104 2283
rect 4408 2277 4424 2283
rect 4456 2277 4520 2283
rect 4600 2277 4856 2283
rect 4968 2277 5016 2283
rect 5048 2277 5059 2283
rect 5112 2277 5144 2283
rect 5528 2277 5560 2283
rect 5576 2277 5720 2283
rect 5421 2268 5427 2272
rect 216 2257 264 2263
rect 568 2257 872 2263
rect 904 2257 1336 2263
rect 1432 2257 2136 2263
rect 2152 2257 2200 2263
rect 2216 2257 2264 2263
rect 2280 2257 2392 2263
rect 2408 2257 2520 2263
rect 2760 2257 2888 2263
rect 2904 2257 2920 2263
rect 3245 2257 3336 2263
rect 392 2237 712 2243
rect 728 2237 1096 2243
rect 1944 2237 2072 2243
rect 2445 2237 2456 2243
rect 2888 2237 2952 2243
rect 2984 2237 3128 2243
rect 3245 2243 3251 2257
rect 3640 2257 3688 2263
rect 3800 2257 3880 2263
rect 3976 2257 4296 2263
rect 4648 2257 4696 2263
rect 5192 2257 5256 2263
rect 3192 2237 3251 2243
rect 3272 2237 3432 2243
rect 3560 2237 3576 2243
rect 4232 2237 4312 2243
rect 4616 2237 4824 2243
rect 5288 2237 5368 2243
rect 5592 2237 5848 2243
rect 88 2217 424 2223
rect 648 2217 680 2223
rect 856 2217 1016 2223
rect 1048 2217 1272 2223
rect 1288 2217 1448 2223
rect 1480 2217 1512 2223
rect 24 2197 536 2203
rect 584 2197 840 2203
rect 856 2197 984 2203
rect 1000 2197 1192 2203
rect 1208 2197 1304 2203
rect 1320 2197 1400 2203
rect 2184 2217 2200 2223
rect 2392 2217 2648 2223
rect 2669 2217 2904 2223
rect 2669 2203 2675 2217
rect 2936 2217 3256 2223
rect 3448 2217 3480 2223
rect 3512 2217 3896 2223
rect 2440 2197 2675 2203
rect 2808 2197 2888 2203
rect 2920 2197 3496 2203
rect 3624 2197 3752 2203
rect 3848 2197 3944 2203
rect 4088 2217 4152 2223
rect 4248 2217 4552 2223
rect 4584 2217 4936 2223
rect 4952 2217 5176 2223
rect 5784 2217 5880 2223
rect 4040 2197 4312 2203
rect 4760 2197 4920 2203
rect 4936 2197 5176 2203
rect 5304 2197 5784 2203
rect 152 2177 488 2183
rect 520 2177 1896 2183
rect 1928 2177 2136 2183
rect 2712 2177 2728 2183
rect 2776 2177 2904 2183
rect 2936 2177 3064 2183
rect 3096 2177 3464 2183
rect 3480 2177 3592 2183
rect 3608 2177 3832 2183
rect 3864 2177 4104 2183
rect 4184 2177 4424 2183
rect 4520 2177 4568 2183
rect 4840 2177 5304 2183
rect 5480 2177 5704 2183
rect -51 2157 8 2163
rect 24 2157 72 2163
rect 88 2157 136 2163
rect 152 2157 360 2163
rect 424 2157 728 2163
rect 792 2157 856 2163
rect 872 2157 952 2163
rect 968 2157 1064 2163
rect 1128 2157 1304 2163
rect 1384 2157 1507 2163
rect 216 2137 232 2143
rect 248 2137 280 2143
rect 296 2137 376 2143
rect 568 2137 600 2143
rect 648 2137 664 2143
rect 712 2137 760 2143
rect 1048 2137 1144 2143
rect 1181 2137 1192 2143
rect 1448 2137 1480 2143
rect 1501 2143 1507 2157
rect 1784 2157 1832 2163
rect 1848 2157 1912 2163
rect 2397 2163 2403 2172
rect 2392 2157 2403 2163
rect 2616 2157 2792 2163
rect 2840 2157 3048 2163
rect 3064 2157 3608 2163
rect 3768 2157 4232 2163
rect 4248 2157 4280 2163
rect 4296 2157 4632 2163
rect 4840 2157 5096 2163
rect 5128 2157 5224 2163
rect 5336 2157 5400 2163
rect 5608 2157 5720 2163
rect 1501 2137 1592 2143
rect 1704 2137 1816 2143
rect 1848 2137 2072 2143
rect 2184 2137 2248 2143
rect 2424 2137 2456 2143
rect 2552 2137 2696 2143
rect 2952 2137 3096 2143
rect 3368 2137 3416 2143
rect 3832 2137 3848 2143
rect 4104 2137 4392 2143
rect 4536 2137 4584 2143
rect 4664 2137 4696 2143
rect 5016 2137 5048 2143
rect 5192 2137 5448 2143
rect 5496 2137 5528 2143
rect 5624 2137 5736 2143
rect 5832 2137 5880 2143
rect 5896 2137 5928 2143
rect 5613 2128 5619 2132
rect -51 2117 184 2123
rect 328 2117 472 2123
rect 488 2117 648 2123
rect 712 2117 1096 2123
rect 1112 2117 1576 2123
rect 1592 2117 1688 2123
rect 1720 2117 1896 2123
rect 1912 2117 2008 2123
rect 2504 2117 2552 2123
rect 2664 2117 2792 2123
rect 2824 2117 3000 2123
rect 3144 2117 3160 2123
rect 3208 2117 3320 2123
rect 3336 2117 3368 2123
rect 3416 2117 3480 2123
rect 3624 2117 3704 2123
rect 3720 2117 3768 2123
rect 3784 2117 3864 2123
rect 3880 2117 4040 2123
rect 4056 2117 4072 2123
rect 4152 2117 4344 2123
rect 4360 2117 4376 2123
rect 4552 2117 4680 2123
rect 4840 2117 4872 2123
rect 4888 2117 4920 2123
rect 4936 2117 5160 2123
rect 5176 2117 5288 2123
rect 5304 2117 5592 2123
rect 5640 2117 5816 2123
rect 5896 2117 5960 2123
rect 168 2097 216 2103
rect 264 2097 504 2103
rect 984 2097 1128 2103
rect 1272 2097 1640 2103
rect 1672 2097 2024 2103
rect 2056 2097 2504 2103
rect 2632 2097 2643 2103
rect 2637 2088 2643 2097
rect 2664 2097 2888 2103
rect 3160 2097 3480 2103
rect 3496 2097 3544 2103
rect 3848 2097 4040 2103
rect 4056 2097 4280 2103
rect 4312 2097 4760 2103
rect 5064 2097 5336 2103
rect 5368 2097 5496 2103
rect 5592 2097 5688 2103
rect 2893 2088 2899 2092
rect 72 2077 120 2083
rect 200 2077 264 2083
rect 280 2077 360 2083
rect 840 2077 1288 2083
rect 1560 2077 1848 2083
rect 1928 2077 2152 2083
rect 2184 2077 2408 2083
rect 2424 2077 2456 2083
rect 3416 2077 3448 2083
rect 3464 2077 3704 2083
rect 3928 2077 4216 2083
rect 4632 2077 4824 2083
rect 4984 2077 5064 2083
rect 5128 2077 5272 2083
rect 5384 2077 5816 2083
rect 696 2057 1560 2063
rect 1848 2057 2200 2063
rect 2232 2057 3288 2063
rect 3400 2057 3816 2063
rect 3832 2057 4120 2063
rect 4152 2057 4184 2063
rect 4248 2057 4259 2063
rect 4376 2057 4696 2063
rect 4936 2057 5368 2063
rect 88 2037 104 2043
rect 152 2037 216 2043
rect 344 2037 408 2043
rect 536 2037 600 2043
rect 1144 2037 1448 2043
rect 1640 2037 1784 2043
rect 2008 2037 2168 2043
rect 2184 2037 3640 2043
rect 3832 2037 5000 2043
rect 5240 2037 5480 2043
rect 5560 2037 5624 2043
rect 216 2017 344 2023
rect 600 2017 824 2023
rect 1336 2017 1384 2023
rect 1592 2017 1891 2023
rect 1032 1997 1864 2003
rect 1885 2003 1891 2017
rect 2152 2017 2184 2023
rect 2200 2017 2344 2023
rect 2584 2017 2872 2023
rect 1885 1997 2184 2003
rect 2264 1997 2824 2003
rect 3080 2017 3272 2023
rect 3288 2017 3464 2023
rect 3480 2017 3800 2023
rect 3816 2017 3848 2023
rect 3928 2017 4296 2023
rect 4504 2017 4792 2023
rect 3192 1997 3288 2003
rect 3304 1997 3320 2003
rect 3352 1997 3624 2003
rect 3640 1997 4200 2003
rect 4264 1997 4280 2003
rect 4328 1997 4504 2003
rect 4536 1997 4712 2003
rect 4904 1997 5000 2003
rect 1016 1977 2216 1983
rect 2360 1977 3224 1983
rect 3240 1977 3256 1983
rect 3272 1977 3304 1983
rect 3624 1977 4136 1983
rect 4168 1977 4312 1983
rect 4376 1977 4808 1983
rect 4952 1977 5976 1983
rect 1016 1957 1704 1963
rect 1768 1957 1912 1963
rect 2056 1957 2088 1963
rect 2152 1957 2440 1963
rect 2632 1957 2712 1963
rect 2728 1957 3192 1963
rect 3208 1957 3240 1963
rect 3256 1957 3272 1963
rect 3672 1957 3800 1963
rect 3944 1957 3955 1963
rect 4184 1957 4472 1963
rect 4488 1957 4600 1963
rect 4664 1957 5144 1963
rect -51 1937 488 1943
rect 504 1937 712 1943
rect 920 1937 1128 1943
rect 1288 1937 1704 1943
rect 1736 1937 1816 1943
rect 1912 1937 2008 1943
rect 2440 1937 2584 1943
rect 2664 1937 2696 1943
rect 2856 1937 2888 1943
rect 2989 1937 3064 1943
rect 56 1917 72 1923
rect 88 1917 168 1923
rect 264 1917 280 1923
rect 856 1917 888 1923
rect 984 1917 1720 1923
rect 1752 1917 1832 1923
rect 2024 1917 2296 1923
rect 2312 1917 2376 1923
rect 2408 1917 2760 1923
rect 2989 1923 2995 1937
rect 3224 1937 3368 1943
rect 3688 1937 4728 1943
rect 4744 1937 4856 1943
rect 4872 1937 5256 1943
rect 5416 1937 5736 1943
rect 2776 1917 2995 1923
rect 3016 1917 3128 1923
rect 3544 1917 3720 1923
rect 3800 1917 4131 1923
rect 477 1908 483 1912
rect 765 1908 771 1912
rect 216 1897 328 1903
rect 488 1897 696 1903
rect 712 1897 744 1903
rect 808 1897 920 1903
rect 1224 1897 1432 1903
rect 1592 1897 1624 1903
rect 1688 1897 1736 1903
rect 1768 1897 2216 1903
rect 2280 1897 2296 1903
rect 2344 1897 2584 1903
rect 2680 1897 2920 1903
rect 3000 1897 3443 1903
rect 56 1877 152 1883
rect 520 1877 584 1883
rect 616 1877 648 1883
rect 792 1877 1064 1883
rect 1368 1877 2184 1883
rect 2216 1877 2280 1883
rect 2472 1877 2504 1883
rect 2584 1877 2648 1883
rect 2712 1877 2824 1883
rect 2840 1877 2856 1883
rect 2952 1877 3016 1883
rect 3064 1877 3112 1883
rect 3240 1877 3416 1883
rect 3437 1883 3443 1897
rect 3464 1897 3496 1903
rect 3656 1897 3752 1903
rect 3768 1897 3832 1903
rect 4125 1903 4131 1917
rect 4312 1917 4840 1923
rect 4856 1917 5224 1923
rect 5272 1917 5528 1923
rect 5544 1917 5640 1923
rect 4125 1897 4184 1903
rect 4264 1897 4275 1903
rect 4285 1897 4296 1903
rect 4472 1897 4648 1903
rect 4728 1897 4744 1903
rect 4760 1897 5016 1903
rect 5256 1897 5464 1903
rect 5480 1897 5576 1903
rect 5592 1897 5624 1903
rect 5656 1897 5768 1903
rect 5869 1888 5875 1892
rect 3437 1877 3496 1883
rect 3704 1877 3715 1883
rect 3736 1877 3800 1883
rect 3832 1877 3864 1883
rect 3944 1877 3960 1883
rect 4248 1877 4376 1883
rect 4424 1877 4504 1883
rect 4568 1877 4616 1883
rect 5224 1877 5320 1883
rect 5384 1877 5416 1883
rect 5432 1877 5576 1883
rect 5640 1877 5672 1883
rect 5768 1877 5864 1883
rect -51 1857 8 1863
rect 24 1857 56 1863
rect 280 1857 376 1863
rect 392 1857 472 1863
rect 648 1857 1288 1863
rect 1432 1857 1768 1863
rect 1896 1857 1912 1863
rect 1960 1857 1971 1863
rect 2168 1857 2232 1863
rect 2472 1857 2696 1863
rect 2856 1857 3048 1863
rect 3144 1857 3224 1863
rect 3352 1857 3368 1863
rect 3608 1857 3640 1863
rect 4024 1857 4248 1863
rect 4264 1857 4424 1863
rect 4488 1857 4536 1863
rect 5496 1857 5848 1863
rect 5864 1857 5944 1863
rect 376 1837 424 1843
rect 456 1837 520 1843
rect 600 1837 952 1843
rect 1608 1837 2760 1843
rect 2808 1837 2888 1843
rect 2920 1837 2936 1843
rect 2952 1837 3176 1843
rect 3224 1837 3272 1843
rect 3288 1837 3528 1843
rect 3592 1837 3928 1843
rect 4072 1837 4424 1843
rect 4568 1837 4856 1843
rect 5144 1837 5176 1843
rect 152 1817 536 1823
rect 584 1817 760 1823
rect 1128 1817 1368 1823
rect -51 1797 8 1803
rect 24 1797 88 1803
rect 264 1797 456 1803
rect 488 1797 584 1803
rect 621 1797 1000 1803
rect 104 1777 152 1783
rect 168 1777 376 1783
rect 408 1777 456 1783
rect 621 1783 627 1797
rect 1624 1797 1736 1803
rect 2072 1817 3560 1823
rect 2024 1797 2248 1803
rect 2568 1797 2632 1803
rect 2664 1797 2968 1803
rect 3032 1797 3064 1803
rect 3128 1797 3368 1803
rect 3432 1797 3688 1803
rect 4136 1817 4824 1823
rect 4872 1817 5000 1823
rect 5016 1817 5224 1823
rect 5240 1817 5304 1823
rect 5320 1817 5720 1823
rect 4040 1797 4232 1803
rect 4248 1797 4808 1803
rect 5160 1797 5192 1803
rect 5400 1797 5528 1803
rect 5544 1797 5560 1803
rect 5608 1797 5640 1803
rect 5848 1797 5896 1803
rect 472 1777 627 1783
rect 637 1777 824 1783
rect -51 1757 8 1763
rect 93 1757 104 1763
rect 360 1757 520 1763
rect 637 1763 643 1777
rect 888 1777 1144 1783
rect 1304 1777 1320 1783
rect 1560 1777 2024 1783
rect 2040 1777 2072 1783
rect 2104 1777 2168 1783
rect 2184 1777 2424 1783
rect 2504 1777 2536 1783
rect 2632 1777 2760 1783
rect 2920 1777 3016 1783
rect 3048 1777 3368 1783
rect 3480 1777 3560 1783
rect 3832 1777 3896 1783
rect 3976 1777 3992 1783
rect 4008 1777 4088 1783
rect 4152 1777 4168 1783
rect 4712 1777 4968 1783
rect 4984 1777 5096 1783
rect 5144 1777 5432 1783
rect 5624 1777 5704 1783
rect 5736 1777 5896 1783
rect 552 1757 643 1763
rect 744 1757 1000 1763
rect 1144 1757 1176 1763
rect 1624 1757 2040 1763
rect 2088 1757 2280 1763
rect 2536 1757 2936 1763
rect 3064 1757 3208 1763
rect 3240 1757 3272 1763
rect 3352 1757 3400 1763
rect 3560 1757 3848 1763
rect 3896 1757 3960 1763
rect 3992 1757 4024 1763
rect 4104 1757 4472 1763
rect 4664 1757 4696 1763
rect 4728 1757 4739 1763
rect 4824 1757 5032 1763
rect 5048 1757 5144 1763
rect 5160 1757 5176 1763
rect 5192 1757 5640 1763
rect 5688 1757 5816 1763
rect 3213 1748 3219 1752
rect 136 1737 344 1743
rect 376 1737 392 1743
rect 408 1737 616 1743
rect 632 1737 680 1743
rect 696 1737 712 1743
rect 824 1737 856 1743
rect 941 1737 952 1743
rect 1064 1737 1128 1743
rect 1192 1737 1240 1743
rect 1272 1737 1320 1743
rect 1544 1737 1592 1743
rect 1816 1737 1912 1743
rect 2328 1737 2440 1743
rect 2488 1737 2552 1743
rect 2680 1737 2856 1743
rect 2888 1737 3027 1743
rect 781 1728 787 1732
rect -51 1703 -45 1723
rect 40 1717 184 1723
rect 264 1717 280 1723
rect 360 1717 408 1723
rect 424 1717 600 1723
rect 909 1723 915 1732
rect 1773 1728 1779 1732
rect 904 1717 915 1723
rect 1192 1717 1256 1723
rect 1416 1717 1432 1723
rect 1496 1717 1560 1723
rect 2216 1717 2227 1723
rect 2392 1717 2424 1723
rect 2440 1717 2488 1723
rect 2616 1717 2664 1723
rect 2685 1708 2691 1723
rect 2712 1717 2872 1723
rect 2952 1717 3000 1723
rect 3021 1723 3027 1737
rect 3128 1737 3160 1743
rect 3288 1737 3304 1743
rect 3688 1737 3768 1743
rect 3805 1737 3816 1743
rect 3960 1737 4008 1743
rect 4024 1737 4120 1743
rect 4152 1737 4280 1743
rect 4296 1737 4696 1743
rect 4712 1737 5016 1743
rect 5032 1737 5096 1743
rect 5144 1737 5336 1743
rect 5352 1737 5384 1743
rect 5464 1737 5496 1743
rect 5640 1737 5880 1743
rect 3021 1717 3432 1723
rect 3480 1717 3512 1723
rect 3560 1717 3832 1723
rect 3944 1717 4136 1723
rect 4312 1717 4632 1723
rect 4648 1717 4792 1723
rect 4808 1717 4824 1723
rect 5176 1717 5256 1723
rect 5384 1717 5608 1723
rect 5624 1717 5768 1723
rect -51 1697 40 1703
rect 328 1697 424 1703
rect 456 1697 536 1703
rect 888 1697 1160 1703
rect 1240 1697 1288 1703
rect 1432 1697 2088 1703
rect 2120 1697 2568 1703
rect 2840 1697 3272 1703
rect 3304 1697 3352 1703
rect 3640 1697 3651 1703
rect 3736 1697 4376 1703
rect 4824 1697 4936 1703
rect 5368 1697 5448 1703
rect 5464 1697 5816 1703
rect 5912 1697 5960 1703
rect -51 1677 344 1683
rect 824 1677 936 1683
rect 952 1677 1320 1683
rect 1336 1677 1832 1683
rect 2056 1677 2232 1683
rect 2248 1677 2392 1683
rect 2600 1677 3656 1683
rect 4280 1677 4328 1683
rect 4344 1677 4664 1683
rect 344 1657 456 1663
rect 584 1657 632 1663
rect 648 1657 744 1663
rect 760 1657 1352 1663
rect 1480 1657 1672 1663
rect 1736 1657 2520 1663
rect 2584 1657 3224 1663
rect 3752 1657 3912 1663
rect 4696 1657 4712 1663
rect 5416 1657 5432 1663
rect 744 1637 968 1643
rect 1176 1637 1272 1643
rect 1480 1637 1496 1643
rect 1768 1637 2040 1643
rect 2456 1637 2552 1643
rect 2568 1637 2616 1643
rect 2632 1637 2808 1643
rect 2968 1637 3384 1643
rect 3416 1637 3800 1643
rect 3816 1637 4056 1643
rect 4200 1637 4888 1643
rect 5112 1637 5304 1643
rect 24 1617 216 1623
rect 232 1617 600 1623
rect 632 1617 760 1623
rect -51 1597 56 1603
rect 216 1597 616 1603
rect 1048 1617 1512 1623
rect 2136 1617 2504 1623
rect 2536 1617 2840 1623
rect 1096 1597 1224 1603
rect 1320 1597 1784 1603
rect 1816 1597 2440 1603
rect 2728 1597 2744 1603
rect 2872 1597 2936 1603
rect 3400 1617 3416 1623
rect 3640 1617 3656 1623
rect 3064 1597 3224 1603
rect 3512 1597 3928 1603
rect 5416 1617 5544 1623
rect 280 1577 584 1583
rect 680 1577 1096 1583
rect 1128 1577 1208 1583
rect 1256 1577 1592 1583
rect 1608 1577 1672 1583
rect 1832 1577 2088 1583
rect 2296 1577 2664 1583
rect 2776 1577 2872 1583
rect 3080 1577 3192 1583
rect 3208 1577 3288 1583
rect 3592 1577 4072 1583
rect 4120 1577 4264 1583
rect 4280 1577 5288 1583
rect -51 1557 8 1563
rect 184 1557 536 1563
rect 776 1557 888 1563
rect 904 1557 1272 1563
rect 1288 1557 1752 1563
rect 2088 1557 2152 1563
rect 2168 1557 2328 1563
rect 2376 1557 2488 1563
rect 2504 1557 2568 1563
rect 2584 1557 2888 1563
rect 2904 1557 3592 1563
rect 3704 1557 3736 1563
rect 3928 1557 4040 1563
rect 4248 1557 4312 1563
rect 4328 1557 4344 1563
rect 4360 1557 4600 1563
rect 4696 1557 4824 1563
rect 200 1537 424 1543
rect 1016 1537 1048 1543
rect 1112 1537 1160 1543
rect 1192 1537 1336 1543
rect 1896 1537 2232 1543
rect 2248 1537 2456 1543
rect 2936 1537 2952 1543
rect 2968 1537 3112 1543
rect 3144 1537 3192 1543
rect 3352 1537 4072 1543
rect 4104 1537 4136 1543
rect 4264 1537 4376 1543
rect 4392 1537 4472 1543
rect 4504 1537 4744 1543
rect -51 1517 744 1523
rect 776 1517 1128 1523
rect 1304 1517 1528 1523
rect 1544 1517 1624 1523
rect 1656 1517 1992 1523
rect 2056 1517 2200 1523
rect 2296 1517 2312 1523
rect 2344 1517 2392 1523
rect 2424 1517 2456 1523
rect 2616 1517 2648 1523
rect 2744 1517 3096 1523
rect 3128 1517 3176 1523
rect 3192 1517 3256 1523
rect 3336 1517 3496 1523
rect 3800 1517 3832 1523
rect 3928 1517 4104 1523
rect 4312 1517 4392 1523
rect 4488 1517 4616 1523
rect 4632 1517 4776 1523
rect 5016 1517 5240 1523
rect 5656 1517 5704 1523
rect 5720 1517 5784 1523
rect 104 1497 152 1503
rect 344 1497 392 1503
rect 456 1497 520 1503
rect 669 1497 680 1503
rect 669 1488 675 1497
rect 760 1497 776 1503
rect 824 1497 904 1503
rect 1000 1497 1064 1503
rect 1112 1497 1240 1503
rect 1320 1497 1432 1503
rect 1464 1497 1912 1503
rect 1992 1497 2312 1503
rect 2360 1497 2584 1503
rect 2696 1497 2728 1503
rect 2936 1497 3288 1503
rect 3320 1497 3480 1503
rect 3512 1497 3544 1503
rect 3624 1497 3816 1503
rect 3832 1497 4008 1503
rect 4152 1497 4456 1503
rect 4616 1497 4728 1503
rect 4744 1497 4808 1503
rect 4856 1497 4872 1503
rect 5096 1497 5144 1503
rect 1293 1488 1299 1492
rect 56 1477 104 1483
rect 504 1477 648 1483
rect 728 1477 824 1483
rect 1096 1477 1192 1483
rect 1384 1477 1416 1483
rect 1448 1477 1608 1483
rect 1752 1477 1848 1483
rect 1864 1477 2472 1483
rect 2520 1477 2664 1483
rect 2680 1477 2872 1483
rect 2888 1477 2920 1483
rect 2936 1477 3128 1483
rect 3272 1477 3832 1483
rect 3880 1477 4024 1483
rect 4088 1477 4184 1483
rect 4232 1477 4280 1483
rect 4440 1477 4504 1483
rect 4664 1477 4712 1483
rect 4792 1477 4904 1483
rect 5496 1477 5560 1483
rect 5624 1477 5704 1483
rect 5720 1477 5752 1483
rect 5800 1477 5960 1483
rect 792 1457 808 1463
rect 824 1457 872 1463
rect 952 1457 1720 1463
rect 1784 1457 1816 1463
rect 1848 1457 2216 1463
rect 2248 1457 2376 1463
rect 2392 1457 2616 1463
rect 3112 1457 3128 1463
rect 3160 1457 3320 1463
rect 3448 1457 3528 1463
rect 3560 1457 3576 1463
rect 3976 1457 3992 1463
rect 4024 1457 4328 1463
rect 4456 1457 4504 1463
rect 4808 1457 4856 1463
rect 5272 1457 5288 1463
rect 5304 1457 5416 1463
rect 5432 1457 5544 1463
rect 5704 1457 5736 1463
rect 5912 1457 5960 1463
rect 712 1437 744 1443
rect 1128 1437 1224 1443
rect 1576 1437 1624 1443
rect 1912 1437 2024 1443
rect 2040 1437 2152 1443
rect 2168 1437 2728 1443
rect 2760 1437 3048 1443
rect 3528 1437 3560 1443
rect 3672 1437 3752 1443
rect 4200 1437 4584 1443
rect 4872 1437 4952 1443
rect 4968 1437 5416 1443
rect 5688 1437 5880 1443
rect 5928 1437 5960 1443
rect 632 1417 728 1423
rect 776 1417 1016 1423
rect 1048 1417 1096 1423
rect 1112 1417 1720 1423
rect 520 1397 552 1403
rect 648 1397 840 1403
rect 856 1397 1256 1403
rect 1272 1397 1368 1403
rect 1384 1397 1480 1403
rect 1496 1397 1560 1403
rect 1576 1397 1640 1403
rect 2184 1417 2232 1423
rect 2312 1417 2344 1423
rect 2365 1417 2632 1423
rect 2365 1403 2371 1417
rect 2680 1417 2808 1423
rect 3064 1417 3096 1423
rect 3112 1417 3240 1423
rect 3400 1417 3864 1423
rect 2328 1397 2371 1403
rect 2440 1397 2888 1403
rect 3096 1397 3400 1403
rect 3464 1397 3896 1403
rect 4232 1417 4728 1423
rect 5416 1417 5496 1423
rect 4344 1397 4536 1403
rect 4632 1397 4904 1403
rect 5096 1397 5288 1403
rect 5533 1388 5539 1392
rect 152 1377 296 1383
rect 424 1377 1048 1383
rect 1208 1377 1224 1383
rect 1720 1377 2008 1383
rect 2024 1377 2216 1383
rect 2232 1377 2424 1383
rect 2600 1377 2648 1383
rect 2680 1377 2776 1383
rect 3128 1377 3368 1383
rect 3880 1377 4040 1383
rect 4104 1377 4376 1383
rect 4392 1377 5176 1383
rect 5560 1377 5752 1383
rect 5832 1377 5848 1383
rect 472 1357 552 1363
rect 808 1357 1064 1363
rect 1080 1357 2200 1363
rect 2296 1357 2344 1363
rect 2424 1357 2600 1363
rect 2712 1357 2776 1363
rect 3016 1357 3064 1363
rect 3240 1357 3304 1363
rect 3496 1357 3592 1363
rect 3624 1357 3688 1363
rect 3864 1357 3880 1363
rect 4216 1357 4227 1363
rect 4344 1357 4440 1363
rect 4456 1357 4504 1363
rect 4776 1357 4872 1363
rect 5160 1357 5352 1363
rect 5592 1357 5656 1363
rect 573 1337 584 1343
rect 712 1337 792 1343
rect 840 1337 872 1343
rect 1192 1337 1208 1343
rect 1240 1337 1304 1343
rect 1320 1337 1448 1343
rect 1464 1337 1544 1343
rect 1688 1337 1768 1343
rect 1789 1337 1848 1343
rect -51 1317 8 1323
rect 248 1317 616 1323
rect 856 1317 904 1323
rect 1160 1317 1192 1323
rect 1496 1317 1507 1323
rect 1528 1317 1576 1323
rect 1597 1317 1608 1323
rect 1789 1323 1795 1337
rect 1960 1337 2040 1343
rect 2296 1337 2360 1343
rect 2408 1337 2424 1343
rect 2472 1337 2488 1343
rect 2504 1337 2744 1343
rect 2792 1337 2824 1343
rect 3096 1337 3176 1343
rect 3304 1337 3336 1343
rect 3480 1337 3512 1343
rect 3544 1337 3672 1343
rect 3752 1337 3768 1343
rect 3928 1337 3944 1343
rect 4056 1337 4104 1343
rect 4456 1337 4467 1343
rect 4493 1337 4504 1343
rect 4776 1337 4808 1343
rect 5224 1337 5272 1343
rect 5400 1337 5448 1343
rect 5720 1337 5896 1343
rect 1704 1317 1795 1323
rect 1816 1317 1864 1323
rect 1880 1317 1896 1323
rect 2088 1317 2312 1323
rect 2344 1317 2392 1323
rect 2472 1317 3144 1323
rect 3176 1317 3736 1323
rect 3800 1317 3816 1323
rect 3944 1317 3960 1323
rect 4280 1317 4360 1323
rect 4712 1317 4776 1323
rect 4920 1317 4984 1323
rect 5000 1317 5160 1323
rect 5192 1317 5224 1323
rect 5464 1317 5592 1323
rect 616 1297 792 1303
rect 984 1297 1208 1303
rect 1544 1297 1704 1303
rect 1720 1297 2376 1303
rect 2488 1297 2584 1303
rect 2600 1297 2760 1303
rect 2776 1297 2872 1303
rect 2968 1297 3336 1303
rect 3512 1297 3608 1303
rect 3656 1297 3752 1303
rect 3768 1297 4104 1303
rect 4392 1297 4403 1303
rect 4584 1297 4696 1303
rect 4904 1297 5048 1303
rect 5192 1297 5368 1303
rect 5480 1297 5512 1303
rect 5528 1297 5544 1303
rect -51 1277 1240 1283
rect 1256 1277 1272 1283
rect 1288 1277 1464 1283
rect 1480 1277 1528 1283
rect 2568 1277 2712 1283
rect 2728 1277 2776 1283
rect 2808 1277 3272 1283
rect 3304 1277 3704 1283
rect 3720 1277 3784 1283
rect 3912 1277 4312 1283
rect 4328 1277 4776 1283
rect 616 1257 1016 1263
rect 1560 1257 1752 1263
rect 1768 1257 2360 1263
rect 2616 1257 2808 1263
rect 2872 1257 2920 1263
rect 2936 1257 3448 1263
rect 4056 1257 4328 1263
rect 4744 1257 5128 1263
rect 5656 1257 5800 1263
rect 552 1237 648 1243
rect 824 1237 3000 1243
rect 3368 1237 3480 1243
rect 3544 1237 3768 1243
rect 4056 1237 4120 1243
rect 4456 1237 4664 1243
rect 4952 1237 5016 1243
rect 5240 1237 5288 1243
rect 5592 1237 5608 1243
rect 568 1217 776 1223
rect 1272 1217 2824 1223
rect 1256 1197 2632 1203
rect 2792 1197 2856 1203
rect 4168 1217 4696 1223
rect 3176 1197 3208 1203
rect 3592 1197 3720 1203
rect 3880 1197 4136 1203
rect 5304 1197 5528 1203
rect 1224 1177 1560 1183
rect 2296 1177 2312 1183
rect 2584 1177 2616 1183
rect 2632 1177 2680 1183
rect 2856 1177 3144 1183
rect 3160 1177 4200 1183
rect 4440 1177 4552 1183
rect 4872 1177 5096 1183
rect -51 1157 104 1163
rect 440 1157 520 1163
rect 936 1157 968 1163
rect 1016 1157 2008 1163
rect 2040 1157 2056 1163
rect 2088 1157 2168 1163
rect 2221 1157 2472 1163
rect 104 1137 424 1143
rect 808 1137 888 1143
rect 1272 1137 1288 1143
rect 2221 1143 2227 1157
rect 2520 1157 2568 1163
rect 2664 1157 3880 1163
rect 4184 1157 4472 1163
rect 4840 1157 4856 1163
rect 5176 1157 5224 1163
rect 5240 1157 5560 1163
rect 5576 1157 5608 1163
rect 1336 1137 2227 1143
rect 2248 1137 2360 1143
rect 2456 1137 2552 1143
rect 2680 1137 3048 1143
rect 3080 1137 4200 1143
rect 4504 1137 4696 1143
rect 5112 1137 5176 1143
rect 5432 1137 5528 1143
rect -51 1117 8 1123
rect 776 1117 824 1123
rect 872 1117 1080 1123
rect 1096 1117 1416 1123
rect 1432 1117 1656 1123
rect 1688 1117 1832 1123
rect 1864 1117 1960 1123
rect 1976 1117 2120 1123
rect 2136 1117 2328 1123
rect 2424 1117 2456 1123
rect 2808 1117 2840 1123
rect 2952 1117 2984 1123
rect 3032 1117 3064 1123
rect 3080 1117 3320 1123
rect 3368 1117 3528 1123
rect 3720 1117 3731 1123
rect 3976 1117 4456 1123
rect 4488 1117 5240 1123
rect 5496 1117 5672 1123
rect 5768 1117 5864 1123
rect 344 1097 392 1103
rect 744 1097 904 1103
rect 1288 1097 1304 1103
rect 1496 1097 1544 1103
rect 2072 1097 2104 1103
rect 2136 1097 2280 1103
rect 2696 1097 2760 1103
rect 2840 1097 3144 1103
rect 3160 1097 3176 1103
rect 3352 1097 3416 1103
rect 3576 1097 3592 1103
rect 3656 1097 3672 1103
rect 3752 1097 3768 1103
rect 3832 1097 3960 1103
rect 4072 1097 4104 1103
rect 4120 1097 4344 1103
rect 4360 1097 4552 1103
rect 4568 1097 4616 1103
rect 4632 1097 4680 1103
rect 4696 1097 4792 1103
rect 4936 1097 4952 1103
rect 5016 1097 5160 1103
rect 5640 1097 5704 1103
rect 1133 1088 1139 1092
rect 632 1077 680 1083
rect 728 1077 936 1083
rect 1192 1077 1336 1083
rect 1816 1077 1864 1083
rect 1880 1077 2008 1083
rect 2024 1077 2200 1083
rect 2216 1077 2280 1083
rect 2509 1083 2515 1092
rect 5869 1088 5875 1092
rect 2509 1077 2520 1083
rect 2728 1077 2984 1083
rect 3256 1077 3368 1083
rect 3432 1077 3448 1083
rect 3592 1077 3603 1083
rect 3656 1077 3752 1083
rect 3768 1077 3960 1083
rect 4264 1077 4392 1083
rect 4728 1077 4744 1083
rect 4760 1077 4872 1083
rect 4904 1077 5176 1083
rect 5192 1077 5224 1083
rect 5256 1077 5400 1083
rect 5704 1077 5816 1083
rect 5896 1077 5912 1083
rect 3549 1068 3555 1072
rect 424 1057 696 1063
rect 744 1057 1032 1063
rect 1224 1057 1336 1063
rect 1416 1057 1496 1063
rect 1768 1057 2200 1063
rect 2232 1057 2440 1063
rect 2888 1057 3160 1063
rect 3192 1057 3208 1063
rect 3224 1057 3320 1063
rect 3784 1057 3800 1063
rect 3848 1057 4040 1063
rect 4056 1057 4120 1063
rect 4168 1057 4184 1063
rect 4264 1057 4408 1063
rect 4424 1057 4632 1063
rect 4712 1057 4760 1063
rect 4776 1057 5208 1063
rect 5432 1057 5576 1063
rect 888 1037 984 1043
rect 1000 1037 1160 1043
rect 1176 1037 1400 1043
rect 1624 1037 1688 1043
rect 1928 1037 2136 1043
rect 2184 1037 2232 1043
rect 2264 1037 2840 1043
rect 3240 1037 3304 1043
rect 3336 1037 3480 1043
rect 3496 1037 3672 1043
rect 3896 1037 3944 1043
rect 3960 1037 4264 1043
rect 4440 1037 5032 1043
rect 5064 1037 5864 1043
rect 813 1028 819 1032
rect 680 1017 728 1023
rect 872 1017 1224 1023
rect 1480 1017 1816 1023
rect 680 997 1096 1003
rect 1592 997 1848 1003
rect 2056 1017 2296 1023
rect 2440 1017 2504 1023
rect 2520 1017 2568 1023
rect 3064 1017 3656 1023
rect 2200 997 2232 1003
rect 2536 997 2568 1003
rect 2600 997 2936 1003
rect 3112 997 3480 1003
rect 4280 1017 4440 1023
rect 4472 1017 4840 1023
rect 5144 1017 5416 1023
rect 5592 1017 5832 1023
rect 4152 997 4472 1003
rect 4552 997 4648 1003
rect 4680 997 4904 1003
rect 5192 997 5224 1003
rect 152 977 424 983
rect 888 977 968 983
rect 1112 977 1480 983
rect 1496 977 1560 983
rect 1736 977 1768 983
rect 1848 977 1928 983
rect 1944 977 2472 983
rect 2808 977 3192 983
rect 3320 977 3336 983
rect 3357 977 3688 983
rect -51 957 56 963
rect 424 957 616 963
rect 648 957 664 963
rect 904 957 968 963
rect 1320 957 1352 963
rect 1368 957 2264 963
rect 2312 957 2328 963
rect 2344 957 2392 963
rect 2904 957 2936 963
rect 3176 957 3192 963
rect 3224 957 3256 963
rect 3357 963 3363 977
rect 3816 977 3832 983
rect 4344 977 4456 983
rect 4488 977 4808 983
rect 5064 977 5080 983
rect 5288 977 5544 983
rect 5736 977 5752 983
rect 5784 977 5944 983
rect 4205 968 4211 972
rect 3288 957 3363 963
rect 3416 957 3448 963
rect 3496 957 3544 963
rect 3560 957 3576 963
rect 4056 957 4072 963
rect 4360 957 4376 963
rect 4536 957 4936 963
rect 5000 957 5144 963
rect 5160 957 5320 963
rect 5352 957 5384 963
rect 5544 957 5560 963
rect 5736 957 5800 963
rect 5816 957 5832 963
rect 1261 948 1267 952
rect 376 937 584 943
rect 936 937 1000 943
rect 1320 937 1544 943
rect 1560 937 1640 943
rect 1688 937 1752 943
rect 1768 937 1832 943
rect 1880 937 1896 943
rect 1928 937 1960 943
rect 1992 937 2008 943
rect 2072 937 2088 943
rect 2104 937 2296 943
rect 2424 937 2440 943
rect 2632 937 2648 943
rect 2680 937 2728 943
rect 2920 937 3080 943
rect 3096 937 3224 943
rect 3448 937 3512 943
rect 3528 937 3560 943
rect 3800 937 4280 943
rect 4312 937 4392 943
rect 4408 937 4456 943
rect 4600 937 4680 943
rect 4808 937 5224 943
rect 5336 937 5448 943
rect 5528 937 5640 943
rect 5752 937 5896 943
rect -51 917 8 923
rect 56 917 152 923
rect 344 917 392 923
rect 568 917 616 923
rect 856 917 904 923
rect 1144 917 1208 923
rect 1416 917 1432 923
rect 1528 917 1608 923
rect 2216 917 2248 923
rect 2504 917 2520 923
rect 2536 917 2632 923
rect 2968 917 3032 923
rect 3176 917 3256 923
rect 3544 917 3624 923
rect 3928 917 4616 923
rect 4664 917 4776 923
rect 4936 917 5208 923
rect 5272 917 5416 923
rect 5464 917 5480 923
rect 5576 917 5592 923
rect 472 897 1064 903
rect 1160 897 1176 903
rect 1240 897 1272 903
rect 1720 897 1944 903
rect 2184 897 2328 903
rect 2344 897 2504 903
rect 3256 897 3352 903
rect 3368 897 3432 903
rect 3496 897 3944 903
rect 5432 897 5448 903
rect 232 877 1080 883
rect 1096 877 1112 883
rect 1128 877 1288 883
rect 1304 877 1560 883
rect 1576 877 1656 883
rect 1704 877 1720 883
rect 1736 877 1848 883
rect 1864 877 1912 883
rect 2488 877 2536 883
rect 2552 877 2600 883
rect 2904 877 3064 883
rect 3080 877 3128 883
rect 3144 877 3208 883
rect 3880 877 4744 883
rect 680 857 696 863
rect 1272 857 1304 863
rect 1640 857 1768 863
rect 2440 857 2520 863
rect 2920 857 3171 863
rect 824 837 1224 843
rect 1640 837 1672 843
rect 2856 837 3048 843
rect 3165 843 3171 857
rect 3192 857 3256 863
rect 3336 857 3368 863
rect 3656 857 4696 863
rect 4712 857 4840 863
rect 3165 837 3640 843
rect 4264 837 4488 843
rect 1064 817 1128 823
rect 1192 817 1304 823
rect 1368 817 1880 823
rect 1896 817 2200 823
rect 2216 817 2472 823
rect 2696 817 2872 823
rect 1720 797 1816 803
rect 1832 797 2056 803
rect 2077 797 2408 803
rect 2077 783 2083 797
rect 2744 797 2888 803
rect 3784 817 4312 823
rect 3448 797 3640 803
rect 3960 797 4584 803
rect 888 777 2083 783
rect 2168 777 2184 783
rect 2216 777 2696 783
rect 2776 777 2840 783
rect 2872 777 3000 783
rect 3128 777 4056 783
rect 4792 777 4808 783
rect 4824 777 4840 783
rect 5384 777 5944 783
rect 968 757 1000 763
rect 1240 757 1528 763
rect 1544 757 2344 763
rect 2360 757 2680 763
rect 2696 757 2744 763
rect 3448 757 3544 763
rect 3576 757 4392 763
rect 4568 757 4776 763
rect 4952 757 5128 763
rect 5400 757 5544 763
rect 5560 757 5640 763
rect 104 737 328 743
rect 1112 737 1192 743
rect 1240 737 1256 743
rect 1272 737 1320 743
rect 1336 737 1368 743
rect 1432 737 1544 743
rect 1560 737 1656 743
rect 1800 737 1848 743
rect 1864 737 1912 743
rect 1928 737 2072 743
rect 2232 737 2280 743
rect 2296 737 2360 743
rect 2440 737 2584 743
rect 3032 737 3080 743
rect 3096 737 3112 743
rect 3128 737 3144 743
rect 3160 737 3176 743
rect 3512 737 3880 743
rect 4056 737 4104 743
rect 4120 737 4904 743
rect 5016 737 5096 743
rect -51 717 8 723
rect 328 717 648 723
rect 840 717 1000 723
rect 1160 717 1240 723
rect 1352 717 1432 723
rect 1608 717 1736 723
rect 1832 717 1864 723
rect 1880 717 2088 723
rect 2120 717 2168 723
rect 2328 717 2376 723
rect 2536 717 2568 723
rect 2840 717 2920 723
rect 2936 717 2984 723
rect 3144 717 3224 723
rect 3784 717 3912 723
rect 3944 717 4200 723
rect 4488 717 4520 723
rect 4648 717 4936 723
rect 4968 717 5112 723
rect 5128 717 5288 723
rect 5832 717 5912 723
rect 2445 708 2451 712
rect 2733 708 2739 712
rect 3629 708 3635 712
rect 248 697 296 703
rect 472 697 552 703
rect 584 697 648 703
rect 664 697 840 703
rect 984 697 1032 703
rect 1272 697 1400 703
rect 1448 697 1480 703
rect 1496 697 1544 703
rect 1768 697 1896 703
rect 2056 697 2136 703
rect 2168 697 2200 703
rect 2216 697 2392 703
rect 2536 697 2547 703
rect 600 677 776 683
rect 1080 677 1112 683
rect 1128 677 1480 683
rect 1496 677 1736 683
rect 1864 677 1896 683
rect 1960 677 2248 683
rect 2509 683 2515 692
rect 2541 688 2547 697
rect 2776 697 2792 703
rect 2856 697 2968 703
rect 3016 697 3112 703
rect 3128 697 3176 703
rect 3224 697 3384 703
rect 3464 697 3475 703
rect 3704 697 3816 703
rect 3912 697 4136 703
rect 4248 697 4264 703
rect 4296 697 4328 703
rect 4456 697 4968 703
rect 5192 697 5288 703
rect 5320 697 5432 703
rect 5448 697 5640 703
rect 5688 697 5896 703
rect 2509 677 2520 683
rect 2760 677 3528 683
rect 3816 677 3848 683
rect 4072 677 4120 683
rect 4328 677 4568 683
rect 4632 677 4648 683
rect 4744 677 4760 683
rect 4840 677 5320 683
rect 5432 677 5464 683
rect 5480 677 5496 683
rect 5672 677 5736 683
rect 5752 677 5832 683
rect 552 657 584 663
rect 760 657 904 663
rect 1016 657 1208 663
rect 1224 657 1448 663
rect 1512 657 1656 663
rect 1672 657 1720 663
rect 1912 657 2200 663
rect 2232 657 2280 663
rect 2536 657 2584 663
rect 2632 657 3656 663
rect 3688 657 3784 663
rect 3928 657 4200 663
rect 4392 657 4584 663
rect 4712 657 4760 663
rect 5000 657 5240 663
rect 5256 657 5288 663
rect 5736 657 5752 663
rect 5832 657 5880 663
rect 648 637 712 643
rect 904 637 1016 643
rect 1048 637 1672 643
rect 2120 637 2707 643
rect 488 617 1000 623
rect 1528 617 1560 623
rect 1656 617 1896 623
rect 648 597 840 603
rect 1752 597 1923 603
rect 2264 617 2680 623
rect 2701 623 2707 637
rect 2872 637 2920 643
rect 3192 637 3272 643
rect 3528 637 3576 643
rect 3592 637 3704 643
rect 3976 637 4120 643
rect 4136 637 4184 643
rect 4200 637 4264 643
rect 4392 637 4456 643
rect 5224 637 5304 643
rect 2701 617 3592 623
rect 520 577 536 583
rect 552 577 600 583
rect 920 577 1032 583
rect 1576 577 1672 583
rect 1752 577 1880 583
rect 1917 583 1923 597
rect 2152 597 2424 603
rect 2728 597 2760 603
rect 3384 597 3400 603
rect 3512 597 3720 603
rect 4136 617 4184 623
rect 4200 617 4312 623
rect 4920 617 4936 623
rect 4952 617 4968 623
rect 4984 617 5064 623
rect 5624 617 5720 623
rect 4648 597 4712 603
rect 4760 597 4872 603
rect 4888 597 5096 603
rect 5112 597 5208 603
rect 5224 597 5240 603
rect 5352 597 5528 603
rect 5720 597 5880 603
rect 1917 577 2616 583
rect 2632 577 2760 583
rect 2824 577 2904 583
rect 3048 577 3192 583
rect 3208 577 3240 583
rect 3320 577 3848 583
rect 3880 577 3976 583
rect 4312 577 4680 583
rect 4696 577 4872 583
rect 4904 577 5112 583
rect 5288 577 5496 583
rect 5560 577 5768 583
rect 5784 577 5800 583
rect 584 557 616 563
rect 632 557 728 563
rect 824 557 872 563
rect 968 557 1160 563
rect 1208 557 1256 563
rect 1304 557 1512 563
rect 1560 557 1624 563
rect 1928 557 1944 563
rect 2696 557 2888 563
rect 3064 557 3096 563
rect 3144 557 3320 563
rect 3640 557 3816 563
rect 3848 557 4056 563
rect 4072 557 4120 563
rect 4141 557 4152 563
rect 4248 557 4376 563
rect 4440 557 4552 563
rect 4696 557 4867 563
rect 232 537 584 543
rect 616 537 632 543
rect 664 537 968 543
rect 984 537 1016 543
rect 1160 537 1320 543
rect 1592 537 1656 543
rect 1672 537 1688 543
rect 1720 537 1848 543
rect 1944 537 1976 543
rect 2312 537 2408 543
rect 2472 537 2552 543
rect 2968 537 3064 543
rect 3096 537 3144 543
rect 3160 537 3256 543
rect 3784 537 3795 543
rect 3832 537 4504 543
rect 4520 537 4840 543
rect 4861 543 4867 557
rect 4952 557 5144 563
rect 5416 557 5512 563
rect 5624 557 5704 563
rect 5736 557 5864 563
rect 5933 563 5939 572
rect 5928 557 5939 563
rect 4861 537 5000 543
rect 5112 537 5224 543
rect 5240 537 5400 543
rect 5432 537 5576 543
rect 5752 537 5848 543
rect -51 517 8 523
rect 328 517 616 523
rect 632 517 696 523
rect 1032 517 2232 523
rect 2248 517 2328 523
rect 2349 508 2355 523
rect 2536 517 2616 523
rect 2872 517 2952 523
rect 2984 517 3016 523
rect 3032 517 3128 523
rect 3160 517 3192 523
rect 3208 517 3400 523
rect 3672 517 3768 523
rect 3784 517 3912 523
rect 4072 517 4328 523
rect 4504 517 4536 523
rect 4568 517 4776 523
rect 4840 517 5064 523
rect 5096 517 5144 523
rect 5160 517 5320 523
rect 5368 517 5379 523
rect 440 497 552 503
rect 760 497 1224 503
rect 1256 497 1432 503
rect 1608 497 1624 503
rect 1640 497 1736 503
rect 1816 497 1880 503
rect 2408 497 2488 503
rect 2520 497 2568 503
rect 2584 497 2600 503
rect 2936 497 2952 503
rect 2968 497 3000 503
rect 3016 497 3080 503
rect 3160 497 3240 503
rect 3656 497 3667 503
rect 4120 497 4520 503
rect 4536 497 4648 503
rect 280 477 488 483
rect 504 477 568 483
rect 1000 477 1048 483
rect 1336 477 3208 483
rect 4296 477 4488 483
rect 4632 477 5224 483
rect 872 457 968 463
rect 1512 457 1576 463
rect 1704 457 1736 463
rect 1768 457 1800 463
rect 1832 457 1848 463
rect 1864 457 1944 463
rect 4568 457 4696 463
rect 232 437 296 443
rect 472 437 520 443
rect 1064 437 2248 443
rect 2264 437 2312 443
rect 2568 437 2600 443
rect 2696 437 3464 443
rect 5576 437 5736 443
rect 1400 417 1528 423
rect 2088 417 2120 423
rect 1320 397 1640 403
rect 1688 397 1768 403
rect 1784 397 1976 403
rect 1992 397 2056 403
rect 2072 397 2216 403
rect 3400 397 4280 403
rect 4552 397 4712 403
rect 4728 397 4856 403
rect 5176 417 5464 423
rect 5480 417 5608 423
rect 5608 397 5624 403
rect 808 377 1064 383
rect 1672 377 1752 383
rect 1768 377 1784 383
rect 1928 377 2024 383
rect 2696 377 3928 383
rect 4456 377 5160 383
rect 5640 377 5864 383
rect 1592 357 2680 363
rect 2744 357 3272 363
rect 3704 357 5016 363
rect 1240 337 1731 343
rect -51 317 8 323
rect 760 317 1304 323
rect 1725 323 1731 337
rect 1960 337 2024 343
rect 2056 337 3352 343
rect 3848 337 4056 343
rect 4072 337 4472 343
rect 4936 337 4968 343
rect 4984 337 5112 343
rect 5784 337 5800 343
rect 5149 328 5155 332
rect 1725 317 2632 323
rect 3064 317 3368 323
rect 3544 317 3784 323
rect 3976 317 4072 323
rect 4328 317 4760 323
rect 4792 317 4824 323
rect 4840 317 4952 323
rect 4968 317 5000 323
rect 5256 317 5432 323
rect 5736 317 5928 323
rect 1709 308 1715 312
rect 680 297 728 303
rect 1112 297 1128 303
rect 1176 297 1352 303
rect 1480 297 1496 303
rect 1736 297 1848 303
rect 2136 297 2360 303
rect 2792 297 2840 303
rect 2872 297 2984 303
rect 3176 297 3224 303
rect 3368 297 3432 303
rect 3512 297 3592 303
rect 3912 297 4248 303
rect 4344 297 4376 303
rect 4392 297 4456 303
rect 4504 297 4552 303
rect 4952 297 5288 303
rect 5336 297 5384 303
rect 5400 297 5496 303
rect 5512 297 5576 303
rect 5624 297 5880 303
rect 5896 297 5944 303
rect 989 277 1000 283
rect 1128 277 1176 283
rect 1496 277 1592 283
rect 1752 277 1800 283
rect 1816 277 1848 283
rect 2296 277 2328 283
rect 2392 277 3384 283
rect 3416 277 3512 283
rect 3912 277 4072 283
rect 4280 277 4344 283
rect 4408 277 4419 283
rect 4808 277 4835 283
rect 616 257 808 263
rect 1560 257 1576 263
rect 1896 257 1960 263
rect 1976 257 2040 263
rect 2056 257 2088 263
rect 2616 257 3192 263
rect 3432 257 3480 263
rect 4344 257 4392 263
rect 4760 257 4808 263
rect 4829 263 4835 277
rect 5128 277 5192 283
rect 5224 277 5448 283
rect 5480 277 5624 283
rect 5640 277 5688 283
rect 5704 277 5752 283
rect 4829 257 5480 263
rect 5608 257 5672 263
rect 552 237 632 243
rect 712 237 744 243
rect 952 237 1000 243
rect 1256 237 1304 243
rect 1640 237 2312 243
rect 2328 237 2344 243
rect 3000 237 3080 243
rect 3288 237 3560 243
rect 3576 237 3752 243
rect 4184 237 5240 243
rect 5336 237 5896 243
rect 888 197 1528 203
rect 1992 217 2136 223
rect 2248 217 2392 223
rect 2136 197 2392 203
rect 2408 197 2776 203
rect 3480 197 3624 203
rect 4632 217 4680 223
rect 4920 217 4952 223
rect 4968 217 5224 223
rect 5464 217 5704 223
rect 4088 197 4216 203
rect 4392 197 5112 203
rect 5288 197 5352 203
rect 5560 197 5576 203
rect 5800 197 5832 203
rect 520 177 840 183
rect 856 177 1272 183
rect 1288 177 2072 183
rect 2088 177 2600 183
rect 3208 177 3864 183
rect 3928 177 4088 183
rect 4152 177 4632 183
rect 5080 177 5128 183
rect 5144 177 5208 183
rect 5224 177 5336 183
rect 5352 177 5592 183
rect 5736 177 5784 183
rect 1432 157 1976 163
rect 2136 157 2152 163
rect 3128 157 3304 163
rect 3320 157 3528 163
rect 3768 157 4264 163
rect 4280 157 4520 163
rect 4536 157 4680 163
rect 4840 157 5320 163
rect 5336 157 5384 163
rect 5400 157 5512 163
rect 5544 157 5608 163
rect 5949 148 5955 152
rect 1416 137 1448 143
rect 1464 137 1512 143
rect 1528 137 2104 143
rect 2376 137 2440 143
rect 2856 137 3352 143
rect 3752 137 4072 143
rect 4936 137 4968 143
rect 5160 137 5352 143
rect 5416 137 5736 143
rect 5768 137 5928 143
rect -51 117 8 123
rect 248 117 296 123
rect 584 117 856 123
rect 1256 117 1400 123
rect 1800 117 1832 123
rect 2056 117 2104 123
rect 2200 117 2696 123
rect 2760 117 2808 123
rect 3336 117 3384 123
rect 3688 117 3720 123
rect 3944 117 4104 123
rect 4248 117 4296 123
rect 4664 117 4712 123
rect 5016 117 5080 123
rect 5112 117 5416 123
rect 5464 117 5544 123
rect 5800 117 5864 123
rect 792 97 840 103
rect 856 97 1480 103
rect 1496 97 3240 103
rect 5544 97 5800 103
rect 2488 57 2536 63
rect 1704 37 1720 43
rect 1832 37 1880 43
rect 1912 37 1976 43
rect 216 17 232 23
rect 1000 17 1016 23
rect 1240 17 1256 23
rect 1720 17 1736 23
rect 1768 17 1816 23
rect 3672 17 3688 23
rect 3720 17 3736 23
rect 4552 17 4568 23
<< m4contact >>
rect 792 4012 808 4028
rect 926 4002 954 4018
rect 2744 4012 2760 4028
rect 2920 4012 2936 4028
rect 2974 4002 3002 4018
rect 3320 4012 3336 4028
rect 3576 4012 3592 4028
rect 3640 4012 3656 4028
rect 4040 4012 4056 4028
rect 4168 4012 4184 4028
rect 3720 3992 3736 4008
rect 5022 4002 5050 4018
rect 712 3972 728 3988
rect 2024 3972 2040 3988
rect 4264 3972 4280 3988
rect 1352 3952 1368 3968
rect 1208 3932 1224 3948
rect 2024 3932 2040 3948
rect 3192 3932 3208 3948
rect 3336 3932 3352 3948
rect 4248 3932 4264 3948
rect 4824 3932 4840 3948
rect 200 3912 216 3928
rect 968 3912 984 3928
rect 2136 3912 2152 3928
rect 2328 3912 2344 3928
rect 648 3892 664 3908
rect 936 3892 952 3908
rect 1176 3892 1192 3908
rect 3608 3892 3624 3908
rect 3720 3892 3736 3908
rect 328 3872 344 3888
rect 392 3872 408 3888
rect 1624 3872 1640 3888
rect 2248 3872 2264 3888
rect 2296 3872 2312 3888
rect 2392 3872 2408 3888
rect 2552 3872 2568 3888
rect 2712 3872 2728 3888
rect 2808 3872 2824 3888
rect 3656 3872 3672 3888
rect 4248 3872 4264 3888
rect 4456 3892 4472 3908
rect 5320 3892 5336 3908
rect 5336 3892 5352 3908
rect 4376 3872 4392 3888
rect 4600 3872 4616 3888
rect 5416 3872 5432 3888
rect 5880 3872 5896 3888
rect 4520 3852 4536 3868
rect 4584 3852 4600 3868
rect 920 3832 936 3848
rect 1720 3832 1736 3848
rect 1288 3812 1304 3828
rect 1934 3802 1962 3818
rect 3448 3812 3464 3828
rect 3224 3792 3240 3808
rect 3304 3792 3320 3808
rect 3720 3792 3736 3808
rect 3982 3802 4010 3818
rect 4168 3812 4184 3828
rect 4568 3812 4584 3828
rect 4856 3812 4872 3828
rect 24 3772 40 3788
rect 1208 3772 1224 3788
rect 2776 3772 2792 3788
rect 4344 3792 4360 3808
rect 4248 3772 4264 3788
rect 2680 3752 2696 3768
rect 3528 3752 3544 3768
rect 4840 3752 4856 3768
rect 24 3732 40 3748
rect 856 3732 872 3748
rect 1944 3732 1960 3748
rect 1048 3712 1064 3728
rect 1560 3712 1576 3728
rect 1896 3712 1912 3728
rect 2440 3732 2456 3748
rect 4344 3732 4360 3748
rect 4824 3732 4840 3748
rect 5784 3732 5800 3748
rect 2168 3712 2184 3728
rect 2296 3712 2312 3728
rect 2472 3712 2488 3728
rect 2936 3712 2952 3728
rect 3256 3712 3272 3728
rect 3304 3712 3336 3728
rect 3448 3712 3480 3728
rect 3512 3712 3528 3728
rect 3944 3712 3960 3728
rect 4648 3712 4664 3728
rect 5688 3712 5704 3728
rect 5752 3712 5768 3728
rect 872 3692 888 3708
rect 1080 3692 1096 3708
rect 1928 3692 1944 3708
rect 2280 3692 2296 3708
rect 2664 3692 2680 3708
rect 2744 3692 2760 3708
rect 1112 3672 1128 3688
rect 2904 3672 2920 3688
rect 3384 3692 3416 3708
rect 3784 3692 3800 3708
rect 3928 3692 3944 3708
rect 3960 3692 3976 3708
rect 3592 3672 3608 3688
rect 3672 3672 3688 3688
rect 5400 3692 5416 3708
rect 4840 3672 4856 3688
rect 3624 3652 3640 3668
rect 4120 3652 4136 3668
rect 5336 3652 5352 3668
rect 728 3632 744 3648
rect 1848 3632 1864 3648
rect 3128 3632 3144 3648
rect 3416 3632 3432 3648
rect 3560 3632 3576 3648
rect 4344 3632 4360 3648
rect 4968 3632 4984 3648
rect 5176 3632 5192 3648
rect 5560 3632 5576 3648
rect 5832 3632 5848 3648
rect 872 3612 888 3628
rect 926 3602 954 3618
rect 1304 3612 1320 3628
rect 2872 3592 2888 3608
rect 2974 3602 3002 3618
rect 3576 3612 3592 3628
rect 5022 3602 5050 3618
rect 5800 3612 5816 3628
rect 5720 3592 5736 3608
rect 2200 3572 2216 3588
rect 2616 3552 2632 3568
rect 4664 3552 4680 3568
rect 4728 3552 4744 3568
rect 5752 3552 5768 3568
rect 2472 3532 2488 3548
rect 5336 3532 5352 3548
rect 472 3512 488 3528
rect 2520 3512 2536 3528
rect 2872 3512 2888 3528
rect 3496 3512 3512 3528
rect 5208 3512 5224 3528
rect 5704 3512 5720 3528
rect 56 3492 72 3508
rect 2232 3492 2248 3508
rect 2712 3492 2728 3508
rect 3432 3492 3448 3508
rect 4200 3492 4216 3508
rect 5864 3492 5880 3508
rect 2984 3472 3000 3488
rect 3528 3472 3544 3488
rect 3896 3472 3912 3488
rect 1656 3452 1672 3468
rect 3336 3452 3352 3468
rect 4152 3472 4168 3488
rect 5240 3472 5256 3488
rect 4792 3452 4808 3468
rect 5368 3452 5384 3468
rect 1128 3432 1144 3448
rect 2232 3432 2248 3448
rect 2568 3432 2584 3448
rect 3112 3432 3128 3448
rect 4584 3432 4600 3448
rect 4872 3432 4888 3448
rect 5448 3432 5464 3448
rect 1288 3392 1304 3408
rect 1934 3402 1962 3418
rect 2952 3412 2968 3428
rect 3512 3412 3528 3428
rect 3528 3412 3544 3428
rect 3544 3412 3560 3428
rect 2552 3392 2568 3408
rect 2680 3392 2696 3408
rect 2744 3392 2760 3408
rect 3176 3392 3192 3408
rect 3982 3402 4010 3418
rect 4856 3412 4872 3428
rect 5544 3392 5560 3408
rect 56 3372 72 3388
rect 2104 3372 2120 3388
rect 2200 3372 2216 3388
rect 4056 3372 4072 3388
rect 3096 3352 3112 3368
rect 3176 3352 3192 3368
rect 3352 3352 3368 3368
rect 4232 3352 4248 3368
rect 4264 3352 4280 3368
rect 4664 3352 4680 3368
rect 728 3332 744 3348
rect 1400 3332 1416 3348
rect 1496 3332 1512 3348
rect 1512 3332 1528 3348
rect 2344 3332 2360 3348
rect 2520 3332 2536 3348
rect 4600 3332 4632 3348
rect 5064 3332 5080 3348
rect 5336 3332 5352 3348
rect 2264 3312 2280 3328
rect 3016 3312 3032 3328
rect 3368 3312 3384 3328
rect 3544 3312 3560 3328
rect 3688 3312 3704 3328
rect 4104 3312 4120 3328
rect 4328 3312 4344 3328
rect 4536 3312 4552 3328
rect 4952 3312 4968 3328
rect 5768 3312 5784 3328
rect 1688 3292 1704 3308
rect 2584 3292 2600 3308
rect 2616 3272 2632 3288
rect 3208 3292 3224 3308
rect 3816 3292 3832 3308
rect 5576 3292 5592 3308
rect 5448 3272 5464 3288
rect 840 3252 856 3268
rect 3736 3252 3752 3268
rect 5896 3252 5912 3268
rect 184 3232 200 3248
rect 456 3232 472 3248
rect 1912 3232 1928 3248
rect 4136 3232 4152 3248
rect 5224 3232 5240 3248
rect 5736 3232 5752 3248
rect 926 3202 954 3218
rect 2920 3212 2936 3228
rect 2974 3202 3002 3218
rect 4216 3192 4232 3208
rect 5022 3202 5050 3218
rect 5752 3212 5768 3228
rect 5112 3192 5128 3208
rect 5432 3192 5448 3208
rect 4568 3172 4584 3188
rect 5688 3152 5704 3168
rect 3256 3132 3272 3148
rect 3960 3132 3976 3148
rect 1128 3112 1144 3128
rect 2392 3112 2408 3128
rect 3080 3112 3096 3128
rect 3480 3112 3496 3128
rect 3624 3112 3640 3128
rect 4456 3112 4472 3128
rect 5640 3112 5656 3128
rect 632 3092 648 3108
rect 1096 3092 1112 3108
rect 3608 3092 3624 3108
rect 4424 3092 4440 3108
rect 4648 3092 4664 3108
rect 5704 3092 5720 3108
rect 1160 3072 1176 3088
rect 1224 3072 1240 3088
rect 2360 3072 2376 3088
rect 3016 3072 3048 3088
rect 3384 3072 3400 3088
rect 3832 3052 3864 3068
rect 4200 3072 4216 3088
rect 4904 3072 4920 3088
rect 5528 3072 5544 3088
rect 5816 3072 5832 3088
rect 4568 3052 4584 3068
rect 4952 3052 4968 3068
rect 4968 3052 4984 3068
rect 2872 3032 2888 3048
rect 2936 3032 2952 3048
rect 3544 3032 3560 3048
rect 3896 3032 3912 3048
rect 696 3012 712 3028
rect 1912 3012 1928 3028
rect 1934 3002 1962 3018
rect 5320 3032 5336 3048
rect 5960 3032 5976 3048
rect 2072 2992 2088 3008
rect 3528 2992 3544 3008
rect 3960 2992 3976 3008
rect 3982 3002 4010 3018
rect 4568 3012 4584 3028
rect 5000 3012 5016 3028
rect 2488 2972 2504 2988
rect 2632 2972 2648 2988
rect 2664 2972 2680 2988
rect 3176 2972 3192 2988
rect 4040 2972 4056 2988
rect 632 2952 648 2968
rect 184 2932 200 2948
rect 1096 2932 1112 2948
rect 2632 2932 2648 2948
rect 2808 2932 2840 2948
rect 2904 2932 2920 2948
rect 3544 2952 3560 2968
rect 3912 2952 3928 2968
rect 4680 2952 4696 2968
rect 5288 2952 5304 2968
rect 5416 2972 5432 2988
rect 3592 2932 3608 2948
rect 5240 2932 5256 2948
rect 5304 2932 5320 2948
rect 5864 2932 5880 2948
rect 696 2912 712 2928
rect 1496 2912 1512 2928
rect 3192 2912 3208 2928
rect 3368 2912 3384 2928
rect 3480 2912 3496 2928
rect 4696 2912 4712 2928
rect 4952 2912 4968 2928
rect 3528 2892 3544 2908
rect 4664 2892 4680 2908
rect 3688 2872 3704 2888
rect 3800 2872 3816 2888
rect 3944 2872 3960 2888
rect 5176 2872 5192 2888
rect 984 2852 1000 2868
rect 2952 2852 2968 2868
rect 760 2832 776 2848
rect 4136 2852 4152 2868
rect 4728 2852 4744 2868
rect 3240 2832 3256 2848
rect 3848 2832 3864 2848
rect 4296 2832 4312 2848
rect 4904 2832 4920 2848
rect 5752 2832 5768 2848
rect 5864 2832 5880 2848
rect 840 2812 856 2828
rect 926 2802 954 2818
rect 2312 2792 2328 2808
rect 2974 2802 3002 2818
rect 3032 2812 3048 2828
rect 3528 2812 3544 2828
rect 4024 2792 4056 2808
rect 5022 2802 5050 2818
rect 5512 2812 5528 2828
rect 5656 2812 5672 2828
rect 5208 2792 5224 2808
rect 4216 2772 4232 2788
rect 5704 2772 5720 2788
rect 3224 2752 3240 2768
rect 3848 2752 3864 2768
rect 4056 2752 4072 2768
rect 4120 2752 4136 2768
rect 5576 2752 5592 2768
rect 1896 2732 1912 2748
rect 4344 2732 4360 2748
rect 4440 2732 4456 2748
rect 5064 2732 5080 2748
rect 2072 2712 2088 2728
rect 2520 2712 2536 2728
rect 3352 2712 3368 2728
rect 3416 2712 3432 2728
rect 4424 2712 4440 2728
rect 4600 2712 4616 2728
rect 72 2692 88 2708
rect 1064 2692 1080 2708
rect 1432 2692 1448 2708
rect 3656 2692 3672 2708
rect 456 2672 472 2688
rect 2712 2672 2728 2688
rect 3240 2672 3256 2688
rect 3560 2672 3576 2688
rect 3592 2672 3608 2688
rect 3640 2672 3656 2688
rect 5496 2692 5512 2708
rect 3912 2672 3928 2688
rect 5544 2672 5560 2688
rect 5672 2672 5688 2688
rect 72 2652 88 2668
rect 4472 2652 4488 2668
rect 5864 2652 5880 2668
rect 808 2632 824 2648
rect 2104 2632 2120 2648
rect 3032 2632 3064 2648
rect 3640 2632 3656 2648
rect 3704 2632 3720 2648
rect 4152 2632 4168 2648
rect 4184 2632 4200 2648
rect 5848 2632 5864 2648
rect 584 2612 600 2628
rect 1934 2602 1962 2618
rect 2168 2612 2184 2628
rect 3208 2612 3224 2628
rect 2904 2592 2920 2608
rect 3864 2592 3880 2608
rect 3982 2602 4010 2618
rect 4904 2612 4920 2628
rect 4968 2612 4984 2628
rect 4104 2592 4120 2608
rect 5240 2592 5256 2608
rect 1560 2572 1576 2588
rect 3640 2572 3656 2588
rect 5928 2572 5944 2588
rect 2440 2552 2456 2568
rect 2520 2552 2536 2568
rect 2904 2552 2920 2568
rect 3240 2552 3256 2568
rect 4440 2552 4456 2568
rect 5912 2552 5928 2568
rect 1896 2532 1912 2548
rect 1976 2532 1992 2548
rect 2200 2532 2216 2548
rect 2312 2532 2328 2548
rect 2424 2532 2440 2548
rect 2744 2532 2760 2548
rect 3224 2532 3240 2548
rect 3400 2532 3416 2548
rect 5112 2532 5128 2548
rect 5224 2532 5240 2548
rect 5864 2532 5880 2548
rect 2040 2512 2056 2528
rect 3224 2512 3240 2528
rect 3320 2512 3336 2528
rect 3432 2512 3448 2528
rect 3960 2512 3976 2528
rect 4152 2512 4168 2528
rect 5400 2512 5416 2528
rect 5720 2512 5736 2528
rect 2056 2492 2072 2508
rect 4856 2492 4872 2508
rect 3112 2472 3128 2488
rect 3896 2472 3912 2488
rect 4296 2472 4312 2488
rect 760 2452 776 2468
rect 3240 2452 3256 2468
rect 3448 2452 3464 2468
rect 4472 2452 4488 2468
rect 4984 2452 5000 2468
rect 376 2432 392 2448
rect 792 2432 808 2448
rect 3048 2432 3064 2448
rect 5896 2432 5912 2448
rect 926 2402 954 2418
rect 2136 2412 2152 2428
rect 2808 2412 2824 2428
rect 2974 2402 3002 2418
rect 3704 2412 3720 2428
rect 4120 2412 4136 2428
rect 4696 2412 4712 2428
rect 4840 2412 4856 2428
rect 3544 2392 3560 2408
rect 4424 2392 4440 2408
rect 5022 2402 5050 2418
rect 5192 2412 5208 2428
rect 5208 2412 5224 2428
rect 5592 2412 5608 2428
rect 1240 2372 1256 2388
rect 2072 2372 2088 2388
rect 4568 2372 4584 2388
rect 5528 2372 5544 2388
rect 808 2352 824 2368
rect 2088 2352 2104 2368
rect 2952 2352 2968 2368
rect 5320 2352 5336 2368
rect 2776 2332 2792 2348
rect 5576 2332 5592 2348
rect 3096 2312 3112 2328
rect 5320 2312 5336 2328
rect 5528 2312 5544 2328
rect 584 2292 600 2308
rect 616 2292 632 2308
rect 984 2292 1000 2308
rect 1512 2292 1528 2308
rect 1816 2292 1832 2308
rect 1912 2292 1928 2308
rect 3096 2292 3112 2308
rect 3224 2292 3240 2308
rect 3336 2292 3352 2308
rect 3720 2292 3752 2308
rect 4968 2292 4984 2308
rect 5496 2292 5512 2308
rect 5752 2292 5784 2308
rect 696 2272 712 2288
rect 792 2272 808 2288
rect 2072 2272 2088 2288
rect 2312 2272 2328 2288
rect 2568 2272 2584 2288
rect 3144 2272 3160 2288
rect 3480 2272 3496 2288
rect 3928 2272 3944 2288
rect 4104 2272 4120 2288
rect 4392 2272 4408 2288
rect 4856 2272 4872 2288
rect 5032 2272 5048 2288
rect 5304 2272 5320 2288
rect 5416 2272 5432 2288
rect 5816 2272 5832 2288
rect 888 2252 904 2268
rect 376 2232 392 2248
rect 2072 2232 2088 2248
rect 2184 2232 2200 2248
rect 2376 2232 2392 2248
rect 2456 2232 2472 2248
rect 2968 2232 2984 2248
rect 3784 2252 3800 2268
rect 5176 2252 5192 2268
rect 3672 2232 3688 2248
rect 3704 2232 3720 2248
rect 5576 2232 5592 2248
rect 680 2212 696 2228
rect 808 2212 824 2228
rect 1016 2212 1032 2228
rect 1934 2202 1962 2218
rect 2168 2212 2184 2228
rect 2120 2192 2136 2208
rect 2424 2192 2440 2208
rect 3896 2212 3912 2228
rect 2792 2192 2808 2208
rect 2904 2192 2920 2208
rect 3832 2192 3848 2208
rect 3982 2202 4010 2218
rect 4056 2212 4072 2228
rect 4568 2212 4584 2228
rect 5768 2212 5784 2228
rect 4024 2192 4040 2208
rect 4632 2192 4648 2208
rect 5288 2192 5304 2208
rect 488 2172 504 2188
rect 1896 2172 1912 2188
rect 2392 2172 2408 2188
rect 2648 2172 2664 2188
rect 2728 2172 2744 2188
rect 2904 2172 2920 2188
rect 3464 2172 3480 2188
rect 3832 2172 3864 2188
rect 4168 2172 4184 2188
rect 5864 2172 5880 2188
rect 360 2152 376 2168
rect 392 2132 408 2148
rect 776 2132 792 2148
rect 808 2132 824 2148
rect 1192 2132 1208 2148
rect 1528 2152 1544 2168
rect 2104 2152 2120 2168
rect 2792 2152 2824 2168
rect 4824 2152 4840 2168
rect 5496 2152 5512 2168
rect 5720 2152 5736 2168
rect 1832 2132 1848 2148
rect 2152 2132 2184 2148
rect 2712 2132 2728 2148
rect 2872 2132 2888 2148
rect 3624 2132 3640 2148
rect 3816 2132 3832 2148
rect 4472 2132 4488 2148
rect 5000 2132 5016 2148
rect 5608 2132 5624 2148
rect 5880 2132 5896 2148
rect 696 2112 712 2128
rect 2488 2112 2504 2128
rect 3192 2112 3208 2128
rect 3368 2112 3384 2128
rect 4136 2112 4152 2128
rect 4344 2112 4360 2128
rect 4872 2112 4888 2128
rect 5624 2112 5640 2128
rect 216 2092 232 2108
rect 968 2092 984 2108
rect 1656 2092 1672 2108
rect 2504 2092 2520 2108
rect 2616 2092 2632 2108
rect 2648 2092 2664 2108
rect 2888 2092 2904 2108
rect 3480 2092 3496 2108
rect 4968 2092 4984 2108
rect 5016 2092 5032 2108
rect 5336 2092 5352 2108
rect 4216 2072 4232 2088
rect 5112 2072 5128 2088
rect 2200 2052 2216 2068
rect 4136 2052 4152 2068
rect 4232 2052 4248 2068
rect 600 2032 616 2048
rect 1448 2032 1464 2048
rect 3784 2032 3800 2048
rect 5544 2032 5560 2048
rect 926 2002 954 2018
rect 2440 2012 2456 2028
rect 2872 2012 2888 2028
rect 2248 1992 2264 2008
rect 2974 2002 3002 2018
rect 3848 2012 3864 2028
rect 4296 2012 4312 2028
rect 4312 1992 4328 2008
rect 4520 1992 4536 2008
rect 5000 1992 5016 2008
rect 5022 2002 5050 2018
rect 4136 1972 4168 1988
rect 1912 1952 1928 1968
rect 2136 1952 2152 1968
rect 2712 1952 2728 1968
rect 3272 1952 3288 1968
rect 3800 1952 3816 1968
rect 3880 1952 3896 1968
rect 3928 1952 3944 1968
rect 4152 1952 4168 1968
rect 4616 1952 4632 1968
rect 1704 1932 1720 1948
rect 2008 1932 2040 1948
rect 2584 1932 2600 1948
rect 2696 1932 2712 1948
rect 2792 1932 2808 1948
rect 1720 1912 1736 1928
rect 2392 1912 2408 1928
rect 5400 1932 5416 1948
rect 3720 1912 3736 1928
rect 472 1892 488 1908
rect 760 1892 776 1908
rect 1736 1892 1752 1908
rect 2216 1892 2248 1908
rect 2664 1892 2680 1908
rect 2920 1892 2936 1908
rect 776 1872 792 1888
rect 2184 1872 2200 1888
rect 2648 1872 2680 1888
rect 2696 1872 2712 1888
rect 2856 1872 2872 1888
rect 3048 1872 3064 1888
rect 3144 1872 3160 1888
rect 3496 1892 3512 1908
rect 4136 1912 4152 1928
rect 4296 1912 4312 1928
rect 4248 1892 4264 1908
rect 4296 1892 4312 1908
rect 5576 1892 5592 1908
rect 5624 1892 5640 1908
rect 3688 1872 3704 1888
rect 3720 1872 3736 1888
rect 3864 1872 3880 1888
rect 3960 1872 3976 1888
rect 4168 1872 4184 1888
rect 4632 1872 4648 1888
rect 5672 1872 5688 1888
rect 5864 1872 5880 1888
rect 472 1852 488 1868
rect 1288 1852 1304 1868
rect 1944 1852 1960 1868
rect 2696 1852 2712 1868
rect 3048 1852 3064 1868
rect 3336 1852 3352 1868
rect 4248 1852 4264 1868
rect 4424 1852 4440 1868
rect 4968 1852 4984 1868
rect 5240 1852 5256 1868
rect 5944 1852 5960 1868
rect 520 1832 536 1848
rect 584 1832 600 1848
rect 2936 1832 2952 1848
rect 3208 1832 3224 1848
rect 4440 1832 4456 1848
rect 5128 1832 5144 1848
rect 536 1812 552 1828
rect 760 1812 776 1828
rect 808 1812 824 1828
rect 88 1792 104 1808
rect 456 1792 472 1808
rect 584 1792 600 1808
rect 1736 1792 1752 1808
rect 1934 1802 1962 1818
rect 2248 1792 2264 1808
rect 3064 1792 3080 1808
rect 3096 1792 3128 1808
rect 3982 1802 4010 1818
rect 4824 1812 4840 1828
rect 5144 1792 5160 1808
rect 5560 1792 5576 1808
rect 5640 1792 5656 1808
rect 5816 1792 5832 1808
rect 8 1752 24 1768
rect 104 1752 120 1768
rect 200 1752 216 1768
rect 1144 1772 1160 1788
rect 2088 1772 2104 1788
rect 2536 1772 2552 1788
rect 2760 1772 2776 1788
rect 3016 1772 3032 1788
rect 3368 1772 3384 1788
rect 4168 1772 4184 1788
rect 4328 1772 4344 1788
rect 5528 1772 5544 1788
rect 5704 1772 5720 1788
rect 1000 1752 1016 1768
rect 1128 1752 1144 1768
rect 1544 1752 1560 1768
rect 3208 1752 3224 1768
rect 3976 1752 3992 1768
rect 4568 1752 4584 1768
rect 4632 1752 4648 1768
rect 4712 1752 4728 1768
rect 344 1732 360 1748
rect 712 1732 728 1748
rect 952 1732 968 1748
rect 1256 1732 1272 1748
rect 2248 1732 2264 1748
rect 2440 1732 2456 1748
rect 2872 1732 2888 1748
rect 776 1712 792 1728
rect 888 1712 904 1728
rect 1768 1712 1784 1728
rect 2200 1712 2216 1728
rect 2376 1712 2392 1728
rect 3256 1732 3272 1748
rect 3816 1732 3832 1748
rect 4120 1732 4152 1748
rect 5624 1732 5640 1748
rect 4152 1712 4168 1728
rect 424 1692 440 1708
rect 1160 1692 1192 1708
rect 1352 1692 1368 1708
rect 2088 1692 2104 1708
rect 2568 1692 2584 1708
rect 2600 1692 2616 1708
rect 2680 1692 2696 1708
rect 3624 1692 3640 1708
rect 5816 1692 5832 1708
rect 5960 1692 5976 1708
rect 808 1672 824 1688
rect 2392 1672 2408 1688
rect 3768 1672 3784 1688
rect 1352 1652 1368 1668
rect 1672 1652 1688 1668
rect 2568 1652 2584 1668
rect 3912 1652 3928 1668
rect 5432 1652 5448 1668
rect 1272 1632 1288 1648
rect 2360 1632 2376 1648
rect 5384 1632 5400 1648
rect 5464 1632 5480 1648
rect 8 1612 24 1628
rect 760 1612 776 1628
rect 200 1592 216 1608
rect 926 1602 954 1618
rect 1784 1592 1800 1608
rect 2568 1592 2584 1608
rect 2744 1592 2760 1608
rect 2974 1602 3002 1618
rect 3272 1612 3288 1628
rect 3048 1592 3064 1608
rect 5022 1602 5050 1618
rect 5544 1612 5560 1628
rect 1096 1572 1112 1588
rect 2248 1572 2264 1588
rect 2712 1572 2728 1588
rect 3288 1572 3304 1588
rect 4088 1572 4120 1588
rect 5288 1572 5304 1588
rect 2152 1552 2168 1568
rect 2328 1552 2344 1568
rect 3736 1552 3752 1568
rect 4040 1552 4056 1568
rect 504 1532 520 1548
rect 1000 1532 1016 1548
rect 1096 1532 1112 1548
rect 1176 1532 1192 1548
rect 1544 1532 1560 1548
rect 1656 1532 1672 1548
rect 2456 1532 2472 1548
rect 2920 1532 2936 1548
rect 3192 1532 3208 1548
rect 4072 1532 4088 1548
rect 4472 1532 4488 1548
rect 760 1512 776 1528
rect 2280 1512 2296 1528
rect 2328 1512 2344 1528
rect 3096 1512 3112 1528
rect 3176 1512 3192 1528
rect 3704 1512 3720 1528
rect 4168 1512 4184 1528
rect 5784 1512 5800 1528
rect 1288 1492 1304 1508
rect 1448 1492 1464 1508
rect 2312 1492 2328 1508
rect 2344 1492 2360 1508
rect 2648 1492 2664 1508
rect 3544 1492 3560 1508
rect 5160 1492 5176 1508
rect 5816 1492 5832 1508
rect 5928 1492 5944 1508
rect 488 1472 504 1488
rect 664 1472 680 1488
rect 1416 1472 1432 1488
rect 2664 1472 2680 1488
rect 3208 1472 3224 1488
rect 3864 1472 3880 1488
rect 4216 1472 4232 1488
rect 4648 1472 4664 1488
rect 472 1452 488 1468
rect 872 1452 888 1468
rect 2216 1452 2232 1468
rect 3048 1452 3064 1468
rect 3144 1452 3160 1468
rect 3432 1452 3448 1468
rect 3544 1452 3560 1468
rect 3944 1452 3976 1468
rect 4328 1452 4344 1468
rect 4440 1452 4456 1468
rect 4568 1452 4584 1468
rect 5688 1452 5704 1468
rect 5896 1452 5912 1468
rect 1112 1432 1128 1448
rect 1848 1432 1864 1448
rect 2744 1432 2760 1448
rect 4856 1432 4872 1448
rect 5416 1432 5432 1448
rect 5960 1432 5976 1448
rect 1934 1402 1962 1418
rect 3864 1412 3880 1428
rect 3880 1412 3896 1428
rect 2408 1392 2424 1408
rect 3400 1392 3416 1408
rect 3448 1392 3464 1408
rect 3982 1402 4010 1418
rect 5736 1412 5752 1428
rect 4616 1392 4632 1408
rect 5288 1392 5304 1408
rect 1224 1372 1240 1388
rect 2504 1372 2520 1388
rect 2584 1372 2600 1388
rect 4088 1372 4104 1388
rect 5176 1372 5192 1388
rect 5336 1372 5352 1388
rect 5528 1372 5544 1388
rect 456 1352 472 1368
rect 2200 1352 2216 1368
rect 2392 1352 2408 1368
rect 3000 1352 3016 1368
rect 3592 1352 3608 1368
rect 3848 1352 3864 1368
rect 4072 1352 4088 1368
rect 4200 1352 4216 1368
rect 584 1332 600 1348
rect 680 1332 696 1348
rect 1208 1332 1224 1348
rect 1144 1312 1160 1328
rect 1480 1312 1496 1328
rect 1608 1312 1624 1328
rect 1912 1332 1928 1348
rect 1944 1332 1960 1348
rect 2424 1332 2440 1348
rect 2456 1332 2472 1348
rect 2776 1332 2792 1348
rect 3032 1332 3048 1348
rect 3080 1332 3096 1348
rect 3528 1332 3544 1348
rect 3784 1332 3800 1348
rect 3912 1332 3928 1348
rect 4440 1332 4456 1348
rect 4504 1332 4520 1348
rect 5336 1332 5352 1348
rect 5496 1332 5512 1348
rect 1896 1312 1912 1328
rect 2312 1312 2328 1328
rect 3144 1312 3160 1328
rect 3736 1312 3752 1328
rect 3784 1312 3800 1328
rect 4776 1312 4792 1328
rect 4984 1312 5000 1328
rect 5176 1312 5192 1328
rect 5272 1312 5288 1328
rect 5416 1312 5432 1328
rect 5448 1312 5464 1328
rect 5768 1312 5784 1328
rect 1704 1292 1720 1308
rect 2376 1292 2392 1308
rect 2408 1292 2424 1308
rect 2888 1292 2904 1308
rect 3336 1292 3352 1308
rect 3432 1292 3448 1308
rect 3640 1292 3656 1308
rect 4104 1292 4120 1308
rect 4280 1292 4296 1308
rect 4376 1292 4392 1308
rect 4696 1292 4712 1308
rect 5880 1292 5896 1308
rect 1880 1272 1896 1288
rect 2792 1272 2808 1288
rect 3288 1272 3304 1288
rect 3800 1272 3816 1288
rect 600 1252 616 1268
rect 2360 1252 2376 1268
rect 2600 1252 2616 1268
rect 2856 1252 2872 1268
rect 5128 1252 5144 1268
rect 5640 1252 5656 1268
rect 5848 1252 5880 1268
rect 3240 1232 3256 1248
rect 4040 1232 4056 1248
rect 5224 1232 5240 1248
rect 5576 1232 5592 1248
rect 5800 1232 5816 1248
rect 926 1202 954 1218
rect 1240 1192 1256 1208
rect 2974 1202 3002 1218
rect 3176 1212 3192 1228
rect 4632 1192 4648 1208
rect 5022 1202 5050 1218
rect 5512 1212 5528 1228
rect 5528 1192 5544 1208
rect 2280 1172 2296 1188
rect 4552 1172 4568 1188
rect 616 1152 632 1168
rect 2072 1152 2088 1168
rect 2648 1152 2664 1168
rect 4472 1152 4488 1168
rect 4856 1152 4872 1168
rect 5160 1152 5176 1168
rect 2232 1132 2248 1148
rect 3064 1132 3080 1148
rect 4328 1132 4344 1148
rect 1672 1112 1688 1128
rect 3016 1112 3032 1128
rect 3528 1112 3544 1128
rect 3704 1112 3720 1128
rect 4472 1112 4488 1128
rect 1272 1092 1288 1108
rect 1336 1092 1352 1108
rect 1992 1092 2008 1108
rect 2104 1092 2120 1108
rect 3176 1092 3192 1108
rect 3560 1092 3576 1108
rect 3624 1092 3640 1108
rect 3672 1092 3688 1108
rect 3768 1092 3784 1108
rect 984 1072 1000 1088
rect 1128 1072 1144 1088
rect 1736 1072 1752 1088
rect 2520 1072 2536 1088
rect 3544 1072 3560 1088
rect 3576 1072 3592 1088
rect 3960 1072 3976 1088
rect 4504 1072 4520 1088
rect 5224 1072 5240 1088
rect 5432 1072 5448 1088
rect 5832 1072 5848 1088
rect 5864 1072 5880 1088
rect 1336 1052 1352 1068
rect 2200 1052 2216 1068
rect 2216 1052 2232 1068
rect 3160 1052 3176 1068
rect 3208 1052 3224 1068
rect 3768 1052 3784 1068
rect 4248 1052 4264 1068
rect 5208 1052 5224 1068
rect 5384 1052 5400 1068
rect 808 1032 824 1048
rect 872 1032 888 1048
rect 2248 1032 2264 1048
rect 3304 1032 3320 1048
rect 1934 1002 1962 1018
rect 2584 992 2600 1008
rect 3096 992 3112 1008
rect 3512 992 3528 1008
rect 3982 1002 4010 1018
rect 4456 1012 4472 1028
rect 968 972 984 988
rect 2472 972 2488 988
rect 1272 952 1288 968
rect 2264 952 2280 968
rect 2328 952 2344 968
rect 4200 972 4216 988
rect 4216 972 4232 988
rect 4456 972 4488 988
rect 3480 952 3496 968
rect 600 932 616 948
rect 1256 932 1272 948
rect 1288 932 1320 948
rect 1864 932 1880 948
rect 1976 932 1992 948
rect 2088 932 2104 948
rect 2296 932 2312 948
rect 5688 932 5704 948
rect 2376 912 2392 928
rect 2632 912 2648 928
rect 5592 912 5608 928
rect 1176 892 1192 908
rect 5416 892 5432 908
rect 216 872 232 888
rect 1560 872 1576 888
rect 1720 872 1736 888
rect 3208 872 3224 888
rect 2904 852 2920 868
rect 4840 852 4856 868
rect 926 802 954 818
rect 1352 812 1368 828
rect 2974 802 3002 818
rect 3640 792 3656 808
rect 5022 802 5050 818
rect 2200 772 2216 788
rect 4056 772 4072 788
rect 4504 772 4520 788
rect 4552 772 4568 788
rect 1224 752 1240 768
rect 3544 752 3560 768
rect 4936 752 4952 768
rect 1256 732 1272 748
rect 1656 732 1672 748
rect 1912 732 1928 748
rect 2376 732 2392 748
rect 2424 732 2440 748
rect 3112 732 3128 748
rect 5656 732 5672 748
rect 1000 712 1016 728
rect 2088 712 2104 728
rect 3928 712 3944 728
rect 4936 712 4952 728
rect 1032 692 1048 708
rect 1544 692 1560 708
rect 1736 692 1752 708
rect 2136 692 2152 708
rect 2440 692 2456 708
rect 2520 692 2536 708
rect 984 672 1000 688
rect 2728 692 2744 708
rect 2760 692 2776 708
rect 2824 692 2840 708
rect 3448 692 3464 708
rect 3624 692 3640 708
rect 3880 692 3896 708
rect 4280 692 4296 708
rect 5640 692 5656 708
rect 2520 672 2536 688
rect 2568 672 2584 688
rect 5912 672 5928 688
rect 3656 652 3672 668
rect 1032 632 1048 648
rect 1976 632 1992 648
rect 472 612 488 628
rect 1736 592 1752 608
rect 1934 602 1962 618
rect 1992 612 2008 628
rect 3832 632 3848 648
rect 504 572 520 588
rect 1880 572 1896 588
rect 2424 592 2440 608
rect 2584 592 2600 608
rect 3400 592 3416 608
rect 3982 602 4010 618
rect 5704 592 5720 608
rect 3304 572 3320 588
rect 728 552 744 568
rect 872 552 888 568
rect 1272 552 1288 568
rect 1880 552 1896 568
rect 2072 552 2088 568
rect 3320 552 3336 568
rect 3512 552 3528 568
rect 3560 552 3576 568
rect 3816 552 3832 568
rect 4152 552 4168 568
rect 648 532 664 548
rect 1416 532 1432 548
rect 1688 532 1704 548
rect 1880 532 1896 548
rect 1976 532 1992 548
rect 2200 532 2216 548
rect 3368 532 3384 548
rect 3768 532 3784 548
rect 5144 552 5160 568
rect 5912 552 5928 568
rect 5400 532 5416 548
rect 5576 532 5592 548
rect 5736 532 5752 548
rect 616 512 632 528
rect 808 512 824 528
rect 2392 512 2408 528
rect 2952 512 2968 528
rect 3144 512 3160 528
rect 3656 512 3672 528
rect 5064 512 5080 528
rect 5352 512 5368 528
rect 1560 492 1576 508
rect 1752 492 1768 508
rect 2344 492 2360 508
rect 2488 492 2504 508
rect 3240 492 3256 508
rect 3640 492 3656 508
rect 1736 452 1752 468
rect 4552 452 4568 468
rect 2248 432 2264 448
rect 2680 432 2696 448
rect 3528 432 3544 448
rect 926 402 954 418
rect 1656 392 1672 408
rect 2974 402 3002 418
rect 5022 402 5050 418
rect 5464 412 5480 428
rect 5624 372 5640 388
rect 2680 352 2696 368
rect 5960 352 5976 368
rect 3352 332 3368 348
rect 3832 332 3848 348
rect 4776 312 4792 328
rect 5144 312 5160 328
rect 5720 312 5736 328
rect 1000 292 1016 308
rect 1704 292 1720 308
rect 2120 292 2136 308
rect 2856 292 2872 308
rect 3896 292 3912 308
rect 5608 292 5624 308
rect 1000 272 1016 288
rect 3384 272 3400 288
rect 3400 272 3416 288
rect 4392 272 4408 288
rect 600 252 616 268
rect 2088 252 2104 268
rect 4216 252 4232 268
rect 5448 272 5464 288
rect 5320 232 5336 248
rect 1934 202 1962 218
rect 1976 212 1992 228
rect 3982 202 4010 218
rect 4904 212 4920 228
rect 5448 212 5464 228
rect 3912 172 3928 188
rect 4632 172 4648 188
rect 1976 152 1992 168
rect 3528 152 3544 168
rect 5752 132 5768 148
rect 5944 132 5960 148
rect 3912 112 3928 128
rect 5784 112 5800 128
rect 1720 32 1736 48
rect 1896 32 1912 48
rect 3672 32 3688 48
rect 926 2 954 18
rect 1176 12 1192 28
rect 1256 12 1272 28
rect 1704 12 1720 28
rect 1912 12 1928 28
rect 2088 12 2104 28
rect 2248 12 2264 28
rect 2376 12 2392 28
rect 2424 12 2440 28
rect 2974 2 3002 18
rect 3112 12 3128 28
rect 3208 12 3224 28
rect 3800 12 3816 28
rect 5022 2 5050 18
<< metal4 >>
rect 652 3976 660 3984
rect 29 3748 35 3772
rect 61 3388 67 3492
rect 189 2948 195 3232
rect 77 2668 83 2692
rect 93 1764 99 1792
rect 205 1768 211 3912
rect 653 3908 659 3976
rect 364 3896 372 3904
rect 316 3883 324 3884
rect 316 3877 328 3883
rect 316 3876 324 3877
rect 365 2168 371 3896
rect 381 2248 387 2432
rect 397 2148 403 3872
rect 461 2688 467 3232
rect 92 1763 100 1764
rect 92 1757 104 1763
rect 92 1756 100 1757
rect 13 1628 19 1752
rect 205 1608 211 1752
rect 221 888 227 2092
rect 477 1908 483 3512
rect 637 2968 643 3092
rect 589 2308 595 2612
rect 604 2303 612 2304
rect 604 2297 616 2303
rect 604 2296 612 2297
rect 461 1368 467 1792
rect 477 1468 483 1852
rect 493 1488 499 2172
rect 525 1784 531 1832
rect 524 1776 532 1784
rect 541 1724 547 1812
rect 589 1808 595 1832
rect 540 1716 548 1724
rect 477 628 483 1452
rect 509 588 515 1532
rect 572 1343 580 1344
rect 572 1337 584 1343
rect 572 1336 580 1337
rect 605 1268 611 2032
rect 605 268 611 932
rect 621 528 627 1152
rect 653 548 659 3892
rect 701 2928 707 3012
rect 668 1496 676 1504
rect 669 1488 675 1496
rect 685 1348 691 2212
rect 701 2128 707 2272
rect 717 1748 723 3972
rect 797 3944 803 4012
rect 954 4006 960 4014
rect 972 3956 980 3964
rect 796 3936 804 3944
rect 973 3928 979 3956
rect 1196 3903 1204 3904
rect 1192 3897 1204 3903
rect 1196 3896 1204 3897
rect 924 3876 932 3884
rect 925 3848 931 3876
rect 861 3724 867 3732
rect 860 3716 868 3724
rect 733 3348 739 3632
rect 877 3628 883 3692
rect 941 3644 947 3892
rect 1084 3876 1092 3884
rect 1036 3723 1044 3724
rect 1036 3717 1048 3723
rect 1036 3716 1044 3717
rect 1085 3708 1091 3876
rect 1213 3788 1219 3932
rect 1117 3664 1123 3672
rect 1116 3656 1124 3664
rect 940 3636 948 3644
rect 765 2468 771 2832
rect 845 2828 851 3252
rect 797 2288 803 2432
rect 813 2368 819 2632
rect 797 2143 803 2272
rect 813 2228 819 2352
rect 797 2137 808 2143
rect 765 1828 771 1892
rect 781 1888 787 2132
rect 780 1736 788 1744
rect 781 1728 787 1736
rect 813 1688 819 1812
rect 765 1528 771 1612
rect 877 1468 883 3612
rect 954 3606 960 3614
rect 954 3206 960 3214
rect 1101 2948 1107 3092
rect 954 2806 960 2814
rect 954 2406 960 2414
rect 989 2308 995 2852
rect 892 2296 900 2304
rect 893 2268 899 2296
rect 954 2006 960 2014
rect 940 1743 948 1744
rect 940 1737 952 1743
rect 940 1736 948 1737
rect 908 1723 916 1724
rect 904 1717 916 1723
rect 908 1716 916 1717
rect 954 1606 960 1614
rect 954 1206 960 1214
rect 813 528 819 1032
rect 877 568 883 1032
rect 973 988 979 2092
rect 1005 1548 1011 1752
rect 954 806 960 814
rect 989 688 995 1072
rect 1021 944 1027 2212
rect 1101 1548 1107 1572
rect 1117 1448 1123 3656
rect 1133 3128 1139 3432
rect 1293 3408 1299 3812
rect 1309 3544 1315 3612
rect 1308 3536 1316 3544
rect 1244 3083 1252 3084
rect 1240 3077 1252 3083
rect 1244 3076 1252 3077
rect 1180 2143 1188 2144
rect 1180 2137 1192 2143
rect 1180 2136 1188 2137
rect 1133 1088 1139 1752
rect 1149 1328 1155 1772
rect 1196 1703 1204 1704
rect 1192 1697 1204 1703
rect 1196 1696 1204 1697
rect 1165 1604 1171 1692
rect 1164 1596 1172 1604
rect 1181 1504 1187 1532
rect 1180 1496 1188 1504
rect 1213 1304 1219 1332
rect 1212 1296 1220 1304
rect 1020 936 1028 944
rect 954 406 960 414
rect 1005 308 1011 712
rect 1037 648 1043 692
rect 988 283 996 284
rect 988 277 1000 283
rect 988 276 996 277
rect 1181 28 1187 892
rect 1229 768 1235 1372
rect 1245 1208 1251 2372
rect 1277 1108 1283 1632
rect 1293 1508 1299 1852
rect 1260 956 1268 964
rect 1261 948 1267 956
rect 1261 28 1267 732
rect 1277 568 1283 952
rect 1309 948 1315 3536
rect 1357 1708 1363 3952
rect 2029 3948 2035 3972
rect 2300 3916 2308 3924
rect 2301 3888 2307 3916
rect 2556 3896 2564 3904
rect 2557 3888 2563 3896
rect 1629 3864 1635 3872
rect 1628 3856 1636 3864
rect 1962 3806 1968 3814
rect 1932 3776 1940 3784
rect 1564 3736 1572 3744
rect 1565 3728 1571 3736
rect 1901 3704 1907 3712
rect 1933 3708 1939 3776
rect 1964 3743 1972 3744
rect 1960 3737 1972 3743
rect 1964 3736 1972 3737
rect 2172 3736 2180 3744
rect 2173 3728 2179 3736
rect 1900 3696 1908 3704
rect 1661 3384 1667 3452
rect 1660 3376 1668 3384
rect 1388 3343 1396 3344
rect 1388 3337 1400 3343
rect 1388 3336 1396 3337
rect 1501 2928 1507 3332
rect 1437 2684 1443 2692
rect 1436 2676 1444 2684
rect 1565 2544 1571 2572
rect 1564 2536 1572 2544
rect 1500 2303 1508 2304
rect 1500 2297 1512 2303
rect 1500 2296 1508 2297
rect 1516 2163 1524 2164
rect 1516 2157 1528 2163
rect 1516 2156 1524 2157
rect 1341 1068 1347 1092
rect 1357 828 1363 1652
rect 1453 1508 1459 2032
rect 1549 1548 1555 1752
rect 1661 1548 1667 2092
rect 1500 1323 1508 1324
rect 1496 1317 1508 1323
rect 1500 1316 1508 1317
rect 1596 1323 1604 1324
rect 1596 1317 1608 1323
rect 1596 1316 1604 1317
rect 1677 1128 1683 1652
rect 1549 644 1555 692
rect 1548 636 1556 644
rect 1421 524 1427 532
rect 1420 516 1428 524
rect 1565 508 1571 872
rect 1661 408 1667 732
rect 1693 548 1699 3292
rect 1821 2284 1827 2292
rect 1820 2276 1828 2284
rect 1836 2156 1844 2164
rect 1837 2148 1843 2156
rect 1708 1956 1716 1964
rect 1709 1948 1715 1956
rect 1741 1864 1747 1892
rect 1740 1856 1748 1864
rect 1709 308 1715 1292
rect 1741 1088 1747 1792
rect 1772 1776 1780 1784
rect 1773 1728 1779 1776
rect 1789 1584 1795 1592
rect 1788 1576 1796 1584
rect 1853 1448 1859 3632
rect 1962 3406 1968 3414
rect 2205 3388 2211 3572
rect 2253 3564 2259 3872
rect 2397 3844 2403 3872
rect 2717 3864 2723 3872
rect 2716 3856 2724 3864
rect 2396 3836 2404 3844
rect 2364 3796 2372 3804
rect 2284 3756 2292 3764
rect 2285 3708 2291 3756
rect 2268 3703 2276 3704
rect 2268 3697 2280 3703
rect 2268 3696 2276 3697
rect 2252 3556 2260 3564
rect 2237 3448 2243 3492
rect 2124 3383 2132 3384
rect 2120 3377 2132 3383
rect 2124 3376 2132 3377
rect 1917 3028 1923 3232
rect 1962 3006 1968 3014
rect 1901 2548 1907 2732
rect 2077 2728 2083 2992
rect 1962 2606 1968 2614
rect 2044 2556 2052 2564
rect 1996 2543 2004 2544
rect 1992 2537 2004 2543
rect 1996 2536 2004 2537
rect 2045 2528 2051 2556
rect 2076 2536 2084 2544
rect 2077 2503 2083 2536
rect 2072 2497 2083 2503
rect 2077 2288 2083 2372
rect 1962 2206 1968 2214
rect 1901 2164 1907 2172
rect 1900 2156 1908 2164
rect 1917 1348 1923 1952
rect 2029 1924 2035 1932
rect 2028 1916 2036 1924
rect 1964 1863 1972 1864
rect 1960 1857 1972 1863
rect 1964 1856 1972 1857
rect 1962 1806 1968 1814
rect 1962 1406 1968 1414
rect 1885 1264 1891 1272
rect 1884 1256 1892 1264
rect 1884 943 1892 944
rect 1880 937 1892 943
rect 1884 936 1892 937
rect 1709 28 1715 292
rect 1725 48 1731 872
rect 1741 608 1747 692
rect 1868 543 1876 544
rect 1868 537 1880 543
rect 1868 536 1876 537
rect 1757 463 1763 492
rect 1752 457 1763 463
rect 1901 48 1907 1312
rect 2077 1168 2083 2232
rect 2093 1788 2099 2352
rect 2109 2168 2115 2632
rect 2108 1116 2116 1124
rect 2109 1108 2115 1116
rect 1962 1006 1968 1014
rect 1917 28 1923 732
rect 1962 606 1968 614
rect 1981 548 1987 632
rect 1997 628 2003 1092
rect 2093 728 2099 932
rect 2076 576 2084 584
rect 2077 568 2083 576
rect 2125 308 2131 2192
rect 2141 1968 2147 2412
rect 2173 2228 2179 2612
rect 2220 2543 2228 2544
rect 2216 2537 2228 2543
rect 2220 2536 2228 2537
rect 2189 2224 2195 2232
rect 2188 2216 2196 2224
rect 2157 1568 2163 2132
rect 2204 2096 2212 2104
rect 2205 2068 2211 2096
rect 2220 2056 2228 2064
rect 2221 1908 2227 2056
rect 2220 1723 2228 1724
rect 2216 1717 2228 1723
rect 2220 1716 2228 1717
rect 2221 1068 2227 1452
rect 2237 1148 2243 1892
rect 2253 1808 2259 1992
rect 2253 1748 2259 1792
rect 2253 964 2259 1032
rect 2269 968 2275 3312
rect 2285 1188 2291 1512
rect 2252 956 2260 964
rect 2301 948 2307 3712
rect 2317 2548 2323 2792
rect 2332 2283 2340 2284
rect 2328 2277 2340 2283
rect 2332 2276 2340 2277
rect 2349 1764 2355 3332
rect 2365 3088 2371 3796
rect 2684 3776 2692 3784
rect 2685 3768 2691 3776
rect 2445 3584 2451 3732
rect 2460 3723 2468 3724
rect 2460 3717 2472 3723
rect 2460 3716 2468 3717
rect 2749 3708 2755 4012
rect 2781 3764 2787 3772
rect 2780 3756 2788 3764
rect 2652 3703 2660 3704
rect 2652 3697 2664 3703
rect 2652 3696 2660 3697
rect 2444 3576 2452 3584
rect 2396 3436 2404 3444
rect 2397 3128 2403 3436
rect 2460 2563 2468 2564
rect 2456 2557 2468 2563
rect 2460 2556 2468 2557
rect 2412 2543 2420 2544
rect 2412 2537 2424 2543
rect 2412 2536 2420 2537
rect 2444 2243 2452 2244
rect 2444 2237 2456 2243
rect 2444 2236 2452 2237
rect 2348 1756 2356 1764
rect 2333 1528 2339 1552
rect 2316 1516 2324 1524
rect 2317 1508 2323 1516
rect 2349 1508 2355 1756
rect 2381 1744 2387 2232
rect 2397 2164 2403 2172
rect 2396 2156 2404 2164
rect 2380 1736 2388 1744
rect 2316 1336 2324 1344
rect 2317 1328 2323 1336
rect 2365 1268 2371 1632
rect 2381 1308 2387 1712
rect 2397 1688 2403 1912
rect 2397 1368 2403 1672
rect 2413 1308 2419 1392
rect 2429 1348 2435 2192
rect 2445 1844 2451 2012
rect 2444 1836 2452 1844
rect 2332 976 2340 984
rect 2333 968 2339 976
rect 2381 928 2387 1292
rect 2205 548 2211 772
rect 2348 516 2356 524
rect 2349 508 2355 516
rect 1962 206 1968 214
rect 1981 168 1987 212
rect 2093 28 2099 252
rect 2253 28 2259 432
rect 2381 28 2387 732
rect 2429 608 2435 732
rect 2445 708 2451 1732
rect 2461 1348 2467 1532
rect 2477 988 2483 3532
rect 2525 3348 2531 3512
rect 2540 3403 2548 3404
rect 2540 3397 2552 3403
rect 2540 3396 2548 3397
rect 2573 3384 2579 3432
rect 2572 3376 2580 3384
rect 2572 3303 2580 3304
rect 2572 3297 2584 3303
rect 2572 3296 2580 3297
rect 2621 3288 2627 3552
rect 2716 3516 2724 3524
rect 2717 3508 2723 3516
rect 2684 3416 2692 3424
rect 2685 3408 2691 3416
rect 2813 3344 2819 3872
rect 2892 3736 2900 3744
rect 2893 3684 2899 3736
rect 2892 3683 2900 3684
rect 2892 3677 2904 3683
rect 2892 3676 2900 3677
rect 2877 3528 2883 3592
rect 2812 3336 2820 3344
rect 2925 3228 2931 4012
rect 3002 4006 3008 4014
rect 2940 3736 2948 3744
rect 2941 3728 2947 3736
rect 3133 3624 3139 3632
rect 3132 3616 3140 3624
rect 3002 3606 3008 3614
rect 2972 3483 2980 3484
rect 2972 3477 2984 3483
rect 2972 3476 2980 3477
rect 3132 3443 3140 3444
rect 3128 3437 3140 3443
rect 3132 3436 3140 3437
rect 3068 3396 3076 3404
rect 3002 3206 3008 3214
rect 3021 3088 3027 3312
rect 2493 2128 2499 2972
rect 2637 2948 2643 2972
rect 2525 2568 2531 2712
rect 2556 2283 2564 2284
rect 2556 2277 2568 2283
rect 2556 2276 2564 2277
rect 2653 2108 2659 2172
rect 2636 2103 2644 2104
rect 2632 2097 2644 2103
rect 2636 2096 2644 2097
rect 2509 1388 2515 2092
rect 2636 2036 2644 2044
rect 2541 1384 2547 1772
rect 2573 1668 2579 1692
rect 2556 1603 2564 1604
rect 2556 1597 2568 1603
rect 2556 1596 2564 1597
rect 2589 1388 2595 1932
rect 2540 1376 2548 1384
rect 2605 1268 2611 1692
rect 2508 1083 2516 1084
rect 2508 1077 2520 1083
rect 2508 1076 2516 1077
rect 2572 736 2580 744
rect 2540 703 2548 704
rect 2536 697 2548 703
rect 2540 696 2548 697
rect 2573 688 2579 736
rect 2508 683 2516 684
rect 2508 677 2520 683
rect 2508 676 2516 677
rect 2589 608 2595 992
rect 2637 928 2643 2036
rect 2669 1908 2675 2972
rect 2828 2956 2836 2964
rect 2829 2948 2835 2956
rect 2717 2148 2723 2672
rect 2749 2524 2755 2532
rect 2748 2516 2756 2524
rect 2652 1896 2660 1904
rect 2653 1888 2659 1896
rect 2701 1888 2707 1932
rect 2653 1168 2659 1492
rect 2669 1488 2675 1872
rect 2701 1868 2707 1872
rect 2684 1716 2692 1724
rect 2685 1708 2691 1716
rect 2717 1588 2723 1952
rect 2733 708 2739 2172
rect 2749 1448 2755 1592
rect 2765 708 2771 1772
rect 2781 1404 2787 2332
rect 2797 2168 2803 2192
rect 2813 2168 2819 2412
rect 2877 2148 2883 3032
rect 2924 2943 2932 2944
rect 2920 2937 2932 2943
rect 2924 2936 2932 2937
rect 2909 2568 2915 2592
rect 2908 2216 2916 2224
rect 2909 2208 2915 2216
rect 2797 1924 2803 1932
rect 2796 1916 2804 1924
rect 2796 1836 2804 1844
rect 2780 1396 2788 1404
rect 2781 1348 2787 1396
rect 2797 1288 2803 1836
rect 2861 1268 2867 1872
rect 2877 1748 2883 2012
rect 2893 1308 2899 2092
rect 2909 868 2915 2172
rect 2925 1548 2931 1892
rect 2941 1848 2947 3032
rect 3037 2964 3043 3072
rect 3036 2956 3044 2964
rect 2957 2368 2963 2852
rect 3002 2806 3008 2814
rect 3037 2648 3043 2812
rect 3053 2544 3059 2632
rect 3052 2536 3060 2544
rect 3002 2406 3008 2414
rect 3002 2006 3008 2014
rect 3053 1888 3059 2432
rect 3020 1796 3028 1804
rect 3021 1788 3027 1796
rect 3002 1606 3008 1614
rect 3053 1608 3059 1852
rect 3069 1808 3075 3396
rect 3181 3368 3187 3392
rect 3181 2988 3187 3352
rect 3197 2928 3203 3932
rect 3308 3896 3316 3904
rect 3309 3808 3315 3896
rect 3212 3803 3220 3804
rect 3212 3797 3224 3803
rect 3212 3796 3220 3797
rect 3325 3728 3331 4012
rect 3261 3148 3267 3712
rect 3309 3484 3315 3712
rect 3308 3476 3316 3484
rect 3309 3324 3315 3476
rect 3341 3468 3347 3932
rect 3453 3728 3459 3812
rect 3388 3596 3396 3604
rect 3372 3363 3380 3364
rect 3368 3357 3380 3363
rect 3372 3356 3380 3357
rect 3308 3316 3316 3324
rect 3373 2928 3379 3312
rect 3389 3088 3395 3596
rect 3117 1808 3123 2472
rect 3149 1888 3155 2272
rect 3084 1803 3092 1804
rect 3084 1797 3096 1803
rect 3084 1796 3092 1797
rect 3084 1376 3092 1384
rect 3085 1348 3091 1376
rect 3037 1324 3043 1332
rect 3036 1316 3044 1324
rect 3020 1256 3028 1264
rect 3002 1206 3008 1214
rect 3021 1128 3027 1256
rect 3069 1084 3075 1132
rect 3068 1076 3076 1084
rect 3101 1008 3107 1512
rect 3149 1468 3155 1872
rect 3197 1548 3203 2112
rect 3213 1848 3219 2612
rect 3229 2548 3235 2752
rect 3245 2688 3251 2832
rect 3245 2468 3251 2552
rect 3228 2316 3236 2324
rect 3229 2308 3235 2316
rect 3212 1776 3220 1784
rect 3213 1768 3219 1776
rect 3260 1756 3268 1764
rect 3261 1748 3267 1756
rect 3277 1628 3283 1952
rect 3149 1328 3155 1452
rect 3181 1228 3187 1512
rect 3213 1464 3219 1472
rect 3212 1456 3220 1464
rect 3164 1103 3172 1104
rect 3164 1097 3176 1103
rect 3164 1096 3172 1097
rect 3164 1076 3172 1084
rect 3165 1068 3171 1076
rect 3213 1068 3219 1456
rect 3293 1288 3299 1572
rect 3002 806 3008 814
rect 2396 536 2404 544
rect 2397 528 2403 536
rect 2429 28 2435 592
rect 2956 536 2964 544
rect 2957 528 2963 536
rect 2685 368 2691 432
rect 3002 406 3008 414
rect 2861 284 2867 292
rect 2860 276 2868 284
rect 3117 28 3123 732
rect 3148 636 3156 644
rect 3149 528 3155 636
rect 3213 28 3219 872
rect 3245 508 3251 1232
rect 3309 588 3315 1032
rect 3325 568 3331 2512
rect 3341 1308 3347 1852
rect 3357 348 3363 2712
rect 3373 2128 3379 2912
rect 3405 2548 3411 3692
rect 3421 2728 3427 3632
rect 3436 3556 3444 3564
rect 3437 3508 3443 3556
rect 3373 548 3379 1772
rect 3405 1408 3411 2532
rect 3437 2528 3443 3492
rect 3453 2468 3459 3712
rect 3469 2188 3475 3712
rect 3500 3576 3508 3584
rect 3501 3528 3507 3576
rect 3484 3436 3492 3444
rect 3485 3128 3491 3436
rect 3517 3428 3523 3712
rect 3533 3488 3539 3752
rect 3565 3524 3571 3632
rect 3581 3628 3587 4012
rect 3645 3924 3651 4012
rect 3644 3916 3652 3924
rect 3725 3908 3731 3992
rect 4045 3984 4051 4012
rect 4044 3976 4052 3984
rect 4173 3964 4179 4012
rect 5050 4006 5056 4014
rect 4172 3956 4180 3964
rect 4269 3944 4275 3972
rect 4268 3943 4276 3944
rect 4264 3937 4276 3943
rect 4268 3936 4276 3937
rect 4444 3903 4452 3904
rect 4444 3897 4456 3903
rect 4444 3896 4452 3897
rect 4524 3896 4532 3904
rect 3613 3744 3619 3892
rect 3725 3884 3731 3892
rect 3724 3876 3732 3884
rect 3612 3736 3620 3744
rect 3564 3516 3572 3524
rect 3500 3416 3508 3424
rect 3437 1308 3443 1452
rect 3485 968 3491 2092
rect 3501 1908 3507 3416
rect 3564 3423 3572 3424
rect 3560 3417 3572 3423
rect 3564 3416 3572 3417
rect 3533 3404 3539 3412
rect 3532 3396 3540 3404
rect 3548 3336 3556 3344
rect 3549 3328 3555 3336
rect 3560 3317 3571 3323
rect 3532 3043 3540 3044
rect 3532 3037 3544 3043
rect 3532 3036 3540 3037
rect 3533 2908 3539 2992
rect 3533 2284 3539 2812
rect 3549 2408 3555 2952
rect 3565 2724 3571 3317
rect 3597 2948 3603 3672
rect 3613 3108 3619 3736
rect 3629 3644 3635 3652
rect 3628 3636 3636 3644
rect 3661 3544 3667 3872
rect 4156 3823 4164 3824
rect 4156 3817 4168 3823
rect 4156 3816 4164 3817
rect 4010 3806 4016 3814
rect 3660 3536 3668 3544
rect 3564 2716 3572 2724
rect 3580 2683 3588 2684
rect 3576 2677 3588 2683
rect 3580 2676 3588 2677
rect 3612 2683 3620 2684
rect 3608 2677 3620 2683
rect 3612 2676 3620 2677
rect 3532 2276 3540 2284
rect 3629 2148 3635 3112
rect 3644 2703 3652 2704
rect 3644 2697 3656 2703
rect 3644 2696 3652 2697
rect 3645 2648 3651 2672
rect 3677 2248 3683 3672
rect 3693 2888 3699 3312
rect 3692 2643 3700 2644
rect 3692 2637 3704 2643
rect 3692 2636 3700 2637
rect 3709 2248 3715 2412
rect 3725 2308 3731 3792
rect 4253 3788 4259 3872
rect 4525 3868 4531 3896
rect 4588 3876 4596 3884
rect 4589 3868 4595 3876
rect 4349 3748 4355 3792
rect 3788 3716 3796 3724
rect 3789 3708 3795 3716
rect 3740 3296 3748 3304
rect 3741 3268 3747 3296
rect 3740 2716 3748 2724
rect 3741 2308 3747 2716
rect 3725 1888 3731 1912
rect 3708 1883 3716 1884
rect 3704 1877 3716 1883
rect 3708 1876 3716 1877
rect 3644 1703 3652 1704
rect 3640 1697 3652 1703
rect 3644 1696 3652 1697
rect 3741 1568 3747 2292
rect 3789 2268 3795 3692
rect 3933 3624 3939 3692
rect 3932 3616 3940 3624
rect 3916 3483 3924 3484
rect 3912 3477 3924 3483
rect 3916 3476 3924 3477
rect 3789 1784 3795 2032
rect 3805 1968 3811 2872
rect 3821 2148 3827 3292
rect 3837 2208 3843 3052
rect 3853 2848 3859 3052
rect 3853 2188 3859 2752
rect 3837 2124 3843 2172
rect 3836 2116 3844 2124
rect 3853 2044 3859 2172
rect 3852 2036 3860 2044
rect 3788 1776 3796 1784
rect 3724 1523 3732 1524
rect 3720 1517 3732 1523
rect 3724 1516 3732 1517
rect 3549 1468 3555 1492
rect 3533 1128 3539 1332
rect 3549 1088 3555 1452
rect 3741 1304 3747 1312
rect 3740 1296 3748 1304
rect 3468 703 3476 704
rect 3464 697 3476 703
rect 3468 696 3476 697
rect 3405 288 3411 592
rect 3517 568 3523 992
rect 3549 768 3555 1072
rect 3565 568 3571 1092
rect 3596 1083 3604 1084
rect 3592 1077 3604 1083
rect 3596 1076 3604 1077
rect 3629 708 3635 1092
rect 3645 808 3651 1292
rect 3724 1123 3732 1124
rect 3720 1117 3732 1123
rect 3724 1116 3732 1117
rect 3773 1108 3779 1672
rect 3789 1348 3795 1776
rect 3804 1743 3812 1744
rect 3804 1737 3816 1743
rect 3804 1736 3812 1737
rect 3853 1368 3859 2012
rect 3869 1924 3875 2592
rect 3901 2488 3907 3032
rect 3917 2688 3923 2952
rect 3933 2288 3939 3616
rect 3949 2888 3955 3712
rect 3965 3664 3971 3692
rect 3964 3656 3972 3664
rect 4060 3516 4068 3524
rect 4010 3406 4016 3414
rect 4061 3388 4067 3516
rect 4108 3356 4116 3364
rect 4109 3328 4115 3356
rect 4060 3316 4068 3324
rect 3965 3008 3971 3132
rect 4044 3036 4052 3044
rect 4010 3006 4016 3014
rect 4045 2988 4051 3036
rect 4010 2606 4016 2614
rect 3885 1944 3891 1952
rect 3884 1936 3892 1944
rect 3868 1916 3876 1924
rect 3869 1888 3875 1916
rect 3869 1428 3875 1472
rect 3661 528 3667 652
rect 3660 503 3668 504
rect 3656 497 3668 503
rect 3660 496 3668 497
rect 3533 168 3539 432
rect 3677 48 3683 1092
rect 3788 1063 3796 1064
rect 3784 1057 3796 1063
rect 3788 1056 3796 1057
rect 3788 543 3796 544
rect 3784 537 3796 543
rect 3788 536 3796 537
rect 3805 28 3811 1272
rect 3885 708 3891 1412
rect 3837 348 3843 632
rect 3901 308 3907 2212
rect 3948 1963 3956 1964
rect 3944 1957 3956 1963
rect 3948 1956 3956 1957
rect 3965 1888 3971 2512
rect 4010 2206 4016 2214
rect 4029 2208 4035 2792
rect 4045 2584 4051 2792
rect 4061 2768 4067 3316
rect 4125 2768 4131 3652
rect 4349 3604 4355 3632
rect 4348 3596 4356 3604
rect 4141 2868 4147 3232
rect 4205 3088 4211 3492
rect 4237 3344 4243 3352
rect 4236 3336 4244 3344
rect 4332 3336 4340 3344
rect 4333 3328 4339 3336
rect 4221 2788 4227 3192
rect 4573 3188 4579 3812
rect 4605 3348 4611 3872
rect 4829 3748 4835 3932
rect 5356 3903 5364 3904
rect 5352 3897 5364 3903
rect 5356 3896 5364 3897
rect 5325 3884 5331 3892
rect 5324 3876 5332 3884
rect 5404 3883 5412 3884
rect 5404 3877 5416 3883
rect 5404 3876 5412 3877
rect 4044 2576 4052 2584
rect 4109 2288 4115 2592
rect 4157 2528 4163 2632
rect 3917 1348 3923 1652
rect 3948 1476 3956 1484
rect 3949 1468 3955 1476
rect 3965 1468 3971 1872
rect 4010 1806 4016 1814
rect 3981 1744 3987 1752
rect 3980 1736 3988 1744
rect 3965 1088 3971 1452
rect 4010 1406 4016 1414
rect 4029 1104 4035 2192
rect 4044 1576 4052 1584
rect 4045 1568 4051 1576
rect 4045 1248 4051 1552
rect 4028 1096 4036 1104
rect 4010 1006 4016 1014
rect 4061 788 4067 2212
rect 4125 1748 4131 2412
rect 4141 1988 4147 2052
rect 4157 1988 4163 2512
rect 4301 2488 4307 2832
rect 4141 1748 4147 1912
rect 4157 1728 4163 1952
rect 4173 1888 4179 2172
rect 4349 2128 4355 2732
rect 4429 2728 4435 3092
rect 4573 3028 4579 3052
rect 4445 2568 4451 2732
rect 4605 2728 4611 3332
rect 4621 3304 4627 3332
rect 4620 3296 4628 3304
rect 4653 3108 4659 3712
rect 4845 3688 4851 3752
rect 4669 3368 4675 3552
rect 4477 2468 4483 2652
rect 4412 2283 4420 2284
rect 4408 2277 4420 2283
rect 4412 2276 4420 2277
rect 4077 1368 4083 1532
rect 4093 1388 4099 1572
rect 4109 1308 4115 1572
rect 4173 1528 4179 1772
rect 4221 1488 4227 2072
rect 4252 2063 4260 2064
rect 4248 2057 4260 2063
rect 4252 2056 4260 2057
rect 4301 1928 4307 2012
rect 4268 1903 4276 1904
rect 4264 1897 4276 1903
rect 4268 1896 4276 1897
rect 4284 1903 4292 1904
rect 4284 1897 4296 1903
rect 4284 1896 4292 1897
rect 4220 1363 4228 1364
rect 4216 1357 4228 1363
rect 4220 1356 4228 1357
rect 4253 1068 4259 1852
rect 4317 1764 4323 1992
rect 4429 1868 4435 2392
rect 4477 2148 4483 2452
rect 4573 2228 4579 2372
rect 4316 1756 4324 1764
rect 4333 1468 4339 1772
rect 4445 1468 4451 1832
rect 4477 1548 4483 2132
rect 4525 1904 4531 1992
rect 4524 1896 4532 1904
rect 4573 1468 4579 1752
rect 4285 1284 4291 1292
rect 4284 1276 4292 1284
rect 4333 1148 4339 1452
rect 4621 1408 4627 1952
rect 4637 1888 4643 2192
rect 4653 1488 4659 3092
rect 4696 2957 4707 2963
rect 4701 2928 4707 2957
rect 4668 2916 4676 2924
rect 4669 2908 4675 2916
rect 4733 2868 4739 3552
rect 4780 3463 4788 3464
rect 4780 3457 4792 3463
rect 4780 3456 4788 3457
rect 4861 2508 4867 3412
rect 4460 1343 4468 1344
rect 4456 1337 4468 1343
rect 4460 1336 4468 1337
rect 4492 1343 4500 1344
rect 4492 1337 4504 1343
rect 4492 1336 4500 1337
rect 4701 1308 4707 2412
rect 4829 1828 4835 2152
rect 4732 1763 4740 1764
rect 4728 1757 4740 1763
rect 4732 1756 4740 1757
rect 4396 1303 4404 1304
rect 4392 1297 4404 1303
rect 4396 1296 4404 1297
rect 4477 1128 4483 1152
rect 4461 988 4467 1012
rect 4205 964 4211 972
rect 4204 956 4212 964
rect 3932 736 3940 744
rect 3933 728 3939 736
rect 4010 606 4016 614
rect 4140 563 4148 564
rect 4140 557 4152 563
rect 4140 556 4148 557
rect 4221 268 4227 972
rect 4477 964 4483 972
rect 4476 956 4484 964
rect 4509 788 4515 1072
rect 4557 788 4563 1172
rect 4285 684 4291 692
rect 4284 676 4292 684
rect 4557 468 4563 772
rect 4412 283 4420 284
rect 4408 277 4420 283
rect 4412 276 4420 277
rect 4010 206 4016 214
rect 4637 188 4643 1192
rect 4781 328 4787 1312
rect 4845 868 4851 2412
rect 4877 2128 4883 3432
rect 4909 2848 4915 3072
rect 4973 3068 4979 3632
rect 5050 3606 5056 3614
rect 5050 3206 5056 3214
rect 4957 2928 4963 3052
rect 4908 2676 4916 2684
rect 4909 2628 4915 2676
rect 4861 1168 4867 1432
rect 4909 228 4915 2612
rect 4973 2308 4979 2612
rect 4973 1868 4979 2092
rect 4989 1328 4995 2452
rect 5005 2148 5011 3012
rect 5050 2806 5056 2814
rect 5069 2748 5075 3332
rect 5117 2548 5123 3192
rect 5181 2888 5187 3632
rect 5341 3548 5347 3652
rect 5213 2808 5219 3512
rect 5229 2548 5235 3232
rect 5245 2948 5251 3472
rect 5341 3348 5347 3532
rect 5050 2406 5056 2414
rect 5052 2283 5060 2284
rect 5048 2277 5060 2283
rect 5052 2276 5060 2277
rect 5005 2008 5011 2132
rect 5036 2103 5044 2104
rect 5032 2097 5044 2103
rect 5036 2096 5044 2097
rect 5117 2088 5123 2532
rect 5050 2006 5056 2014
rect 5050 1606 5056 1614
rect 5133 1268 5139 1832
rect 5050 1206 5056 1214
rect 5050 806 5056 814
rect 4941 728 4947 752
rect 5149 568 5155 1792
rect 5165 1168 5171 1492
rect 5181 1388 5187 2252
rect 5197 1584 5203 2412
rect 5196 1576 5204 1584
rect 5180 1336 5188 1344
rect 5181 1328 5187 1336
rect 5213 1068 5219 2412
rect 5245 1868 5251 2592
rect 5293 2208 5299 2952
rect 5309 2288 5315 2932
rect 5325 2368 5331 3032
rect 5405 2528 5411 3692
rect 5453 3288 5459 3432
rect 5293 1588 5299 2192
rect 5293 1408 5299 1572
rect 5260 1323 5268 1324
rect 5260 1317 5272 1323
rect 5260 1316 5268 1317
rect 5229 1088 5235 1232
rect 5050 406 5056 414
rect 5149 328 5155 552
rect 5325 248 5331 2312
rect 5421 2288 5427 2972
rect 5340 2116 5348 2124
rect 5341 2108 5347 2116
rect 5341 1348 5347 1372
rect 5389 1068 5395 1632
rect 5405 548 5411 1932
rect 5437 1668 5443 3192
rect 5516 3083 5524 3084
rect 5516 3077 5528 3083
rect 5516 3076 5524 3077
rect 5501 2308 5507 2692
rect 5421 1328 5427 1432
rect 5421 908 5427 1312
rect 5437 1088 5443 1652
rect 5372 523 5380 524
rect 5368 517 5380 523
rect 5372 516 5380 517
rect 5469 428 5475 1632
rect 5501 1348 5507 2152
rect 5517 1228 5523 2812
rect 5533 2388 5539 3072
rect 5549 2688 5555 3392
rect 5533 1788 5539 2312
rect 5549 1628 5555 2032
rect 5565 1808 5571 3632
rect 5581 2768 5587 3292
rect 5693 3168 5699 3712
rect 5581 2348 5587 2752
rect 5581 1908 5587 2232
rect 5533 1208 5539 1372
rect 5581 548 5587 1232
rect 5597 928 5603 2412
rect 5613 2104 5619 2132
rect 5612 2096 5620 2104
rect 5613 308 5619 2096
rect 5629 1748 5635 1892
rect 5645 1808 5651 3112
rect 5709 3108 5715 3512
rect 5629 388 5635 1732
rect 5645 708 5651 1252
rect 5661 748 5667 2812
rect 5709 2788 5715 3092
rect 5677 1888 5683 2672
rect 5725 2528 5731 3592
rect 5757 3568 5763 3712
rect 5693 948 5699 1452
rect 5709 608 5715 1772
rect 5725 328 5731 2152
rect 5741 1428 5747 3232
rect 5757 3228 5763 3552
rect 5757 2824 5763 2832
rect 5756 2816 5764 2824
rect 5773 2308 5779 3312
rect 5740 1356 5748 1364
rect 5741 548 5747 1356
rect 5453 228 5459 272
rect 3917 128 3923 172
rect 5757 148 5763 2292
rect 5773 1328 5779 2212
rect 5789 1528 5795 3732
rect 5789 128 5795 1512
rect 5805 1248 5811 3612
rect 5821 2288 5827 3072
rect 5821 1708 5827 1792
rect 5821 1508 5827 1692
rect 5837 1088 5843 3632
rect 5869 3084 5875 3492
rect 5868 3076 5876 3084
rect 5869 2948 5875 3076
rect 5853 2837 5864 2843
rect 5853 1268 5859 2632
rect 5869 2548 5875 2652
rect 5869 1888 5875 2172
rect 5885 2148 5891 3872
rect 5901 2464 5907 3252
rect 5900 2456 5908 2464
rect 5884 2116 5892 2124
rect 5885 1308 5891 2116
rect 5901 1468 5907 2432
rect 5869 1088 5875 1252
rect 5917 688 5923 2552
rect 5933 1508 5939 2572
rect 5932 563 5940 564
rect 5928 557 5940 563
rect 5932 556 5940 557
rect 5949 148 5955 1852
rect 5965 1708 5971 3032
rect 5965 368 5971 1432
rect 954 6 960 14
rect 3002 6 3008 14
rect 5050 6 5056 14
use AND2X2  AND2X2_506
timestamp 1516238463
transform -1 0 72 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_528
timestamp 1516238463
transform 1 0 72 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_505
timestamp 1516238463
transform -1 0 200 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_482
timestamp 1516238463
transform 1 0 200 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_481
timestamp 1516238463
transform -1 0 328 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_4
timestamp 1516238463
transform -1 0 424 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_104
timestamp 1516238463
transform -1 0 520 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_3
timestamp 1516238463
transform 1 0 520 0 1 3810
box 0 0 96 200
use AND2X2  AND2X2_494
timestamp 1516238463
transform 1 0 616 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_347
timestamp 1516238463
transform 1 0 680 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_493
timestamp 1516238463
transform -1 0 808 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_472
timestamp 1516238463
transform 1 0 808 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_103
timestamp 1516238463
transform -1 0 968 0 1 3810
box 0 0 96 200
use FILL  FILL_19_0_0
timestamp 1516238463
transform -1 0 984 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_1
timestamp 1516238463
transform -1 0 1000 0 1 3810
box 0 0 16 200
use AND2X2  AND2X2_471
timestamp 1516238463
transform -1 0 1064 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_370
timestamp 1516238463
transform -1 0 1128 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_84
timestamp 1516238463
transform -1 0 1224 0 1 3810
box 0 0 96 200
use AND2X2  AND2X2_386
timestamp 1516238463
transform 1 0 1224 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_261
timestamp 1516238463
transform -1 0 1352 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_458
timestamp 1516238463
transform -1 0 1416 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_387
timestamp 1516238463
transform -1 0 1480 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_402
timestamp 1516238463
transform -1 0 1544 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_431
timestamp 1516238463
transform -1 0 1608 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_456
timestamp 1516238463
transform -1 0 1672 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_110
timestamp 1516238463
transform -1 0 1736 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_112
timestamp 1516238463
transform 1 0 1736 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_413
timestamp 1516238463
transform -1 0 1864 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_303
timestamp 1516238463
transform -1 0 1928 0 1 3810
box 0 0 64 200
use FILL  FILL_19_1_0
timestamp 1516238463
transform -1 0 1944 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_1
timestamp 1516238463
transform -1 0 1960 0 1 3810
box 0 0 16 200
use AND2X2  AND2X2_443
timestamp 1516238463
transform -1 0 2024 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_442
timestamp 1516238463
transform -1 0 2088 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_100
timestamp 1516238463
transform -1 0 2184 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_99
timestamp 1516238463
transform -1 0 2280 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_101
timestamp 1516238463
transform -1 0 2376 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_102
timestamp 1516238463
transform -1 0 2472 0 1 3810
box 0 0 96 200
use BUFX4  BUFX4_37
timestamp 1516238463
transform -1 0 2536 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_39
timestamp 1516238463
transform -1 0 2600 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_109
timestamp 1516238463
transform -1 0 2664 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_86
timestamp 1516238463
transform -1 0 2760 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_90
timestamp 1516238463
transform -1 0 2856 0 1 3810
box 0 0 96 200
use BUFX4  BUFX4_90
timestamp 1516238463
transform -1 0 2920 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_92
timestamp 1516238463
transform -1 0 2984 0 1 3810
box 0 0 64 200
use FILL  FILL_19_2_0
timestamp 1516238463
transform 1 0 2984 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_1
timestamp 1516238463
transform 1 0 3000 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_114
timestamp 1516238463
transform 1 0 3016 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_34
timestamp 1516238463
transform 1 0 3080 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_187
timestamp 1516238463
transform -1 0 3208 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_43
timestamp 1516238463
transform -1 0 3272 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_121
timestamp 1516238463
transform -1 0 3336 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_122
timestamp 1516238463
transform -1 0 3400 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_59
timestamp 1516238463
transform -1 0 3464 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_49
timestamp 1516238463
transform -1 0 3560 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_69
timestamp 1516238463
transform -1 0 3656 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_11
timestamp 1516238463
transform -1 0 3752 0 1 3810
box 0 0 96 200
use BUFX4  BUFX4_84
timestamp 1516238463
transform -1 0 3816 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_87
timestamp 1516238463
transform 1 0 3816 0 1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_19
timestamp 1516238463
transform 1 0 3880 0 1 3810
box 0 0 96 200
use FILL  FILL_19_3_0
timestamp 1516238463
transform 1 0 3976 0 1 3810
box 0 0 16 200
use FILL  FILL_19_3_1
timestamp 1516238463
transform 1 0 3992 0 1 3810
box 0 0 16 200
use MUX2X1  MUX2X1_12
timestamp 1516238463
transform 1 0 4008 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_21
timestamp 1516238463
transform 1 0 4104 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_13
timestamp 1516238463
transform 1 0 4200 0 1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_20
timestamp 1516238463
transform 1 0 4296 0 1 3810
box 0 0 96 200
use AND2X2  AND2X2_368
timestamp 1516238463
transform -1 0 4456 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_379
timestamp 1516238463
transform -1 0 4520 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_45
timestamp 1516238463
transform -1 0 4584 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_20
timestamp 1516238463
transform -1 0 4648 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_85
timestamp 1516238463
transform -1 0 4712 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_84
timestamp 1516238463
transform -1 0 4776 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_620
timestamp 1516238463
transform -1 0 4840 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_621
timestamp 1516238463
transform -1 0 4904 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_38
timestamp 1516238463
transform -1 0 4968 0 1 3810
box 0 0 64 200
use BUFX4  BUFX4_115
timestamp 1516238463
transform 1 0 4968 0 1 3810
box 0 0 64 200
use FILL  FILL_19_4_0
timestamp 1516238463
transform 1 0 5032 0 1 3810
box 0 0 16 200
use FILL  FILL_19_4_1
timestamp 1516238463
transform 1 0 5048 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_36
timestamp 1516238463
transform 1 0 5064 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_50
timestamp 1516238463
transform -1 0 5192 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_65
timestamp 1516238463
transform -1 0 5256 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_66
timestamp 1516238463
transform -1 0 5320 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_631
timestamp 1516238463
transform -1 0 5384 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_568
timestamp 1516238463
transform 1 0 5384 0 1 3810
box 0 0 64 200
use OR2X2  OR2X2_346
timestamp 1516238463
transform -1 0 5512 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_579
timestamp 1516238463
transform -1 0 5576 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_57
timestamp 1516238463
transform -1 0 5640 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_3
timestamp 1516238463
transform -1 0 5704 0 1 3810
box 0 0 64 200
use AND2X2  AND2X2_46
timestamp 1516238463
transform -1 0 5768 0 1 3810
box 0 0 64 200
use BUFX2  BUFX2_35
timestamp 1516238463
transform 1 0 5768 0 1 3810
box 0 0 48 200
use BUFX2  BUFX2_70
timestamp 1516238463
transform 1 0 5816 0 1 3810
box 0 0 48 200
use XOR2X1  XOR2X1_4
timestamp 1516238463
transform -1 0 5976 0 1 3810
box 0 0 112 200
use FILL  FILL_20_1
timestamp 1516238463
transform 1 0 5976 0 1 3810
box 0 0 16 200
use OR2X2  OR2X2_358
timestamp 1516238463
transform 1 0 8 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_376
timestamp 1516238463
transform -1 0 136 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_529
timestamp 1516238463
transform -1 0 200 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_337
timestamp 1516238463
transform -1 0 264 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_370
timestamp 1516238463
transform -1 0 328 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_520
timestamp 1516238463
transform -1 0 392 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_519
timestamp 1516238463
transform -1 0 456 0 -1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_5
timestamp 1516238463
transform -1 0 552 0 -1 3810
box 0 0 96 200
use AND2X2  AND2X2_544
timestamp 1516238463
transform 1 0 552 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_389
timestamp 1516238463
transform 1 0 616 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_391
timestamp 1516238463
transform 1 0 680 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_543
timestamp 1516238463
transform -1 0 808 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_322
timestamp 1516238463
transform -1 0 872 0 -1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_6
timestamp 1516238463
transform -1 0 968 0 -1 3810
box 0 0 96 200
use FILL  FILL_18_0_0
timestamp 1516238463
transform -1 0 984 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_1
timestamp 1516238463
transform -1 0 1000 0 -1 3810
box 0 0 16 200
use MUX2X1  MUX2X1_7
timestamp 1516238463
transform -1 0 1096 0 -1 3810
box 0 0 96 200
use NAND3X1  NAND3X1_60
timestamp 1516238463
transform -1 0 1160 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_311
timestamp 1516238463
transform -1 0 1224 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_418
timestamp 1516238463
transform -1 0 1288 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_398
timestamp 1516238463
transform -1 0 1352 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_272
timestamp 1516238463
transform -1 0 1416 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_403
timestamp 1516238463
transform -1 0 1480 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_294
timestamp 1516238463
transform -1 0 1544 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_430
timestamp 1516238463
transform -1 0 1608 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_282
timestamp 1516238463
transform -1 0 1672 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_414
timestamp 1516238463
transform -1 0 1736 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_304
timestamp 1516238463
transform -1 0 1800 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_447
timestamp 1516238463
transform -1 0 1864 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_448
timestamp 1516238463
transform -1 0 1928 0 -1 3810
box 0 0 64 200
use FILL  FILL_18_1_0
timestamp 1516238463
transform -1 0 1944 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_1
timestamp 1516238463
transform -1 0 1960 0 -1 3810
box 0 0 16 200
use OR2X2  OR2X2_283
timestamp 1516238463
transform -1 0 2024 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_416
timestamp 1516238463
transform -1 0 2088 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_417
timestamp 1516238463
transform -1 0 2152 0 -1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_81
timestamp 1516238463
transform -1 0 2248 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_96
timestamp 1516238463
transform -1 0 2344 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_87
timestamp 1516238463
transform -1 0 2440 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_82
timestamp 1516238463
transform -1 0 2536 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_77
timestamp 1516238463
transform -1 0 2632 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_98
timestamp 1516238463
transform 1 0 2632 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_95
timestamp 1516238463
transform 1 0 2728 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_80
timestamp 1516238463
transform -1 0 2920 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_73
timestamp 1516238463
transform -1 0 3016 0 -1 3810
box 0 0 96 200
use FILL  FILL_18_2_0
timestamp 1516238463
transform -1 0 3032 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_1
timestamp 1516238463
transform -1 0 3048 0 -1 3810
box 0 0 16 200
use OR2X2  OR2X2_92
timestamp 1516238463
transform -1 0 3112 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_186
timestamp 1516238463
transform -1 0 3176 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_250
timestamp 1516238463
transform -1 0 3240 0 -1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_74
timestamp 1516238463
transform -1 0 3336 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_76
timestamp 1516238463
transform -1 0 3432 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_64
timestamp 1516238463
transform -1 0 3528 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_16
timestamp 1516238463
transform -1 0 3624 0 -1 3810
box 0 0 96 200
use BUFX4  BUFX4_86
timestamp 1516238463
transform -1 0 3688 0 -1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_94
timestamp 1516238463
transform 1 0 3688 0 -1 3810
box 0 0 96 200
use BUFX4  BUFX4_91
timestamp 1516238463
transform -1 0 3848 0 -1 3810
box 0 0 64 200
use MUX2X1  MUX2X1_83
timestamp 1516238463
transform -1 0 3944 0 -1 3810
box 0 0 96 200
use MUX2X1  MUX2X1_10
timestamp 1516238463
transform 1 0 3944 0 -1 3810
box 0 0 96 200
use FILL  FILL_18_3_0
timestamp 1516238463
transform 1 0 4040 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_1
timestamp 1516238463
transform 1 0 4056 0 -1 3810
box 0 0 16 200
use MUX2X1  MUX2X1_22
timestamp 1516238463
transform 1 0 4072 0 -1 3810
box 0 0 96 200
use INVX4  INVX4_4
timestamp 1516238463
transform -1 0 4216 0 -1 3810
box 0 0 48 200
use OR2X2  OR2X2_453
timestamp 1516238463
transform -1 0 4280 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_44
timestamp 1516238463
transform -1 0 4344 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_235
timestamp 1516238463
transform -1 0 4408 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_157
timestamp 1516238463
transform -1 0 4472 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_257
timestamp 1516238463
transform -1 0 4536 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_268
timestamp 1516238463
transform -1 0 4600 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_33
timestamp 1516238463
transform -1 0 4664 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_113
timestamp 1516238463
transform -1 0 4728 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_416
timestamp 1516238463
transform -1 0 4792 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_455
timestamp 1516238463
transform -1 0 4856 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_49
timestamp 1516238463
transform -1 0 4920 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_111
timestamp 1516238463
transform 1 0 4920 0 -1 3810
box 0 0 64 200
use INVX1  INVX1_1
timestamp 1516238463
transform 1 0 4984 0 -1 3810
box 0 0 32 200
use FILL  FILL_18_4_0
timestamp 1516238463
transform 1 0 5016 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_4_1
timestamp 1516238463
transform 1 0 5032 0 -1 3810
box 0 0 16 200
use OR2X2  OR2X2_414
timestamp 1516238463
transform 1 0 5048 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_335
timestamp 1516238463
transform -1 0 5176 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_8
timestamp 1516238463
transform -1 0 5240 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_426
timestamp 1516238463
transform -1 0 5304 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_632
timestamp 1516238463
transform -1 0 5368 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_116
timestamp 1516238463
transform -1 0 5432 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_4
timestamp 1516238463
transform -1 0 5496 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_428
timestamp 1516238463
transform 1 0 5496 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_35
timestamp 1516238463
transform -1 0 5624 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_120
timestamp 1516238463
transform 1 0 5624 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_445
timestamp 1516238463
transform 1 0 5688 0 -1 3810
box 0 0 64 200
use AND2X2  AND2X2_556
timestamp 1516238463
transform 1 0 5752 0 -1 3810
box 0 0 64 200
use OR2X2  OR2X2_452
timestamp 1516238463
transform 1 0 5816 0 -1 3810
box 0 0 64 200
use BUFX4  BUFX4_42
timestamp 1516238463
transform 1 0 5880 0 -1 3810
box 0 0 64 200
use FILL  FILL_19_1
timestamp 1516238463
transform -1 0 5960 0 -1 3810
box 0 0 16 200
use FILL  FILL_19_2
timestamp 1516238463
transform -1 0 5976 0 -1 3810
box 0 0 16 200
use FILL  FILL_19_3
timestamp 1516238463
transform -1 0 5992 0 -1 3810
box 0 0 16 200
use AND2X2  AND2X2_504
timestamp 1516238463
transform -1 0 72 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_530
timestamp 1516238463
transform 1 0 72 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_531
timestamp 1516238463
transform -1 0 200 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_459
timestamp 1516238463
transform -1 0 264 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_521
timestamp 1516238463
transform 1 0 264 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_483
timestamp 1516238463
transform 1 0 328 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_455
timestamp 1516238463
transform -1 0 456 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_404
timestamp 1516238463
transform 1 0 456 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_400
timestamp 1516238463
transform -1 0 584 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_484
timestamp 1516238463
transform -1 0 648 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_371
timestamp 1516238463
transform 1 0 648 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_546
timestamp 1516238463
transform -1 0 776 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_392
timestamp 1516238463
transform -1 0 840 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_432
timestamp 1516238463
transform 1 0 840 0 1 3410
box 0 0 64 200
use FILL  FILL_17_0_0
timestamp 1516238463
transform -1 0 920 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_1
timestamp 1516238463
transform -1 0 936 0 1 3410
box 0 0 16 200
use OR2X2  OR2X2_245
timestamp 1516238463
transform -1 0 1000 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_429
timestamp 1516238463
transform -1 0 1064 0 1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_63
timestamp 1516238463
transform -1 0 1112 0 1 3410
box 0 0 48 200
use AND2X2  AND2X2_369
timestamp 1516238463
transform -1 0 1176 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_284
timestamp 1516238463
transform -1 0 1240 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_551
timestamp 1516238463
transform -1 0 1304 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_415
timestamp 1516238463
transform -1 0 1368 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_325
timestamp 1516238463
transform -1 0 1432 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_10
timestamp 1516238463
transform -1 0 1496 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_449
timestamp 1516238463
transform -1 0 1560 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_339
timestamp 1516238463
transform 1 0 1560 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_338
timestamp 1516238463
transform -1 0 1688 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_302
timestamp 1516238463
transform -1 0 1752 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_300
timestamp 1516238463
transform -1 0 1816 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_267
timestamp 1516238463
transform -1 0 1880 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_266
timestamp 1516238463
transform -1 0 1944 0 1 3410
box 0 0 64 200
use FILL  FILL_17_1_0
timestamp 1516238463
transform 1 0 1944 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_1
timestamp 1516238463
transform 1 0 1960 0 1 3410
box 0 0 16 200
use MUX2X1  MUX2X1_88
timestamp 1516238463
transform 1 0 1976 0 1 3410
box 0 0 96 200
use AND2X2  AND2X2_352
timestamp 1516238463
transform -1 0 2136 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_353
timestamp 1516238463
transform -1 0 2200 0 1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_97
timestamp 1516238463
transform -1 0 2296 0 1 3410
box 0 0 96 200
use MUX2X1  MUX2X1_93
timestamp 1516238463
transform -1 0 2392 0 1 3410
box 0 0 96 200
use AND2X2  AND2X2_316
timestamp 1516238463
transform -1 0 2456 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_233
timestamp 1516238463
transform -1 0 2520 0 1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_85
timestamp 1516238463
transform -1 0 2616 0 1 3410
box 0 0 96 200
use AND2X2  AND2X2_317
timestamp 1516238463
transform -1 0 2680 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_284
timestamp 1516238463
transform 1 0 2680 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_232
timestamp 1516238463
transform -1 0 2808 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_155
timestamp 1516238463
transform -1 0 2872 0 1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_75
timestamp 1516238463
transform 1 0 2872 0 1 3410
box 0 0 96 200
use FILL  FILL_17_2_0
timestamp 1516238463
transform -1 0 2984 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_1
timestamp 1516238463
transform -1 0 3000 0 1 3410
box 0 0 16 200
use AND2X2  AND2X2_154
timestamp 1516238463
transform -1 0 3064 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_97
timestamp 1516238463
transform 1 0 3064 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_137
timestamp 1516238463
transform -1 0 3192 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_285
timestamp 1516238463
transform -1 0 3256 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_249
timestamp 1516238463
transform -1 0 3320 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_346
timestamp 1516238463
transform -1 0 3384 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_224
timestamp 1516238463
transform -1 0 3448 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_335
timestamp 1516238463
transform -1 0 3512 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_4
timestamp 1516238463
transform 1 0 3512 0 1 3410
box 0 0 48 200
use NAND2X1  NAND2X1_52
timestamp 1516238463
transform -1 0 3608 0 1 3410
box 0 0 48 200
use BUFX4  BUFX4_88
timestamp 1516238463
transform -1 0 3672 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_89
timestamp 1516238463
transform 1 0 3672 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_177
timestamp 1516238463
transform -1 0 3800 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_51
timestamp 1516238463
transform 1 0 3800 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_468
timestamp 1516238463
transform -1 0 3928 0 1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_15
timestamp 1516238463
transform 1 0 3928 0 1 3410
box 0 0 96 200
use FILL  FILL_17_3_0
timestamp 1516238463
transform -1 0 4040 0 1 3410
box 0 0 16 200
use FILL  FILL_17_3_1
timestamp 1516238463
transform -1 0 4056 0 1 3410
box 0 0 16 200
use MUX2X1  MUX2X1_14
timestamp 1516238463
transform -1 0 4152 0 1 3410
box 0 0 96 200
use AND2X2  AND2X2_120
timestamp 1516238463
transform -1 0 4216 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_119
timestamp 1516238463
transform -1 0 4280 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_268
timestamp 1516238463
transform -1 0 4344 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_446
timestamp 1516238463
transform -1 0 4408 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_457
timestamp 1516238463
transform -1 0 4472 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_52
timestamp 1516238463
transform 1 0 4472 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_36
timestamp 1516238463
transform 1 0 4536 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_257
timestamp 1516238463
transform -1 0 4664 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_412
timestamp 1516238463
transform -1 0 4728 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_423
timestamp 1516238463
transform -1 0 4792 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_40
timestamp 1516238463
transform -1 0 4856 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_32
timestamp 1516238463
transform 1 0 4856 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_415
timestamp 1516238463
transform -1 0 4984 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_618
timestamp 1516238463
transform -1 0 5048 0 1 3410
box 0 0 64 200
use FILL  FILL_17_4_0
timestamp 1516238463
transform -1 0 5064 0 1 3410
box 0 0 16 200
use FILL  FILL_17_4_1
timestamp 1516238463
transform -1 0 5080 0 1 3410
box 0 0 16 200
use AND2X2  AND2X2_619
timestamp 1516238463
transform -1 0 5144 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_39
timestamp 1516238463
transform -1 0 5208 0 1 3410
box 0 0 64 200
use OR2X2  OR2X2_425
timestamp 1516238463
transform -1 0 5272 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_88
timestamp 1516238463
transform -1 0 5336 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_13
timestamp 1516238463
transform 1 0 5336 0 1 3410
box 0 0 64 200
use XNOR2X1  XNOR2X1_1
timestamp 1516238463
transform -1 0 5512 0 1 3410
box 0 0 112 200
use AND2X2  AND2X2_70
timestamp 1516238463
transform -1 0 5576 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_90
timestamp 1516238463
transform 1 0 5576 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_101
timestamp 1516238463
transform -1 0 5704 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_6
timestamp 1516238463
transform 1 0 5704 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_7
timestamp 1516238463
transform -1 0 5832 0 1 3410
box 0 0 64 200
use BUFX4  BUFX4_119
timestamp 1516238463
transform 1 0 5832 0 1 3410
box 0 0 64 200
use AND2X2  AND2X2_203
timestamp 1516238463
transform -1 0 5960 0 1 3410
box 0 0 64 200
use FILL  FILL_18_1
timestamp 1516238463
transform 1 0 5960 0 1 3410
box 0 0 16 200
use FILL  FILL_18_2
timestamp 1516238463
transform 1 0 5976 0 1 3410
box 0 0 16 200
use OR2X2  OR2X2_359
timestamp 1516238463
transform 1 0 8 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_507
timestamp 1516238463
transform -1 0 136 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_377
timestamp 1516238463
transform 1 0 136 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_313
timestamp 1516238463
transform -1 0 264 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_371
timestamp 1516238463
transform -1 0 328 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_518
timestamp 1516238463
transform -1 0 392 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_554
timestamp 1516238463
transform 1 0 392 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_273
timestamp 1516238463
transform -1 0 520 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_338
timestamp 1516238463
transform -1 0 584 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_399
timestamp 1516238463
transform -1 0 648 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_247
timestamp 1516238463
transform -1 0 712 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_367
timestamp 1516238463
transform -1 0 776 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_303
timestamp 1516238463
transform 1 0 776 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_185
timestamp 1516238463
transform -1 0 904 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_0_0
timestamp 1516238463
transform -1 0 920 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_1
timestamp 1516238463
transform -1 0 936 0 -1 3410
box 0 0 16 200
use OR2X2  OR2X2_295
timestamp 1516238463
transform -1 0 1000 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_348
timestamp 1516238463
transform -1 0 1064 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_299
timestamp 1516238463
transform -1 0 1128 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_552
timestamp 1516238463
transform 1 0 1128 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_553
timestamp 1516238463
transform -1 0 1256 0 -1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_91
timestamp 1516238463
transform -1 0 1352 0 -1 3410
box 0 0 96 200
use OR2X2  OR2X2_218
timestamp 1516238463
transform -1 0 1416 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_337
timestamp 1516238463
transform -1 0 1480 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_17
timestamp 1516238463
transform -1 0 1544 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_340
timestamp 1516238463
transform -1 0 1608 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_217
timestamp 1516238463
transform -1 0 1672 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_184
timestamp 1516238463
transform -1 0 1736 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_131
timestamp 1516238463
transform -1 0 1800 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_152
timestamp 1516238463
transform -1 0 1864 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_128
timestamp 1516238463
transform -1 0 1928 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_1_0
timestamp 1516238463
transform -1 0 1944 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_1
timestamp 1516238463
transform -1 0 1960 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_134
timestamp 1516238463
transform -1 0 2024 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_234
timestamp 1516238463
transform -1 0 2088 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_74
timestamp 1516238463
transform 1 0 2088 0 -1 3410
box 0 0 48 200
use OR2X2  OR2X2_421
timestamp 1516238463
transform -1 0 2200 0 -1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_79
timestamp 1516238463
transform -1 0 2296 0 -1 3410
box 0 0 96 200
use AND2X2  AND2X2_318
timestamp 1516238463
transform -1 0 2360 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_198
timestamp 1516238463
transform -1 0 2424 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_122
timestamp 1516238463
transform -1 0 2488 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_66
timestamp 1516238463
transform -1 0 2552 0 -1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_78
timestamp 1516238463
transform 1 0 2552 0 -1 3410
box 0 0 96 200
use OR2X2  OR2X2_170
timestamp 1516238463
transform -1 0 2712 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_28
timestamp 1516238463
transform -1 0 2776 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_96
timestamp 1516238463
transform -1 0 2840 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_133
timestamp 1516238463
transform 1 0 2840 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_462
timestamp 1516238463
transform -1 0 2968 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_2_0
timestamp 1516238463
transform -1 0 2984 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_1
timestamp 1516238463
transform -1 0 3000 0 -1 3410
box 0 0 16 200
use AND2X2  AND2X2_58
timestamp 1516238463
transform -1 0 3064 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_461
timestamp 1516238463
transform -1 0 3128 0 -1 3410
box 0 0 64 200
use INVX1  INVX1_44
timestamp 1516238463
transform -1 0 3160 0 -1 3410
box 0 0 32 200
use AND2X2  AND2X2_176
timestamp 1516238463
transform 1 0 3160 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_84
timestamp 1516238463
transform -1 0 3288 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_451
timestamp 1516238463
transform -1 0 3352 0 -1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_48
timestamp 1516238463
transform -1 0 3448 0 -1 3410
box 0 0 96 200
use NOR2X1  NOR2X1_10
timestamp 1516238463
transform -1 0 3496 0 -1 3410
box 0 0 48 200
use MUX2X1  MUX2X1_18
timestamp 1516238463
transform -1 0 3592 0 -1 3410
box 0 0 96 200
use MUX2X1  MUX2X1_2
timestamp 1516238463
transform -1 0 3688 0 -1 3410
box 0 0 96 200
use MUX2X1  MUX2X1_23
timestamp 1516238463
transform 1 0 3688 0 -1 3410
box 0 0 96 200
use OR2X2  OR2X2_457
timestamp 1516238463
transform -1 0 3848 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_54
timestamp 1516238463
transform -1 0 3912 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_87
timestamp 1516238463
transform -1 0 3976 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_3_0
timestamp 1516238463
transform -1 0 3992 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_3_1
timestamp 1516238463
transform -1 0 4008 0 -1 3410
box 0 0 16 200
use AND2X2  AND2X2_180
timestamp 1516238463
transform -1 0 4072 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_181
timestamp 1516238463
transform -1 0 4136 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_41
timestamp 1516238463
transform -1 0 4200 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_448
timestamp 1516238463
transform -1 0 4264 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_38
timestamp 1516238463
transform -1 0 4328 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_41
timestamp 1516238463
transform -1 0 4392 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_184
timestamp 1516238463
transform -1 0 4456 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_456
timestamp 1516238463
transform -1 0 4520 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_53
timestamp 1516238463
transform -1 0 4584 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_446
timestamp 1516238463
transform -1 0 4648 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_37
timestamp 1516238463
transform -1 0 4712 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_168
timestamp 1516238463
transform -1 0 4776 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_290
timestamp 1516238463
transform -1 0 4840 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_301
timestamp 1516238463
transform -1 0 4904 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_40
timestamp 1516238463
transform 1 0 4904 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_447
timestamp 1516238463
transform -1 0 5032 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_4_0
timestamp 1516238463
transform 1 0 5032 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_4_1
timestamp 1516238463
transform 1 0 5048 0 -1 3410
box 0 0 16 200
use AND2X2  AND2X2_89
timestamp 1516238463
transform 1 0 5064 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_22
timestamp 1516238463
transform -1 0 5192 0 -1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_65
timestamp 1516238463
transform -1 0 5288 0 -1 3410
box 0 0 96 200
use AND2X2  AND2X2_24
timestamp 1516238463
transform 1 0 5288 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_24
timestamp 1516238463
transform -1 0 5416 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_10
timestamp 1516238463
transform -1 0 5480 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_71
timestamp 1516238463
transform -1 0 5544 0 -1 3410
box 0 0 64 200
use AND2X2  AND2X2_133
timestamp 1516238463
transform -1 0 5608 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_57
timestamp 1516238463
transform 1 0 5608 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_7
timestamp 1516238463
transform -1 0 5736 0 -1 3410
box 0 0 64 200
use OR2X2  OR2X2_429
timestamp 1516238463
transform -1 0 5800 0 -1 3410
box 0 0 64 200
use BUFX4  BUFX4_8
timestamp 1516238463
transform 1 0 5800 0 -1 3410
box 0 0 64 200
use MUX2X1  MUX2X1_51
timestamp 1516238463
transform 1 0 5864 0 -1 3410
box 0 0 96 200
use FILL  FILL_17_1
timestamp 1516238463
transform -1 0 5976 0 -1 3410
box 0 0 16 200
use FILL  FILL_17_2
timestamp 1516238463
transform -1 0 5992 0 -1 3410
box 0 0 16 200
use AND2X2  AND2X2_555
timestamp 1516238463
transform -1 0 72 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_508
timestamp 1516238463
transform 1 0 72 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_532
timestamp 1516238463
transform -1 0 200 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_372
timestamp 1516238463
transform 1 0 200 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_522
timestamp 1516238463
transform 1 0 264 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_373
timestamp 1516238463
transform -1 0 392 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_324
timestamp 1516238463
transform 1 0 392 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_485
timestamp 1516238463
transform -1 0 520 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_474
timestamp 1516238463
transform -1 0 584 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_473
timestamp 1516238463
transform -1 0 648 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_393
timestamp 1516238463
transform 1 0 648 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_470
timestamp 1516238463
transform -1 0 776 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_62
timestamp 1516238463
transform 1 0 776 0 1 3010
box 0 0 48 200
use AOI21X1  AOI21X1_30
timestamp 1516238463
transform 1 0 824 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_419
timestamp 1516238463
transform 1 0 888 0 1 3010
box 0 0 64 200
use FILL  FILL_15_0_0
timestamp 1516238463
transform -1 0 968 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_1
timestamp 1516238463
transform -1 0 984 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_496
timestamp 1516238463
transform -1 0 1048 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_495
timestamp 1516238463
transform -1 0 1112 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_234
timestamp 1516238463
transform -1 0 1176 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_231
timestamp 1516238463
transform -1 0 1240 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_349
timestamp 1516238463
transform -1 0 1304 0 1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_89
timestamp 1516238463
transform -1 0 1400 0 1 3010
box 0 0 96 200
use BUFX4  BUFX4_18
timestamp 1516238463
transform -1 0 1464 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_444
timestamp 1516238463
transform -1 0 1528 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_156
timestamp 1516238463
transform 1 0 1528 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_269
timestamp 1516238463
transform 1 0 1592 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_265
timestamp 1516238463
transform 1 0 1656 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_153
timestamp 1516238463
transform 1 0 1720 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_270
timestamp 1516238463
transform 1 0 1784 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_354
timestamp 1516238463
transform -1 0 1912 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_355
timestamp 1516238463
transform -1 0 1976 0 1 3010
box 0 0 64 200
use FILL  FILL_15_1_0
timestamp 1516238463
transform 1 0 1976 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_1
timestamp 1516238463
transform 1 0 1992 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_381
timestamp 1516238463
transform 1 0 2008 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_319
timestamp 1516238463
transform -1 0 2136 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_252
timestamp 1516238463
transform -1 0 2200 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_251
timestamp 1516238463
transform -1 0 2264 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_123
timestamp 1516238463
transform -1 0 2328 0 1 3010
box 0 0 64 200
use AOI21X1  AOI21X1_39
timestamp 1516238463
transform -1 0 2392 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_171
timestamp 1516238463
transform -1 0 2456 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_286
timestamp 1516238463
transform -1 0 2520 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_287
timestamp 1516238463
transform -1 0 2584 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_188
timestamp 1516238463
transform 1 0 2584 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_189
timestamp 1516238463
transform -1 0 2712 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_3
timestamp 1516238463
transform -1 0 2776 0 1 3010
box 0 0 64 200
use INVX1  INVX1_45
timestamp 1516238463
transform 1 0 2776 0 1 3010
box 0 0 32 200
use NAND2X1  NAND2X1_67
timestamp 1516238463
transform -1 0 2856 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_15
timestamp 1516238463
transform 1 0 2856 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_41
timestamp 1516238463
transform -1 0 2952 0 1 3010
box 0 0 48 200
use FILL  FILL_15_2_0
timestamp 1516238463
transform 1 0 2952 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_1
timestamp 1516238463
transform 1 0 2968 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_11
timestamp 1516238463
transform 1 0 2984 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_47
timestamp 1516238463
transform -1 0 3112 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_390
timestamp 1516238463
transform -1 0 3176 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_130
timestamp 1516238463
transform 1 0 3176 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_117
timestamp 1516238463
transform 1 0 3240 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_116
timestamp 1516238463
transform -1 0 3368 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_434
timestamp 1516238463
transform -1 0 3432 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_14
timestamp 1516238463
transform -1 0 3496 0 1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_8
timestamp 1516238463
transform -1 0 3592 0 1 3010
box 0 0 96 200
use MUX2X1  MUX2X1_39
timestamp 1516238463
transform 1 0 3592 0 1 3010
box 0 0 96 200
use AND2X2  AND2X2_185
timestamp 1516238463
transform -1 0 3752 0 1 3010
box 0 0 64 200
use INVX4  INVX4_3
timestamp 1516238463
transform 1 0 3752 0 1 3010
box 0 0 48 200
use OR2X2  OR2X2_21
timestamp 1516238463
transform -1 0 3864 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_135
timestamp 1516238463
transform 1 0 3864 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_132
timestamp 1516238463
transform 1 0 3928 0 1 3010
box 0 0 64 200
use FILL  FILL_15_3_0
timestamp 1516238463
transform 1 0 3992 0 1 3010
box 0 0 16 200
use FILL  FILL_15_3_1
timestamp 1516238463
transform 1 0 4008 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_214
timestamp 1516238463
transform 1 0 4024 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_34
timestamp 1516238463
transform -1 0 4152 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_279
timestamp 1516238463
transform -1 0 4216 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_88
timestamp 1516238463
transform -1 0 4280 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_183
timestamp 1516238463
transform -1 0 4344 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_445
timestamp 1516238463
transform -1 0 4408 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_30
timestamp 1516238463
transform -1 0 4472 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_443
timestamp 1516238463
transform -1 0 4536 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_29
timestamp 1516238463
transform -1 0 4600 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_4
timestamp 1516238463
transform 1 0 4600 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_28
timestamp 1516238463
transform -1 0 4728 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_545
timestamp 1516238463
transform -1 0 4792 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_124
timestamp 1516238463
transform -1 0 4856 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_179
timestamp 1516238463
transform -1 0 4920 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_190
timestamp 1516238463
transform -1 0 4984 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_33
timestamp 1516238463
transform -1 0 5048 0 1 3010
box 0 0 64 200
use FILL  FILL_15_4_0
timestamp 1516238463
transform -1 0 5064 0 1 3010
box 0 0 16 200
use FILL  FILL_15_4_1
timestamp 1516238463
transform -1 0 5080 0 1 3010
box 0 0 16 200
use OR2X2  OR2X2_444
timestamp 1516238463
transform -1 0 5144 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_32
timestamp 1516238463
transform -1 0 5208 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_112
timestamp 1516238463
transform -1 0 5272 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_408
timestamp 1516238463
transform 1 0 5272 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_6
timestamp 1516238463
transform 1 0 5336 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_12
timestamp 1516238463
transform 1 0 5400 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_132
timestamp 1516238463
transform -1 0 5528 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_124
timestamp 1516238463
transform -1 0 5592 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_11
timestamp 1516238463
transform 1 0 5592 0 1 3010
box 0 0 64 200
use BUFX4  BUFX4_121
timestamp 1516238463
transform -1 0 5720 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_15
timestamp 1516238463
transform 1 0 5720 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_22
timestamp 1516238463
transform 1 0 5784 0 1 3010
box 0 0 64 200
use AND2X2  AND2X2_19
timestamp 1516238463
transform 1 0 5848 0 1 3010
box 0 0 64 200
use OR2X2  OR2X2_390
timestamp 1516238463
transform 1 0 5912 0 1 3010
box 0 0 64 200
use FILL  FILL_16_1
timestamp 1516238463
transform 1 0 5976 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_460
timestamp 1516238463
transform 1 0 8 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_314
timestamp 1516238463
transform -1 0 136 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_378
timestamp 1516238463
transform -1 0 200 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_360
timestamp 1516238463
transform -1 0 264 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_461
timestamp 1516238463
transform -1 0 328 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_527
timestamp 1516238463
transform -1 0 392 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_374
timestamp 1516238463
transform 1 0 392 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_339
timestamp 1516238463
transform 1 0 456 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_326
timestamp 1516238463
transform 1 0 520 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_433
timestamp 1516238463
transform 1 0 584 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_296
timestamp 1516238463
transform 1 0 648 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_327
timestamp 1516238463
transform 1 0 712 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_435
timestamp 1516238463
transform -1 0 840 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_340
timestamp 1516238463
transform 1 0 840 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_0_0
timestamp 1516238463
transform -1 0 920 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_1
timestamp 1516238463
transform -1 0 936 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_20
timestamp 1516238463
transform -1 0 1000 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_350
timestamp 1516238463
transform 1 0 1000 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_123
timestamp 1516238463
transform -1 0 1128 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_183
timestamp 1516238463
transform -1 0 1192 0 -1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_92
timestamp 1516238463
transform 1 0 1192 0 -1 3010
box 0 0 96 200
use OR2X2  OR2X2_395
timestamp 1516238463
transform -1 0 1352 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_351
timestamp 1516238463
transform 1 0 1352 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_394
timestamp 1516238463
transform -1 0 1480 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_21
timestamp 1516238463
transform 1 0 1480 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_67
timestamp 1516238463
transform -1 0 1608 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_153
timestamp 1516238463
transform -1 0 1672 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_492
timestamp 1516238463
transform -1 0 1736 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_236
timestamp 1516238463
transform -1 0 1800 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_22
timestamp 1516238463
transform -1 0 1864 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_422
timestamp 1516238463
transform 1 0 1864 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_1_0
timestamp 1516238463
transform 1 0 1928 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_1
timestamp 1516238463
transform 1 0 1944 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_394
timestamp 1516238463
transform 1 0 1960 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_199
timestamp 1516238463
transform -1 0 2088 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_138
timestamp 1516238463
transform -1 0 2152 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_269
timestamp 1516238463
transform -1 0 2216 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_44
timestamp 1516238463
transform -1 0 2280 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_395
timestamp 1516238463
transform -1 0 2344 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_172
timestamp 1516238463
transform 1 0 2344 0 -1 3010
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1516238463
transform -1 0 2536 0 -1 3010
box 0 0 128 200
use OR2X2  OR2X2_37
timestamp 1516238463
transform -1 0 2600 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_93
timestamp 1516238463
transform -1 0 2664 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_48
timestamp 1516238463
transform 1 0 2664 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_83
timestamp 1516238463
transform -1 0 2792 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_454
timestamp 1516238463
transform -1 0 2856 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_43
timestamp 1516238463
transform -1 0 2920 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_458
timestamp 1516238463
transform 1 0 2920 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_2_0
timestamp 1516238463
transform -1 0 3000 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_1
timestamp 1516238463
transform -1 0 3016 0 -1 3010
box 0 0 16 200
use OR2X2  OR2X2_246
timestamp 1516238463
transform -1 0 3080 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_357
timestamp 1516238463
transform -1 0 3144 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_282
timestamp 1516238463
transform -1 0 3208 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_55
timestamp 1516238463
transform -1 0 3272 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_38
timestamp 1516238463
transform -1 0 3336 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_279
timestamp 1516238463
transform -1 0 3400 0 -1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_17
timestamp 1516238463
transform 1 0 3400 0 -1 3010
box 0 0 96 200
use MUX2X1  MUX2X1_25
timestamp 1516238463
transform 1 0 3496 0 -1 3010
box 0 0 96 200
use OR2X2  OR2X2_232
timestamp 1516238463
transform -1 0 3656 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_89
timestamp 1516238463
transform -1 0 3720 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_182
timestamp 1516238463
transform -1 0 3784 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1516238463
transform 1 0 3784 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_42
timestamp 1516238463
transform 1 0 3848 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_449
timestamp 1516238463
transform -1 0 3976 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_3_0
timestamp 1516238463
transform -1 0 3992 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_3_1
timestamp 1516238463
transform -1 0 4008 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_12
timestamp 1516238463
transform -1 0 4072 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_179
timestamp 1516238463
transform -1 0 4136 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_312
timestamp 1516238463
transform -1 0 4200 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_110
timestamp 1516238463
transform 1 0 4200 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_215
timestamp 1516238463
transform -1 0 4328 0 -1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_1
timestamp 1516238463
transform -1 0 4424 0 -1 3010
box 0 0 96 200
use AND2X2  AND2X2_91
timestamp 1516238463
transform -1 0 4488 0 -1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_68
timestamp 1516238463
transform 1 0 4488 0 -1 3010
box 0 0 96 200
use OR2X2  OR2X2_146
timestamp 1516238463
transform -1 0 4648 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_201
timestamp 1516238463
transform -1 0 4712 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_235
timestamp 1516238463
transform -1 0 4776 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_135
timestamp 1516238463
transform -1 0 4840 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_212
timestamp 1516238463
transform -1 0 4904 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_224
timestamp 1516238463
transform -1 0 4968 0 -1 3010
box 0 0 64 200
use MUX2X1  MUX2X1_28
timestamp 1516238463
transform -1 0 5064 0 -1 3010
box 0 0 96 200
use FILL  FILL_14_4_0
timestamp 1516238463
transform 1 0 5064 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_4_1
timestamp 1516238463
transform 1 0 5080 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_31
timestamp 1516238463
transform 1 0 5096 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_23
timestamp 1516238463
transform 1 0 5160 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_334
timestamp 1516238463
transform 1 0 5224 0 -1 3010
box 0 0 64 200
use INVX1  INVX1_19
timestamp 1516238463
transform -1 0 5320 0 -1 3010
box 0 0 32 200
use MUX2X1  MUX2X1_61
timestamp 1516238463
transform 1 0 5320 0 -1 3010
box 0 0 96 200
use OR2X2  OR2X2_51
timestamp 1516238463
transform 1 0 5416 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_68
timestamp 1516238463
transform -1 0 5544 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_135
timestamp 1516238463
transform -1 0 5608 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_433
timestamp 1516238463
transform 1 0 5608 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_16
timestamp 1516238463
transform 1 0 5672 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_434
timestamp 1516238463
transform 1 0 5736 0 -1 3010
box 0 0 64 200
use OR2X2  OR2X2_437
timestamp 1516238463
transform 1 0 5800 0 -1 3010
box 0 0 64 200
use AND2X2  AND2X2_599
timestamp 1516238463
transform 1 0 5864 0 -1 3010
box 0 0 64 200
use FILL  FILL_15_1
timestamp 1516238463
transform -1 0 5944 0 -1 3010
box 0 0 16 200
use FILL  FILL_15_2
timestamp 1516238463
transform -1 0 5960 0 -1 3010
box 0 0 16 200
use FILL  FILL_15_3
timestamp 1516238463
transform -1 0 5976 0 -1 3010
box 0 0 16 200
use FILL  FILL_15_4
timestamp 1516238463
transform -1 0 5992 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_550
timestamp 1516238463
transform 1 0 8 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_400
timestamp 1516238463
transform 1 0 72 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_558
timestamp 1516238463
transform 1 0 136 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_503
timestamp 1516238463
transform -1 0 264 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_372
timestamp 1516238463
transform -1 0 328 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_405
timestamp 1516238463
transform 1 0 328 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_399
timestamp 1516238463
transform -1 0 456 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_304
timestamp 1516238463
transform 1 0 456 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_524
timestamp 1516238463
transform 1 0 520 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_298
timestamp 1516238463
transform -1 0 648 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_436
timestamp 1516238463
transform -1 0 712 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_547
timestamp 1516238463
transform 1 0 712 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_341
timestamp 1516238463
transform -1 0 840 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_13
timestamp 1516238463
transform 1 0 840 0 1 2610
box 0 0 64 200
use FILL  FILL_13_0_0
timestamp 1516238463
transform 1 0 904 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_1
timestamp 1516238463
transform 1 0 920 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_35
timestamp 1516238463
transform 1 0 936 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_285
timestamp 1516238463
transform 1 0 1000 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_420
timestamp 1516238463
transform 1 0 1064 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_411
timestamp 1516238463
transform -1 0 1192 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_48
timestamp 1516238463
transform 1 0 1192 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_388
timestamp 1516238463
transform 1 0 1256 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_320
timestamp 1516238463
transform -1 0 1384 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_497
timestamp 1516238463
transform -1 0 1448 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_68
timestamp 1516238463
transform 1 0 1448 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_356
timestamp 1516238463
transform -1 0 1576 0 1 2610
box 0 0 64 200
use AOI21X1  AOI21X1_25
timestamp 1516238463
transform 1 0 1576 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_65
timestamp 1516238463
transform 1 0 1640 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_154
timestamp 1516238463
transform -1 0 1768 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_264
timestamp 1516238463
transform -1 0 1832 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_174
timestamp 1516238463
transform -1 0 1896 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_256
timestamp 1516238463
transform 1 0 1896 0 1 2610
box 0 0 64 200
use FILL  FILL_13_1_0
timestamp 1516238463
transform -1 0 1976 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_1
timestamp 1516238463
transform -1 0 1992 0 1 2610
box 0 0 16 200
use AND2X2  AND2X2_382
timestamp 1516238463
transform -1 0 2056 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_258
timestamp 1516238463
transform 1 0 2056 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_139
timestamp 1516238463
transform 1 0 2120 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_396
timestamp 1516238463
transform 1 0 2184 0 1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_9
timestamp 1516238463
transform 1 0 2248 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_288
timestamp 1516238463
transform -1 0 2360 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_72
timestamp 1516238463
transform 1 0 2360 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_4
timestamp 1516238463
transform -1 0 2488 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_169
timestamp 1516238463
transform -1 0 2552 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_175
timestamp 1516238463
transform 1 0 2552 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_85
timestamp 1516238463
transform 1 0 2616 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_178
timestamp 1516238463
transform -1 0 2744 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_351
timestamp 1516238463
transform -1 0 2808 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_231
timestamp 1516238463
transform -1 0 2872 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_46
timestamp 1516238463
transform -1 0 2936 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_247
timestamp 1516238463
transform -1 0 3000 0 1 2610
box 0 0 64 200
use FILL  FILL_13_2_0
timestamp 1516238463
transform -1 0 3016 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_1
timestamp 1516238463
transform -1 0 3032 0 1 2610
box 0 0 16 200
use AND2X2  AND2X2_479
timestamp 1516238463
transform -1 0 3096 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_118
timestamp 1516238463
transform -1 0 3160 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_44
timestamp 1516238463
transform 1 0 3160 0 1 2610
box 0 0 48 200
use NOR2X1  NOR2X1_2
timestamp 1516238463
transform -1 0 3256 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_324
timestamp 1516238463
transform 1 0 3256 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_283
timestamp 1516238463
transform -1 0 3384 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_248
timestamp 1516238463
transform -1 0 3448 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_69
timestamp 1516238463
transform 1 0 3448 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_323
timestamp 1516238463
transform -1 0 3576 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_345
timestamp 1516238463
transform -1 0 3640 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_369
timestamp 1516238463
transform -1 0 3704 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_322
timestamp 1516238463
transform -1 0 3768 0 1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_7
timestamp 1516238463
transform -1 0 3816 0 1 2610
box 0 0 48 200
use AND2X2  AND2X2_86
timestamp 1516238463
transform 1 0 3816 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_47
timestamp 1516238463
transform 1 0 3880 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_246
timestamp 1516238463
transform -1 0 4008 0 1 2610
box 0 0 64 200
use FILL  FILL_13_3_0
timestamp 1516238463
transform 1 0 4008 0 1 2610
box 0 0 16 200
use FILL  FILL_13_3_1
timestamp 1516238463
transform 1 0 4024 0 1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_50
timestamp 1516238463
transform 1 0 4040 0 1 2610
box 0 0 96 200
use BUFX4  BUFX4_15
timestamp 1516238463
transform -1 0 4200 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_16
timestamp 1516238463
transform 1 0 4200 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_150
timestamp 1516238463
transform -1 0 4328 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_67
timestamp 1516238463
transform -1 0 4392 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_622
timestamp 1516238463
transform -1 0 4456 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_623
timestamp 1516238463
transform -1 0 4520 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_626
timestamp 1516238463
transform 1 0 4520 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_92
timestamp 1516238463
transform 1 0 4584 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_23
timestamp 1516238463
transform -1 0 4712 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_93
timestamp 1516238463
transform -1 0 4776 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_9
timestamp 1516238463
transform -1 0 4840 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_196
timestamp 1516238463
transform 1 0 4840 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_427
timestamp 1516238463
transform -1 0 4968 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_630
timestamp 1516238463
transform -1 0 5032 0 1 2610
box 0 0 64 200
use FILL  FILL_13_4_0
timestamp 1516238463
transform -1 0 5048 0 1 2610
box 0 0 16 200
use FILL  FILL_13_4_1
timestamp 1516238463
transform -1 0 5064 0 1 2610
box 0 0 16 200
use OR2X2  OR2X2_367
timestamp 1516238463
transform -1 0 5128 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_633
timestamp 1516238463
transform -1 0 5192 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_163
timestamp 1516238463
transform 1 0 5192 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_35
timestamp 1516238463
transform -1 0 5320 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_334
timestamp 1516238463
transform 1 0 5320 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_134
timestamp 1516238463
transform -1 0 5448 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_68
timestamp 1516238463
transform -1 0 5512 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_104
timestamp 1516238463
transform -1 0 5576 0 1 2610
box 0 0 64 200
use MUX2X1  MUX2X1_66
timestamp 1516238463
transform -1 0 5672 0 1 2610
box 0 0 96 200
use AND2X2  AND2X2_20
timestamp 1516238463
transform 1 0 5672 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_613
timestamp 1516238463
transform 1 0 5736 0 1 2610
box 0 0 64 200
use OR2X2  OR2X2_436
timestamp 1516238463
transform 1 0 5800 0 1 2610
box 0 0 64 200
use AND2X2  AND2X2_602
timestamp 1516238463
transform -1 0 5928 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_117
timestamp 1516238463
transform -1 0 5992 0 1 2610
box 0 0 64 200
use BUFX4  BUFX4_71
timestamp 1516238463
transform 1 0 8 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_70
timestamp 1516238463
transform 1 0 72 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_361
timestamp 1516238463
transform -1 0 200 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_366
timestamp 1516238463
transform -1 0 264 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_248
timestamp 1516238463
transform 1 0 264 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_125
timestamp 1516238463
transform 1 0 328 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_274
timestamp 1516238463
transform 1 0 392 0 -1 2610
box 0 0 64 200
use INVX4  INVX4_2
timestamp 1516238463
transform -1 0 504 0 -1 2610
box 0 0 48 200
use OR2X2  OR2X2_186
timestamp 1516238463
transform 1 0 504 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_297
timestamp 1516238463
transform 1 0 568 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_298
timestamp 1516238463
transform 1 0 632 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_437
timestamp 1516238463
transform -1 0 760 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_219
timestamp 1516238463
transform -1 0 824 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_336
timestamp 1516238463
transform -1 0 888 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_69
timestamp 1516238463
transform -1 0 952 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_0_0
timestamp 1516238463
transform 1 0 952 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_1
timestamp 1516238463
transform 1 0 968 0 -1 2610
box 0 0 16 200
use OR2X2  OR2X2_286
timestamp 1516238463
transform 1 0 984 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_421
timestamp 1516238463
transform -1 0 1112 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_287
timestamp 1516238463
transform 1 0 1112 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_45
timestamp 1516238463
transform -1 0 1240 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_321
timestamp 1516238463
transform 1 0 1240 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_200
timestamp 1516238463
transform 1 0 1304 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_358
timestamp 1516238463
transform -1 0 1432 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_237
timestamp 1516238463
transform -1 0 1496 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_305
timestamp 1516238463
transform 1 0 1496 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_306
timestamp 1516238463
transform 1 0 1560 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_450
timestamp 1516238463
transform -1 0 1688 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_94
timestamp 1516238463
transform -1 0 1752 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_205
timestamp 1516238463
transform -1 0 1816 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_115
timestamp 1516238463
transform 1 0 1816 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_239
timestamp 1516238463
transform 1 0 1880 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_1_0
timestamp 1516238463
transform 1 0 1944 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_1
timestamp 1516238463
transform 1 0 1960 0 -1 2610
box 0 0 16 200
use OR2X2  OR2X2_262
timestamp 1516238463
transform 1 0 1976 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_15
timestamp 1516238463
transform 1 0 2040 0 -1 2610
box 0 0 64 200
use INVX1  INVX1_26
timestamp 1516238463
transform -1 0 2136 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_11
timestamp 1516238463
transform -1 0 2200 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_270
timestamp 1516238463
transform 1 0 2200 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_233
timestamp 1516238463
transform -1 0 2328 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_67
timestamp 1516238463
transform 1 0 2328 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_134
timestamp 1516238463
transform 1 0 2392 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_39
timestamp 1516238463
transform 1 0 2456 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_136
timestamp 1516238463
transform 1 0 2520 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_1
timestamp 1516238463
transform -1 0 2648 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1516238463
transform 1 0 2648 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_204
timestamp 1516238463
transform -1 0 2776 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_167
timestamp 1516238463
transform -1 0 2840 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_166
timestamp 1516238463
transform -1 0 2904 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_401
timestamp 1516238463
transform 1 0 2904 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_2_0
timestamp 1516238463
transform 1 0 2968 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_1
timestamp 1516238463
transform 1 0 2984 0 -1 2610
box 0 0 16 200
use OR2X2  OR2X2_290
timestamp 1516238463
transform 1 0 3000 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_56
timestamp 1516238463
transform -1 0 3128 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_7
timestamp 1516238463
transform 1 0 3128 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_460
timestamp 1516238463
transform -1 0 3256 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_203
timestamp 1516238463
transform -1 0 3320 0 -1 2610
box 0 0 64 200
use MUX2X1  MUX2X1_26
timestamp 1516238463
transform -1 0 3416 0 -1 2610
box 0 0 96 200
use OR2X2  OR2X2_450
timestamp 1516238463
transform 1 0 3416 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_190
timestamp 1516238463
transform -1 0 3544 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_62
timestamp 1516238463
transform -1 0 3608 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_42
timestamp 1516238463
transform 1 0 3608 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_10
timestamp 1516238463
transform -1 0 3736 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_271
timestamp 1516238463
transform 1 0 3736 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_156
timestamp 1516238463
transform -1 0 3864 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_272
timestamp 1516238463
transform -1 0 3928 0 -1 2610
box 0 0 64 200
use MUX2X1  MUX2X1_45
timestamp 1516238463
transform -1 0 4024 0 -1 2610
box 0 0 96 200
use FILL  FILL_12_3_0
timestamp 1516238463
transform -1 0 4040 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_3_1
timestamp 1516238463
transform -1 0 4056 0 -1 2610
box 0 0 16 200
use OR2X2  OR2X2_63
timestamp 1516238463
transform -1 0 4120 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_151
timestamp 1516238463
transform -1 0 4184 0 -1 2610
box 0 0 64 200
use MUX2X1  MUX2X1_46
timestamp 1516238463
transform 1 0 4184 0 -1 2610
box 0 0 96 200
use NAND2X1  NAND2X1_18
timestamp 1516238463
transform 1 0 4280 0 -1 2610
box 0 0 48 200
use OR2X2  OR2X2_417
timestamp 1516238463
transform -1 0 4392 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_25
timestamp 1516238463
transform -1 0 4456 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_94
timestamp 1516238463
transform -1 0 4520 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_418
timestamp 1516238463
transform -1 0 4584 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_625
timestamp 1516238463
transform -1 0 4648 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_217
timestamp 1516238463
transform 1 0 4648 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_50
timestamp 1516238463
transform -1 0 4776 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_557
timestamp 1516238463
transform 1 0 4776 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_357
timestamp 1516238463
transform -1 0 4904 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_74
timestamp 1516238463
transform -1 0 4968 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_98
timestamp 1516238463
transform 1 0 4968 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_4_0
timestamp 1516238463
transform -1 0 5048 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_4_1
timestamp 1516238463
transform -1 0 5064 0 -1 2610
box 0 0 16 200
use AND2X2  AND2X2_197
timestamp 1516238463
transform -1 0 5128 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_590
timestamp 1516238463
transform -1 0 5192 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_46
timestamp 1516238463
transform -1 0 5256 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_43
timestamp 1516238463
transform -1 0 5320 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_52
timestamp 1516238463
transform -1 0 5384 0 -1 2610
box 0 0 64 200
use AND2X2  AND2X2_131
timestamp 1516238463
transform -1 0 5448 0 -1 2610
box 0 0 64 200
use MUX2X1  MUX2X1_72
timestamp 1516238463
transform 1 0 5448 0 -1 2610
box 0 0 96 200
use MUX2X1  MUX2X1_67
timestamp 1516238463
transform 1 0 5544 0 -1 2610
box 0 0 96 200
use BUFX4  BUFX4_45
timestamp 1516238463
transform -1 0 5704 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_9
timestamp 1516238463
transform -1 0 5768 0 -1 2610
box 0 0 64 200
use BUFX4  BUFX4_41
timestamp 1516238463
transform 1 0 5768 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_2
timestamp 1516238463
transform 1 0 5832 0 -1 2610
box 0 0 64 200
use OR2X2  OR2X2_54
timestamp 1516238463
transform 1 0 5896 0 -1 2610
box 0 0 64 200
use FILL  FILL_13_1
timestamp 1516238463
transform -1 0 5976 0 -1 2610
box 0 0 16 200
use FILL  FILL_13_2
timestamp 1516238463
transform -1 0 5992 0 -1 2610
box 0 0 16 200
use AND2X2  AND2X2_462
timestamp 1516238463
transform -1 0 72 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_533
timestamp 1516238463
transform -1 0 136 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_509
timestamp 1516238463
transform -1 0 200 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_403
timestamp 1516238463
transform 1 0 200 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_402
timestamp 1516238463
transform -1 0 328 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_559
timestamp 1516238463
transform -1 0 392 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_29
timestamp 1516238463
transform 1 0 392 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_406
timestamp 1516238463
transform 1 0 456 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_356
timestamp 1516238463
transform -1 0 584 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_525
timestamp 1516238463
transform 1 0 584 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_423
timestamp 1516238463
transform 1 0 648 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_19
timestamp 1516238463
transform 1 0 712 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_396
timestamp 1516238463
transform 1 0 776 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_486
timestamp 1516238463
transform -1 0 904 0 1 2210
box 0 0 64 200
use FILL  FILL_11_0_0
timestamp 1516238463
transform -1 0 920 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1516238463
transform -1 0 936 0 1 2210
box 0 0 16 200
use OR2X2  OR2X2_336
timestamp 1516238463
transform -1 0 1000 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_21
timestamp 1516238463
transform 1 0 1000 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_47
timestamp 1516238463
transform 1 0 1064 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_498
timestamp 1516238463
transform -1 0 1192 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_491
timestamp 1516238463
transform -1 0 1256 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_344
timestamp 1516238463
transform -1 0 1320 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_363
timestamp 1516238463
transform 1 0 1320 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_22
timestamp 1516238463
transform 1 0 1384 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_202
timestamp 1516238463
transform 1 0 1448 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_173
timestamp 1516238463
transform 1 0 1512 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_30
timestamp 1516238463
transform 1 0 1576 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_364
timestamp 1516238463
transform -1 0 1704 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_292
timestamp 1516238463
transform 1 0 1704 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_206
timestamp 1516238463
transform 1 0 1768 0 1 2210
box 0 0 64 200
use INVX8  INVX8_1
timestamp 1516238463
transform 1 0 1832 0 1 2210
box 0 0 80 200
use AND2X2  AND2X2_326
timestamp 1516238463
transform 1 0 1912 0 1 2210
box 0 0 64 200
use FILL  FILL_11_1_0
timestamp 1516238463
transform 1 0 1976 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1516238463
transform 1 0 1992 0 1 2210
box 0 0 16 200
use AND2X2  AND2X2_327
timestamp 1516238463
transform 1 0 2008 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_328
timestamp 1516238463
transform 1 0 2072 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_155
timestamp 1516238463
transform 1 0 2136 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_95
timestamp 1516238463
transform 1 0 2200 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_362
timestamp 1516238463
transform 1 0 2264 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_293
timestamp 1516238463
transform 1 0 2328 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_5
timestamp 1516238463
transform 1 0 2392 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_192
timestamp 1516238463
transform 1 0 2456 0 1 2210
box 0 0 64 200
use AOI22X1  AOI22X1_1
timestamp 1516238463
transform -1 0 2600 0 1 2210
box 0 0 80 200
use NAND2X1  NAND2X1_76
timestamp 1516238463
transform -1 0 2648 0 1 2210
box 0 0 48 200
use AND2X2  AND2X2_258
timestamp 1516238463
transform 1 0 2648 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_397
timestamp 1516238463
transform 1 0 2712 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_393
timestamp 1516238463
transform -1 0 2840 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_267
timestamp 1516238463
transform -1 0 2904 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_221
timestamp 1516238463
transform -1 0 2968 0 1 2210
box 0 0 64 200
use FILL  FILL_11_2_0
timestamp 1516238463
transform -1 0 2984 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1516238463
transform -1 0 3000 0 1 2210
box 0 0 16 200
use AND2X2  AND2X2_193
timestamp 1516238463
transform -1 0 3064 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_12
timestamp 1516238463
transform 1 0 3064 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_60
timestamp 1516238463
transform 1 0 3128 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_14
timestamp 1516238463
transform 1 0 3192 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_459
timestamp 1516238463
transform 1 0 3256 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_61
timestamp 1516238463
transform 1 0 3320 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_91
timestamp 1516238463
transform -1 0 3448 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_62
timestamp 1516238463
transform 1 0 3448 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_66
timestamp 1516238463
transform 1 0 3512 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_149
timestamp 1516238463
transform 1 0 3576 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_64
timestamp 1516238463
transform -1 0 3704 0 1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_30
timestamp 1516238463
transform 1 0 3704 0 1 2210
box 0 0 96 200
use OR2X2  OR2X2_420
timestamp 1516238463
transform 1 0 3800 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_627
timestamp 1516238463
transform 1 0 3864 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_24
timestamp 1516238463
transform 1 0 3928 0 1 2210
box 0 0 64 200
use FILL  FILL_11_3_0
timestamp 1516238463
transform -1 0 4008 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_1
timestamp 1516238463
transform -1 0 4024 0 1 2210
box 0 0 16 200
use AND2X2  AND2X2_152
timestamp 1516238463
transform -1 0 4088 0 1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_47
timestamp 1516238463
transform -1 0 4184 0 1 2210
box 0 0 96 200
use OR2X2  OR2X2_214
timestamp 1516238463
transform 1 0 4184 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_35
timestamp 1516238463
transform -1 0 4296 0 1 2210
box 0 0 48 200
use AOI21X1  AOI21X1_5
timestamp 1516238463
transform -1 0 4360 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_19
timestamp 1516238463
transform -1 0 4408 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_75
timestamp 1516238463
transform 1 0 4408 0 1 2210
box 0 0 48 200
use AND2X2  AND2X2_147
timestamp 1516238463
transform 1 0 4456 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_148
timestamp 1516238463
transform -1 0 4584 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_612
timestamp 1516238463
transform 1 0 4584 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_411
timestamp 1516238463
transform -1 0 4712 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_616
timestamp 1516238463
transform -1 0 4776 0 1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_41
timestamp 1516238463
transform 1 0 4776 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_410
timestamp 1516238463
transform -1 0 4904 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_615
timestamp 1516238463
transform -1 0 4968 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_222
timestamp 1516238463
transform -1 0 5032 0 1 2210
box 0 0 64 200
use FILL  FILL_11_4_0
timestamp 1516238463
transform -1 0 5048 0 1 2210
box 0 0 16 200
use FILL  FILL_11_4_1
timestamp 1516238463
transform -1 0 5064 0 1 2210
box 0 0 16 200
use OR2X2  OR2X2_409
timestamp 1516238463
transform -1 0 5128 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_610
timestamp 1516238463
transform -1 0 5192 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_103
timestamp 1516238463
transform -1 0 5256 0 1 2210
box 0 0 64 200
use OR2X2  OR2X2_441
timestamp 1516238463
transform 1 0 5256 0 1 2210
box 0 0 64 200
use XOR2X1  XOR2X1_5
timestamp 1516238463
transform -1 0 5432 0 1 2210
box 0 0 112 200
use MUX2X1  MUX2X1_24
timestamp 1516238463
transform -1 0 5528 0 1 2210
box 0 0 96 200
use BUFX4  BUFX4_5
timestamp 1516238463
transform 1 0 5528 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_73
timestamp 1516238463
transform 1 0 5592 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_74
timestamp 1516238463
transform -1 0 5720 0 1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_27
timestamp 1516238463
transform -1 0 5816 0 1 2210
box 0 0 96 200
use BUFX4  BUFX4_4
timestamp 1516238463
transform 1 0 5816 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_139
timestamp 1516238463
transform 1 0 5880 0 1 2210
box 0 0 64 200
use FILL  FILL_12_1
timestamp 1516238463
transform 1 0 5944 0 1 2210
box 0 0 16 200
use FILL  FILL_12_2
timestamp 1516238463
transform 1 0 5960 0 1 2210
box 0 0 16 200
use FILL  FILL_12_3
timestamp 1516238463
transform 1 0 5976 0 1 2210
box 0 0 16 200
use INVX1  INVX1_17
timestamp 1516238463
transform 1 0 8 0 -1 2210
box 0 0 32 200
use NAND3X1  NAND3X1_40
timestamp 1516238463
transform -1 0 104 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_38
timestamp 1516238463
transform -1 0 168 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_49
timestamp 1516238463
transform -1 0 232 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_58
timestamp 1516238463
transform 1 0 232 0 -1 2210
box 0 0 48 200
use OR2X2  OR2X2_321
timestamp 1516238463
transform 1 0 280 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_50
timestamp 1516238463
transform -1 0 408 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_380
timestamp 1516238463
transform 1 0 408 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_381
timestamp 1516238463
transform 1 0 472 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_316
timestamp 1516238463
transform 1 0 536 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_315
timestamp 1516238463
transform -1 0 664 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_463
timestamp 1516238463
transform -1 0 728 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_526
timestamp 1516238463
transform -1 0 792 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_328
timestamp 1516238463
transform 1 0 792 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_187
timestamp 1516238463
transform 1 0 856 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_0_0
timestamp 1516238463
transform 1 0 920 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1516238463
transform 1 0 936 0 -1 2210
box 0 0 16 200
use OR2X2  OR2X2_70
timestamp 1516238463
transform 1 0 952 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_475
timestamp 1516238463
transform 1 0 1016 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_126
timestamp 1516238463
transform 1 0 1080 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_329
timestamp 1516238463
transform -1 0 1208 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_489
timestamp 1516238463
transform -1 0 1272 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_249
timestamp 1516238463
transform 1 0 1272 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_517
timestamp 1516238463
transform -1 0 1400 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_385
timestamp 1516238463
transform 1 0 1400 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_238
timestamp 1516238463
transform 1 0 1464 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_220
timestamp 1516238463
transform 1 0 1528 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_516
timestamp 1516238463
transform -1 0 1656 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_342
timestamp 1516238463
transform -1 0 1720 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_291
timestamp 1516238463
transform -1 0 1784 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_175
timestamp 1516238463
transform -1 0 1848 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_386
timestamp 1516238463
transform -1 0 1912 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_240
timestamp 1516238463
transform 1 0 1912 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_1_0
timestamp 1516238463
transform 1 0 1976 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1516238463
transform 1 0 1992 0 -1 2210
box 0 0 16 200
use AND2X2  AND2X2_360
timestamp 1516238463
transform 1 0 2008 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_361
timestamp 1516238463
transform 1 0 2072 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_201
timestamp 1516238463
transform 1 0 2136 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_253
timestamp 1516238463
transform 1 0 2200 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_140
timestamp 1516238463
transform 1 0 2264 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_256
timestamp 1516238463
transform 1 0 2328 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_275
timestamp 1516238463
transform 1 0 2392 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_16
timestamp 1516238463
transform -1 0 2520 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_2
timestamp 1516238463
transform 1 0 2520 0 -1 2210
box 0 0 32 200
use AOI22X1  AOI22X1_2
timestamp 1516238463
transform -1 0 2632 0 -1 2210
box 0 0 80 200
use NAND3X1  NAND3X1_3
timestamp 1516238463
transform 1 0 2632 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_302
timestamp 1516238463
transform -1 0 2760 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_86
timestamp 1516238463
transform 1 0 2760 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_141
timestamp 1516238463
transform -1 0 2888 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_23
timestamp 1516238463
transform -1 0 2952 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_2_0
timestamp 1516238463
transform 1 0 2952 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1516238463
transform 1 0 2968 0 -1 2210
box 0 0 16 200
use AND2X2  AND2X2_194
timestamp 1516238463
transform 1 0 2984 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_11
timestamp 1516238463
transform -1 0 3096 0 -1 2210
box 0 0 48 200
use AND2X2  AND2X2_98
timestamp 1516238463
transform -1 0 3160 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_18
timestamp 1516238463
transform 1 0 3160 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_106
timestamp 1516238463
transform 1 0 3224 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_20
timestamp 1516238463
transform -1 0 3352 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_274
timestamp 1516238463
transform 1 0 3352 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_159
timestamp 1516238463
transform -1 0 3480 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_275
timestamp 1516238463
transform 1 0 3480 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_64
timestamp 1516238463
transform -1 0 3608 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_32
timestamp 1516238463
transform 1 0 3608 0 -1 2210
box 0 0 96 200
use OR2X2  OR2X2_158
timestamp 1516238463
transform -1 0 3768 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_33
timestamp 1516238463
transform 1 0 3768 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_31
timestamp 1516238463
transform 1 0 3864 0 -1 2210
box 0 0 96 200
use FILL  FILL_10_3_0
timestamp 1516238463
transform -1 0 3976 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_3_1
timestamp 1516238463
transform -1 0 3992 0 -1 2210
box 0 0 16 200
use MUX2X1  MUX2X1_38
timestamp 1516238463
transform -1 0 4088 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_37
timestamp 1516238463
transform 1 0 4088 0 -1 2210
box 0 0 96 200
use OR2X2  OR2X2_111
timestamp 1516238463
transform -1 0 4248 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_39
timestamp 1516238463
transform -1 0 4312 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_34
timestamp 1516238463
transform -1 0 4408 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_35
timestamp 1516238463
transform 1 0 4408 0 -1 2210
box 0 0 96 200
use AND2X2  AND2X2_333
timestamp 1516238463
transform -1 0 4568 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_61
timestamp 1516238463
transform 1 0 4568 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_215
timestamp 1516238463
transform 1 0 4632 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_13
timestamp 1516238463
transform 1 0 4696 0 -1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_33
timestamp 1516238463
transform 1 0 4744 0 -1 2210
box 0 0 48 200
use OR2X2  OR2X2_116
timestamp 1516238463
transform -1 0 4856 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_614
timestamp 1516238463
transform 1 0 4856 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_57
timestamp 1516238463
transform 1 0 4920 0 -1 2210
box 0 0 96 200
use FILL  FILL_10_4_0
timestamp 1516238463
transform 1 0 5016 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_4_1
timestamp 1516238463
transform 1 0 5032 0 -1 2210
box 0 0 16 200
use MUX2X1  MUX2X1_59
timestamp 1516238463
transform 1 0 5048 0 -1 2210
box 0 0 96 200
use AND2X2  AND2X2_611
timestamp 1516238463
transform -1 0 5208 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_58
timestamp 1516238463
transform -1 0 5304 0 -1 2210
box 0 0 96 200
use AND2X2  AND2X2_220
timestamp 1516238463
transform -1 0 5368 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_112
timestamp 1516238463
transform -1 0 5432 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_219
timestamp 1516238463
transform 1 0 5432 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_115
timestamp 1516238463
transform -1 0 5560 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_218
timestamp 1516238463
transform -1 0 5624 0 -1 2210
box 0 0 64 200
use OR2X2  OR2X2_11
timestamp 1516238463
transform -1 0 5688 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_29
timestamp 1516238463
transform 1 0 5688 0 -1 2210
box 0 0 96 200
use NAND2X1  NAND2X1_45
timestamp 1516238463
transform 1 0 5784 0 -1 2210
box 0 0 48 200
use XOR2X1  XOR2X1_2
timestamp 1516238463
transform 1 0 5832 0 -1 2210
box 0 0 112 200
use FILL  FILL_11_1
timestamp 1516238463
transform -1 0 5960 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_2
timestamp 1516238463
transform -1 0 5976 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_3
timestamp 1516238463
transform -1 0 5992 0 -1 2210
box 0 0 16 200
use INVX1  INVX1_18
timestamp 1516238463
transform 1 0 8 0 1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_36
timestamp 1516238463
transform 1 0 40 0 1 1810
box 0 0 48 200
use AND2X2  AND2X2_373
timestamp 1516238463
transform 1 0 88 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_8
timestamp 1516238463
transform 1 0 152 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_13
timestamp 1516238463
transform 1 0 216 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_59
timestamp 1516238463
transform -1 0 328 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_28
timestamp 1516238463
transform 1 0 328 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_466
timestamp 1516238463
transform 1 0 392 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_57
timestamp 1516238463
transform 1 0 456 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_561
timestamp 1516238463
transform 1 0 520 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_499
timestamp 1516238463
transform 1 0 584 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_355
timestamp 1516238463
transform -1 0 712 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_66
timestamp 1516238463
transform -1 0 760 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_24
timestamp 1516238463
transform 1 0 760 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_464
timestamp 1516238463
transform 1 0 824 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_454
timestamp 1516238463
transform -1 0 952 0 1 1810
box 0 0 64 200
use FILL  FILL_9_0_0
timestamp 1516238463
transform -1 0 968 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1516238463
transform -1 0 984 0 1 1810
box 0 0 16 200
use AND2X2  AND2X2_476
timestamp 1516238463
transform -1 0 1048 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_31
timestamp 1516238463
transform -1 0 1112 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_310
timestamp 1516238463
transform 1 0 1112 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_549
timestamp 1516238463
transform -1 0 1240 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_548
timestamp 1516238463
transform -1 0 1304 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_126
timestamp 1516238463
transform 1 0 1304 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_376
timestamp 1516238463
transform 1 0 1368 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_542
timestamp 1516238463
transform -1 0 1496 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_541
timestamp 1516238463
transform -1 0 1560 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_438
timestamp 1516238463
transform 1 0 1560 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_428
timestamp 1516238463
transform -1 0 1688 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_63
timestamp 1516238463
transform -1 0 1752 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_377
timestamp 1516238463
transform 1 0 1752 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_56
timestamp 1516238463
transform 1 0 1816 0 1 1810
box 0 0 48 200
use AND2X2  AND2X2_469
timestamp 1516238463
transform -1 0 1928 0 1 1810
box 0 0 64 200
use FILL  FILL_9_1_0
timestamp 1516238463
transform -1 0 1944 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1516238463
transform -1 0 1960 0 1 1810
box 0 0 16 200
use OR2X2  OR2X2_293
timestamp 1516238463
transform -1 0 2024 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_309
timestamp 1516238463
transform -1 0 2088 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_105
timestamp 1516238463
transform -1 0 2152 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_65
timestamp 1516238463
transform 1 0 2152 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_159
timestamp 1516238463
transform 1 0 2216 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_160
timestamp 1516238463
transform 1 0 2280 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_103
timestamp 1516238463
transform 1 0 2344 0 1 1810
box 0 0 64 200
use INVX2  INVX2_4
timestamp 1516238463
transform -1 0 2440 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_451
timestamp 1516238463
transform 1 0 2440 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_441
timestamp 1516238463
transform -1 0 2568 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_161
timestamp 1516238463
transform 1 0 2568 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_2
timestamp 1516238463
transform -1 0 2696 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_490
timestamp 1516238463
transform 1 0 2696 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_191
timestamp 1516238463
transform -1 0 2824 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_16
timestamp 1516238463
transform 1 0 2824 0 1 1810
box 0 0 64 200
use INVX1  INVX1_23
timestamp 1516238463
transform -1 0 2920 0 1 1810
box 0 0 32 200
use AND2X2  AND2X2_512
timestamp 1516238463
transform 1 0 2920 0 1 1810
box 0 0 64 200
use FILL  FILL_9_2_0
timestamp 1516238463
transform -1 0 3000 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1516238463
transform -1 0 3016 0 1 1810
box 0 0 16 200
use OR2X2  OR2X2_312
timestamp 1516238463
transform -1 0 3080 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_255
timestamp 1516238463
transform -1 0 3144 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_2
timestamp 1516238463
transform 1 0 3144 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_104
timestamp 1516238463
transform -1 0 3272 0 1 1810
box 0 0 64 200
use INVX1  INVX1_25
timestamp 1516238463
transform 1 0 3272 0 1 1810
box 0 0 32 200
use BUFX4  BUFX4_108
timestamp 1516238463
transform 1 0 3304 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_332
timestamp 1516238463
transform -1 0 3432 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_212
timestamp 1516238463
transform 1 0 3432 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_523
timestamp 1516238463
transform 1 0 3496 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_216
timestamp 1516238463
transform -1 0 3624 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_18
timestamp 1516238463
transform 1 0 3624 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_127
timestamp 1516238463
transform 1 0 3688 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_276
timestamp 1516238463
transform -1 0 3816 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_87
timestamp 1516238463
transform 1 0 3816 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_319
timestamp 1516238463
transform -1 0 3944 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_388
timestamp 1516238463
transform -1 0 4008 0 1 1810
box 0 0 64 200
use FILL  FILL_9_3_0
timestamp 1516238463
transform -1 0 4024 0 1 1810
box 0 0 16 200
use FILL  FILL_9_3_1
timestamp 1516238463
transform -1 0 4040 0 1 1810
box 0 0 16 200
use INVX2  INVX2_2
timestamp 1516238463
transform -1 0 4072 0 1 1810
box 0 0 32 200
use XOR2X1  XOR2X1_7
timestamp 1516238463
transform 1 0 4072 0 1 1810
box 0 0 112 200
use OR2X2  OR2X2_151
timestamp 1516238463
transform -1 0 4248 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_34
timestamp 1516238463
transform -1 0 4312 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_145
timestamp 1516238463
transform -1 0 4376 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_150
timestamp 1516238463
transform -1 0 4440 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_221
timestamp 1516238463
transform -1 0 4504 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_263
timestamp 1516238463
transform -1 0 4568 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_617
timestamp 1516238463
transform -1 0 4632 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_42
timestamp 1516238463
transform -1 0 4728 0 1 1810
box 0 0 96 200
use AND2X2  AND2X2_228
timestamp 1516238463
transform 1 0 4728 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_227
timestamp 1516238463
transform -1 0 4856 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_226
timestamp 1516238463
transform -1 0 4920 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_117
timestamp 1516238463
transform -1 0 4984 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_225
timestamp 1516238463
transform -1 0 5048 0 1 1810
box 0 0 64 200
use FILL  FILL_9_4_0
timestamp 1516238463
transform 1 0 5048 0 1 1810
box 0 0 16 200
use FILL  FILL_9_4_1
timestamp 1516238463
transform 1 0 5064 0 1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_36
timestamp 1516238463
transform 1 0 5080 0 1 1810
box 0 0 96 200
use OR2X2  OR2X2_73
timestamp 1516238463
transform -1 0 5240 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_70
timestamp 1516238463
transform 1 0 5240 0 1 1810
box 0 0 96 200
use AND2X2  AND2X2_164
timestamp 1516238463
transform -1 0 5400 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_105
timestamp 1516238463
transform 1 0 5400 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_52
timestamp 1516238463
transform 1 0 5464 0 1 1810
box 0 0 96 200
use AND2X2  AND2X2_204
timestamp 1516238463
transform -1 0 5624 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_207
timestamp 1516238463
transform 1 0 5624 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_208
timestamp 1516238463
transform -1 0 5752 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_603
timestamp 1516238463
transform 1 0 5752 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_206
timestamp 1516238463
transform -1 0 5880 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_141
timestamp 1516238463
transform 1 0 5880 0 1 1810
box 0 0 64 200
use FILL  FILL_10_1
timestamp 1516238463
transform 1 0 5944 0 1 1810
box 0 0 16 200
use FILL  FILL_10_2
timestamp 1516238463
transform 1 0 5960 0 1 1810
box 0 0 16 200
use FILL  FILL_10_3
timestamp 1516238463
transform 1 0 5976 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_71
timestamp 1516238463
transform 1 0 8 0 -1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_7
timestamp 1516238463
transform -1 0 104 0 -1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_37
timestamp 1516238463
transform -1 0 168 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_42
timestamp 1516238463
transform -1 0 200 0 -1 1810
box 0 0 32 200
use OR2X2  OR2X2_343
timestamp 1516238463
transform 1 0 200 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_488
timestamp 1516238463
transform 1 0 264 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_47
timestamp 1516238463
transform -1 0 392 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_310
timestamp 1516238463
transform 1 0 392 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_330
timestamp 1516238463
transform 1 0 456 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_453
timestamp 1516238463
transform 1 0 520 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_48
timestamp 1516238463
transform -1 0 648 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_55
timestamp 1516238463
transform -1 0 696 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_55
timestamp 1516238463
transform -1 0 760 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_32
timestamp 1516238463
transform 1 0 760 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_560
timestamp 1516238463
transform -1 0 888 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1516238463
transform 1 0 888 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_0_0
timestamp 1516238463
transform -1 0 968 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1516238463
transform -1 0 984 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_85
timestamp 1516238463
transform -1 0 1048 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_48
timestamp 1516238463
transform -1 0 1112 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_125
timestamp 1516238463
transform 1 0 1112 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_27
timestamp 1516238463
transform 1 0 1176 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_33
timestamp 1516238463
transform 1 0 1240 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_375
timestamp 1516238463
transform 1 0 1304 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_309
timestamp 1516238463
transform -1 0 1432 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_308
timestamp 1516238463
transform -1 0 1496 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_354
timestamp 1516238463
transform -1 0 1560 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_192
timestamp 1516238463
transform -1 0 1624 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_19
timestamp 1516238463
transform -1 0 1688 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_28
timestamp 1516238463
transform 1 0 1688 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_25
timestamp 1516238463
transform 1 0 1752 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_64
timestamp 1516238463
transform -1 0 1880 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_467
timestamp 1516238463
transform -1 0 1944 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_1_0
timestamp 1516238463
transform -1 0 1960 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1516238463
transform -1 0 1976 0 -1 1810
box 0 0 16 200
use OR2X2  OR2X2_320
timestamp 1516238463
transform -1 0 2040 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_301
timestamp 1516238463
transform -1 0 2104 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_383
timestamp 1516238463
transform 1 0 2104 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_259
timestamp 1516238463
transform 1 0 2168 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_142
timestamp 1516238463
transform 1 0 2232 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_255
timestamp 1516238463
transform 1 0 2296 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_1
timestamp 1516238463
transform -1 0 2424 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_1
timestamp 1516238463
transform 1 0 2424 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_52
timestamp 1516238463
transform 1 0 2488 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_36
timestamp 1516238463
transform -1 0 2616 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_20
timestamp 1516238463
transform -1 0 2680 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_384
timestamp 1516238463
transform 1 0 2680 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_501
timestamp 1516238463
transform 1 0 2744 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_13
timestamp 1516238463
transform -1 0 2872 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_380
timestamp 1516238463
transform -1 0 2936 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_24
timestamp 1516238463
transform 1 0 2936 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_2_0
timestamp 1516238463
transform 1 0 3000 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1516238463
transform 1 0 3016 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_24
timestamp 1516238463
transform 1 0 3032 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_273
timestamp 1516238463
transform 1 0 3096 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_160
timestamp 1516238463
transform -1 0 3224 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_216
timestamp 1516238463
transform -1 0 3288 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_389
timestamp 1516238463
transform 1 0 3288 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_264
timestamp 1516238463
transform -1 0 3416 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_32
timestamp 1516238463
transform -1 0 3448 0 -1 1810
box 0 0 32 200
use AND2X2  AND2X2_99
timestamp 1516238463
transform 1 0 3448 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_27
timestamp 1516238463
transform -1 0 3576 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_114
timestamp 1516238463
transform 1 0 3576 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_189
timestamp 1516238463
transform -1 0 3704 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_121
timestamp 1516238463
transform 1 0 3704 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_188
timestamp 1516238463
transform -1 0 3832 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_26
timestamp 1516238463
transform -1 0 3896 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_305
timestamp 1516238463
transform -1 0 3960 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_95
timestamp 1516238463
transform -1 0 4024 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_3_0
timestamp 1516238463
transform -1 0 4040 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_3_1
timestamp 1516238463
transform -1 0 4056 0 -1 1810
box 0 0 16 200
use AND2X2  AND2X2_306
timestamp 1516238463
transform -1 0 4120 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_82
timestamp 1516238463
transform 1 0 4120 0 -1 1810
box 0 0 64 200
use INVX2  INVX2_3
timestamp 1516238463
transform 1 0 4184 0 -1 1810
box 0 0 32 200
use MUX2X1  MUX2X1_43
timestamp 1516238463
transform -1 0 4312 0 -1 1810
box 0 0 96 200
use OR2X2  OR2X2_60
timestamp 1516238463
transform 1 0 4312 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_120
timestamp 1516238463
transform -1 0 4440 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_230
timestamp 1516238463
transform -1 0 4504 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_119
timestamp 1516238463
transform -1 0 4568 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_229
timestamp 1516238463
transform -1 0 4632 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_60
timestamp 1516238463
transform 1 0 4632 0 -1 1810
box 0 0 96 200
use OR2X2  OR2X2_118
timestamp 1516238463
transform -1 0 4792 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_62
timestamp 1516238463
transform 1 0 4792 0 -1 1810
box 0 0 96 200
use OR2X2  OR2X2_223
timestamp 1516238463
transform -1 0 4952 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_54
timestamp 1516238463
transform -1 0 5048 0 -1 1810
box 0 0 96 200
use FILL  FILL_8_4_0
timestamp 1516238463
transform -1 0 5064 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_4_1
timestamp 1516238463
transform -1 0 5080 0 -1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_40
timestamp 1516238463
transform -1 0 5176 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_55
timestamp 1516238463
transform -1 0 5272 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_71
timestamp 1516238463
transform -1 0 5368 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_41
timestamp 1516238463
transform -1 0 5464 0 -1 1810
box 0 0 96 200
use OR2X2  OR2X2_30
timestamp 1516238463
transform -1 0 5528 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_53
timestamp 1516238463
transform -1 0 5624 0 -1 1810
box 0 0 96 200
use AND2X2  AND2X2_209
timestamp 1516238463
transform 1 0 5624 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_105
timestamp 1516238463
transform 1 0 5688 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_99
timestamp 1516238463
transform -1 0 5816 0 -1 1810
box 0 0 64 200
use OR2X2  OR2X2_103
timestamp 1516238463
transform 1 0 5816 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_604
timestamp 1516238463
transform 1 0 5880 0 -1 1810
box 0 0 64 200
use FILL  FILL_9_1
timestamp 1516238463
transform -1 0 5960 0 -1 1810
box 0 0 16 200
use FILL  FILL_9_2
timestamp 1516238463
transform -1 0 5976 0 -1 1810
box 0 0 16 200
use FILL  FILL_9_3
timestamp 1516238463
transform -1 0 5992 0 -1 1810
box 0 0 16 200
use BUFX2  BUFX2_61
timestamp 1516238463
transform -1 0 56 0 1 1410
box 0 0 48 200
use BUFX2  BUFX2_59
timestamp 1516238463
transform -1 0 104 0 1 1410
box 0 0 48 200
use BUFX2  BUFX2_26
timestamp 1516238463
transform -1 0 152 0 1 1410
box 0 0 48 200
use BUFX2  BUFX2_24
timestamp 1516238463
transform -1 0 200 0 1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_18
timestamp 1516238463
transform -1 0 392 0 1 1410
box 0 0 192 200
use INVX1  INVX1_34
timestamp 1516238463
transform -1 0 424 0 1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_72
timestamp 1516238463
transform -1 0 472 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_36
timestamp 1516238463
transform -1 0 536 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_73
timestamp 1516238463
transform -1 0 584 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_53
timestamp 1516238463
transform -1 0 648 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_510
timestamp 1516238463
transform 1 0 648 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_511
timestamp 1516238463
transform -1 0 776 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_5
timestamp 1516238463
transform -1 0 824 0 1 1410
box 0 0 48 200
use AND2X2  AND2X2_514
timestamp 1516238463
transform 1 0 824 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_365
timestamp 1516238463
transform 1 0 888 0 1 1410
box 0 0 64 200
use FILL  FILL_7_0_0
timestamp 1516238463
transform 1 0 952 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1516238463
transform 1 0 968 0 1 1410
box 0 0 16 200
use AOI21X1  AOI21X1_32
timestamp 1516238463
transform 1 0 984 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_68
timestamp 1516238463
transform -1 0 1096 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_27
timestamp 1516238463
transform -1 0 1160 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_57
timestamp 1516238463
transform -1 0 1208 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_11
timestamp 1516238463
transform -1 0 1272 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_28
timestamp 1516238463
transform 1 0 1272 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_502
timestamp 1516238463
transform -1 0 1400 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_500
timestamp 1516238463
transform -1 0 1464 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_74
timestamp 1516238463
transform -1 0 1528 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_30
timestamp 1516238463
transform -1 0 1592 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_7
timestamp 1516238463
transform 1 0 1592 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_77
timestamp 1516238463
transform -1 0 1720 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_515
timestamp 1516238463
transform 1 0 1720 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_366
timestamp 1516238463
transform -1 0 1848 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_80
timestamp 1516238463
transform -1 0 1912 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_237
timestamp 1516238463
transform 1 0 1912 0 1 1410
box 0 0 64 200
use FILL  FILL_7_1_0
timestamp 1516238463
transform 1 0 1976 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1516238463
transform 1 0 1992 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_75
timestamp 1516238463
transform 1 0 2008 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_345
timestamp 1516238463
transform -1 0 2136 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_344
timestamp 1516238463
transform -1 0 2200 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_23
timestamp 1516238463
transform 1 0 2200 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_251
timestamp 1516238463
transform -1 0 2328 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_37
timestamp 1516238463
transform 1 0 2328 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_45
timestamp 1516238463
transform 1 0 2376 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_1
timestamp 1516238463
transform -1 0 2488 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_41
timestamp 1516238463
transform 1 0 2488 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_61
timestamp 1516238463
transform -1 0 2616 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_31
timestamp 1516238463
transform 1 0 2616 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_83
timestamp 1516238463
transform 1 0 2680 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_79
timestamp 1516238463
transform 1 0 2744 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_1
timestamp 1516238463
transform 1 0 2808 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_62
timestamp 1516238463
transform 1 0 2856 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_12
timestamp 1516238463
transform 1 0 2920 0 1 1410
box 0 0 48 200
use FILL  FILL_7_2_0
timestamp 1516238463
transform -1 0 2984 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1516238463
transform -1 0 3000 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_23
timestamp 1516238463
transform -1 0 3048 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_1
timestamp 1516238463
transform -1 0 3112 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_56
timestamp 1516238463
transform 1 0 3112 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_42
timestamp 1516238463
transform -1 0 3224 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_43
timestamp 1516238463
transform -1 0 3272 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_10
timestamp 1516238463
transform -1 0 3336 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_392
timestamp 1516238463
transform -1 0 3400 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_54
timestamp 1516238463
transform -1 0 3448 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_53
timestamp 1516238463
transform -1 0 3496 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_47
timestamp 1516238463
transform -1 0 3544 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_46
timestamp 1516238463
transform -1 0 3592 0 1 1410
box 0 0 48 200
use INVX2  INVX2_5
timestamp 1516238463
transform -1 0 3624 0 1 1410
box 0 0 32 200
use AND2X2  AND2X2_239
timestamp 1516238463
transform -1 0 3688 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_238
timestamp 1516238463
transform -1 0 3752 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_277
timestamp 1516238463
transform -1 0 3816 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_223
timestamp 1516238463
transform 1 0 3816 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_100
timestamp 1516238463
transform -1 0 3944 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_353
timestamp 1516238463
transform -1 0 4008 0 1 1410
box 0 0 64 200
use FILL  FILL_7_3_0
timestamp 1516238463
transform -1 0 4024 0 1 1410
box 0 0 16 200
use FILL  FILL_7_3_1
timestamp 1516238463
transform -1 0 4040 0 1 1410
box 0 0 16 200
use OR2X2  OR2X2_430
timestamp 1516238463
transform -1 0 4104 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_19
timestamp 1516238463
transform -1 0 4168 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_8
timestamp 1516238463
transform -1 0 4216 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_6
timestamp 1516238463
transform -1 0 4280 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_628
timestamp 1516238463
transform 1 0 4280 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_2
timestamp 1516238463
transform -1 0 4392 0 1 1410
box 0 0 48 200
use OR2X2  OR2X2_413
timestamp 1516238463
transform -1 0 4456 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_18
timestamp 1516238463
transform -1 0 4520 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_412
timestamp 1516238463
transform -1 0 4584 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_609
timestamp 1516238463
transform -1 0 4648 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_44
timestamp 1516238463
transform -1 0 4744 0 1 1410
box 0 0 96 200
use AND2X2  AND2X2_83
timestamp 1516238463
transform -1 0 4808 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_63
timestamp 1516238463
transform 1 0 4808 0 1 1410
box 0 0 96 200
use XOR2X1  XOR2X1_1
timestamp 1516238463
transform 1 0 4904 0 1 1410
box 0 0 112 200
use FILL  FILL_7_4_0
timestamp 1516238463
transform -1 0 5032 0 1 1410
box 0 0 16 200
use FILL  FILL_7_4_1
timestamp 1516238463
transform -1 0 5048 0 1 1410
box 0 0 16 200
use AND2X2  AND2X2_138
timestamp 1516238463
transform -1 0 5112 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_80
timestamp 1516238463
transform -1 0 5176 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_56
timestamp 1516238463
transform -1 0 5272 0 1 1410
box 0 0 96 200
use AND2X2  AND2X2_72
timestamp 1516238463
transform 1 0 5272 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_75
timestamp 1516238463
transform -1 0 5400 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_200
timestamp 1516238463
transform 1 0 5400 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_102
timestamp 1516238463
transform 1 0 5464 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_5
timestamp 1516238463
transform 1 0 5528 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_100
timestamp 1516238463
transform -1 0 5656 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_101
timestamp 1516238463
transform -1 0 5720 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_142
timestamp 1516238463
transform -1 0 5784 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_601
timestamp 1516238463
transform 1 0 5784 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_605
timestamp 1516238463
transform -1 0 5912 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_379
timestamp 1516238463
transform 1 0 5912 0 1 1410
box 0 0 64 200
use FILL  FILL_8_1
timestamp 1516238463
transform 1 0 5976 0 1 1410
box 0 0 16 200
use BUFX2  BUFX2_64
timestamp 1516238463
transform -1 0 56 0 -1 1410
box 0 0 48 200
use BUFX2  BUFX2_29
timestamp 1516238463
transform -1 0 104 0 -1 1410
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_24
timestamp 1516238463
transform -1 0 296 0 -1 1410
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_20
timestamp 1516238463
transform -1 0 488 0 -1 1410
box 0 0 192 200
use OR2X2  OR2X2_404
timestamp 1516238463
transform 1 0 488 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_252
timestamp 1516238463
transform 1 0 552 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_39
timestamp 1516238463
transform -1 0 648 0 -1 1410
box 0 0 32 200
use OR2X2  OR2X2_375
timestamp 1516238463
transform -1 0 712 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_362
timestamp 1516238463
transform -1 0 776 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_33
timestamp 1516238463
transform -1 0 808 0 -1 1410
box 0 0 32 200
use AND2X2  AND2X2_513
timestamp 1516238463
transform -1 0 872 0 -1 1410
box 0 0 64 200
use XNOR2X1  XNOR2X1_3
timestamp 1516238463
transform -1 0 984 0 -1 1410
box 0 0 112 200
use FILL  FILL_6_0_0
timestamp 1516238463
transform -1 0 1000 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1516238463
transform -1 0 1016 0 -1 1410
box 0 0 16 200
use AND2X2  AND2X2_581
timestamp 1516238463
transform -1 0 1080 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_317
timestamp 1516238463
transform -1 0 1144 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_465
timestamp 1516238463
transform -1 0 1208 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_58
timestamp 1516238463
transform 1 0 1208 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_69
timestamp 1516238463
transform -1 0 1320 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_37
timestamp 1516238463
transform -1 0 1384 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_359
timestamp 1516238463
transform 1 0 1384 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_387
timestamp 1516238463
transform 1 0 1448 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_59
timestamp 1516238463
transform -1 0 1576 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_540
timestamp 1516238463
transform 1 0 1576 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_22
timestamp 1516238463
transform 1 0 1640 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_98
timestamp 1516238463
transform -1 0 1768 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_427
timestamp 1516238463
transform -1 0 1832 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_3
timestamp 1516238463
transform 1 0 1832 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_3
timestamp 1516238463
transform 1 0 1880 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_1_0
timestamp 1516238463
transform -1 0 1960 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1516238463
transform -1 0 1976 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_81
timestamp 1516238463
transform -1 0 2040 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_378
timestamp 1516238463
transform -1 0 2104 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_82
timestamp 1516238463
transform -1 0 2168 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_73
timestamp 1516238463
transform -1 0 2232 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_343
timestamp 1516238463
transform -1 0 2296 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_383
timestamp 1516238463
transform -1 0 2360 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_222
timestamp 1516238463
transform -1 0 2424 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_76
timestamp 1516238463
transform 1 0 2424 0 -1 1410
box 0 0 64 200
use INVX2  INVX2_1
timestamp 1516238463
transform -1 0 2520 0 -1 1410
box 0 0 32 200
use OR2X2  OR2X2_250
timestamp 1516238463
transform 1 0 2520 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_374
timestamp 1516238463
transform 1 0 2584 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_1
timestamp 1516238463
transform -1 0 2712 0 -1 1410
box 0 0 64 200
use INVX2  INVX2_7
timestamp 1516238463
transform 1 0 2712 0 -1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_1
timestamp 1516238463
transform 1 0 2744 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_288
timestamp 1516238463
transform 1 0 2808 0 -1 1410
box 0 0 64 200
use INVX2  INVX2_6
timestamp 1516238463
transform 1 0 2872 0 -1 1410
box 0 0 32 200
use BUFX4  BUFX4_78
timestamp 1516238463
transform 1 0 2904 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_2_0
timestamp 1516238463
transform -1 0 2984 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1516238463
transform -1 0 3000 0 -1 1410
box 0 0 16 200
use OR2X2  OR2X2_323
timestamp 1516238463
transform -1 0 3064 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_307
timestamp 1516238463
transform -1 0 3128 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_452
timestamp 1516238463
transform -1 0 3192 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_17
timestamp 1516238463
transform 1 0 3192 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_265
timestamp 1516238463
transform -1 0 3320 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_93
timestamp 1516238463
transform 1 0 3320 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_26
timestamp 1516238463
transform -1 0 3448 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_14
timestamp 1516238463
transform 1 0 3448 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_21
timestamp 1516238463
transform -1 0 3544 0 -1 1410
box 0 0 32 200
use AOI21X1  AOI21X1_19
timestamp 1516238463
transform 1 0 3544 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_14
timestamp 1516238463
transform 1 0 3608 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_38
timestamp 1516238463
transform -1 0 3704 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_20
timestamp 1516238463
transform -1 0 3752 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_25
timestamp 1516238463
transform 1 0 3752 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_534
timestamp 1516238463
transform -1 0 3880 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_40
timestamp 1516238463
transform 1 0 3880 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_128
timestamp 1516238463
transform 1 0 3944 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_3_0
timestamp 1516238463
transform -1 0 4024 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_3_1
timestamp 1516238463
transform -1 0 4040 0 -1 1410
box 0 0 16 200
use AND2X2  AND2X2_391
timestamp 1516238463
transform -1 0 4104 0 -1 1410
box 0 0 64 200
use XOR2X1  XOR2X1_3
timestamp 1516238463
transform -1 0 4216 0 -1 1410
box 0 0 112 200
use AOI21X1  AOI21X1_23
timestamp 1516238463
transform -1 0 4280 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_308
timestamp 1516238463
transform -1 0 4344 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_3
timestamp 1516238463
transform -1 0 4392 0 -1 1410
box 0 0 48 200
use OR2X2  OR2X2_300
timestamp 1516238463
transform -1 0 4456 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_244
timestamp 1516238463
transform -1 0 4520 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_629
timestamp 1516238463
transform 1 0 4520 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_424
timestamp 1516238463
transform 1 0 4584 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_118
timestamp 1516238463
transform -1 0 4712 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1516238463
transform 1 0 4712 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_99
timestamp 1516238463
transform -1 0 4840 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_198
timestamp 1516238463
transform -1 0 4904 0 -1 1410
box 0 0 64 200
use XOR2X1  XOR2X1_6
timestamp 1516238463
transform 1 0 4904 0 -1 1410
box 0 0 112 200
use FILL  FILL_6_4_0
timestamp 1516238463
transform -1 0 5032 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_4_1
timestamp 1516238463
transform -1 0 5048 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_34
timestamp 1516238463
transform -1 0 5096 0 -1 1410
box 0 0 48 200
use OR2X2  OR2X2_15
timestamp 1516238463
transform -1 0 5160 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_364
timestamp 1516238463
transform 1 0 5160 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_243
timestamp 1516238463
transform -1 0 5288 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_12
timestamp 1516238463
transform -1 0 5352 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_78
timestamp 1516238463
transform -1 0 5416 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_64
timestamp 1516238463
transform 1 0 5416 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_419
timestamp 1516238463
transform 1 0 5480 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_365
timestamp 1516238463
transform 1 0 5544 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_431
timestamp 1516238463
transform -1 0 5672 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_8
timestamp 1516238463
transform -1 0 5736 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_44
timestamp 1516238463
transform -1 0 5800 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_401
timestamp 1516238463
transform -1 0 5864 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_243
timestamp 1516238463
transform -1 0 5928 0 -1 1410
box 0 0 64 200
use FILL  FILL_7_1
timestamp 1516238463
transform -1 0 5944 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_2
timestamp 1516238463
transform -1 0 5960 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_3
timestamp 1516238463
transform -1 0 5976 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_4
timestamp 1516238463
transform -1 0 5992 0 -1 1410
box 0 0 16 200
use BUFX2  BUFX2_58
timestamp 1516238463
transform -1 0 56 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_23
timestamp 1516238463
transform -1 0 104 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_63
timestamp 1516238463
transform -1 0 152 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_28
timestamp 1516238463
transform -1 0 200 0 1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_22
timestamp 1516238463
transform -1 0 392 0 1 1010
box 0 0 192 200
use INVX1  INVX1_38
timestamp 1516238463
transform -1 0 424 0 1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_17
timestamp 1516238463
transform -1 0 616 0 1 1010
box 0 0 192 200
use AND2X2  AND2X2_589
timestamp 1516238463
transform 1 0 616 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_384
timestamp 1516238463
transform -1 0 744 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_64
timestamp 1516238463
transform 1 0 744 0 1 1010
box 0 0 48 200
use INVX1  INVX1_46
timestamp 1516238463
transform 1 0 792 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_65
timestamp 1516238463
transform -1 0 872 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_54
timestamp 1516238463
transform -1 0 936 0 1 1010
box 0 0 64 200
use FILL  FILL_5_0_0
timestamp 1516238463
transform -1 0 952 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1516238463
transform -1 0 968 0 1 1010
box 0 0 16 200
use AND2X2  AND2X2_538
timestamp 1516238463
transform -1 0 1032 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_539
timestamp 1516238463
transform -1 0 1096 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_397
timestamp 1516238463
transform -1 0 1160 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_35
timestamp 1516238463
transform -1 0 1224 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_70
timestamp 1516238463
transform 1 0 1224 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_311
timestamp 1516238463
transform -1 0 1336 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_241
timestamp 1516238463
transform 1 0 1336 0 1 1010
box 0 0 64 200
use INVX1  INVX1_30
timestamp 1516238463
transform 1 0 1400 0 1 1010
box 0 0 32 200
use BUFX4  BUFX4_95
timestamp 1516238463
transform -1 0 1496 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_97
timestamp 1516238463
transform -1 0 1560 0 1 1010
box 0 0 64 200
use XNOR2X1  XNOR2X1_2
timestamp 1516238463
transform 1 0 1560 0 1 1010
box 0 0 112 200
use AND2X2  AND2X2_440
timestamp 1516238463
transform 1 0 1672 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_439
timestamp 1516238463
transform 1 0 1736 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_4
timestamp 1516238463
transform 1 0 1800 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_29
timestamp 1516238463
transform 1 0 1864 0 1 1010
box 0 0 64 200
use FILL  FILL_5_1_0
timestamp 1516238463
transform -1 0 1944 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1516238463
transform -1 0 1960 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_37
timestamp 1516238463
transform -1 0 2024 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_537
timestamp 1516238463
transform -1 0 2088 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_536
timestamp 1516238463
transform -1 0 2152 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_5
timestamp 1516238463
transform -1 0 2216 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_225
timestamp 1516238463
transform 1 0 2216 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_38
timestamp 1516238463
transform 1 0 2280 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_35
timestamp 1516238463
transform -1 0 2408 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_34
timestamp 1516238463
transform 1 0 2408 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_182
timestamp 1516238463
transform -1 0 2536 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_12
timestamp 1516238463
transform -1 0 2600 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_2
timestamp 1516238463
transform 1 0 2600 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_18
timestamp 1516238463
transform -1 0 2728 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_424
timestamp 1516238463
transform -1 0 2792 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_5
timestamp 1516238463
transform -1 0 2840 0 1 1010
box 0 0 48 200
use AND2X2  AND2X2_480
timestamp 1516238463
transform -1 0 2904 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_478
timestamp 1516238463
transform -1 0 2968 0 1 1010
box 0 0 64 200
use FILL  FILL_5_2_0
timestamp 1516238463
transform 1 0 2968 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1516238463
transform 1 0 2984 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_17
timestamp 1516238463
transform 1 0 3000 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_94
timestamp 1516238463
transform 1 0 3064 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1516238463
transform -1 0 3192 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_38
timestamp 1516238463
transform 1 0 3192 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_410
timestamp 1516238463
transform 1 0 3256 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_39
timestamp 1516238463
transform 1 0 3320 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_15
timestamp 1516238463
transform -1 0 3432 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_40
timestamp 1516238463
transform 1 0 3432 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_6
timestamp 1516238463
transform -1 0 3544 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_21
timestamp 1516238463
transform 1 0 3544 0 1 1010
box 0 0 48 200
use OR2X2  OR2X2_331
timestamp 1516238463
transform -1 0 3656 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_408
timestamp 1516238463
transform 1 0 3656 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_382
timestamp 1516238463
transform -1 0 3784 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_292
timestamp 1516238463
transform -1 0 3848 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_199
timestamp 1516238463
transform -1 0 3912 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_137
timestamp 1516238463
transform -1 0 3976 0 1 1010
box 0 0 64 200
use FILL  FILL_5_3_0
timestamp 1516238463
transform -1 0 3992 0 1 1010
box 0 0 16 200
use FILL  FILL_5_3_1
timestamp 1516238463
transform -1 0 4008 0 1 1010
box 0 0 16 200
use OR2X2  OR2X2_318
timestamp 1516238463
transform -1 0 4072 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_79
timestamp 1516238463
transform -1 0 4136 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_113
timestamp 1516238463
transform -1 0 4200 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_297
timestamp 1516238463
transform -1 0 4264 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_178
timestamp 1516238463
transform -1 0 4328 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_69
timestamp 1516238463
transform 1 0 4328 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_181
timestamp 1516238463
transform -1 0 4456 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_53
timestamp 1516238463
transform -1 0 4520 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_130
timestamp 1516238463
transform -1 0 4584 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_166
timestamp 1516238463
transform -1 0 4648 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_330
timestamp 1516238463
transform -1 0 4712 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_136
timestamp 1516238463
transform -1 0 4776 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_62
timestamp 1516238463
transform -1 0 4840 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_76
timestamp 1516238463
transform -1 0 4904 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_56
timestamp 1516238463
transform -1 0 4968 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_143
timestamp 1516238463
transform -1 0 5032 0 1 1010
box 0 0 64 200
use FILL  FILL_5_4_0
timestamp 1516238463
transform -1 0 5048 0 1 1010
box 0 0 16 200
use FILL  FILL_5_4_1
timestamp 1516238463
transform -1 0 5064 0 1 1010
box 0 0 16 200
use OR2X2  OR2X2_180
timestamp 1516238463
transform -1 0 5128 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_295
timestamp 1516238463
transform -1 0 5192 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_296
timestamp 1516238463
transform -1 0 5256 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_624
timestamp 1516238463
transform -1 0 5320 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_12
timestamp 1516238463
transform -1 0 5384 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_113
timestamp 1516238463
transform -1 0 5448 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_146
timestamp 1516238463
transform -1 0 5512 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_108
timestamp 1516238463
transform 1 0 5512 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_244
timestamp 1516238463
transform -1 0 5640 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_109
timestamp 1516238463
transform -1 0 5704 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_130
timestamp 1516238463
transform -1 0 5768 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_242
timestamp 1516238463
transform -1 0 5832 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_104
timestamp 1516238463
transform -1 0 5896 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_25
timestamp 1516238463
transform 1 0 5896 0 1 1010
box 0 0 64 200
use FILL  FILL_6_1
timestamp 1516238463
transform 1 0 5960 0 1 1010
box 0 0 16 200
use FILL  FILL_6_2
timestamp 1516238463
transform 1 0 5976 0 1 1010
box 0 0 16 200
use BUFX2  BUFX2_65
timestamp 1516238463
transform -1 0 56 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_66
timestamp 1516238463
transform -1 0 104 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_31
timestamp 1516238463
transform -1 0 152 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_30
timestamp 1516238463
transform -1 0 200 0 -1 1010
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_25
timestamp 1516238463
transform -1 0 392 0 -1 1010
box 0 0 192 200
use INVX1  INVX1_40
timestamp 1516238463
transform -1 0 424 0 -1 1010
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_26
timestamp 1516238463
transform -1 0 616 0 -1 1010
box 0 0 192 200
use INVX1  INVX1_41
timestamp 1516238463
transform -1 0 648 0 -1 1010
box 0 0 32 200
use AND2X2  AND2X2_588
timestamp 1516238463
transform 1 0 648 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_591
timestamp 1516238463
transform 1 0 712 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_592
timestamp 1516238463
transform 1 0 776 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_352
timestamp 1516238463
transform -1 0 904 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_0_0
timestamp 1516238463
transform 1 0 904 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1516238463
transform 1 0 920 0 -1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_31
timestamp 1516238463
transform 1 0 936 0 -1 1010
box 0 0 64 200
use XNOR2X1  XNOR2X1_4
timestamp 1516238463
transform 1 0 1000 0 -1 1010
box 0 0 112 200
use NAND3X1  NAND3X1_36
timestamp 1516238463
transform 1 0 1112 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_31
timestamp 1516238463
transform -1 0 1224 0 -1 1010
box 0 0 48 200
use AND2X2  AND2X2_487
timestamp 1516238463
transform -1 0 1288 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_29
timestamp 1516238463
transform 1 0 1288 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_193
timestamp 1516238463
transform 1 0 1352 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_307
timestamp 1516238463
transform 1 0 1416 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_535
timestamp 1516238463
transform -1 0 1544 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_33
timestamp 1516238463
transform 1 0 1544 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_6
timestamp 1516238463
transform -1 0 1656 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_22
timestamp 1516238463
transform 1 0 1656 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_16
timestamp 1516238463
transform -1 0 1768 0 -1 1010
box 0 0 48 200
use OR2X2  OR2X2_299
timestamp 1516238463
transform 1 0 1768 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_143
timestamp 1516238463
transform 1 0 1832 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_21
timestamp 1516238463
transform -1 0 1960 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_1_0
timestamp 1516238463
transform 1 0 1960 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1516238463
transform 1 0 1976 0 -1 1010
box 0 0 16 200
use AND2X2  AND2X2_254
timestamp 1516238463
transform 1 0 1992 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_6
timestamp 1516238463
transform 1 0 2056 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_342
timestamp 1516238463
transform 1 0 2120 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_325
timestamp 1516238463
transform 1 0 2184 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_207
timestamp 1516238463
transform -1 0 2312 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_63
timestamp 1516238463
transform -1 0 2376 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_158
timestamp 1516238463
transform -1 0 2440 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_71
timestamp 1516238463
transform -1 0 2504 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_14
timestamp 1516238463
transform 1 0 2504 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_25
timestamp 1516238463
transform -1 0 2632 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_425
timestamp 1516238463
transform 1 0 2632 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_422
timestamp 1516238463
transform -1 0 2760 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_6
timestamp 1516238463
transform 1 0 2760 0 -1 1010
box 0 0 48 200
use AND2X2  AND2X2_191
timestamp 1516238463
transform -1 0 2872 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_42
timestamp 1516238463
transform -1 0 2936 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_407
timestamp 1516238463
transform 1 0 2936 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_2_0
timestamp 1516238463
transform -1 0 3016 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1516238463
transform -1 0 3032 0 -1 1010
box 0 0 16 200
use OR2X2  OR2X2_278
timestamp 1516238463
transform -1 0 3096 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_48
timestamp 1516238463
transform 1 0 3096 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_49
timestamp 1516238463
transform -1 0 3192 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_43
timestamp 1516238463
transform -1 0 3256 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_20
timestamp 1516238463
transform 1 0 3256 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_280
timestamp 1516238463
transform 1 0 3320 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_260
timestamp 1516238463
transform 1 0 3384 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_385
timestamp 1516238463
transform -1 0 3512 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_4
timestamp 1516238463
transform 1 0 3512 0 -1 1010
box 0 0 48 200
use OR2X2  OR2X2_7
timestamp 1516238463
transform 1 0 3560 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_34
timestamp 1516238463
transform 1 0 3624 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_409
timestamp 1516238463
transform -1 0 3752 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_276
timestamp 1516238463
transform -1 0 3816 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_108
timestamp 1516238463
transform -1 0 3880 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_58
timestamp 1516238463
transform -1 0 3944 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_254
timestamp 1516238463
transform -1 0 4008 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_3_0
timestamp 1516238463
transform 1 0 4008 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_1
timestamp 1516238463
transform 1 0 4024 0 -1 1010
box 0 0 16 200
use OR2X2  OR2X2_101
timestamp 1516238463
transform 1 0 4040 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_168
timestamp 1516238463
transform 1 0 4104 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_16
timestamp 1516238463
transform -1 0 4232 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_77
timestamp 1516238463
transform -1 0 4296 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_14
timestamp 1516238463
transform -1 0 4360 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_227
timestamp 1516238463
transform -1 0 4424 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_129
timestamp 1516238463
transform -1 0 4488 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_211
timestamp 1516238463
transform -1 0 4552 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_75
timestamp 1516238463
transform -1 0 4616 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_144
timestamp 1516238463
transform -1 0 4680 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_165
timestamp 1516238463
transform -1 0 4744 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_213
timestamp 1516238463
transform -1 0 4808 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_81
timestamp 1516238463
transform -1 0 4872 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_58
timestamp 1516238463
transform -1 0 4936 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_210
timestamp 1516238463
transform -1 0 5000 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_4_0
timestamp 1516238463
transform -1 0 5016 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_4_1
timestamp 1516238463
transform -1 0 5032 0 -1 1010
box 0 0 16 200
use AND2X2  AND2X2_331
timestamp 1516238463
transform -1 0 5096 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_131
timestamp 1516238463
transform -1 0 5160 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_56
timestamp 1516238463
transform -1 0 5224 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_107
timestamp 1516238463
transform -1 0 5288 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_79
timestamp 1516238463
transform -1 0 5352 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_607
timestamp 1516238463
transform -1 0 5416 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_205
timestamp 1516238463
transform -1 0 5480 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_32
timestamp 1516238463
transform -1 0 5544 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_211
timestamp 1516238463
transform -1 0 5608 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_210
timestamp 1516238463
transform -1 0 5672 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_106
timestamp 1516238463
transform -1 0 5736 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_438
timestamp 1516238463
transform -1 0 5800 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_21
timestamp 1516238463
transform -1 0 5864 0 -1 1010
box 0 0 64 200
use OR2X2  OR2X2_55
timestamp 1516238463
transform -1 0 5928 0 -1 1010
box 0 0 64 200
use FILL  FILL_5_1
timestamp 1516238463
transform -1 0 5944 0 -1 1010
box 0 0 16 200
use FILL  FILL_5_2
timestamp 1516238463
transform -1 0 5960 0 -1 1010
box 0 0 16 200
use FILL  FILL_5_3
timestamp 1516238463
transform -1 0 5976 0 -1 1010
box 0 0 16 200
use FILL  FILL_5_4
timestamp 1516238463
transform -1 0 5992 0 -1 1010
box 0 0 16 200
use BUFX2  BUFX2_62
timestamp 1516238463
transform -1 0 56 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_27
timestamp 1516238463
transform -1 0 104 0 1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_27
timestamp 1516238463
transform -1 0 296 0 1 610
box 0 0 192 200
use INVX1  INVX1_43
timestamp 1516238463
transform -1 0 328 0 1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_21
timestamp 1516238463
transform -1 0 520 0 1 610
box 0 0 192 200
use INVX1  INVX1_36
timestamp 1516238463
transform -1 0 552 0 1 610
box 0 0 32 200
use INVX1  INVX1_37
timestamp 1516238463
transform -1 0 584 0 1 610
box 0 0 32 200
use AND2X2  AND2X2_577
timestamp 1516238463
transform 1 0 584 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_578
timestamp 1516238463
transform 1 0 648 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_580
timestamp 1516238463
transform 1 0 712 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_341
timestamp 1516238463
transform -1 0 840 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_242
timestamp 1516238463
transform -1 0 904 0 1 610
box 0 0 64 200
use FILL  FILL_3_0_0
timestamp 1516238463
transform -1 0 920 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1516238463
transform -1 0 936 0 1 610
box 0 0 16 200
use AND2X2  AND2X2_583
timestamp 1516238463
transform -1 0 1000 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_11
timestamp 1516238463
transform -1 0 1064 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_32
timestamp 1516238463
transform 1 0 1064 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_26
timestamp 1516238463
transform 1 0 1112 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_8
timestamp 1516238463
transform 1 0 1160 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_25
timestamp 1516238463
transform -1 0 1272 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_137
timestamp 1516238463
transform -1 0 1336 0 1 610
box 0 0 64 200
use INVX2  INVX2_8
timestamp 1516238463
transform -1 0 1368 0 1 610
box 0 0 32 200
use NAND3X1  NAND3X1_28
timestamp 1516238463
transform -1 0 1432 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_136
timestamp 1516238463
transform 1 0 1432 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_3
timestamp 1516238463
transform 1 0 1496 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_17
timestamp 1516238463
transform 1 0 1560 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_4
timestamp 1516238463
transform 1 0 1608 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_582
timestamp 1516238463
transform -1 0 1736 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_30
timestamp 1516238463
transform 1 0 1736 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_29
timestamp 1516238463
transform -1 0 1832 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_33
timestamp 1516238463
transform -1 0 1896 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_10
timestamp 1516238463
transform 1 0 1896 0 1 610
box 0 0 64 200
use FILL  FILL_3_1_0
timestamp 1516238463
transform -1 0 1976 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1516238463
transform -1 0 1992 0 1 610
box 0 0 16 200
use AND2X2  AND2X2_347
timestamp 1516238463
transform -1 0 2056 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_35
timestamp 1516238463
transform -1 0 2120 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_32
timestamp 1516238463
transform -1 0 2184 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_30
timestamp 1516238463
transform 1 0 2184 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_9
timestamp 1516238463
transform -1 0 2312 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_28
timestamp 1516238463
transform -1 0 2360 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_27
timestamp 1516238463
transform -1 0 2408 0 1 610
box 0 0 48 200
use AND2X2  AND2X2_363
timestamp 1516238463
transform -1 0 2472 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_230
timestamp 1516238463
transform -1 0 2536 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_213
timestamp 1516238463
transform -1 0 2600 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_8
timestamp 1516238463
transform -1 0 2648 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_9
timestamp 1516238463
transform -1 0 2696 0 1 610
box 0 0 48 200
use AND2X2  AND2X2_259
timestamp 1516238463
transform -1 0 2760 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_162
timestamp 1516238463
transform -1 0 2824 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_44
timestamp 1516238463
transform 1 0 2824 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_289
timestamp 1516238463
transform -1 0 2952 0 1 610
box 0 0 64 200
use FILL  FILL_3_2_0
timestamp 1516238463
transform 1 0 2952 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1516238463
transform 1 0 2968 0 1 610
box 0 0 16 200
use NAND3X1  NAND3X1_16
timestamp 1516238463
transform 1 0 2984 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_96
timestamp 1516238463
transform -1 0 3112 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_10
timestamp 1516238463
transform 1 0 3112 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_15
timestamp 1516238463
transform -1 0 3224 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_11
timestamp 1516238463
transform -1 0 3272 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_42
timestamp 1516238463
transform 1 0 3272 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_126
timestamp 1516238463
transform -1 0 3400 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_127
timestamp 1516238463
transform 1 0 3400 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_59
timestamp 1516238463
transform -1 0 3528 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_133
timestamp 1516238463
transform -1 0 3592 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_240
timestamp 1516238463
transform -1 0 3656 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_109
timestamp 1516238463
transform -1 0 3720 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_277
timestamp 1516238463
transform -1 0 3784 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_29
timestamp 1516238463
transform 1 0 3784 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_102
timestamp 1516238463
transform -1 0 3912 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_149
timestamp 1516238463
transform -1 0 3976 0 1 610
box 0 0 64 200
use FILL  FILL_3_3_0
timestamp 1516238463
transform -1 0 3992 0 1 610
box 0 0 16 200
use FILL  FILL_3_3_1
timestamp 1516238463
transform -1 0 4008 0 1 610
box 0 0 16 200
use OR2X2  OR2X2_253
timestamp 1516238463
transform -1 0 4072 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_90
timestamp 1516238463
transform -1 0 4136 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_17
timestamp 1516238463
transform -1 0 4200 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_332
timestamp 1516238463
transform -1 0 4264 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_209
timestamp 1516238463
transform -1 0 4328 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_350
timestamp 1516238463
transform -1 0 4392 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_245
timestamp 1516238463
transform -1 0 4456 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_407
timestamp 1516238463
transform 1 0 4456 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_406
timestamp 1516238463
transform -1 0 4584 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_262
timestamp 1516238463
transform -1 0 4648 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_145
timestamp 1516238463
transform -1 0 4712 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_348
timestamp 1516238463
transform -1 0 4776 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_608
timestamp 1516238463
transform -1 0 4840 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_61
timestamp 1516238463
transform 1 0 4840 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_157
timestamp 1516238463
transform -1 0 4968 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_132
timestamp 1516238463
transform -1 0 5032 0 1 610
box 0 0 64 200
use FILL  FILL_3_4_0
timestamp 1516238463
transform -1 0 5048 0 1 610
box 0 0 16 200
use FILL  FILL_3_4_1
timestamp 1516238463
transform -1 0 5064 0 1 610
box 0 0 16 200
use AND2X2  AND2X2_241
timestamp 1516238463
transform -1 0 5128 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_148
timestamp 1516238463
transform -1 0 5192 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_147
timestamp 1516238463
transform -1 0 5256 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_261
timestamp 1516238463
transform -1 0 5320 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_405
timestamp 1516238463
transform -1 0 5384 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_606
timestamp 1516238463
transform -1 0 5448 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_60
timestamp 1516238463
transform 1 0 5448 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_111
timestamp 1516238463
transform -1 0 5576 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_172
timestamp 1516238463
transform -1 0 5640 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_14
timestamp 1516238463
transform 1 0 5640 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_171
timestamp 1516238463
transform -1 0 5768 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_169
timestamp 1516238463
transform -1 0 5832 0 1 610
box 0 0 64 200
use OR2X2  OR2X2_77
timestamp 1516238463
transform 1 0 5832 0 1 610
box 0 0 64 200
use MUX2X1  MUX2X1_9
timestamp 1516238463
transform 1 0 5896 0 1 610
box 0 0 96 200
use BUFX2  BUFX2_67
timestamp 1516238463
transform -1 0 56 0 -1 610
box 0 0 48 200
use BUFX2  BUFX2_32
timestamp 1516238463
transform -1 0 104 0 -1 610
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1516238463
transform -1 0 296 0 -1 610
box 0 0 192 200
use INVX1  INVX1_20
timestamp 1516238463
transform -1 0 328 0 -1 610
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1516238463
transform -1 0 520 0 -1 610
box 0 0 192 200
use INVX1  INVX1_35
timestamp 1516238463
transform -1 0 552 0 -1 610
box 0 0 32 200
use INVX1  INVX1_15
timestamp 1516238463
transform -1 0 584 0 -1 610
box 0 0 32 200
use INVX1  INVX1_16
timestamp 1516238463
transform -1 0 616 0 -1 610
box 0 0 32 200
use AND2X2  AND2X2_565
timestamp 1516238463
transform 1 0 616 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_566
timestamp 1516238463
transform 1 0 680 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_584
timestamp 1516238463
transform 1 0 744 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_29
timestamp 1516238463
transform -1 0 872 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_61
timestamp 1516238463
transform 1 0 872 0 -1 610
box 0 0 48 200
use FILL  FILL_2_0_0
timestamp 1516238463
transform 1 0 920 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1516238463
transform 1 0 936 0 -1 610
box 0 0 16 200
use NAND3X1  NAND3X1_51
timestamp 1516238463
transform 1 0 952 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_60
timestamp 1516238463
transform 1 0 1016 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_125
timestamp 1516238463
transform -1 0 1128 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_122
timestamp 1516238463
transform 1 0 1128 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_567
timestamp 1516238463
transform -1 0 1256 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_194
timestamp 1516238463
transform 1 0 1256 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_123
timestamp 1516238463
transform 1 0 1320 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_177
timestamp 1516238463
transform -1 0 1448 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_7
timestamp 1516238463
transform -1 0 1512 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_24
timestamp 1516238463
transform 1 0 1512 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_27
timestamp 1516238463
transform 1 0 1560 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_22
timestamp 1516238463
transform -1 0 1672 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_14
timestamp 1516238463
transform 1 0 1672 0 -1 610
box 0 0 48 200
use AOI21X1  AOI21X1_2
timestamp 1516238463
transform -1 0 1784 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_17
timestamp 1516238463
transform 1 0 1784 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_13
timestamp 1516238463
transform -1 0 1896 0 -1 610
box 0 0 48 200
use OR2X2  OR2X2_226
timestamp 1516238463
transform -1 0 1960 0 -1 610
box 0 0 64 200
use FILL  FILL_2_1_0
timestamp 1516238463
transform -1 0 1976 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1516238463
transform -1 0 1992 0 -1 610
box 0 0 16 200
use AND2X2  AND2X2_236
timestamp 1516238463
transform -1 0 2056 0 -1 610
box 0 0 64 200
use INVX1  INVX1_31
timestamp 1516238463
transform 1 0 2056 0 -1 610
box 0 0 32 200
use OR2X2  OR2X2_128
timestamp 1516238463
transform 1 0 2088 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_144
timestamp 1516238463
transform -1 0 2216 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_52
timestamp 1516238463
transform 1 0 2216 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1516238463
transform -1 0 2344 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_294
timestamp 1516238463
transform -1 0 2408 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_477
timestamp 1516238463
transform 1 0 2408 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_13
timestamp 1516238463
transform 1 0 2472 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_333
timestamp 1516238463
transform 1 0 2536 0 -1 610
box 0 0 64 200
use INVX1  INVX1_29
timestamp 1516238463
transform -1 0 2632 0 -1 610
box 0 0 32 200
use AOI21X1  AOI21X1_40
timestamp 1516238463
transform 1 0 2632 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_72
timestamp 1516238463
transform 1 0 2696 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_291
timestamp 1516238463
transform -1 0 2824 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_426
timestamp 1516238463
transform -1 0 2888 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_21
timestamp 1516238463
transform -1 0 2952 0 -1 610
box 0 0 64 200
use FILL  FILL_2_2_0
timestamp 1516238463
transform -1 0 2968 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1516238463
transform -1 0 2984 0 -1 610
box 0 0 16 200
use NAND3X1  NAND3X1_46
timestamp 1516238463
transform -1 0 3048 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_51
timestamp 1516238463
transform -1 0 3096 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_50
timestamp 1516238463
transform -1 0 3144 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_139
timestamp 1516238463
transform -1 0 3208 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_124
timestamp 1516238463
transform 1 0 3208 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_97
timestamp 1516238463
transform -1 0 3336 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_195
timestamp 1516238463
transform -1 0 3400 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_138
timestamp 1516238463
transform 1 0 3400 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_161
timestamp 1516238463
transform -1 0 3528 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_271
timestamp 1516238463
transform -1 0 3592 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_398
timestamp 1516238463
transform -1 0 3656 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_165
timestamp 1516238463
transform -1 0 3720 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_27
timestamp 1516238463
transform -1 0 3784 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_281
timestamp 1516238463
transform -1 0 3848 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_49
timestamp 1516238463
transform 1 0 3848 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_26
timestamp 1516238463
transform 1 0 3912 0 -1 610
box 0 0 64 200
use FILL  FILL_2_3_0
timestamp 1516238463
transform -1 0 3992 0 -1 610
box 0 0 16 200
use FILL  FILL_2_3_1
timestamp 1516238463
transform -1 0 4008 0 -1 610
box 0 0 16 200
use AND2X2  AND2X2_129
timestamp 1516238463
transform -1 0 4072 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_263
timestamp 1516238463
transform -1 0 4136 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_266
timestamp 1516238463
transform -1 0 4200 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_23
timestamp 1516238463
transform 1 0 4200 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_13
timestamp 1516238463
transform 1 0 4264 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_36
timestamp 1516238463
transform -1 0 4392 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_34
timestamp 1516238463
transform -1 0 4456 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_107
timestamp 1516238463
transform -1 0 4520 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_598
timestamp 1516238463
transform 1 0 4520 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_229
timestamp 1516238463
transform -1 0 4648 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_368
timestamp 1516238463
transform -1 0 4712 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_596
timestamp 1516238463
transform -1 0 4776 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_114
timestamp 1516238463
transform -1 0 4840 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_31
timestamp 1516238463
transform -1 0 4904 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_12
timestamp 1516238463
transform -1 0 4952 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_129
timestamp 1516238463
transform 1 0 4952 0 -1 610
box 0 0 64 200
use FILL  FILL_2_4_0
timestamp 1516238463
transform -1 0 5032 0 -1 610
box 0 0 16 200
use FILL  FILL_2_4_1
timestamp 1516238463
transform -1 0 5048 0 -1 610
box 0 0 16 200
use AND2X2  AND2X2_597
timestamp 1516238463
transform -1 0 5112 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_106
timestamp 1516238463
transform -1 0 5176 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_260
timestamp 1516238463
transform -1 0 5240 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_228
timestamp 1516238463
transform -1 0 5304 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_55
timestamp 1516238463
transform 1 0 5304 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_33
timestamp 1516238463
transform -1 0 5432 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_110
timestamp 1516238463
transform -1 0 5496 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_349
timestamp 1516238463
transform -1 0 5560 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_78
timestamp 1516238463
transform -1 0 5624 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_435
timestamp 1516238463
transform -1 0 5688 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_17
timestamp 1516238463
transform -1 0 5752 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_26
timestamp 1516238463
transform 1 0 5752 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_76
timestamp 1516238463
transform -1 0 5880 0 -1 610
box 0 0 64 200
use OR2X2  OR2X2_100
timestamp 1516238463
transform -1 0 5944 0 -1 610
box 0 0 64 200
use FILL  FILL_3_1
timestamp 1516238463
transform -1 0 5960 0 -1 610
box 0 0 16 200
use FILL  FILL_3_2
timestamp 1516238463
transform -1 0 5976 0 -1 610
box 0 0 16 200
use FILL  FILL_3_3
timestamp 1516238463
transform -1 0 5992 0 -1 610
box 0 0 16 200
use BUFX2  BUFX2_50
timestamp 1516238463
transform -1 0 56 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_15
timestamp 1516238463
transform -1 0 104 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1516238463
transform -1 0 296 0 1 210
box 0 0 192 200
use BUFX2  BUFX2_14
timestamp 1516238463
transform -1 0 344 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_19
timestamp 1516238463
transform -1 0 536 0 1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1516238463
transform -1 0 728 0 1 210
box 0 0 192 200
use INVX1  INVX1_13
timestamp 1516238463
transform -1 0 760 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1516238463
transform 1 0 760 0 1 210
box 0 0 192 200
use FILL  FILL_1_0_0
timestamp 1516238463
transform 1 0 952 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1516238463
transform 1 0 968 0 1 210
box 0 0 16 200
use AND2X2  AND2X2_593
timestamp 1516238463
transform 1 0 984 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_594
timestamp 1516238463
transform 1 0 1048 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_595
timestamp 1516238463
transform 1 0 1112 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_576
timestamp 1516238463
transform -1 0 1240 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1516238463
transform -1 0 1432 0 1 210
box 0 0 192 200
use AND2X2  AND2X2_564
timestamp 1516238463
transform -1 0 1496 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_563
timestamp 1516238463
transform -1 0 1560 0 1 210
box 0 0 64 200
use INVX1  INVX1_11
timestamp 1516238463
transform -1 0 1592 0 1 210
box 0 0 32 200
use AND2X2  AND2X2_562
timestamp 1516238463
transform -1 0 1656 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_96
timestamp 1516238463
transform -1 0 1720 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_26
timestamp 1516238463
transform -1 0 1784 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_176
timestamp 1516238463
transform 1 0 1784 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_289
timestamp 1516238463
transform 1 0 1848 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_127
timestamp 1516238463
transform -1 0 1976 0 1 210
box 0 0 64 200
use FILL  FILL_1_1_0
timestamp 1516238463
transform -1 0 1992 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1516238463
transform -1 0 2008 0 1 210
box 0 0 16 200
use NAND3X1  NAND3X1_19
timestamp 1516238463
transform -1 0 2072 0 1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1516238463
transform 1 0 2072 0 1 210
box 0 0 192 200
use OR2X2  OR2X2_208
timestamp 1516238463
transform 1 0 2264 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_329
timestamp 1516238463
transform -1 0 2392 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_21
timestamp 1516238463
transform -1 0 2440 0 1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1516238463
transform -1 0 2632 0 1 210
box 0 0 192 200
use AND2X2  AND2X2_575
timestamp 1516238463
transform -1 0 2696 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_573
timestamp 1516238463
transform -1 0 2760 0 1 210
box 0 0 64 200
use INVX1  INVX1_7
timestamp 1516238463
transform 1 0 2760 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_31
timestamp 1516238463
transform 1 0 2792 0 1 210
box 0 0 192 200
use FILL  FILL_1_2_0
timestamp 1516238463
transform -1 0 3000 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1516238463
transform -1 0 3016 0 1 210
box 0 0 16 200
use AND2X2  AND2X2_587
timestamp 1516238463
transform -1 0 3080 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_585
timestamp 1516238463
transform -1 0 3144 0 1 210
box 0 0 64 200
use INVX1  INVX1_24
timestamp 1516238463
transform 1 0 3144 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1516238463
transform 1 0 3176 0 1 210
box 0 0 192 200
use AND2X2  AND2X2_586
timestamp 1516238463
transform -1 0 3432 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_18
timestamp 1516238463
transform 1 0 3432 0 1 210
box 0 0 48 200
use INVX1  INVX1_22
timestamp 1516238463
transform 1 0 3480 0 1 210
box 0 0 32 200
use INVX1  INVX1_28
timestamp 1516238463
transform 1 0 3512 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_10
timestamp 1516238463
transform 1 0 3544 0 1 210
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_14
timestamp 1516238463
transform 1 0 3736 0 1 210
box 0 0 192 200
use AND2X2  AND2X2_571
timestamp 1516238463
transform -1 0 3992 0 1 210
box 0 0 64 200
use FILL  FILL_1_3_0
timestamp 1516238463
transform -1 0 4008 0 1 210
box 0 0 16 200
use FILL  FILL_1_3_1
timestamp 1516238463
transform -1 0 4024 0 1 210
box 0 0 16 200
use AND2X2  AND2X2_569
timestamp 1516238463
transform -1 0 4088 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_570
timestamp 1516238463
transform -1 0 4152 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_6
timestamp 1516238463
transform -1 0 4216 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_63
timestamp 1516238463
transform -1 0 4280 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_82
timestamp 1516238463
transform -1 0 4344 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_442
timestamp 1516238463
transform -1 0 4408 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_197
timestamp 1516238463
transform -1 0 4472 0 1 210
box 0 0 64 200
use INVX1  INVX1_5
timestamp 1516238463
transform 1 0 4472 0 1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_29
timestamp 1516238463
transform 1 0 4504 0 1 210
box 0 0 192 200
use AND2X2  AND2X2_167
timestamp 1516238463
transform 1 0 4696 0 1 210
box 0 0 64 200
use OR2X2  OR2X2_81
timestamp 1516238463
transform -1 0 4824 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_2
timestamp 1516238463
transform 1 0 4824 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_15
timestamp 1516238463
transform 1 0 4888 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_57
timestamp 1516238463
transform 1 0 4936 0 1 210
box 0 0 64 200
use FILL  FILL_1_4_0
timestamp 1516238463
transform 1 0 5000 0 1 210
box 0 0 16 200
use FILL  FILL_1_4_1
timestamp 1516238463
transform 1 0 5016 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_107
timestamp 1516238463
transform 1 0 5032 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_31
timestamp 1516238463
transform -1 0 5160 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_315
timestamp 1516238463
transform -1 0 5224 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_634
timestamp 1516238463
transform 1 0 5224 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_59
timestamp 1516238463
transform 1 0 5288 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_9
timestamp 1516238463
transform -1 0 5416 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_278
timestamp 1516238463
transform 1 0 5416 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_314
timestamp 1516238463
transform 1 0 5480 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_280
timestamp 1516238463
transform -1 0 5608 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_313
timestamp 1516238463
transform 1 0 5608 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_18
timestamp 1516238463
transform 1 0 5672 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_173
timestamp 1516238463
transform 1 0 5736 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_170
timestamp 1516238463
transform 1 0 5800 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_140
timestamp 1516238463
transform 1 0 5864 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_202
timestamp 1516238463
transform 1 0 5928 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_68
timestamp 1516238463
transform -1 0 56 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_33
timestamp 1516238463
transform -1 0 104 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_16
timestamp 1516238463
transform 1 0 104 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_51
timestamp 1516238463
transform 1 0 152 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_60
timestamp 1516238463
transform -1 0 248 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_49
timestamp 1516238463
transform -1 0 296 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_25
timestamp 1516238463
transform -1 0 344 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_46
timestamp 1516238463
transform -1 0 392 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_11
timestamp 1516238463
transform -1 0 440 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1516238463
transform -1 0 632 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_12
timestamp 1516238463
transform 1 0 632 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_47
timestamp 1516238463
transform 1 0 680 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_53
timestamp 1516238463
transform -1 0 792 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_50
timestamp 1516238463
transform -1 0 856 0 -1 210
box 0 0 64 200
use INVX1  INVX1_12
timestamp 1516238463
transform -1 0 888 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_36
timestamp 1516238463
transform -1 0 936 0 -1 210
box 0 0 48 200
use FILL  FILL_0_0_0
timestamp 1516238463
transform -1 0 952 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1516238463
transform -1 0 968 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_1
timestamp 1516238463
transform -1 0 1016 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_43
timestamp 1516238463
transform -1 0 1064 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_8
timestamp 1516238463
transform -1 0 1112 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_33
timestamp 1516238463
transform -1 0 1304 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_34
timestamp 1516238463
transform 1 0 1304 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_69
timestamp 1516238463
transform 1 0 1352 0 -1 210
box 0 0 48 200
use INVX1  INVX1_9
timestamp 1516238463
transform -1 0 1432 0 -1 210
box 0 0 32 200
use BUFX4  BUFX4_51
timestamp 1516238463
transform -1 0 1496 0 -1 210
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1516238463
transform 1 0 1496 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_10
timestamp 1516238463
transform 1 0 1688 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_45
timestamp 1516238463
transform 1 0 1736 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_44
timestamp 1516238463
transform 1 0 1784 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_9
timestamp 1516238463
transform -1 0 1880 0 -1 210
box 0 0 48 200
use FILL  FILL_0_1_0
timestamp 1516238463
transform -1 0 1896 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1516238463
transform -1 0 1912 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1516238463
transform -1 0 2104 0 -1 210
box 0 0 192 200
use INVX1  INVX1_10
timestamp 1516238463
transform -1 0 2136 0 -1 210
box 0 0 32 200
use AND2X2  AND2X2_572
timestamp 1516238463
transform 1 0 2136 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_56
timestamp 1516238463
transform -1 0 2248 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_22
timestamp 1516238463
transform 1 0 2248 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_57
timestamp 1516238463
transform 1 0 2296 0 -1 210
box 0 0 48 200
use INVX1  INVX1_14
timestamp 1516238463
transform 1 0 2344 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1516238463
transform 1 0 2376 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_13
timestamp 1516238463
transform 1 0 2568 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_48
timestamp 1516238463
transform 1 0 2616 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_574
timestamp 1516238463
transform -1 0 2728 0 -1 210
box 0 0 64 200
use INVX1  INVX1_8
timestamp 1516238463
transform 1 0 2728 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_32
timestamp 1516238463
transform 1 0 2760 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_7
timestamp 1516238463
transform 1 0 2952 0 -1 210
box 0 0 48 200
use FILL  FILL_0_2_0
timestamp 1516238463
transform 1 0 3000 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1516238463
transform 1 0 3016 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_42
timestamp 1516238463
transform 1 0 3032 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_6
timestamp 1516238463
transform 1 0 3080 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_41
timestamp 1516238463
transform 1 0 3128 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_49
timestamp 1516238463
transform -1 0 3240 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_54
timestamp 1516238463
transform 1 0 3240 0 -1 210
box 0 0 64 200
use INVX1  INVX1_27
timestamp 1516238463
transform 1 0 3304 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1516238463
transform 1 0 3336 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_19
timestamp 1516238463
transform 1 0 3528 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_54
timestamp 1516238463
transform 1 0 3576 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_53
timestamp 1516238463
transform 1 0 3624 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_38
timestamp 1516238463
transform 1 0 3672 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_3
timestamp 1516238463
transform -1 0 3768 0 -1 210
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_28
timestamp 1516238463
transform -1 0 3960 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_52
timestamp 1516238463
transform -1 0 4008 0 -1 210
box 0 0 48 200
use FILL  FILL_0_3_0
timestamp 1516238463
transform -1 0 4024 0 -1 210
box 0 0 16 200
use FILL  FILL_0_3_1
timestamp 1516238463
transform -1 0 4040 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_17
timestamp 1516238463
transform -1 0 4088 0 -1 210
box 0 0 48 200
use INVX1  INVX1_4
timestamp 1516238463
transform -1 0 4120 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_20
timestamp 1516238463
transform 1 0 4120 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_55
timestamp 1516238463
transform 1 0 4168 0 -1 210
box 0 0 48 200
use INVX1  INVX1_6
timestamp 1516238463
transform 1 0 4216 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_30
timestamp 1516238463
transform 1 0 4248 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_5
timestamp 1516238463
transform 1 0 4440 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_40
timestamp 1516238463
transform 1 0 4488 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_39
timestamp 1516238463
transform -1 0 4584 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_4
timestamp 1516238463
transform -1 0 4632 0 -1 210
box 0 0 48 200
use INVX1  INVX1_3
timestamp 1516238463
transform 1 0 4632 0 -1 210
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_23
timestamp 1516238463
transform 1 0 4664 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_2
timestamp 1516238463
transform 1 0 4856 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_37
timestamp 1516238463
transform 1 0 4904 0 -1 210
box 0 0 48 200
use OR2X2  OR2X2_162
timestamp 1516238463
transform 1 0 4952 0 -1 210
box 0 0 64 200
use FILL  FILL_0_4_0
timestamp 1516238463
transform -1 0 5032 0 -1 210
box 0 0 16 200
use FILL  FILL_0_4_1
timestamp 1516238463
transform -1 0 5048 0 -1 210
box 0 0 16 200
use AND2X2  AND2X2_281
timestamp 1516238463
transform -1 0 5112 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_440
timestamp 1516238463
transform -1 0 5176 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_10
timestamp 1516238463
transform -1 0 5240 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_432
timestamp 1516238463
transform -1 0 5304 0 -1 210
box 0 0 64 200
use INVX4  INVX4_1
timestamp 1516238463
transform -1 0 5352 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_27
timestamp 1516238463
transform -1 0 5416 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_164
timestamp 1516238463
transform -1 0 5480 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_174
timestamp 1516238463
transform -1 0 5544 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_163
timestamp 1516238463
transform -1 0 5608 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_195
timestamp 1516238463
transform 1 0 5608 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_196
timestamp 1516238463
transform 1 0 5672 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_439
timestamp 1516238463
transform -1 0 5800 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_80
timestamp 1516238463
transform -1 0 5864 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_102
timestamp 1516238463
transform 1 0 5864 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_600
timestamp 1516238463
transform 1 0 5928 0 -1 210
box 0 0 64 200
<< labels >>
flabel space 1156 42 1164 136 6 FreeSans 48 0 0 0 vdd
port 0 nsew
flabel space 2164 42 2172 136 6 FreeSans 48 0 0 0 gnd
port 1 nsew
flabel metal2 3136 4060 3136 4060 3 FreeSans 48 90 0 0 ULA_A<0>
port 2 nsew
flabel metal2 3488 4060 3488 4060 3 FreeSans 48 90 0 0 ULA_A<1>
port 3 nsew
flabel metal2 3536 4060 3536 4060 3 FreeSans 48 90 0 0 ULA_A<2>
port 4 nsew
flabel metal2 3616 4060 3616 4060 3 FreeSans 48 90 0 0 ULA_A<3>
port 5 nsew
flabel metal2 3664 4060 3664 4060 3 FreeSans 48 90 0 0 ULA_A<4>
port 6 nsew
flabel metal2 3024 4060 3024 4060 3 FreeSans 48 90 0 0 ULA_A<5>
port 7 nsew
flabel metal2 3312 4060 3312 4060 3 FreeSans 48 90 0 0 ULA_A<6>
port 8 nsew
flabel metal2 2096 -40 2096 -40 7 FreeSans 48 270 0 0 ULA_A<7>
port 9 nsew
flabel metal2 3408 4060 3408 4060 3 FreeSans 48 90 0 0 ULA_A<8>
port 10 nsew
flabel metal2 2624 4060 2624 4060 3 FreeSans 48 90 0 0 ULA_A<9>
port 11 nsew
flabel metal2 1824 -40 1824 -40 7 FreeSans 48 270 0 0 ULA_A<10>
port 12 nsew
flabel metal2 2880 4060 2880 4060 3 FreeSans 48 90 0 0 ULA_A<11>
port 13 nsew
flabel metal2 3712 4060 3712 4060 3 FreeSans 48 90 0 0 ULA_A<12>
port 14 nsew
flabel metal2 2256 4060 2256 4060 3 FreeSans 48 90 0 0 ULA_A<13>
port 15 nsew
flabel metal2 1200 4060 1200 4060 3 FreeSans 48 90 0 0 ULA_A<14>
port 16 nsew
flabel metal3 -48 2160 -48 2160 7 FreeSans 48 0 0 0 ULA_A<15>
port 17 nsew
flabel metal2 2800 4060 2800 4060 3 FreeSans 48 90 0 0 ULA_A<16>
port 18 nsew
flabel metal2 2832 4060 2832 4060 3 FreeSans 48 90 0 0 ULA_A<17>
port 19 nsew
flabel metal2 2752 4060 2752 4060 3 FreeSans 48 90 0 0 ULA_A<18>
port 20 nsew
flabel metal2 2208 4060 2208 4060 3 FreeSans 48 90 0 0 ULA_A<19>
port 21 nsew
flabel metal2 2112 4060 2112 4060 3 FreeSans 48 90 0 0 ULA_A<20>
port 22 nsew
flabel metal2 4000 4060 4000 4060 3 FreeSans 48 90 0 0 ULA_A<21>
port 23 nsew
flabel metal2 2400 4060 2400 4060 3 FreeSans 48 90 0 0 ULA_A<22>
port 24 nsew
flabel metal2 896 4060 896 4060 3 FreeSans 48 90 0 0 ULA_A<23>
port 25 nsew
flabel metal2 448 4060 448 4060 3 FreeSans 48 90 0 0 ULA_A<24>
port 26 nsew
flabel metal2 4048 4060 4048 4060 3 FreeSans 48 90 0 0 ULA_A<25>
port 27 nsew
flabel metal2 4176 4060 4176 4060 3 FreeSans 48 90 0 0 ULA_A<26>
port 28 nsew
flabel metal2 496 4060 496 4060 3 FreeSans 48 90 0 0 ULA_A<27>
port 29 nsew
flabel metal2 4368 4060 4368 4060 3 FreeSans 48 90 0 0 ULA_A<28>
port 30 nsew
flabel metal2 3760 4060 3760 4060 3 FreeSans 48 90 0 0 ULA_A<29>
port 31 nsew
flabel metal2 3888 4060 3888 4060 3 FreeSans 48 90 0 0 ULA_A<30>
port 32 nsew
flabel metal3 -48 1800 -48 1800 7 FreeSans 48 0 0 0 ULA_A<31>
port 33 nsew
flabel metal2 2976 4060 2976 4060 3 FreeSans 48 90 0 0 ULA_B<0>
port 34 nsew
flabel metal2 4864 4060 4864 4060 3 FreeSans 48 90 0 0 ULA_B<1>
port 35 nsew
flabel metal2 1488 4060 1488 4060 3 FreeSans 48 90 0 0 ULA_B<2>
port 36 nsew
flabel metal3 -48 2520 -48 2520 7 FreeSans 48 0 0 0 ULA_B<3>
port 37 nsew
flabel metal3 -48 2320 -48 2320 7 FreeSans 48 0 0 0 ULA_B<4>
port 38 nsew
flabel metal2 2576 -40 2576 -40 7 FreeSans 48 270 0 0 ULA_B<5>
port 39 nsew
flabel metal2 3120 -40 3120 -40 7 FreeSans 48 270 0 0 ULA_B<6>
port 40 nsew
flabel metal2 2048 -40 2048 -40 7 FreeSans 48 270 0 0 ULA_B<7>
port 41 nsew
flabel metal2 1696 -40 1696 -40 7 FreeSans 48 270 0 0 ULA_B<8>
port 42 nsew
flabel metal2 3792 -40 3792 -40 7 FreeSans 48 270 0 0 ULA_B<9>
port 43 nsew
flabel metal2 1856 -40 1856 -40 7 FreeSans 48 270 0 0 ULA_B<10>
port 44 nsew
flabel metal2 1232 -40 1232 -40 7 FreeSans 48 270 0 0 ULA_B<11>
port 45 nsew
flabel metal2 2384 -40 2384 -40 7 FreeSans 48 270 0 0 ULA_B<12>
port 46 nsew
flabel metal2 1936 -40 1936 -40 7 FreeSans 48 270 0 0 ULA_B<13>
port 47 nsew
flabel metal2 1184 -40 1184 -40 7 FreeSans 48 270 0 0 ULA_B<14>
port 48 nsew
flabel metal3 -48 1860 -48 1860 7 FreeSans 48 0 0 0 ULA_B<15>
port 49 nsew
flabel metal2 3664 -40 3664 -40 7 FreeSans 48 270 0 0 ULA_B<16>
port 50 nsew
flabel metal2 2928 4060 2928 4060 3 FreeSans 48 90 0 0 ULA_B<17>
port 51 nsew
flabel metal2 3200 4060 3200 4060 3 FreeSans 48 90 0 0 ULA_B<18>
port 52 nsew
flabel metal2 3216 -40 3216 -40 7 FreeSans 48 270 0 0 ULA_B<19>
port 53 nsew
flabel metal2 2976 -40 2976 -40 7 FreeSans 48 270 0 0 ULA_B<20>
port 54 nsew
flabel metal2 1984 -40 1984 -40 7 FreeSans 48 270 0 0 ULA_B<21>
port 55 nsew
flabel metal2 3584 4060 3584 4060 3 FreeSans 48 90 0 0 ULA_B<22>
port 56 nsew
flabel metal3 -48 1680 -48 1680 7 FreeSans 48 0 0 0 ULA_B<23>
port 57 nsew
flabel metal3 -48 2120 -48 2120 7 FreeSans 48 0 0 0 ULA_B<24>
port 58 nsew
flabel metal2 2256 -40 2256 -40 7 FreeSans 48 270 0 0 ULA_B<25>
port 59 nsew
flabel metal3 -48 1760 -48 1760 7 FreeSans 48 0 0 0 ULA_B<26>
port 60 nsew
flabel metal3 -48 1940 -48 1940 7 FreeSans 48 0 0 0 ULA_B<27>
port 61 nsew
flabel metal3 -48 1520 -48 1520 7 FreeSans 48 0 0 0 ULA_B<28>
port 62 nsew
flabel metal2 1616 -40 1616 -40 7 FreeSans 48 270 0 0 ULA_B<29>
port 63 nsew
flabel metal3 -48 1280 -48 1280 7 FreeSans 48 0 0 0 ULA_B<30>
port 64 nsew
flabel metal3 -48 1720 -48 1720 7 FreeSans 48 0 0 0 ULA_B<31>
port 65 nsew
flabel metal2 1136 -40 1136 -40 7 FreeSans 48 270 0 0 ULA_ctrl<0>
port 66 nsew
flabel metal2 1744 -40 1744 -40 7 FreeSans 48 270 0 0 ULA_ctrl<1>
port 67 nsew
flabel metal2 2432 -40 2432 -40 7 FreeSans 48 270 0 0 ULA_ctrl<2>
port 68 nsew
flabel metal2 2480 -40 2480 -40 7 FreeSans 48 270 0 0 ULA_ctrl<3>
port 69 nsew
flabel metal2 3264 -40 3264 -40 7 FreeSans 48 270 0 0 clk
port 70 nsew
flabel metal2 896 -40 896 -40 7 FreeSans 48 270 0 0 ULA_OUT<0>
port 71 nsew
flabel metal2 4944 -40 4944 -40 7 FreeSans 48 270 0 0 ULA_OUT<1>
port 72 nsew
flabel metal2 3744 -40 3744 -40 7 FreeSans 48 270 0 0 ULA_OUT<2>
port 73 nsew
flabel metal2 4576 -40 4576 -40 7 FreeSans 48 270 0 0 ULA_OUT<3>
port 74 nsew
flabel metal2 4528 -40 4528 -40 7 FreeSans 48 270 0 0 ULA_OUT<4>
port 75 nsew
flabel metal2 3168 -40 3168 -40 7 FreeSans 48 270 0 0 ULA_OUT<5>
port 76 nsew
flabel metal2 3072 -40 3072 -40 7 FreeSans 48 270 0 0 ULA_OUT<6>
port 77 nsew
flabel metal2 992 -40 992 -40 7 FreeSans 48 270 0 0 ULA_OUT<7>
port 78 nsew
flabel metal2 1904 -40 1904 -40 7 FreeSans 48 270 0 0 ULA_OUT<8>
port 79 nsew
flabel metal2 1776 -40 1776 -40 7 FreeSans 48 270 0 0 ULA_OUT<9>
port 80 nsew
flabel metal2 352 -40 352 -40 7 FreeSans 48 270 0 0 ULA_OUT<10>
port 81 nsew
flabel metal2 720 -40 720 -40 7 FreeSans 48 270 0 0 ULA_OUT<11>
port 82 nsew
flabel metal2 2656 -40 2656 -40 7 FreeSans 48 270 0 0 ULA_OUT<12>
port 83 nsew
flabel metal2 272 -40 272 -40 7 FreeSans 48 270 0 0 ULA_OUT<13>
port 84 nsew
flabel metal3 -48 320 -48 320 7 FreeSans 48 0 0 0 ULA_OUT<14>
port 85 nsew
flabel metal2 192 -40 192 -40 7 FreeSans 48 270 0 0 ULA_OUT<15>
port 86 nsew
flabel metal2 3968 -40 3968 -40 7 FreeSans 48 270 0 0 ULA_OUT<16>
port 87 nsew
flabel metal2 3712 -40 3712 -40 7 FreeSans 48 270 0 0 ULA_OUT<17>
port 88 nsew
flabel metal2 3616 -40 3616 -40 7 FreeSans 48 270 0 0 ULA_OUT<18>
port 89 nsew
flabel metal2 4208 -40 4208 -40 7 FreeSans 48 270 0 0 ULA_OUT<19>
port 90 nsew
flabel metal2 2208 -40 2208 -40 7 FreeSans 48 270 0 0 ULA_OUT<20>
port 91 nsew
flabel metal2 2336 -40 2336 -40 7 FreeSans 48 270 0 0 ULA_OUT<21>
port 92 nsew
flabel metal3 -48 1120 -48 1120 7 FreeSans 48 0 0 0 ULA_OUT<22>
port 93 nsew
flabel metal3 -48 1600 -48 1600 7 FreeSans 48 0 0 0 ULA_OUT<23>
port 94 nsew
flabel metal2 240 -40 240 -40 7 FreeSans 48 270 0 0 ULA_OUT<24>
port 95 nsew
flabel metal3 -48 1560 -48 1560 7 FreeSans 48 0 0 0 ULA_OUT<25>
port 96 nsew
flabel metal3 -48 720 -48 720 7 FreeSans 48 0 0 0 ULA_OUT<26>
port 97 nsew
flabel metal3 -48 1160 -48 1160 7 FreeSans 48 0 0 0 ULA_OUT<27>
port 98 nsew
flabel metal3 -48 1320 -48 1320 7 FreeSans 48 0 0 0 ULA_OUT<28>
port 99 nsew
flabel metal3 -48 920 -48 920 7 FreeSans 48 0 0 0 ULA_OUT<29>
port 100 nsew
flabel metal3 -48 960 -48 960 7 FreeSans 48 0 0 0 ULA_OUT<30>
port 101 nsew
flabel metal3 -48 520 -48 520 7 FreeSans 48 0 0 0 ULA_OUT<31>
port 102 nsew
flabel metal3 -48 120 -48 120 7 FreeSans 48 0 0 0 ULA_flags<0>
port 103 nsew
flabel metal2 1392 -40 1392 -40 7 FreeSans 48 270 0 0 ULA_flags<1>
port 104 nsew
flabel metal2 5856 4060 5856 4060 3 FreeSans 48 90 0 0 ULA_flags<2>
port 105 nsew
<< end >>
