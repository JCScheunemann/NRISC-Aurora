module NRISC_InstructionDecoder ( gnd, vdd, CORE_InstructionIN, CORE_ctrl, CORE_ULA_flags, clk, rst, CORE_InstructionToULAMux, CORE_Status_ctrl, CORE_ULA_ctrl, CORE_ULAMux_inc_dec, CORE_REG_RF1, CORE_REG_RF2, CORE_REG_RD, CORE_REG_write, CORE_DATA_write, CORE_DATA_load, CORE_DATA_ctrl, CORE_DATA_ADDR_mux, CORE_DATA_REGMux, CORE_STACK_ctrl, CORE_PC_ctrl, CORE_PC_clk, CORE_INT_CHA, CORE_INT_ctrl);

input gnd, vdd;
input clk;
input rst;
output CORE_ULAMux_inc_dec;
output CORE_REG_write;
output CORE_DATA_write;
output CORE_DATA_load;
output CORE_DATA_ADDR_mux;
output CORE_DATA_REGMux;
output CORE_PC_clk;
input [15:0] CORE_InstructionIN;
input [2:0] CORE_ctrl;
input [2:0] CORE_ULA_flags;
output [1:0] CORE_InstructionToULAMux;
output [4:0] CORE_Status_ctrl;
output [3:0] CORE_ULA_ctrl;
output [3:0] CORE_REG_RF1;
output [3:0] CORE_REG_RF2;
output [3:0] CORE_REG_RD;
output [2:0] CORE_DATA_ctrl;
output [1:0] CORE_STACK_ctrl;
output [1:0] CORE_PC_ctrl;
output [7:0] CORE_INT_CHA;
output [1:0] CORE_INT_ctrl;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_16__bF_buf4) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_16__bF_buf3) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_16__bF_buf2) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_16__bF_buf1) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_16__bF_buf0) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf3) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf2) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf1) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[15]), .Y(CORE_InstructionIN_15_bF_buf0) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf0), .Y(_16_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .Y(_17_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[13]), .Y(_18_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(CORE_InstructionIN[12]), .Y(_19_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_18_), .Y(_20_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf2), .B(_17_), .C(_20_), .Y(_21_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_211__0_), .B(CORE_InstructionIN[14]), .Y(_22_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[10]), .Y(_23_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[9]), .Y(_24_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .B(_24_), .C(_23_), .Y(_25_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_211__0_), .B(_23_), .C(_25_), .Y(_26_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf2), .B(_22_), .C(_26_), .D(_21_), .Y(_6__0_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .Y(_27_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf3), .B(_27_), .Y(_28_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_211__1_), .B(_28_), .Y(_29_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[9]), .C(CORE_InstructionIN[10]), .Y(_30_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_31_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_211__1_), .C(_31_), .Y(_32_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_21_), .C(_29_), .Y(_6__1_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_210__0_), .Y(_33_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[0]), .Y(_34_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[9]), .B(_23_), .Y(_35_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_21_), .Y(_36_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_33_), .S(_36_), .Y(_5__0_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_210__1_), .Y(_37_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[1]), .Y(_38_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_37_), .S(_36_), .Y(_5__1_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_210__2_), .Y(_39_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[2]), .Y(_40_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_39_), .S(_36_), .Y(_5__2_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_210__3_), .Y(_41_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[3]), .Y(_42_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_41_), .S(_36_), .Y(_5__3_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_210__4_), .Y(_43_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[4]), .Y(_44_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_43_), .S(_36_), .Y(_5__4_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_210__5_), .Y(_45_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[5]), .Y(_46_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_45_), .S(_36_), .Y(_5__5_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_210__6_), .Y(_47_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[6]), .Y(_48_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_47_), .S(_36_), .Y(_5__6_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_210__7_), .Y(_49_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[7]), .Y(_50_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_49_), .S(_36_), .Y(_5__7_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .B(CORE_ULA_flags[1]), .C(_24_), .Y(_51_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[9]), .C(CORE_ULA_flags[0]), .Y(_52_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .Y(_53_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(CORE_ULA_flags[2]), .B(_24_), .C(_53_), .Y(_54_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_52_), .C(_54_), .Y(_55_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_213__0_), .Y(_56_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[12]), .B(_27_), .C(_18_), .Y(_57_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_56_), .C(_57_), .Y(_58_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_55_), .C(_58_), .Y(_59_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(CORE_InstructionIN[11]), .C(_19_), .Y(_60_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_60_), .Y(_61_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_24_), .Y(_62_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_62_), .C(_31_), .Y(_63_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_213__0_), .C(_61_), .D(_63_), .Y(_64_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_59_), .C(CORE_InstructionIN_15_bF_buf1), .Y(_8__0_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_213__1_), .Y(_65_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_61_), .Y(_66_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_57_), .Y(_67_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_60_), .C(_27_), .Y(_68_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_68_), .C(_16__bF_buf4), .Y(_69_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(_69_), .Y(_8__1_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_24_), .C(_218__0_), .Y(_70_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_31_), .Y(_71_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_218__0_), .C(_61_), .D(_71_), .Y(_72_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf1), .B(_72_), .Y(_13__0_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_218__1_), .Y(_73_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_60_), .Y(_74_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_74_), .C(_16__bF_buf4), .Y(_75_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_66_), .C(_75_), .Y(_13__1_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[2]), .B(_38_), .C(_42_), .Y(_76_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[0]), .B(CORE_InstructionIN[1]), .Y(_77_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[2]), .B(CORE_InstructionIN[3]), .Y(_78_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_79_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_79_), .C(_76_), .Y(_80_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_78_), .Y(_81_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_81_), .C(_80_), .Y(_82_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[13]), .B(_19_), .Y(_83_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_84_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf2), .B(_84_), .Y(_85_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_28_), .Y(_86_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_82_), .C(_86_), .Y(_1_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_18_), .Y(_87_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf3), .B(_88_), .C(_207__0_), .Y(_89_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[13]), .B(CORE_InstructionIN[12]), .Y(_90_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_90_), .Y(_91_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_207__0_), .Y(_92_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[0]), .B(CORE_InstructionIN[1]), .C(_78_), .Y(_93_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_76_), .C(_93_), .Y(_94_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[1]), .B(_34_), .Y(_95_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[13]), .B(_19_), .C(_76_), .Y(_96_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_95_), .C(_96_), .Y(_97_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_17_), .Y(_98_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_17_), .C(_92_), .D(_98_), .Y(_99_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_99_), .C(_94_), .D(_97_), .Y(_100_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf3), .B(_100_), .C(_89_), .Y(_2__0_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .Y(_101_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf3), .B(_88_), .Y(_102_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_35_), .C(_101_), .D(_98_), .Y(_103_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_101_), .C(_83_), .Y(_104_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_91_), .C(_93_), .D(_104_), .Y(_105_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_102_), .C(CORE_InstructionIN_15_bF_buf3), .D(_105_), .Y(_2__1_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf2), .B(_88_), .C(_207__2_), .Y(_106_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_207__2_), .Y(_107_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_76_), .C(_93_), .Y(_108_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[3]), .B(_40_), .Y(_109_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[0]), .B(_40_), .C(_42_), .Y(_110_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[13]), .B(_19_), .C(_110_), .Y(_111_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_95_), .C(_111_), .Y(_112_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[10]), .B(CORE_InstructionIN[11]), .Y(_113_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_107_), .C(_113_), .Y(_114_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_114_), .C(_108_), .D(_112_), .Y(_115_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf2), .B(_115_), .C(_106_), .Y(_2__2_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[12]), .Y(_116_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_116_), .C(_27_), .Y(_117_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_27_), .C(_16__bF_buf3), .Y(_119_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_118_), .Y(_0_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_208_), .Y(_120_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_208_), .Y(_121_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_121_), .C(_84_), .Y(_122_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_120_), .C(CORE_InstructionIN_15_bF_buf2), .Y(_3_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_27_), .C(_16__bF_buf3), .Y(_123_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_118_), .Y(_4_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_116_), .C(_16__bF_buf1), .Y(_124_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_30_), .C(_124_), .Y(_125_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_30_), .Y(_126_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_126_), .C(CORE_InstructionIN[14]), .Y(_127_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_216__0_), .B(_16__bF_buf1), .Y(_128_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_128_), .C(_34_), .D(_125_), .Y(_11__0_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_216__1_), .B(_16__bF_buf1), .Y(_129_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_129_), .C(_38_), .D(_125_), .Y(_11__1_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_216__2_), .B(_16__bF_buf3), .Y(_130_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_130_), .C(_40_), .D(_125_), .Y(_11__2_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_216__3_), .B(_16__bF_buf1), .Y(_131_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_131_), .C(_42_), .D(_125_), .Y(_11__3_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_17_), .Y(_132_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_30_), .C(CORE_InstructionIN_15_bF_buf0), .Y(_133_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_215__0_), .Y(_134_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_19_), .Y(_135_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_134_), .C(_135_), .Y(_136_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[4]), .B(_133_), .C(_136_), .Y(_137_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf1), .B(_87_), .C(CORE_InstructionIN[4]), .Y(_138_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_134_), .C(_57_), .Y(_139_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf1), .B(_113_), .C(_44_), .Y(_140_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_215__0_), .B(_28_), .C(_140_), .D(_139_), .Y(_141_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_141_), .C(_137_), .Y(_10__0_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_57_), .C(_127_), .Y(_142_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf4), .B(_215__1_), .Y(_143_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_142_), .Y(_144_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .B(_30_), .Y(_145_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_60_), .Y(_146_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_147_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_18_), .C(_16__bF_buf2), .Y(_148_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_149_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_57_), .C(_149_), .Y(_150_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_150_), .C(CORE_InstructionIN[5]), .Y(_151_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_144_), .Y(_10__1_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf4), .B(_215__2_), .Y(_152_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_142_), .Y(_153_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_150_), .C(CORE_InstructionIN[6]), .Y(_154_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_153_), .Y(_10__2_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf4), .B(_215__3_), .Y(_155_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_142_), .Y(_156_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_150_), .C(CORE_InstructionIN[7]), .Y(_157_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_156_), .Y(_10__3_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_214__0_), .B(_148_), .Y(_158_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_148_), .C(_158_), .Y(_9__0_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_214__1_), .B(_148_), .Y(_159_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_148_), .C(_159_), .Y(_9__1_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_214__2_), .B(_148_), .Y(_160_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_148_), .C(_160_), .Y(_9__2_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_214__3_), .Y(_161_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_149_), .C(_17_), .D(_102_), .Y(_9__3_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_126_), .C(_117_), .Y(_162_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(_163_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(CORE_InstructionIN[11]), .C(_163_), .Y(_164_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_220__0_), .B(_16__bF_buf3), .Y(_165_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_165_), .C(_16__bF_buf3), .D(_164_), .Y(_15__0_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_116_), .C(_83_), .Y(_166_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_91_), .C(_166_), .Y(_167_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_220__1_), .B(_16__bF_buf0), .Y(_168_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_168_), .C(_16__bF_buf0), .D(_167_), .Y(_15__1_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(CORE_InstructionIN[12]), .C(CORE_InstructionIN[13]), .Y(_169_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_220__2_), .B(_16__bF_buf3), .Y(_170_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf1), .B(_169_), .C(_170_), .D(_162_), .Y(_15__2_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_220__3_), .B(_16__bF_buf0), .Y(_171_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf0), .B(_27_), .C(_171_), .D(_162_), .Y(_15__3_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf2), .B(_20_), .Y(_172_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(CORE_InstructionIN[8]), .Y(_173_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf2), .B(_87_), .C(_173_), .D(_172_), .Y(_174_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_174_), .Y(_175_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[11]), .B(_163_), .Y(_176_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_176_), .Y(_177_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_212__0_), .B(_16__bF_buf0), .Y(_178_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_175_), .Y(_7__0_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_212__1_), .B(_117_), .Y(_179_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_212__1_), .Y(_180_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_126_), .C(_180_), .Y(_181_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_67_), .C(_181_), .Y(_182_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_179_), .C(CORE_InstructionIN_15_bF_buf0), .Y(_7__1_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[1]), .B(_110_), .Y(_183_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[4]), .B(CORE_InstructionIN[5]), .Y(_184_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[6]), .B(CORE_InstructionIN[7]), .Y(_185_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_185_), .Y(_186_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_145_), .Y(_187_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_187_), .Y(_188_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_188_), .C(_219__0_), .Y(_189_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_78_), .C(_187_), .Y(_190_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_190_), .C(_189_), .Y(_14__0_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_219__1_), .Y(_191_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[0]), .B(CORE_InstructionIN[1]), .Y(_192_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_79_), .Y(_193_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN_15_bF_buf0), .B(_135_), .Y(_194_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_24_), .C(_113_), .Y(_195_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_195_), .Y(_196_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_196_), .Y(_197_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_197_), .Y(_198_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[0]), .B(CORE_InstructionIN[1]), .C(_93_), .Y(_199_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_199_), .C(_196_), .Y(_200_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_191_), .C(_193_), .D(_198_), .Y(_14__1_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_219__2_), .B(_200_), .Y(_201_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_197_), .C(_201_), .Y(_14__2_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[8]), .B(CORE_InstructionIN[9]), .C(_98_), .Y(_202_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_172_), .C(_219__3_), .Y(_203_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(_14__3_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(CORE_InstructionIN[14]), .B(_74_), .C(_217_), .Y(_204_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_16__bF_buf4), .B(_83_), .C(_204_), .Y(_12_) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_205_), .Y(CORE_DATA_ADDR_mux) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_206_), .Y(CORE_DATA_REGMux) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_207__0_), .Y(CORE_DATA_ctrl[0]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .Y(CORE_DATA_ctrl[1]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_207__2_), .Y(CORE_DATA_ctrl[2]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_208_), .Y(CORE_DATA_load) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_209_), .Y(CORE_DATA_write) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_210__0_), .Y(CORE_INT_CHA[0]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_210__1_), .Y(CORE_INT_CHA[1]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_210__2_), .Y(CORE_INT_CHA[2]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_210__3_), .Y(CORE_INT_CHA[3]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_210__4_), .Y(CORE_INT_CHA[4]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_210__5_), .Y(CORE_INT_CHA[5]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_210__6_), .Y(CORE_INT_CHA[6]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_210__7_), .Y(CORE_INT_CHA[7]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_211__0_), .Y(CORE_INT_ctrl[0]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_211__1_), .Y(CORE_INT_ctrl[1]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_212__0_), .Y(CORE_InstructionToULAMux[0]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_212__1_), .Y(CORE_InstructionToULAMux[1]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(CORE_PC_clk) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_213__0_), .Y(CORE_PC_ctrl[0]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_213__1_), .Y(CORE_PC_ctrl[1]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_214__0_), .Y(CORE_REG_RD[0]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_214__1_), .Y(CORE_REG_RD[1]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_214__2_), .Y(CORE_REG_RD[2]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_214__3_), .Y(CORE_REG_RD[3]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_215__0_), .Y(CORE_REG_RF1[0]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_215__1_), .Y(CORE_REG_RF1[1]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_215__2_), .Y(CORE_REG_RF1[2]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_215__3_), .Y(CORE_REG_RF1[3]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_216__0_), .Y(CORE_REG_RF2[0]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_216__1_), .Y(CORE_REG_RF2[1]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_216__2_), .Y(CORE_REG_RF2[2]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_216__3_), .Y(CORE_REG_RF2[3]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(CORE_REG_write) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_218__0_), .Y(CORE_STACK_ctrl[0]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_218__1_), .Y(CORE_STACK_ctrl[1]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_219__0_), .Y(CORE_Status_ctrl[0]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_219__1_), .Y(CORE_Status_ctrl[1]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_219__2_), .Y(CORE_Status_ctrl[2]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_219__3_), .Y(CORE_Status_ctrl[3]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(CORE_Status_ctrl[4]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(CORE_ULAMux_inc_dec) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_220__0_), .Y(CORE_ULA_ctrl[0]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_220__1_), .Y(CORE_ULA_ctrl[1]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_220__2_), .Y(CORE_ULA_ctrl[2]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_220__3_), .Y(CORE_ULA_ctrl[3]) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_14__0_), .Q(_219__0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_14__1_), .Q(_219__1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_14__2_), .Q(_219__2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_14__3_), .Q(_219__3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_7__0_), .Q(_212__0_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_7__1_), .Q(_212__1_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_15__0_), .Q(_220__0_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_15__1_), .Q(_220__1_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_15__2_), .Q(_220__2_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_15__3_), .Q(_220__3_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_9__0_), .Q(_214__0_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_9__1_), .Q(_214__1_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_9__2_), .Q(_214__2_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_9__3_), .Q(_214__3_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_10__0_), .Q(_215__0_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_10__1_), .Q(_215__1_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_10__2_), .Q(_215__2_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_10__3_), .Q(_215__3_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_11__0_), .Q(_216__0_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_11__1_), .Q(_216__1_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_11__2_), .Q(_216__2_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_11__3_), .Q(_216__3_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_12_), .Q(_217_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_4_), .Q(_209_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3_), .Q(_208_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0_), .Q(_205_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2__0_), .Q(_207__0_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2__1_), .Q(_207__1_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2__2_), .Q(_207__2_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_1_), .Q(_206_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_13__0_), .Q(_218__0_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_13__1_), .Q(_218__1_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_8__0_), .Q(_213__0_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8__1_), .Q(_213__1_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_5__0_), .Q(_210__0_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_5__1_), .Q(_210__1_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_5__2_), .Q(_210__2_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_5__3_), .Q(_210__3_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_5__4_), .Q(_210__4_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_5__5_), .Q(_210__5_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_5__6_), .Q(_210__6_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_5__7_), .Q(_210__7_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__0_), .Q(_211__0_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6__1_), .Q(_211__1_) );
endmodule
