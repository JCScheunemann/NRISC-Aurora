module NRISC_ULA ( gnd, vdd, ULA_A, ULA_B, ULA_ctrl, clk, ULA_OUT, ULA_flags);

input gnd, vdd;
input clk;
input [31:0] ULA_A;
input [31:0] ULA_B;
input [3:0] ULA_ctrl;
output [31:0] ULA_OUT;
output [2:0] ULA_flags;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(ULA_ctrl_1_bF_buf5) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(ULA_ctrl_1_bF_buf4) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(ULA_ctrl_1_bF_buf3) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(ULA_ctrl_1_bF_buf2) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(ULA_ctrl_1_bF_buf1) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[1]), .Y(ULA_ctrl_1_bF_buf0) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_447_), .Y(_447__bF_buf3) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_447_), .Y(_447__bF_buf2) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_447_), .Y(_447__bF_buf1) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_447_), .Y(_447__bF_buf0) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_212__bF_buf5) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_212__bF_buf4) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_212__bF_buf3) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_212__bF_buf2) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_212__bF_buf1) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_212__bF_buf0) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_664_), .Y(_664__bF_buf4) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_664_), .Y(_664__bF_buf3) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_664_), .Y(_664__bF_buf2) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_664_), .Y(_664__bF_buf1) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_664_), .Y(_664__bF_buf0) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_244_), .Y(_244__bF_buf3) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_244_), .Y(_244__bF_buf2) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_244_), .Y(_244__bF_buf1) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_244_), .Y(_244__bF_buf0) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf7) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf6) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf5) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf4) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf3) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf2) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf1) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[3]), .Y(ULA_B_3_bF_buf0) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_74__bF_buf4) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_74__bF_buf3) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_74__bF_buf2) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_74__bF_buf1) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_74__bF_buf0) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_106__bF_buf4) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_106__bF_buf3) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_106__bF_buf2) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_106__bF_buf1) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_106__bF_buf0) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf7) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf6) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf5) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf4) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf3) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf2) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf1) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[0]), .Y(ULA_B_0_bF_buf0) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_138__bF_buf4) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_138__bF_buf3) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_138__bF_buf2) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_138__bF_buf1) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_138__bF_buf0) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_458_), .Y(_458__bF_buf3) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_458_), .Y(_458__bF_buf2) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_458_), .Y(_458__bF_buf1) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_458_), .Y(_458__bF_buf0) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_705__bF_buf4) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_705__bF_buf3) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_705__bF_buf2) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_705__bF_buf1) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(_705_), .Y(_705__bF_buf0) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf6) );
BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf5) );
BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf4) );
BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf3) );
BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf2) );
BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf1) );
BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(_684_), .Y(_684__bF_buf0) );
BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_490__bF_buf4) );
BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_490__bF_buf3) );
BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_490__bF_buf2) );
BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_490__bF_buf1) );
BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_490__bF_buf0) );
BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf5) );
BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf4) );
BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf3) );
BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf2) );
BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf1) );
BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf0) );
BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf6) );
BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf5) );
BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf4) );
BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf3) );
BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf2) );
BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf1) );
BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_255__bF_buf0) );
BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_149__bF_buf4) );
BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_149__bF_buf3) );
BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_149__bF_buf2) );
BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_149__bF_buf1) );
BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_149__bF_buf0) );
BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_340__bF_buf5) );
BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_340__bF_buf4) );
BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_340__bF_buf3) );
BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_340__bF_buf2) );
BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_340__bF_buf1) );
BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_340__bF_buf0) );
BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf7) );
BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf6) );
BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf5) );
BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf4) );
BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf3) );
BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf2) );
BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf1) );
BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[2]), .Y(ULA_B_2_bF_buf0) );
BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(_842_), .Y(_842__bF_buf3) );
BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(_842_), .Y(_842__bF_buf2) );
BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(_842_), .Y(_842__bF_buf1) );
BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(_842_), .Y(_842__bF_buf0) );
BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(_639_), .Y(_639__bF_buf3) );
BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(_639_), .Y(_639__bF_buf2) );
BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(_639_), .Y(_639__bF_buf1) );
BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(_639_), .Y(_639__bF_buf0) );
BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[4]), .Y(ULA_B_4_bF_buf3) );
BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[4]), .Y(ULA_B_4_bF_buf2) );
BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[4]), .Y(ULA_B_4_bF_buf1) );
BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[4]), .Y(ULA_B_4_bF_buf0) );
BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf7) );
BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf6) );
BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf5) );
BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf4) );
BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf3) );
BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf2) );
BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf1) );
BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[1]), .Y(ULA_B_1_bF_buf0) );
BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_277__bF_buf4) );
BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_277__bF_buf3) );
BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_277__bF_buf2) );
BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_277__bF_buf1) );
BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_277__bF_buf0) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf3), .Y(_30_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(ULA_ctrl[2]), .C(ULA_ctrl[3]), .Y(_41_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .B(ULA_ctrl_1_bF_buf3), .C(ULA_ctrl[3]), .Y(_42_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_42_), .Y(_52_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_52_), .Y(_63_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .Y(_74_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf3), .B(ULA_ctrl[3]), .C(_30_), .Y(_94_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf2), .B(ULA_ctrl_1_bF_buf3), .C(ULA_ctrl[3]), .Y(_105_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[3]), .Y(_106_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .B(_106__bF_buf4), .Y(_127_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_105_), .C(_127_), .Y(_137_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_137_), .Y(_138_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .Y(_149_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .B(ULA_B_0_bF_buf1), .Y(_169_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf1), .B(_169_), .Y(_180_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(ULA_A[0]), .C(ULA_B_0_bF_buf1), .Y(_181_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .C(_138__bF_buf3), .Y(_201_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf2), .Y(_212_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(ULA_B_1_bF_buf0), .Y(_213_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf3), .B(_213_), .Y(_223_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(_223_), .Y(_234_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf4), .B(_234_), .Y(_244_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf5), .Y(_255_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(_213_), .Y(_266_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_255__bF_buf3), .B(_266_), .Y(_277_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_A[2]), .S(ULA_B_0_bF_buf3), .Y(_287_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(ULA_B_1_bF_buf0), .Y(_298_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_298_), .Y(_308_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(ULA_B_1_bF_buf0), .Y(_319_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(ULA_ctrl_0_bF_buf0), .Y(_330_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_330_), .Y(_340_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_A[0]), .S(ULA_B_0_bF_buf3), .Y(_351_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_287_), .S(_340__bF_buf3), .Y(_362_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_A[4]), .S(ULA_B_0_bF_buf4), .Y(_372_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_A[6]), .S(ULA_B_0_bF_buf4), .Y(_383_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_383_), .S(_340__bF_buf3), .Y(_394_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_362_), .S(_277__bF_buf4), .Y(_404_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_244__bF_buf0), .B(_404_), .Y(_415_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf6), .B(_223_), .Y(_426_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(ULA_ctrl_0_bF_buf3), .Y(_436_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_4_bF_buf3), .B(_436_), .Y(_447_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf3), .B(_266_), .Y(_458_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(ULA_B_1_bF_buf0), .Y(_468_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf2), .B(_468_), .Y(_479_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_298_), .Y(_490_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .B(ULA_A[14]), .S(ULA_B_0_bF_buf5), .Y(_500_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf1), .B(_500_), .Y(_511_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_A[12]), .S(ULA_B_0_bF_buf6), .Y(_522_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf1), .B(_522_), .Y(_532_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_511_), .Y(_543_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_A[10]), .S(ULA_B_0_bF_buf6), .Y(_554_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf3), .B(_554_), .Y(_564_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_A[8]), .S(ULA_B_0_bF_buf4), .Y(_575_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf0), .B(_575_), .Y(_585_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_564_), .Y(_596_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_543_), .S(_458__bF_buf2), .Y(_607_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_244__bF_buf0), .B(_607_), .C(_447__bF_buf1), .Y(_617_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_415_), .Y(_638_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_42_), .Y(_639_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf1), .B(_447__bF_buf0), .Y(_649_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .B(ULA_A[30]), .S(ULA_B_0_bF_buf7), .Y(_650_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf4), .B(_650_), .Y(_651_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[29]), .B(ULA_A[28]), .S(ULA_B_0_bF_buf7), .Y(_652_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf2), .B(_652_), .Y(_653_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_651_), .Y(_654_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_277__bF_buf2), .Y(_655_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[25]), .B(ULA_A[24]), .S(ULA_B_0_bF_buf5), .Y(_656_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf1), .B(_656_), .Y(_657_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[27]), .B(ULA_A[26]), .S(ULA_B_0_bF_buf7), .Y(_658_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf1), .B(_658_), .Y(_659_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_659_), .Y(_660_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_458__bF_buf0), .Y(_661_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_661_), .Y(_662_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_244__bF_buf1), .Y(_663_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf6), .B(_234_), .Y(_664_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[23]), .B(ULA_A[22]), .S(ULA_B_0_bF_buf3), .Y(_665_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf1), .B(_665_), .Y(_666_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[21]), .B(ULA_A[20]), .S(ULA_B_0_bF_buf4), .Y(_667_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf1), .B(_667_), .Y(_668_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_666_), .Y(_669_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_277__bF_buf1), .Y(_670_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[19]), .B(ULA_A[18]), .S(ULA_B_0_bF_buf6), .Y(_671_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf0), .B(_671_), .Y(_672_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[17]), .B(ULA_A[16]), .S(ULA_B_0_bF_buf6), .Y(_673_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf0), .B(_673_), .Y(_674_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_672_), .Y(_675_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_458__bF_buf2), .Y(_676_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_676_), .Y(_677_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_664__bF_buf2), .Y(_678_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf1), .B(_678_), .Y(_679_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_679_), .Y(_680_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_649_), .Y(_681_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_638_), .Y(_682_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(ULA_B_1_bF_buf4), .Y(_683_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf6), .Y(_684_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_684__bF_buf4), .Y(_685_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_685_), .Y(_686_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(ULA_B_2_bF_buf2), .Y(_687_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_684__bF_buf4), .Y(_688_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(ULA_B_1_bF_buf4), .Y(_689_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_688_), .B(_689_), .Y(_690_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_255__bF_buf3), .Y(_691_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_691_), .Y(_692_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_212__bF_buf1), .Y(_693_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(ULA_B_1_bF_buf6), .Y(_694_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_684__bF_buf2), .Y(_695_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_695_), .Y(_696_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(ULA_B_2_bF_buf5), .Y(_697_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(ULA_B_1_bF_buf4), .Y(_698_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_684__bF_buf2), .Y(_699_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_699_), .Y(_700_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_255__bF_buf3), .Y(_701_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_701_), .Y(_702_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(ULA_B_3_bF_buf3), .Y(_703_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_703_), .Y(_704_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_4_bF_buf2), .B(_105_), .Y(_705_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf3), .B(_704_), .Y(_706_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_684__bF_buf1), .Y(_707_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(ULA_B_1_bF_buf5), .Y(_708_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_708_), .Y(_709_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(ULA_B_2_bF_buf6), .Y(_710_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(ULA_B_1_bF_buf2), .Y(_711_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_684__bF_buf0), .Y(_712_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_712_), .Y(_713_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_255__bF_buf5), .Y(_714_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_714_), .Y(_715_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(ULA_B_3_bF_buf3), .Y(_716_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(ULA_B_1_bF_buf4), .Y(_717_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_684__bF_buf2), .Y(_718_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_717_), .B(_718_), .Y(_719_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(ULA_B_2_bF_buf4), .Y(_720_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(ULA_B_1_bF_buf6), .Y(_721_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_684__bF_buf2), .Y(_722_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_722_), .Y(_723_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_255__bF_buf2), .Y(_724_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_724_), .Y(_725_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_212__bF_buf2), .Y(_726_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_726_), .Y(_727_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_4_bF_buf1), .Y(_728_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_105_), .Y(_729_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_727_), .Y(_730_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_426_), .Y(_731_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(ULA_B_4_bF_buf3), .Y(_732_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(ULA_A[0]), .C(_731_), .Y(_733_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_106__bF_buf3), .B(ULA_ctrl[2]), .C(ULA_ctrl_1_bF_buf1), .Y(_734_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(ULA_ctrl[2]), .C(_106__bF_buf3), .Y(_735_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_735_), .Y(_736_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .Y(_737_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .Y(_738_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(_738_), .Y(_739_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .B(ULA_B_0_bF_buf1), .C(ULA_ctrl_1_bF_buf5), .Y(_740_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_739_), .C(_740_), .Y(_741_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_138__bF_buf3), .Y(_742_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_733_), .Y(_743_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_730_), .Y(_744_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_706_), .Y(_745_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_745_), .Y(_746_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_746_), .Y(_747_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_747_), .Y(_0__0_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_B_1_bF_buf0), .Y(_748_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf2), .B(_748_), .Y(_749_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_138__bF_buf4), .B(_749_), .Y(_750_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(ULA_B_1_bF_buf0), .C(ULA_A[31]), .Y(_751_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[30]), .B(ULA_A[29]), .S(ULA_B_0_bF_buf7), .Y(_752_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_490__bF_buf4), .Y(_753_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_751_), .Y(_754_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_277__bF_buf2), .Y(_755_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[28]), .B(ULA_A[27]), .S(ULA_B_0_bF_buf7), .Y(_756_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf4), .B(_756_), .Y(_757_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[26]), .B(ULA_A[25]), .S(ULA_B_0_bF_buf7), .Y(_758_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf2), .B(_758_), .Y(_759_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_757_), .Y(_760_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_458__bF_buf0), .Y(_761_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_761_), .Y(_762_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_244__bF_buf2), .Y(_763_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[22]), .B(ULA_A[21]), .S(ULA_B_0_bF_buf5), .Y(_764_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[24]), .B(ULA_A[23]), .S(ULA_B_0_bF_buf3), .Y(_765_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_765_), .S(_340__bF_buf4), .Y(_766_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[18]), .B(ULA_A[17]), .S(ULA_B_0_bF_buf3), .Y(_767_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[20]), .B(ULA_A[19]), .S(ULA_B_0_bF_buf3), .Y(_768_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_768_), .S(_340__bF_buf4), .Y(_769_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_766_), .S(_458__bF_buf3), .Y(_770_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_664__bF_buf0), .Y(_771_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_771_), .Y(_772_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_447__bF_buf0), .Y(_773_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf3), .Y(_774_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[16]), .B(ULA_A[15]), .S(ULA_B_0_bF_buf4), .Y(_775_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf2), .B(_775_), .Y(_776_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_A[13]), .S(ULA_B_0_bF_buf4), .Y(_777_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf4), .B(_777_), .Y(_778_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_776_), .Y(_779_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_277__bF_buf4), .Y(_780_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_A[11]), .S(ULA_B_0_bF_buf4), .Y(_781_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf3), .B(_781_), .Y(_782_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_A[9]), .S(ULA_B_0_bF_buf4), .Y(_783_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf5), .B(_783_), .Y(_784_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_782_), .Y(_785_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_458__bF_buf1), .Y(_786_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_786_), .Y(_787_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_244__bF_buf3), .Y(_788_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_A[3]), .S(ULA_B_0_bF_buf3), .Y(_789_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_A[1]), .S(ULA_B_0_bF_buf3), .Y(_790_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_789_), .S(_340__bF_buf3), .Y(_791_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_A[5]), .S(ULA_B_0_bF_buf3), .Y(_792_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_A[7]), .S(ULA_B_0_bF_buf4), .Y(_793_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_793_), .S(_340__bF_buf5), .Y(_794_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_791_), .S(_277__bF_buf4), .Y(_795_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_795_), .B(_664__bF_buf4), .Y(_796_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_796_), .Y(_797_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_774_), .Y(_798_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_798_), .Y(_799_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf3), .B(_799_), .Y(_800_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_789_), .S(_684__bF_buf4), .Y(_801_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_792_), .S(ULA_B_1_bF_buf7), .Y(_802_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_801_), .S(ULA_B_2_bF_buf3), .Y(_803_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_803_), .B(_212__bF_buf4), .Y(_804_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(ULA_B_1_bF_buf7), .Y(_805_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_684__bF_buf4), .Y(_806_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_806_), .Y(_807_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(ULA_B_2_bF_buf2), .Y(_808_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(ULA_B_1_bF_buf7), .Y(_809_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_684__bF_buf4), .Y(_810_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_810_), .Y(_811_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_255__bF_buf0), .Y(_812_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_812_), .Y(_813_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(ULA_B_3_bF_buf6), .Y(_814_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_814_), .B(_804_), .Y(_815_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf0), .B(_815_), .Y(_816_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_684__bF_buf0), .Y(_817_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .Y(_818_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(_818_), .Y(_819_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_819_), .B(ULA_B_1_bF_buf0), .Y(_820_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_820_), .Y(_821_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_756_), .B(ULA_B_1_bF_buf2), .Y(_822_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_684__bF_buf0), .Y(_823_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(_823_), .Y(_824_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_824_), .S(ULA_B_2_bF_buf3), .Y(_825_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(ULA_B_1_bF_buf0), .Y(_826_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_684__bF_buf0), .Y(_827_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_827_), .Y(_828_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(ULA_B_1_bF_buf7), .Y(_829_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_684__bF_buf0), .Y(_830_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(_830_), .Y(_831_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_828_), .S(_255__bF_buf0), .Y(_832_) );
MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_832_), .S(ULA_B_3_bF_buf6), .Y(_833_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_833_), .Y(_834_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf4), .B(ULA_A[1]), .C(ULA_B_1_bF_buf2), .Y(_835_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_B_1_bF_buf2), .C(_835_), .Y(_836_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[2]), .B(_836_), .Y(_837_) );
MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .B(ULA_A[1]), .S(ULA_B_0_bF_buf7), .Y(_838_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf5), .B(_838_), .Y(_839_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf0), .B(_839_), .Y(_840_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(ULA_B_3_bF_buf0), .Y(_841_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_4_bF_buf2), .B(_52_), .Y(_842_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf0), .Y(_843_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_106__bF_buf0), .B(_837_), .C(_841_), .D(_843_), .Y(_844_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_844_), .Y(_845_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_816_), .Y(_846_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_846_), .Y(_847_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_847_), .Y(_848_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_848_), .Y(_0__1_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_B_2_bF_buf3), .Y(_849_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf2), .B(_849_), .Y(_850_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(ULA_A[2]), .C(ULA_B_2_bF_buf3), .Y(_851_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_851_), .C(_138__bF_buf4), .Y(_852_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_490__bF_buf4), .Y(_853_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_277__bF_buf2), .B(_853_), .Y(_854_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf2), .B(_658_), .Y(_855_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf4), .B(_652_), .Y(_856_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_856_), .Y(_857_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_857_), .B(_458__bF_buf0), .Y(_858_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_858_), .Y(_859_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_244__bF_buf2), .Y(_860_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf1), .B(_656_), .Y(_861_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf1), .B(_665_), .Y(_862_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_861_), .Y(_863_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_277__bF_buf1), .Y(_864_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf2), .B(_667_), .Y(_865_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf1), .B(_671_), .Y(_866_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_865_), .Y(_867_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_458__bF_buf2), .Y(_868_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_868_), .Y(_869_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_664__bF_buf0), .Y(_870_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_870_), .Y(_871_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_871_), .B(_447__bF_buf3), .Y(_872_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf0), .B(_673_), .Y(_873_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf3), .B(_500_), .Y(_874_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_873_), .Y(_875_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_277__bF_buf3), .Y(_876_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf0), .B(_522_), .Y(_877_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf0), .B(_554_), .Y(_878_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_877_), .Y(_879_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_458__bF_buf1), .Y(_880_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_880_), .Y(_881_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_244__bF_buf3), .Y(_882_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf0), .B(_575_), .Y(_883_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf0), .B(_383_), .Y(_884_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_883_), .Y(_885_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_277__bF_buf3), .Y(_886_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf0), .B(_372_), .Y(_887_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf3), .B(_287_), .Y(_888_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_887_), .Y(_889_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_889_), .B(_458__bF_buf1), .Y(_890_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_890_), .Y(_891_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_664__bF_buf4), .Y(_892_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_882_), .B(_892_), .Y(_893_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_774_), .Y(_894_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_894_), .Y(_895_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf3), .B(_895_), .Y(_896_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(ULA_B_1_bF_buf4), .Y(_897_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_684__bF_buf2), .Y(_898_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_897_), .B(_898_), .Y(_899_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(ULA_B_2_bF_buf5), .Y(_900_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_684__bF_buf4), .Y(_901_) );
AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(ULA_B_1_bF_buf4), .Y(_902_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_902_), .Y(_903_) );
AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_255__bF_buf3), .Y(_904_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_904_), .Y(_905_) );
AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_212__bF_buf1), .Y(_906_) );
AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(ULA_B_1_bF_buf6), .Y(_907_) );
AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_684__bF_buf2), .Y(_908_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_908_), .Y(_909_) );
AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(ULA_B_2_bF_buf5), .Y(_910_) );
AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(ULA_B_1_bF_buf4), .Y(_911_) );
AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_684__bF_buf2), .Y(_912_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_912_), .Y(_913_) );
AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_913_), .B(_255__bF_buf2), .Y(_914_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_914_), .Y(_915_) );
AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_915_), .B(ULA_B_3_bF_buf0), .Y(_916_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(_916_), .Y(_917_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf1), .B(_917_), .Y(_918_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_1_bF_buf5), .B(_650_), .Y(_919_) );
AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(ULA_B_2_bF_buf6), .Y(_920_) );
AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(ULA_B_1_bF_buf2), .Y(_921_) );
AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_684__bF_buf0), .Y(_922_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_921_), .B(_922_), .Y(_923_) );
AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_255__bF_buf5), .Y(_924_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_920_), .B(_924_), .Y(_925_) );
AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(ULA_B_3_bF_buf7), .Y(_926_) );
AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_684__bF_buf2), .Y(_927_) );
AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(ULA_B_1_bF_buf4), .Y(_928_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_928_), .Y(_929_) );
AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(ULA_B_2_bF_buf5), .Y(_930_) );
AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(ULA_B_1_bF_buf6), .Y(_931_) );
AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_684__bF_buf2), .Y(_932_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_932_), .Y(_933_) );
AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_255__bF_buf2), .Y(_934_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_934_), .Y(_935_) );
AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_212__bF_buf2), .Y(_936_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_936_), .Y(_937_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_937_), .Y(_938_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_B_2_bF_buf4), .Y(_939_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf4), .B(ULA_A[2]), .C(ULA_B_2_bF_buf4), .Y(_940_) );
AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_939_), .Y(_941_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf2), .B(_941_), .C(_106__bF_buf0), .Y(_942_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf1), .B(_737_), .Y(_943_) );
AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(ULA_B_1_bF_buf2), .Y(_944_) );
MUX2X1 MUX2X1_49 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[1]), .B(ULA_A[2]), .S(ULA_B_0_bF_buf5), .Y(_945_) );
AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_684__bF_buf1), .Y(_946_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_944_), .Y(_947_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf6), .B(_947_), .Y(_948_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf0), .B(_948_), .Y(_949_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf0), .B(_949_), .Y(_950_) );
AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_942_), .Y(_951_) );
AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_951_), .Y(_952_) );
AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_918_), .Y(_953_) );
AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_953_), .Y(_954_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_954_), .Y(_955_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_955_), .Y(_0__2_) );
AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_B_3_bF_buf6), .Y(_956_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(_956_), .Y(_957_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(_956_), .Y(_958_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_958_), .C(_138__bF_buf4), .Y(_959_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_0_bF_buf7), .B(ULA_B_1_bF_buf2), .Y(_960_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(ULA_B_2_bF_buf4), .C(ULA_A[31]), .Y(_961_) );
AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf4), .B(_752_), .Y(_962_) );
AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf2), .B(_756_), .Y(_963_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_962_), .Y(_964_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_277__bF_buf0), .B(_964_), .Y(_965_) );
AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_965_), .B(_961_), .Y(_966_) );
AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_244__bF_buf1), .Y(_967_) );
AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf1), .B(_758_), .Y(_968_) );
AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf1), .B(_765_), .Y(_969_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_968_), .Y(_970_) );
AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_277__bF_buf1), .Y(_971_) );
AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf2), .B(_764_), .Y(_972_) );
AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf4), .B(_768_), .Y(_973_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_972_), .Y(_974_) );
AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(_458__bF_buf3), .Y(_975_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_975_), .Y(_976_) );
AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_664__bF_buf1), .Y(_977_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_977_), .Y(_978_) );
AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_447__bF_buf2), .Y(_979_) );
MUX2X1 MUX2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_767_), .S(_340__bF_buf4), .Y(_980_) );
MUX2X1 MUX2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_777_), .S(_340__bF_buf5), .Y(_981_) );
MUX2X1 MUX2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(_980_), .S(_458__bF_buf3), .Y(_982_) );
AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_244__bF_buf0), .Y(_983_) );
MUX2X1 MUX2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_792_), .S(_340__bF_buf3), .Y(_984_) );
MUX2X1 MUX2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_783_), .S(_340__bF_buf5), .Y(_985_) );
MUX2X1 MUX2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(_984_), .S(_277__bF_buf1), .Y(_986_) );
AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(_664__bF_buf3), .Y(_987_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_987_), .Y(_988_) );
AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_988_), .B(_774_), .Y(_989_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_979_), .B(_989_), .Y(_990_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf1), .B(_990_), .Y(_991_) );
MUX2X1 MUX2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_775_), .S(ULA_B_1_bF_buf7), .Y(_992_) );
MUX2X1 MUX2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_781_), .S(ULA_B_1_bF_buf7), .Y(_993_) );
MUX2X1 MUX2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_992_), .S(_255__bF_buf3), .Y(_994_) );
AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(ULA_B_3_bF_buf6), .Y(_995_) );
MUX2X1 MUX2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_789_), .S(ULA_B_1_bF_buf7), .Y(_996_) );
MUX2X1 MUX2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_793_), .S(ULA_B_1_bF_buf7), .Y(_997_) );
MUX2X1 MUX2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_996_), .S(ULA_B_2_bF_buf3), .Y(_998_) );
AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_212__bF_buf4), .Y(_999_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf0), .B(_999_), .Y(_1000_) );
OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_995_), .B(_1000_), .Y(_1001_) );
AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(ULA_B_1_bF_buf2), .Y(_1002_) );
AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_756_), .B(_684__bF_buf0), .Y(_1003_) );
OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_1002_), .B(_1003_), .Y(_1004_) );
OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf4), .B(_1004_), .Y(_1005_) );
AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .B(_961_), .Y(_1006_) );
AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(ULA_B_3_bF_buf5), .Y(_1007_) );
AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(ULA_B_1_bF_buf0), .Y(_1008_) );
AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_684__bF_buf0), .Y(_1009_) );
OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_1009_), .Y(_1010_) );
AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(ULA_B_2_bF_buf2), .Y(_1011_) );
AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(ULA_B_1_bF_buf2), .Y(_1012_) );
AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_684__bF_buf0), .Y(_1013_) );
OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_1012_), .B(_1013_), .Y(_1014_) );
AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(_255__bF_buf0), .Y(_1015_) );
OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1015_), .Y(_1016_) );
AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_212__bF_buf4), .Y(_1017_) );
OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .B(_1007_), .Y(_1018_) );
OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1018_), .Y(_1019_) );
AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(ULA_B_1_bF_buf5), .Y(_1020_) );
MUX2X1 MUX2X1_62 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[2]), .B(ULA_A[3]), .S(ULA_B_0_bF_buf7), .Y(_1021_) );
AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .B(_684__bF_buf1), .Y(_1022_) );
OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(_1022_), .Y(_1023_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(ULA_B_2_bF_buf6), .C(ULA_B_3_bF_buf0), .Y(_1024_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_B_3_bF_buf5), .Y(_1025_) );
AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(ULA_ctrl_1_bF_buf4), .Y(_1026_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1025_), .C(ULA_ctrl[2]), .Y(_1027_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_106__bF_buf0), .B(_1027_), .C(_843_), .D(_1024_), .Y(_1028_) );
AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1019_), .Y(_1029_) );
AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(_1001_), .Y(_1030_) );
AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_1030_), .Y(_1031_) );
OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_1031_), .Y(_1032_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .Y(_0__3_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_B_4_bF_buf3), .Y(_1033_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf0), .B(_1033_), .Y(_1034_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(ULA_A[4]), .C(ULA_B_4_bF_buf3), .Y(_1035_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1035_), .C(_138__bF_buf3), .Y(_1036_) );
MUX2X1 MUX2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_650_), .S(_340__bF_buf2), .Y(_1037_) );
AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_458__bF_buf0), .Y(_1038_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_664__bF_buf2), .Y(_1039_) );
AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_277__bF_buf0), .Y(_1040_) );
AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_458__bF_buf3), .Y(_1041_) );
OR2X2 OR2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .B(_1041_), .Y(_1042_) );
AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_664__bF_buf0), .Y(_1043_) );
OR2X2 OR2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .B(_1039_), .Y(_1044_) );
AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_447__bF_buf0), .Y(_1045_) );
AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_277__bF_buf1), .Y(_1046_) );
AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_458__bF_buf2), .Y(_1047_) );
OR2X2 OR2X2_127 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1047_), .Y(_1048_) );
AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_244__bF_buf3), .Y(_1049_) );
MUX2X1 MUX2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_554_), .S(_340__bF_buf0), .Y(_1050_) );
MUX2X1 MUX2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_394_), .S(_277__bF_buf4), .Y(_1051_) );
AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_664__bF_buf4), .Y(_1052_) );
OR2X2 OR2X2_128 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1052_), .Y(_1053_) );
AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_774_), .Y(_1054_) );
OR2X2 OR2X2_129 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1054_), .Y(_1055_) );
OR2X2 OR2X2_130 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf3), .B(_1055_), .Y(_1056_) );
OR2X2 OR2X2_131 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf6), .B(_709_), .Y(_1057_) );
AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(ULA_B_3_bF_buf4), .Y(_1058_) );
AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(ULA_B_2_bF_buf4), .Y(_1059_) );
AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_255__bF_buf5), .Y(_1060_) );
OR2X2 OR2X2_132 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1060_), .Y(_1061_) );
AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_212__bF_buf2), .Y(_1062_) );
OR2X2 OR2X2_133 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1062_), .Y(_1063_) );
OR2X2 OR2X2_134 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1063_), .Y(_1064_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf0), .Y(_1065_) );
AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(ULA_B_2_bF_buf5), .Y(_1066_) );
AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_255__bF_buf2), .Y(_1067_) );
OR2X2 OR2X2_135 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1067_), .Y(_1068_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf0), .B(_1068_), .Y(_1069_) );
MUX2X1 MUX2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_686_), .S(ULA_B_2_bF_buf5), .Y(_1070_) );
OR2X2 OR2X2_136 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf5), .B(_1070_), .Y(_1071_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1065_), .C(_1071_), .Y(_1072_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[0]), .B(_960_), .C(_255__bF_buf5), .Y(_1073_) );
MUX2X1 MUX2X1_67 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[3]), .B(ULA_A[4]), .S(ULA_B_0_bF_buf5), .Y(_1074_) );
AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_684__bF_buf1), .Y(_1075_) );
AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(ULA_B_1_bF_buf5), .Y(_1076_) );
OR2X2 OR2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1076_), .Y(_1077_) );
AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_255__bF_buf5), .Y(_1078_) );
OR2X2 OR2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1078_), .Y(_1079_) );
OR2X2 OR2X2_139 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf4), .B(_1079_), .Y(_1080_) );
OR2X2 OR2X2_140 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf3), .B(_1080_), .Y(_1081_) );
OR2X2 OR2X2_141 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_B_4_bF_buf0), .Y(_1082_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf2), .B(ULA_A[4]), .C(ULA_B_4_bF_buf0), .Y(_1083_) );
AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1082_), .Y(_1084_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf1), .B(_1084_), .C(_106__bF_buf2), .Y(_1085_) );
AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_1085_), .Y(_1086_) );
AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1086_), .Y(_1087_) );
AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(_1064_), .Y(_1088_) );
AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_1056_), .B(_1088_), .Y(_1089_) );
OR2X2 OR2X2_142 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .B(_1089_), .Y(_1090_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .Y(_0__4_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_B[5]), .Y(_1091_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf0), .B(_1091_), .Y(_1092_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .B(ULA_A[5]), .C(ULA_B[5]), .Y(_1093_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_1093_), .C(_138__bF_buf0), .Y(_1094_) );
OR2X2 OR2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_277__bF_buf2), .B(_754_), .Y(_1095_) );
AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_244__bF_buf1), .Y(_1096_) );
AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_277__bF_buf0), .Y(_1097_) );
AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf2), .B(_765_), .Y(_1098_) );
AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf2), .B(_764_), .Y(_1099_) );
OR2X2 OR2X2_144 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1098_), .Y(_1100_) );
AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .B(_458__bF_buf0), .Y(_1101_) );
OR2X2 OR2X2_145 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .B(_1101_), .Y(_1102_) );
AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_664__bF_buf1), .Y(_1103_) );
OR2X2 OR2X2_146 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1103_), .Y(_1104_) );
AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_447__bF_buf2), .Y(_1105_) );
MUX2X1 MUX2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_781_), .S(_340__bF_buf5), .Y(_1106_) );
MUX2X1 MUX2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1106_), .B(_794_), .S(_277__bF_buf4), .Y(_1107_) );
AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .B(_664__bF_buf3), .Y(_1108_) );
AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf3), .B(_768_), .Y(_1109_) );
AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf5), .B(_767_), .Y(_1110_) );
OR2X2 OR2X2_147 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .B(_1109_), .Y(_1111_) );
AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(_1111_), .B(_277__bF_buf4), .Y(_1112_) );
AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_458__bF_buf2), .Y(_1113_) );
OR2X2 OR2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1113_), .Y(_1114_) );
AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_244__bF_buf0), .Y(_1115_) );
OR2X2 OR2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1108_), .Y(_1116_) );
AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .B(_774_), .Y(_1117_) );
OR2X2 OR2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_1117_), .Y(_1118_) );
OR2X2 OR2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf0), .B(_1118_), .Y(_1119_) );
OR2X2 OR2X2_152 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf3), .B(_802_), .Y(_1120_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf2), .B(_811_), .C(ULA_B_3_bF_buf6), .Y(_1121_) );
AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1120_), .Y(_1122_) );
AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(ULA_B_2_bF_buf2), .Y(_1123_) );
AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_255__bF_buf0), .Y(_1124_) );
OR2X2 OR2X2_153 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1124_), .Y(_1125_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .B(_212__bF_buf1), .Y(_1126_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1126_), .C(_1065_), .Y(_1127_) );
OR2X2 OR2X2_154 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf4), .B(_821_), .Y(_1128_) );
AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(ULA_B_3_bF_buf3), .Y(_1129_) );
AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(ULA_B_2_bF_buf2), .Y(_1130_) );
AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_255__bF_buf0), .Y(_1131_) );
OR2X2 OR2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1131_), .Y(_1132_) );
AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_212__bF_buf1), .Y(_1133_) );
OR2X2 OR2X2_156 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_1133_), .Y(_1134_) );
OR2X2 OR2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1134_), .Y(_1135_) );
AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(ULA_B_2_bF_buf0), .Y(_1136_) );
AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .B(ULA_B_1_bF_buf5), .Y(_1137_) );
MUX2X1 MUX2X1_70 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[4]), .B(ULA_A[5]), .S(ULA_B_0_bF_buf5), .Y(_1138_) );
AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_684__bF_buf1), .Y(_1139_) );
OR2X2 OR2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1139_), .Y(_1140_) );
AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_255__bF_buf6), .Y(_1141_) );
OR2X2 OR2X2_159 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1141_), .Y(_1142_) );
OR2X2 OR2X2_160 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf1), .B(_1142_), .Y(_1143_) );
OR2X2 OR2X2_161 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf3), .B(_1143_), .Y(_1144_) );
OR2X2 OR2X2_162 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_B[5]), .Y(_1145_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf3), .B(ULA_A[5]), .C(ULA_B[5]), .Y(_1146_) );
AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .B(_1145_), .Y(_1147_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf2), .B(_1147_), .C(_106__bF_buf1), .Y(_1148_) );
AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1148_), .Y(_1149_) );
AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1149_), .Y(_1150_) );
AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1150_), .Y(_1151_) );
AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_1119_), .B(_1151_), .Y(_1152_) );
OR2X2 OR2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_1094_), .B(_1152_), .Y(_1153_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .Y(_0__5_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_B[6]), .Y(_1154_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf1), .B(_1154_), .Y(_1155_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(ULA_A[6]), .C(ULA_B[6]), .Y(_1156_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1156_), .C(_138__bF_buf3), .Y(_1157_) );
AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_857_), .B(_277__bF_buf0), .Y(_1158_) );
AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_458__bF_buf3), .Y(_1159_) );
OR2X2 OR2X2_164 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .B(_1159_), .Y(_1160_) );
AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_664__bF_buf1), .Y(_1161_) );
OR2X2 OR2X2_165 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_277__bF_buf2), .Y(_1162_) );
AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_244__bF_buf1), .Y(_1163_) );
OR2X2 OR2X2_166 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1161_), .Y(_1164_) );
AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_1164_), .B(_447__bF_buf0), .Y(_1165_) );
OR2X2 OR2X2_167 ( .gnd(gnd), .vdd(vdd), .A(_458__bF_buf1), .B(_879_), .Y(_1166_) );
OR2X2 OR2X2_168 ( .gnd(gnd), .vdd(vdd), .A(_277__bF_buf3), .B(_885_), .Y(_1167_) );
AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_664__bF_buf4), .Y(_1168_) );
AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1166_), .Y(_1169_) );
AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_277__bF_buf3), .Y(_1170_) );
AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_458__bF_buf1), .Y(_1171_) );
OR2X2 OR2X2_169 ( .gnd(gnd), .vdd(vdd), .A(_1170_), .B(_1171_), .Y(_1172_) );
AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(_244__bF_buf3), .Y(_1173_) );
OR2X2 OR2X2_170 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1173_), .Y(_1174_) );
AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_774_), .Y(_1175_) );
OR2X2 OR2X2_171 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1175_), .Y(_1176_) );
OR2X2 OR2X2_172 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf3), .B(_1176_), .Y(_1177_) );
OR2X2 OR2X2_173 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf6), .B(_919_), .Y(_1178_) );
AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(ULA_B_3_bF_buf7), .Y(_1179_) );
AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(ULA_B_2_bF_buf6), .Y(_1180_) );
AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_255__bF_buf2), .Y(_1181_) );
OR2X2 OR2X2_174 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(_1181_), .Y(_1182_) );
AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_212__bF_buf2), .Y(_1183_) );
OR2X2 OR2X2_175 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_1183_), .Y(_1184_) );
OR2X2 OR2X2_176 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1184_), .Y(_1185_) );
AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(ULA_B_2_bF_buf5), .Y(_1186_) );
AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_255__bF_buf2), .Y(_1187_) );
OR2X2 OR2X2_177 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1187_), .Y(_1188_) );
AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(ULA_B_3_bF_buf0), .Y(_1189_) );
AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_255__bF_buf3), .Y(_1190_) );
AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_913_), .B(ULA_B_2_bF_buf5), .Y(_1191_) );
OR2X2 OR2X2_178 ( .gnd(gnd), .vdd(vdd), .A(_1190_), .B(_1191_), .Y(_1192_) );
AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_212__bF_buf1), .Y(_1193_) );
OR2X2 OR2X2_179 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1193_), .Y(_1194_) );
OR2X2 OR2X2_180 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf1), .B(_1194_), .Y(_1195_) );
MUX2X1 MUX2X1_71 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[5]), .B(ULA_A[6]), .S(ULA_B_0_bF_buf5), .Y(_1196_) );
AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_684__bF_buf1), .Y(_1197_) );
AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(ULA_B_1_bF_buf5), .Y(_1198_) );
OR2X2 OR2X2_181 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_1198_), .Y(_1199_) );
AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(_255__bF_buf5), .Y(_1200_) );
AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(ULA_B_2_bF_buf6), .Y(_1201_) );
OR2X2 OR2X2_182 ( .gnd(gnd), .vdd(vdd), .A(_1200_), .B(_1201_), .Y(_1202_) );
OR2X2 OR2X2_183 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf4), .B(_1202_), .Y(_1203_) );
OR2X2 OR2X2_184 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf0), .B(_1203_), .Y(_1204_) );
OR2X2 OR2X2_185 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_B[6]), .Y(_1205_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf5), .B(ULA_A[6]), .C(ULA_B[6]), .Y(_1206_) );
AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_1205_), .Y(_1207_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf0), .B(_1207_), .C(_106__bF_buf4), .Y(_1208_) );
AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1208_), .Y(_1209_) );
AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1209_), .Y(_1210_) );
AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(_1185_), .Y(_1211_) );
AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1211_), .Y(_1212_) );
OR2X2 OR2X2_186 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1212_), .Y(_1213_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .Y(_0__6_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_B[7]), .Y(_1214_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf3), .B(_1214_), .Y(_1215_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(ULA_A[7]), .C(ULA_B[7]), .Y(_1216_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_1216_), .C(_138__bF_buf1), .Y(_1217_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_1218_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .B(_1218_), .C(_664__bF_buf1), .Y(_1219_) );
AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_964_), .B(_277__bF_buf0), .Y(_1220_) );
AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_458__bF_buf0), .Y(_1221_) );
OR2X2 OR2X2_187 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_1221_), .Y(_1222_) );
AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_664__bF_buf1), .Y(_1223_) );
OR2X2 OR2X2_188 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1219_), .Y(_1224_) );
AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_447__bF_buf2), .Y(_1225_) );
AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(_277__bF_buf1), .Y(_1226_) );
AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf2), .B(_767_), .Y(_1227_) );
AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf4), .B(_775_), .Y(_1228_) );
OR2X2 OR2X2_189 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1227_), .Y(_1229_) );
AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .B(_458__bF_buf3), .Y(_1230_) );
OR2X2 OR2X2_190 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1230_), .Y(_1231_) );
AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_244__bF_buf3), .Y(_1232_) );
AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf3), .B(_777_), .Y(_1233_) );
AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf0), .B(_781_), .Y(_1234_) );
OR2X2 OR2X2_191 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1233_), .Y(_1235_) );
OR2X2 OR2X2_192 ( .gnd(gnd), .vdd(vdd), .A(_458__bF_buf1), .B(_1235_), .Y(_1236_) );
AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(_490__bF_buf3), .B(_783_), .Y(_1237_) );
AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_340__bF_buf5), .B(_793_), .Y(_1238_) );
OR2X2 OR2X2_193 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1237_), .Y(_1239_) );
OR2X2 OR2X2_194 ( .gnd(gnd), .vdd(vdd), .A(_277__bF_buf3), .B(_1239_), .Y(_1240_) );
AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_664__bF_buf4), .Y(_1241_) );
AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1236_), .Y(_1242_) );
OR2X2 OR2X2_195 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .B(_1232_), .Y(_1243_) );
AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_1243_), .B(_774_), .Y(_1244_) );
OR2X2 OR2X2_196 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1225_), .Y(_1245_) );
OR2X2 OR2X2_197 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf0), .B(_1245_), .Y(_1246_) );
AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(ULA_B_2_bF_buf4), .Y(_1247_) );
AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_255__bF_buf0), .Y(_1248_) );
OR2X2 OR2X2_198 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_1248_), .Y(_1249_) );
OR2X2 OR2X2_199 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf5), .B(_1249_), .Y(_1250_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1218_), .B(ULA_B_3_bF_buf5), .C(ULA_A[31]), .Y(_1251_) );
AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1251_), .Y(_1252_) );
OR2X2 OR2X2_200 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1252_), .Y(_1253_) );
AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_1014_), .B(ULA_B_2_bF_buf2), .Y(_1254_) );
AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(ULA_B_1_bF_buf7), .Y(_1255_) );
AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_684__bF_buf4), .Y(_1256_) );
OR2X2 OR2X2_201 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(_1256_), .Y(_1257_) );
AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_1257_), .B(_255__bF_buf3), .Y(_1258_) );
OR2X2 OR2X2_202 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1258_), .Y(_1259_) );
AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(_1259_), .B(ULA_B_3_bF_buf6), .Y(_1260_) );
AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(ULA_B_1_bF_buf4), .Y(_1261_) );
AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_684__bF_buf4), .Y(_1262_) );
OR2X2 OR2X2_203 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1262_), .Y(_1263_) );
AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_255__bF_buf3), .Y(_1264_) );
AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(ULA_B_1_bF_buf7), .Y(_1265_) );
AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_684__bF_buf4), .Y(_1266_) );
OR2X2 OR2X2_204 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1266_), .Y(_1267_) );
AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(ULA_B_2_bF_buf3), .Y(_1268_) );
OR2X2 OR2X2_205 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1268_), .Y(_1269_) );
AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(_1269_), .B(_212__bF_buf4), .Y(_1270_) );
OR2X2 OR2X2_206 ( .gnd(gnd), .vdd(vdd), .A(_1260_), .B(_1270_), .Y(_1271_) );
OR2X2 OR2X2_207 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf3), .B(_1271_), .Y(_1272_) );
AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(ULA_B_2_bF_buf0), .Y(_1273_) );
AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(ULA_B_1_bF_buf6), .Y(_1274_) );
MUX2X1 MUX2X1_72 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[6]), .B(ULA_A[7]), .S(ULA_B_0_bF_buf6), .Y(_1275_) );
AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_684__bF_buf6), .Y(_1276_) );
OR2X2 OR2X2_208 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1276_), .Y(_1277_) );
AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_1277_), .B(_255__bF_buf6), .Y(_1278_) );
OR2X2 OR2X2_209 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_1278_), .Y(_1279_) );
OR2X2 OR2X2_210 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf1), .B(_1279_), .Y(_1280_) );
OR2X2 OR2X2_211 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf3), .B(_1280_), .Y(_1281_) );
OR2X2 OR2X2_212 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_B[7]), .Y(_1282_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf0), .B(ULA_A[7]), .C(ULA_B[7]), .Y(_1283_) );
AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1282_), .Y(_1284_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf4), .B(_1284_), .C(_106__bF_buf1), .Y(_1285_) );
AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(_1281_), .B(_1285_), .Y(_1286_) );
AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1286_), .Y(_1287_) );
AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .B(_1253_), .Y(_1288_) );
AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1288_), .Y(_1289_) );
OR2X2 OR2X2_213 ( .gnd(gnd), .vdd(vdd), .A(_1217_), .B(_1289_), .Y(_1290_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .Y(_0__7_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf0), .B(_664__bF_buf2), .Y(_1291_) );
OR2X2 OR2X2_214 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_1291_), .Y(_1292_) );
AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_244__bF_buf2), .Y(_1293_) );
AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_277__bF_buf3), .Y(_1294_) );
AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_458__bF_buf2), .Y(_1295_) );
OR2X2 OR2X2_215 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1295_), .Y(_1296_) );
AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_664__bF_buf3), .Y(_1297_) );
OR2X2 OR2X2_216 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf1), .B(_1297_), .Y(_1298_) );
OR2X2 OR2X2_217 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1298_), .Y(_1299_) );
AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(_1299_), .B(_1292_), .Y(_1300_) );
OR2X2 OR2X2_218 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf0), .B(_1300_), .Y(_1301_) );
AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(ULA_B_3_bF_buf3), .Y(_1302_) );
AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_212__bF_buf2), .Y(_1303_) );
OR2X2 OR2X2_219 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf4), .B(_1303_), .Y(_1304_) );
OR2X2 OR2X2_220 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1304_), .Y(_1305_) );
MUX2X1 MUX2X1_73 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[7]), .B(ULA_A[8]), .S(ULA_B_0_bF_buf5), .Y(_1306_) );
AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_684__bF_buf1), .Y(_1307_) );
AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(ULA_B_1_bF_buf6), .Y(_1308_) );
OR2X2 OR2X2_221 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1308_), .Y(_1309_) );
AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_255__bF_buf5), .Y(_1310_) );
AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(ULA_B_2_bF_buf0), .Y(_1311_) );
OR2X2 OR2X2_222 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .B(_1311_), .Y(_1312_) );
OR2X2 OR2X2_223 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf7), .B(_1312_), .Y(_1313_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1218_), .B(ULA_A[0]), .C(ULA_B_3_bF_buf3), .Y(_1314_) );
AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .B(_1314_), .Y(_1315_) );
OR2X2 OR2X2_224 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf0), .B(_1315_), .Y(_1316_) );
OR2X2 OR2X2_225 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf3), .B(_715_), .Y(_1317_) );
OR2X2 OR2X2_226 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1317_), .Y(_1318_) );
OR2X2 OR2X2_227 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_B[8]), .Y(_1319_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf0), .B(ULA_A[8]), .C(ULA_B[8]), .Y(_1320_) );
AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1319_), .Y(_1321_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf4), .B(_1321_), .C(_106__bF_buf1), .Y(_1322_) );
AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1322_), .Y(_1323_) );
AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1323_), .Y(_1324_) );
AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(_1305_), .Y(_1325_) );
AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_1301_), .B(_1325_), .Y(_1326_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_B[8]), .Y(_1327_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf3), .B(_1327_), .Y(_1328_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_A[8]), .C(ULA_B[8]), .Y(_1329_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(_1329_), .C(_138__bF_buf1), .Y(_1330_) );
OR2X2 OR2X2_228 ( .gnd(gnd), .vdd(vdd), .A(_1330_), .B(_1326_), .Y(_1331_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .Y(_0__8_) );
OR2X2 OR2X2_229 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_1291_), .Y(_1332_) );
AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_244__bF_buf2), .Y(_1333_) );
AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_664__bF_buf3), .Y(_1334_) );
OR2X2 OR2X2_230 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf1), .B(_1334_), .Y(_1335_) );
OR2X2 OR2X2_231 ( .gnd(gnd), .vdd(vdd), .A(_1335_), .B(_1333_), .Y(_1336_) );
AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1332_), .Y(_1337_) );
OR2X2 OR2X2_232 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf1), .B(_1337_), .Y(_1338_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf2), .B(_828_), .Y(_1339_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_255__bF_buf0), .B(_831_), .Y(_1340_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1339_), .B(_1340_), .C(_212__bF_buf4), .Y(_1341_) );
AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_212__bF_buf4), .Y(_1342_) );
OR2X2 OR2X2_233 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf0), .B(_1342_), .Y(_1343_) );
OR2X2 OR2X2_234 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1341_), .Y(_1344_) );
AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(ULA_B_3_bF_buf7), .Y(_1345_) );
AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(ULA_B_2_bF_buf0), .Y(_1346_) );
AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(ULA_B_1_bF_buf1), .Y(_1347_) );
MUX2X1 MUX2X1_74 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[8]), .B(ULA_A[9]), .S(ULA_B_0_bF_buf6), .Y(_1348_) );
AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_684__bF_buf3), .Y(_1349_) );
OR2X2 OR2X2_235 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_1349_), .Y(_1350_) );
AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_255__bF_buf6), .Y(_1351_) );
OR2X2 OR2X2_236 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1351_), .Y(_1352_) );
AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_212__bF_buf0), .Y(_1353_) );
OR2X2 OR2X2_237 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1353_), .Y(_1354_) );
OR2X2 OR2X2_238 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf0), .B(_1354_), .Y(_1355_) );
AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(ULA_B_2_bF_buf4), .Y(_1356_) );
AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_255__bF_buf0), .Y(_1357_) );
OR2X2 OR2X2_239 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1356_), .Y(_1358_) );
OR2X2 OR2X2_240 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf5), .B(_1358_), .Y(_1359_) );
OR2X2 OR2X2_241 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1359_), .Y(_1360_) );
OR2X2 OR2X2_242 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_B[9]), .Y(_1361_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf4), .B(ULA_A[9]), .C(ULA_B[9]), .Y(_1362_) );
AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1361_), .Y(_1363_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf2), .B(_1363_), .C(_106__bF_buf0), .Y(_1364_) );
AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1364_), .Y(_1365_) );
AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_1365_), .B(_1355_), .Y(_1366_) );
AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1344_), .Y(_1367_) );
AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1367_), .Y(_1368_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_B[9]), .Y(_1369_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf2), .B(_1369_), .Y(_1370_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf0), .B(ULA_A[9]), .C(ULA_B[9]), .Y(_1371_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1371_), .C(_138__bF_buf4), .Y(_1372_) );
OR2X2 OR2X2_243 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1368_), .Y(_1373_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .Y(_0__9_) );
OR2X2 OR2X2_244 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_1291_), .Y(_1374_) );
AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_244__bF_buf2), .Y(_1375_) );
AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_664__bF_buf0), .Y(_1376_) );
OR2X2 OR2X2_245 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf3), .B(_1376_), .Y(_1377_) );
OR2X2 OR2X2_246 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .B(_1377_), .Y(_1378_) );
AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .B(_1374_), .Y(_1379_) );
OR2X2 OR2X2_247 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf0), .B(_1379_), .Y(_1380_) );
AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(ULA_B_3_bF_buf0), .Y(_1381_) );
AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_915_), .B(_212__bF_buf2), .Y(_1382_) );
OR2X2 OR2X2_248 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf1), .B(_1382_), .Y(_1383_) );
OR2X2 OR2X2_249 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .B(_1383_), .Y(_1384_) );
OR2X2 OR2X2_250 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf2), .B(_948_), .Y(_1385_) );
MUX2X1 MUX2X1_75 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[9]), .B(ULA_A[10]), .S(ULA_B_0_bF_buf6), .Y(_1386_) );
AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_684__bF_buf1), .Y(_1387_) );
AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(ULA_B_1_bF_buf6), .Y(_1388_) );
OR2X2 OR2X2_251 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .B(_1388_), .Y(_1389_) );
AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_255__bF_buf5), .Y(_1390_) );
AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(ULA_B_2_bF_buf6), .Y(_1391_) );
OR2X2 OR2X2_252 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1391_), .Y(_1392_) );
OR2X2 OR2X2_253 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf7), .B(_1392_), .Y(_1393_) );
AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1385_), .Y(_1394_) );
OR2X2 OR2X2_254 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf1), .B(_1394_), .Y(_1395_) );
OR2X2 OR2X2_255 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf4), .B(_925_), .Y(_1396_) );
OR2X2 OR2X2_256 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1396_), .Y(_1397_) );
OR2X2 OR2X2_257 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_B[10]), .Y(_1398_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf0), .B(ULA_A[10]), .C(ULA_B[10]), .Y(_1399_) );
AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1398_), .Y(_1400_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf4), .B(_1400_), .C(_106__bF_buf2), .Y(_1401_) );
AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1401_), .Y(_1402_) );
AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_1402_), .Y(_1403_) );
AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_1384_), .Y(_1404_) );
AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_1380_), .B(_1404_), .Y(_1405_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_B[10]), .Y(_1406_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf3), .B(_1406_), .Y(_1407_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_A[10]), .C(ULA_B[10]), .Y(_1408_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1408_), .C(_138__bF_buf2), .Y(_1409_) );
OR2X2 OR2X2_258 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_1405_), .Y(_1410_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .Y(_0__10_) );
OR2X2 OR2X2_259 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_1291_), .Y(_1411_) );
AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_244__bF_buf0), .Y(_1412_) );
AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_664__bF_buf3), .Y(_1413_) );
OR2X2 OR2X2_260 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1413_), .Y(_1414_) );
OR2X2 OR2X2_261 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf2), .B(_1414_), .Y(_1415_) );
AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_1415_), .B(_1411_), .Y(_1416_) );
OR2X2 OR2X2_262 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf2), .B(_1416_), .Y(_1417_) );
OR2X2 OR2X2_263 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf0), .B(_1023_), .Y(_1418_) );
AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(ULA_B_3_bF_buf2), .Y(_1419_) );
AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_1277_), .B(ULA_B_2_bF_buf1), .Y(_1420_) );
AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(ULA_B_1_bF_buf1), .Y(_1421_) );
MUX2X1 MUX2X1_76 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[10]), .B(ULA_A[11]), .S(ULA_B_0_bF_buf6), .Y(_1422_) );
AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_684__bF_buf3), .Y(_1423_) );
OR2X2 OR2X2_264 ( .gnd(gnd), .vdd(vdd), .A(_1421_), .B(_1423_), .Y(_1424_) );
AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(_255__bF_buf4), .Y(_1425_) );
OR2X2 OR2X2_265 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1425_), .Y(_1426_) );
AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_212__bF_buf3), .Y(_1427_) );
OR2X2 OR2X2_266 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_1427_), .Y(_1428_) );
OR2X2 OR2X2_267 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf3), .B(_1428_), .Y(_1429_) );
AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(ULA_B_3_bF_buf6), .Y(_1430_) );
AND2X2 AND2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_212__bF_buf4), .Y(_1431_) );
OR2X2 OR2X2_268 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(_1431_), .Y(_1432_) );
OR2X2 OR2X2_269 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf3), .B(_1432_), .Y(_1433_) );
OR2X2 OR2X2_270 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf5), .B(_1006_), .Y(_1434_) );
OR2X2 OR2X2_271 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1434_), .Y(_1435_) );
OR2X2 OR2X2_272 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_B[11]), .Y(_1436_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf0), .B(ULA_A[11]), .C(ULA_B[11]), .Y(_1437_) );
AND2X2 AND2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_1437_), .B(_1436_), .Y(_1438_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf4), .B(_1438_), .C(_106__bF_buf1), .Y(_1439_) );
AND2X2 AND2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_1439_), .Y(_1440_) );
AND2X2 AND2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1440_), .Y(_1441_) );
AND2X2 AND2X2_378 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1429_), .Y(_1442_) );
AND2X2 AND2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1442_), .Y(_1443_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_B[11]), .Y(_1444_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf4), .B(_1444_), .Y(_1445_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_A[11]), .C(ULA_B[11]), .Y(_1446_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1445_), .B(_1446_), .C(_138__bF_buf2), .Y(_1447_) );
OR2X2 OR2X2_273 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1443_), .Y(_1448_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .Y(_0__11_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_B[12]), .Y(_1449_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf0), .B(_1449_), .Y(_1450_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .B(ULA_A[12]), .C(ULA_B[12]), .Y(_1451_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1451_), .C(_138__bF_buf0), .Y(_1452_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1038_), .B(_447__bF_buf3), .C(_664__bF_buf2), .Y(_1453_) );
AND2X2 AND2X2_380 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_244__bF_buf3), .Y(_1454_) );
AND2X2 AND2X2_381 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_664__bF_buf0), .Y(_1455_) );
OR2X2 OR2X2_274 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf3), .B(_1455_), .Y(_1456_) );
OR2X2 OR2X2_275 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_1456_), .Y(_1457_) );
AND2X2 AND2X2_382 ( .gnd(gnd), .vdd(vdd), .A(_1457_), .B(_1453_), .Y(_1458_) );
OR2X2 OR2X2_276 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf3), .B(_1458_), .Y(_1459_) );
MUX2X1 MUX2X1_77 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[11]), .B(ULA_A[12]), .S(ULA_B_0_bF_buf5), .Y(_1460_) );
AND2X2 AND2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_684__bF_buf6), .Y(_1461_) );
AND2X2 AND2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(ULA_B_1_bF_buf6), .Y(_1462_) );
OR2X2 OR2X2_277 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_1462_), .Y(_1463_) );
AND2X2 AND2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_255__bF_buf2), .Y(_1464_) );
AND2X2 AND2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(ULA_B_2_bF_buf0), .Y(_1465_) );
OR2X2 OR2X2_278 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1465_), .Y(_1466_) );
AND2X2 AND2X2_387 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_212__bF_buf0), .Y(_1467_) );
AND2X2 AND2X2_388 ( .gnd(gnd), .vdd(vdd), .A(_1079_), .B(ULA_B_3_bF_buf4), .Y(_1468_) );
OR2X2 OR2X2_279 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1467_), .Y(_1469_) );
OR2X2 OR2X2_280 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf1), .B(_1469_), .Y(_1470_) );
AND2X2 AND2X2_389 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_212__bF_buf1), .Y(_1471_) );
AND2X2 AND2X2_390 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(ULA_B_3_bF_buf3), .Y(_1472_) );
OR2X2 OR2X2_281 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1472_), .Y(_1473_) );
OR2X2 OR2X2_282 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf1), .B(_1473_), .Y(_1474_) );
OR2X2 OR2X2_283 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf4), .B(_1057_), .Y(_1475_) );
OR2X2 OR2X2_284 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_1475_), .Y(_1_) );
OR2X2 OR2X2_285 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_B[12]), .Y(_2_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf3), .B(ULA_A[12]), .C(ULA_B[12]), .Y(_3_) );
AND2X2 AND2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_2_), .Y(_4_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf4), .B(_4_), .C(_106__bF_buf1), .Y(_5_) );
AND2X2 AND2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_5_), .Y(_6_) );
AND2X2 AND2X2_393 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_6_), .Y(_7_) );
AND2X2 AND2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_1470_), .Y(_8_) );
AND2X2 AND2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_8_), .Y(_9_) );
OR2X2 OR2X2_286 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_9_), .Y(_10_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_0__12_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_B[13]), .Y(_11_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf4), .B(_11_), .Y(_12_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .B(ULA_A[13]), .C(ULA_B[13]), .Y(_13_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .C(_138__bF_buf0), .Y(_14_) );
OR2X2 OR2X2_287 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1291_), .Y(_15_) );
AND2X2 AND2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_244__bF_buf1), .Y(_16_) );
AND2X2 AND2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_664__bF_buf2), .Y(_17_) );
OR2X2 OR2X2_288 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf1), .B(_17_), .Y(_18_) );
OR2X2 OR2X2_289 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_18_), .Y(_19_) );
AND2X2 AND2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_15_), .Y(_20_) );
OR2X2 OR2X2_290 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf2), .B(_20_), .Y(_21_) );
OR2X2 OR2X2_291 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf1), .B(_1132_), .Y(_22_) );
OR2X2 OR2X2_292 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf5), .B(_1125_), .Y(_23_) );
AND2X2 AND2X2_399 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_23_), .Y(_24_) );
OR2X2 OR2X2_293 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf3), .B(_24_), .Y(_25_) );
AND2X2 AND2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(ULA_B_3_bF_buf1), .Y(_26_) );
AND2X2 AND2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(ULA_B_2_bF_buf1), .Y(_27_) );
AND2X2 AND2X2_402 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(ULA_B_1_bF_buf1), .Y(_28_) );
MUX2X1 MUX2X1_78 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[12]), .B(ULA_A[13]), .S(ULA_B_0_bF_buf0), .Y(_29_) );
AND2X2 AND2X2_403 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_684__bF_buf3), .Y(_31_) );
OR2X2 OR2X2_294 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_31_), .Y(_32_) );
AND2X2 AND2X2_404 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_255__bF_buf4), .Y(_33_) );
OR2X2 OR2X2_295 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_33_), .Y(_34_) );
AND2X2 AND2X2_405 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_212__bF_buf5), .Y(_35_) );
OR2X2 OR2X2_296 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_35_), .Y(_36_) );
OR2X2 OR2X2_297 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf1), .B(_36_), .Y(_37_) );
OR2X2 OR2X2_298 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf3), .B(_1128_), .Y(_38_) );
OR2X2 OR2X2_299 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_38_), .Y(_39_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf3), .B(ULA_A[13]), .C(ULA_B[13]), .Y(_40_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_B[13]), .C(_40_), .Y(_43_) );
AND2X2 AND2X2_406 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(ULA_ctrl[2]), .Y(_44_) );
OR2X2 OR2X2_300 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[3]), .B(_44_), .Y(_45_) );
AND2X2 AND2X2_407 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_45_), .Y(_46_) );
AND2X2 AND2X2_408 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_46_), .Y(_47_) );
AND2X2 AND2X2_409 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_25_), .Y(_48_) );
AND2X2 AND2X2_410 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_48_), .Y(_49_) );
OR2X2 OR2X2_301 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_49_), .Y(_50_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_50_), .Y(_0__13_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_B[14]), .Y(_51_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf4), .B(_51_), .Y(_53_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_A[14]), .C(ULA_B[14]), .Y(_54_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_54_), .C(_138__bF_buf2), .Y(_55_) );
OR2X2 OR2X2_302 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_1291_), .Y(_56_) );
AND2X2 AND2X2_411 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_244__bF_buf2), .Y(_57_) );
AND2X2 AND2X2_412 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(_664__bF_buf4), .Y(_58_) );
OR2X2 OR2X2_303 ( .gnd(gnd), .vdd(vdd), .A(_447__bF_buf1), .B(_58_), .Y(_59_) );
OR2X2 OR2X2_304 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_59_), .Y(_60_) );
AND2X2 AND2X2_413 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_56_), .Y(_61_) );
OR2X2 OR2X2_305 ( .gnd(gnd), .vdd(vdd), .A(_639__bF_buf2), .B(_61_), .Y(_62_) );
OR2X2 OR2X2_306 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf2), .B(_1182_), .Y(_64_) );
OR2X2 OR2X2_307 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf0), .B(_1188_), .Y(_65_) );
AND2X2 AND2X2_414 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_65_), .Y(_66_) );
OR2X2 OR2X2_308 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf4), .B(_66_), .Y(_67_) );
MUX2X1 MUX2X1_79 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[13]), .B(ULA_A[14]), .S(ULA_B_0_bF_buf0), .Y(_68_) );
AND2X2 AND2X2_415 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_684__bF_buf6), .Y(_69_) );
AND2X2 AND2X2_416 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(ULA_B_1_bF_buf3), .Y(_70_) );
OR2X2 OR2X2_309 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_70_), .Y(_71_) );
AND2X2 AND2X2_417 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_255__bF_buf6), .Y(_72_) );
AND2X2 AND2X2_418 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(ULA_B_2_bF_buf0), .Y(_73_) );
OR2X2 OR2X2_310 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_73_), .Y(_75_) );
AND2X2 AND2X2_419 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_212__bF_buf0), .Y(_76_) );
AND2X2 AND2X2_420 ( .gnd(gnd), .vdd(vdd), .A(_1202_), .B(ULA_B_3_bF_buf4), .Y(_77_) );
OR2X2 OR2X2_311 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .Y(_78_) );
OR2X2 OR2X2_312 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf1), .B(_78_), .Y(_79_) );
OR2X2 OR2X2_313 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf4), .B(_1178_), .Y(_80_) );
OR2X2 OR2X2_314 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_80_), .Y(_81_) );
OR2X2 OR2X2_315 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_B[14]), .Y(_82_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf2), .B(ULA_A[14]), .C(ULA_B[14]), .Y(_83_) );
AND2X2 AND2X2_421 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_82_), .Y(_84_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf1), .B(_84_), .C(_106__bF_buf2), .Y(_85_) );
AND2X2 AND2X2_422 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_85_), .Y(_86_) );
AND2X2 AND2X2_423 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_86_), .Y(_87_) );
AND2X2 AND2X2_424 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_67_), .Y(_88_) );
AND2X2 AND2X2_425 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_88_), .Y(_89_) );
OR2X2 OR2X2_316 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_89_), .Y(_90_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(_0__14_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .Y(_91_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(ULA_B[15]), .Y(_92_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .C(_149__bF_buf4), .Y(_93_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_A[15]), .C(ULA_B[15]), .Y(_95_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_95_), .C(_138__bF_buf2), .Y(_96_) );
AND2X2 AND2X2_426 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_244__bF_buf0), .Y(_97_) );
AND2X2 AND2X2_427 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .B(_664__bF_buf3), .Y(_98_) );
OR2X2 OR2X2_317 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_99_) );
OR2X2 OR2X2_318 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_99_), .Y(_100_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf1), .B(_1259_), .Y(_101_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf5), .B(_1249_), .Y(_102_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_1065_), .C(_102_), .Y(_103_) );
AND2X2 AND2X2_428 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(ULA_B_3_bF_buf1), .Y(_104_) );
AND2X2 AND2X2_429 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(ULA_B_2_bF_buf1), .Y(_107_) );
AND2X2 AND2X2_430 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(ULA_B_1_bF_buf3), .Y(_108_) );
MUX2X1 MUX2X1_80 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[14]), .B(ULA_A[15]), .S(ULA_B_0_bF_buf2), .Y(_109_) );
AND2X2 AND2X2_431 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_684__bF_buf5), .Y(_110_) );
OR2X2 OR2X2_319 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_110_), .Y(_111_) );
AND2X2 AND2X2_432 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_255__bF_buf1), .Y(_112_) );
OR2X2 OR2X2_320 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_112_), .Y(_113_) );
AND2X2 AND2X2_433 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_212__bF_buf5), .Y(_114_) );
OR2X2 OR2X2_321 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_114_), .Y(_115_) );
OR2X2 OR2X2_322 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf1), .B(_115_), .Y(_116_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .Y(_117_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf1), .B(ULA_A[15]), .C(ULA_B[15]), .Y(_118_) );
AND2X2 AND2X2_434 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_118_), .Y(_119_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf3), .B(_119_), .C(_106__bF_buf3), .Y(_120_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .B(_731_), .Y(_121_) );
OR2X2 OR2X2_323 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_639__bF_buf2), .Y(_122_) );
AND2X2 AND2X2_435 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_729_), .Y(_123_) );
OR2X2 OR2X2_324 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_121_), .Y(_124_) );
AND2X2 AND2X2_436 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_120_), .Y(_125_) );
AND2X2 AND2X2_437 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_116_), .Y(_126_) );
AND2X2 AND2X2_438 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_126_), .Y(_128_) );
AND2X2 AND2X2_439 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_100_), .Y(_129_) );
OR2X2 OR2X2_325 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_129_), .Y(_130_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_130_), .Y(_0__15_) );
OR2X2 OR2X2_326 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_678_), .Y(_131_) );
OR2X2 OR2X2_327 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_131_), .Y(_132_) );
OR2X2 OR2X2_328 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf3), .B(_727_), .Y(_133_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[16]), .B(ULA_B[16]), .Y(_134_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[16]), .B(ULA_B[16]), .Y(_135_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_136_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf5), .B(_136_), .C(_134_), .Y(_139_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf2), .B(_139_), .C(_106__bF_buf0), .Y(_140_) );
AND2X2 AND2X2_440 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_133_), .Y(_141_) );
MUX2X1 MUX2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_1386_), .S(_684__bF_buf6), .Y(_142_) );
MUX2X1 MUX2X1_82 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[15]), .B(ULA_A[16]), .S(ULA_B_0_bF_buf0), .Y(_143_) );
MUX2X1 MUX2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_68_), .S(_684__bF_buf6), .Y(_144_) );
MUX2X1 MUX2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_142_), .S(_255__bF_buf1), .Y(_145_) );
AND2X2 AND2X2_441 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_212__bF_buf0), .Y(_146_) );
AND2X2 AND2X2_442 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(ULA_B_3_bF_buf7), .Y(_147_) );
OR2X2 OR2X2_329 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_4_bF_buf1), .B(_147_), .Y(_148_) );
OR2X2 OR2X2_330 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_146_), .Y(_150_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(ULA_A[0]), .C(ULA_B_4_bF_buf3), .Y(_151_) );
AND2X2 AND2X2_443 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .Y(_152_) );
OR2X2 OR2X2_331 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_152_), .Y(_153_) );
AND2X2 AND2X2_444 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_141_), .Y(_154_) );
AND2X2 AND2X2_445 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_132_), .Y(_155_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf1), .B(_135_), .Y(_156_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(_136_), .Y(_157_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .C(_138__bF_buf3), .Y(_158_) );
OR2X2 OR2X2_332 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_155_), .Y(_159_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_159_), .Y(_0__16_) );
MUX2X1 MUX2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1140_), .S(_255__bF_buf6), .Y(_160_) );
AND2X2 AND2X2_446 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(ULA_B_1_bF_buf3), .Y(_161_) );
MUX2X1 MUX2X1_86 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[16]), .B(ULA_A[17]), .S(ULA_B_0_bF_buf0), .Y(_162_) );
AND2X2 AND2X2_447 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_684__bF_buf3), .Y(_163_) );
OR2X2 OR2X2_333 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_163_), .Y(_164_) );
MUX2X1 MUX2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_32_), .S(_255__bF_buf4), .Y(_165_) );
MUX2X1 MUX2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_160_), .S(_212__bF_buf3), .Y(_166_) );
AND2X2 AND2X2_448 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_728_), .Y(_167_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_841_), .C(_63_), .Y(_168_) );
OR2X2 OR2X2_334 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_167_), .Y(_170_) );
OR2X2 OR2X2_335 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_772_), .Y(_171_) );
OR2X2 OR2X2_336 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf0), .B(_833_), .Y(_172_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[17]), .B(ULA_B[17]), .Y(_173_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[17]), .B(ULA_B[17]), .Y(_174_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_174_), .Y(_175_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf5), .B(_175_), .C(_173_), .Y(_176_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf0), .B(_176_), .C(_106__bF_buf4), .Y(_177_) );
AND2X2 AND2X2_449 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_177_), .Y(_178_) );
AND2X2 AND2X2_450 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_171_), .Y(_179_) );
AND2X2 AND2X2_451 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_170_), .Y(_182_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf1), .B(_174_), .Y(_183_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(_175_), .Y(_184_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .C(_138__bF_buf3), .Y(_185_) );
OR2X2 OR2X2_337 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_182_), .Y(_186_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_186_), .Y(_0__17_) );
OR2X2 OR2X2_338 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_871_), .Y(_187_) );
OR2X2 OR2X2_339 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf1), .B(_937_), .Y(_188_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[18]), .B(ULA_B[18]), .Y(_189_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[18]), .B(ULA_B[18]), .Y(_190_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_191_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf4), .B(_191_), .C(_189_), .Y(_192_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf2), .B(_192_), .C(_106__bF_buf0), .Y(_193_) );
AND2X2 AND2X2_452 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_188_), .Y(_194_) );
MUX2X1 MUX2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_1460_), .S(_684__bF_buf6), .Y(_195_) );
MUX2X1 MUX2X1_90 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[17]), .B(ULA_A[18]), .S(ULA_B_0_bF_buf6), .Y(_196_) );
MUX2X1 MUX2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_143_), .S(_684__bF_buf6), .Y(_197_) );
MUX2X1 MUX2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_195_), .S(_255__bF_buf2), .Y(_198_) );
AND2X2 AND2X2_453 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_212__bF_buf0), .Y(_199_) );
AND2X2 AND2X2_454 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .B(ULA_B_3_bF_buf7), .Y(_200_) );
OR2X2 OR2X2_340 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_199_), .Y(_202_) );
AND2X2 AND2X2_455 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_728_), .Y(_203_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_949_), .Y(_204_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_204_), .C(_63_), .Y(_205_) );
OR2X2 OR2X2_341 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_205_), .Y(_206_) );
AND2X2 AND2X2_456 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_194_), .Y(_207_) );
AND2X2 AND2X2_457 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_187_), .Y(_208_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf2), .B(_190_), .Y(_209_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(_191_), .Y(_210_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_210_), .C(_138__bF_buf4), .Y(_211_) );
OR2X2 OR2X2_342 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_208_), .Y(_214_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_214_), .Y(_0__18_) );
AND2X2 AND2X2_458 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(ULA_B_3_bF_buf2), .Y(_215_) );
AND2X2 AND2X2_459 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(ULA_B_2_bF_buf7), .Y(_216_) );
AND2X2 AND2X2_460 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(ULA_B_1_bF_buf1), .Y(_217_) );
MUX2X1 MUX2X1_93 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[18]), .B(ULA_A[19]), .S(ULA_B_0_bF_buf0), .Y(_218_) );
AND2X2 AND2X2_461 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_684__bF_buf3), .Y(_219_) );
OR2X2 OR2X2_343 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_219_), .Y(_220_) );
AND2X2 AND2X2_462 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_255__bF_buf1), .Y(_221_) );
OR2X2 OR2X2_344 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_221_), .Y(_222_) );
AND2X2 AND2X2_463 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_212__bF_buf3), .Y(_224_) );
OR2X2 OR2X2_345 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_224_), .Y(_225_) );
AND2X2 AND2X2_464 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_728_), .Y(_226_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_1024_), .C(_63_), .Y(_227_) );
OR2X2 OR2X2_346 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_227_), .Y(_228_) );
OR2X2 OR2X2_347 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_978_), .Y(_229_) );
OR2X2 OR2X2_348 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf0), .B(_1018_), .Y(_230_) );
OR2X2 OR2X2_349 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[19]), .B(ULA_B[19]), .Y(_231_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf5), .B(ULA_A[19]), .C(ULA_B[19]), .Y(_232_) );
AND2X2 AND2X2_465 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_231_), .Y(_233_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf0), .B(_233_), .C(_106__bF_buf4), .Y(_235_) );
AND2X2 AND2X2_466 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_235_), .Y(_236_) );
AND2X2 AND2X2_467 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_236_), .Y(_237_) );
AND2X2 AND2X2_468 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_228_), .Y(_238_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[19]), .B(ULA_B[19]), .Y(_239_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf1), .B(_239_), .Y(_240_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(ULA_A[19]), .C(ULA_B[19]), .Y(_241_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(_138__bF_buf4), .Y(_242_) );
OR2X2 OR2X2_350 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_238_), .Y(_243_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_0__19_) );
OR2X2 OR2X2_351 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_1044_), .Y(_245_) );
AND2X2 AND2X2_469 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(ULA_B_3_bF_buf1), .Y(_246_) );
MUX2X1 MUX2X1_94 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[19]), .B(ULA_A[20]), .S(ULA_B_0_bF_buf0), .Y(_247_) );
AND2X2 AND2X2_470 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_684__bF_buf3), .Y(_248_) );
AND2X2 AND2X2_471 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(ULA_B_1_bF_buf1), .Y(_249_) );
OR2X2 OR2X2_352 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_249_), .Y(_250_) );
AND2X2 AND2X2_472 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_255__bF_buf1), .Y(_251_) );
AND2X2 AND2X2_473 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_684__bF_buf6), .Y(_252_) );
AND2X2 AND2X2_474 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(ULA_B_1_bF_buf3), .Y(_253_) );
OR2X2 OR2X2_353 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .Y(_254_) );
AND2X2 AND2X2_475 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(ULA_B_2_bF_buf7), .Y(_256_) );
OR2X2 OR2X2_354 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_256_), .Y(_257_) );
AND2X2 AND2X2_476 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_212__bF_buf5), .Y(_258_) );
OR2X2 OR2X2_355 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_258_), .Y(_259_) );
AND2X2 AND2X2_477 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_728_), .Y(_260_) );
AND2X2 AND2X2_478 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(ULA_B_4_bF_buf2), .Y(_261_) );
OR2X2 OR2X2_356 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_261_), .Y(_262_) );
OR2X2 OR2X2_357 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_262_), .Y(_263_) );
OR2X2 OR2X2_358 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf2), .B(_1063_), .Y(_264_) );
OR2X2 OR2X2_359 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[20]), .B(ULA_B[20]), .Y(_265_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf5), .B(ULA_A[20]), .C(ULA_B[20]), .Y(_267_) );
AND2X2 AND2X2_479 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_265_), .Y(_268_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf0), .B(_268_), .C(_106__bF_buf4), .Y(_269_) );
AND2X2 AND2X2_480 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_269_), .Y(_270_) );
AND2X2 AND2X2_481 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_270_), .Y(_271_) );
AND2X2 AND2X2_482 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_245_), .Y(_272_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[20]), .B(ULA_B[20]), .Y(_273_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf1), .B(_273_), .Y(_274_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf3), .B(ULA_A[20]), .C(ULA_B[20]), .Y(_275_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_275_), .C(_138__bF_buf0), .Y(_276_) );
OR2X2 OR2X2_360 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_272_), .Y(_278_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_278_), .Y(_0__20_) );
OR2X2 OR2X2_361 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_1104_), .Y(_279_) );
OR2X2 OR2X2_362 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf4), .B(_1134_), .Y(_280_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[21]), .B(ULA_B[21]), .Y(_281_) );
AND2X2 AND2X2_483 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[21]), .B(ULA_B[21]), .Y(_282_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf2), .B(_282_), .C(_281_), .Y(_283_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf1), .B(_283_), .C(_106__bF_buf2), .Y(_284_) );
AND2X2 AND2X2_484 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_284_), .Y(_285_) );
AND2X2 AND2X2_485 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(ULA_B_2_bF_buf7), .Y(_286_) );
AND2X2 AND2X2_486 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(ULA_B_1_bF_buf1), .Y(_288_) );
MUX2X1 MUX2X1_95 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[20]), .B(ULA_A[21]), .S(ULA_B_0_bF_buf0), .Y(_289_) );
AND2X2 AND2X2_487 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_684__bF_buf3), .Y(_290_) );
OR2X2 OR2X2_363 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_290_), .Y(_291_) );
AND2X2 AND2X2_488 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_255__bF_buf1), .Y(_292_) );
OR2X2 OR2X2_364 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_292_), .Y(_293_) );
AND2X2 AND2X2_489 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_212__bF_buf5), .Y(_294_) );
AND2X2 AND2X2_490 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(ULA_B_3_bF_buf1), .Y(_295_) );
OR2X2 OR2X2_365 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .Y(_296_) );
AND2X2 AND2X2_491 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_728_), .Y(_297_) );
AND2X2 AND2X2_492 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(ULA_B_4_bF_buf2), .Y(_299_) );
OR2X2 OR2X2_366 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_299_), .Y(_300_) );
OR2X2 OR2X2_367 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_300_), .Y(_301_) );
AND2X2 AND2X2_493 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_285_), .Y(_302_) );
AND2X2 AND2X2_494 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_279_), .Y(_303_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_138__bF_buf1), .Y(_304_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(_282_), .Y(_305_) );
AND2X2 AND2X2_495 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_305_), .Y(_306_) );
OR2X2 OR2X2_368 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_303_), .Y(_307_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_307_), .Y(_0__21_) );
OR2X2 OR2X2_369 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_1164_), .Y(_309_) );
OR2X2 OR2X2_370 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf1), .B(_1184_), .Y(_310_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[22]), .B(ULA_B[22]), .Y(_311_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[22]), .B(ULA_B[22]), .Y(_312_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_312_), .Y(_313_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf4), .B(_313_), .C(_311_), .Y(_314_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf0), .B(_314_), .C(_106__bF_buf4), .Y(_315_) );
AND2X2 AND2X2_496 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_310_), .Y(_316_) );
MUX2X1 MUX2X1_96 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[21]), .B(ULA_A[22]), .S(ULA_B_0_bF_buf0), .Y(_317_) );
AND2X2 AND2X2_497 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_684__bF_buf6), .Y(_318_) );
AND2X2 AND2X2_498 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(ULA_B_1_bF_buf1), .Y(_320_) );
OR2X2 OR2X2_371 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_320_), .Y(_321_) );
AND2X2 AND2X2_499 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_255__bF_buf6), .Y(_322_) );
AND2X2 AND2X2_500 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_684__bF_buf3), .Y(_323_) );
AND2X2 AND2X2_501 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(ULA_B_1_bF_buf1), .Y(_324_) );
OR2X2 OR2X2_372 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_324_), .Y(_325_) );
AND2X2 AND2X2_502 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(ULA_B_2_bF_buf7), .Y(_326_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_326_), .C(_212__bF_buf0), .Y(_327_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_73_), .C(ULA_B_3_bF_buf7), .Y(_328_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_328_), .C(ULA_B_4_bF_buf1), .Y(_329_) );
AND2X2 AND2X2_503 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(ULA_B_4_bF_buf1), .Y(_331_) );
OR2X2 OR2X2_373 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_331_), .Y(_332_) );
OR2X2 OR2X2_374 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_329_), .Y(_333_) );
AND2X2 AND2X2_504 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_316_), .Y(_334_) );
AND2X2 AND2X2_505 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_309_), .Y(_335_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf2), .B(_312_), .Y(_336_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf1), .B(_313_), .Y(_337_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_337_), .C(_138__bF_buf4), .Y(_338_) );
OR2X2 OR2X2_375 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_335_), .Y(_339_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_339_), .Y(_0__22_) );
OR2X2 OR2X2_376 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_1224_), .Y(_341_) );
OR2X2 OR2X2_377 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf2), .B(_1252_), .Y(_342_) );
OR2X2 OR2X2_378 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[23]), .B(ULA_B[23]), .Y(_343_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf1), .B(ULA_A[23]), .C(ULA_B[23]), .Y(_344_) );
AND2X2 AND2X2_506 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_343_), .Y(_345_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf3), .B(_345_), .C(_106__bF_buf3), .Y(_346_) );
AND2X2 AND2X2_507 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_346_), .Y(_347_) );
AND2X2 AND2X2_508 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(ULA_B_2_bF_buf7), .Y(_348_) );
AND2X2 AND2X2_509 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(ULA_B_1_bF_buf1), .Y(_349_) );
MUX2X1 MUX2X1_97 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[22]), .B(ULA_A[23]), .S(ULA_B_0_bF_buf0), .Y(_350_) );
AND2X2 AND2X2_510 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_684__bF_buf3), .Y(_352_) );
OR2X2 OR2X2_379 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_352_), .Y(_353_) );
AND2X2 AND2X2_511 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_255__bF_buf1), .Y(_354_) );
OR2X2 OR2X2_380 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_354_), .Y(_355_) );
AND2X2 AND2X2_512 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_212__bF_buf5), .Y(_356_) );
AND2X2 AND2X2_513 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(ULA_B_3_bF_buf2), .Y(_357_) );
OR2X2 OR2X2_381 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_357_), .Y(_358_) );
AND2X2 AND2X2_514 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_728_), .Y(_359_) );
AND2X2 AND2X2_515 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(ULA_B_4_bF_buf0), .Y(_360_) );
OR2X2 OR2X2_382 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_360_), .Y(_361_) );
OR2X2 OR2X2_383 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_361_), .Y(_363_) );
AND2X2 AND2X2_516 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_347_), .Y(_364_) );
AND2X2 AND2X2_517 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_341_), .Y(_365_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[23]), .B(ULA_B[23]), .Y(_366_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf0), .B(_366_), .Y(_367_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .B(ULA_A[23]), .C(ULA_B[23]), .Y(_368_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_368_), .C(_138__bF_buf0), .Y(_369_) );
OR2X2 OR2X2_384 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_365_), .Y(_370_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_370_), .Y(_0__23_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[24]), .B(ULA_B[24]), .Y(_371_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf4), .B(_371_), .Y(_373_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf2), .B(ULA_A[24]), .C(ULA_B[24]), .Y(_374_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_374_), .C(_138__bF_buf2), .Y(_375_) );
OR2X2 OR2X2_385 ( .gnd(gnd), .vdd(vdd), .A(_244__bF_buf1), .B(_649_), .Y(_376_) );
OR2X2 OR2X2_386 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_662_), .Y(_377_) );
OR2X2 OR2X2_387 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf2), .B(_1317_), .Y(_378_) );
OR2X2 OR2X2_388 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[24]), .B(ULA_B[24]), .Y(_379_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf1), .B(ULA_A[24]), .C(ULA_B[24]), .Y(_380_) );
AND2X2 AND2X2_518 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_379_), .Y(_381_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf3), .B(_381_), .C(_106__bF_buf4), .Y(_382_) );
AND2X2 AND2X2_519 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_382_), .Y(_384_) );
AND2X2 AND2X2_520 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_377_), .Y(_385_) );
AND2X2 AND2X2_521 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(ULA_B_3_bF_buf2), .Y(_386_) );
AND2X2 AND2X2_522 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(ULA_B_1_bF_buf3), .Y(_387_) );
MUX2X1 MUX2X1_98 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[23]), .B(ULA_A[24]), .S(ULA_B_0_bF_buf2), .Y(_388_) );
AND2X2 AND2X2_523 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_684__bF_buf5), .Y(_389_) );
OR2X2 OR2X2_389 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_389_), .Y(_390_) );
OR2X2 OR2X2_390 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .B(_390_), .Y(_391_) );
OR2X2 OR2X2_391 ( .gnd(gnd), .vdd(vdd), .A(_255__bF_buf1), .B(_250_), .Y(_392_) );
AND2X2 AND2X2_524 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_212__bF_buf3), .Y(_393_) );
AND2X2 AND2X2_525 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_391_), .Y(_395_) );
OR2X2 OR2X2_392 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf2), .B(_395_), .Y(_396_) );
OR2X2 OR2X2_393 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_386_), .Y(_397_) );
OR2X2 OR2X2_394 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_52_), .Y(_398_) );
OR2X2 OR2X2_395 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_1315_), .Y(_399_) );
AND2X2 AND2X2_526 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_399_), .Y(_400_) );
AND2X2 AND2X2_527 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_385_), .Y(_401_) );
OR2X2 OR2X2_396 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_401_), .Y(_402_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_402_), .Y(_0__24_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[25]), .B(ULA_B[25]), .Y(_403_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf3), .B(_403_), .Y(_405_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(ULA_A[25]), .C(ULA_B[25]), .Y(_406_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_406_), .C(_138__bF_buf1), .Y(_407_) );
OR2X2 OR2X2_397 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_762_), .Y(_408_) );
OR2X2 OR2X2_398 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf3), .B(_1359_), .Y(_409_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf0), .B(ULA_A[25]), .C(ULA_B[25]), .Y(_410_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[25]), .B(ULA_B[25]), .C(_410_), .Y(_411_) );
AND2X2 AND2X2_528 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(ULA_ctrl[2]), .Y(_412_) );
OR2X2 OR2X2_399 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[3]), .B(_412_), .Y(_413_) );
AND2X2 AND2X2_529 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_413_), .Y(_414_) );
AND2X2 AND2X2_530 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_408_), .Y(_416_) );
OR2X2 OR2X2_400 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_1354_), .Y(_417_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .B(_32_), .Y(_418_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_255__bF_buf4), .B(_164_), .Y(_419_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_419_), .C(_212__bF_buf3), .Y(_420_) );
AND2X2 AND2X2_531 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(ULA_B_1_bF_buf3), .Y(_421_) );
MUX2X1 MUX2X1_99 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[24]), .B(ULA_A[25]), .S(ULA_B_0_bF_buf2), .Y(_422_) );
AND2X2 AND2X2_532 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_684__bF_buf5), .Y(_423_) );
OR2X2 OR2X2_401 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_423_), .Y(_424_) );
AND2X2 AND2X2_533 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_255__bF_buf4), .Y(_425_) );
AND2X2 AND2X2_534 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(ULA_B_2_bF_buf7), .Y(_427_) );
OR2X2 OR2X2_402 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_427_), .Y(_428_) );
AND2X2 AND2X2_535 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_212__bF_buf3), .Y(_429_) );
OR2X2 OR2X2_403 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf2), .B(_429_), .Y(_430_) );
OR2X2 OR2X2_404 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_420_), .Y(_431_) );
AND2X2 AND2X2_536 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_417_), .Y(_432_) );
AND2X2 AND2X2_537 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_416_), .Y(_433_) );
OR2X2 OR2X2_405 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_433_), .Y(_434_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_434_), .Y(_0__25_) );
OR2X2 OR2X2_406 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf4), .B(_1396_), .Y(_435_) );
OR2X2 OR2X2_407 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[26]), .B(ULA_B[26]), .Y(_437_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf2), .B(ULA_A[26]), .C(ULA_B[26]), .Y(_438_) );
AND2X2 AND2X2_538 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_437_), .Y(_439_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf1), .B(_439_), .C(_106__bF_buf2), .Y(_440_) );
AND2X2 AND2X2_539 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_440_), .Y(_441_) );
OR2X2 OR2X2_408 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_1394_), .Y(_442_) );
AND2X2 AND2X2_540 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_441_), .Y(_443_) );
OR2X2 OR2X2_409 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_859_), .Y(_444_) );
AND2X2 AND2X2_541 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(ULA_B_3_bF_buf7), .Y(_445_) );
AND2X2 AND2X2_542 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(ULA_B_1_bF_buf3), .Y(_446_) );
MUX2X1 MUX2X1_100 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[25]), .B(ULA_A[26]), .S(ULA_B_0_bF_buf2), .Y(_448_) );
AND2X2 AND2X2_543 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_684__bF_buf5), .Y(_449_) );
OR2X2 OR2X2_410 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_449_), .Y(_450_) );
OR2X2 OR2X2_411 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf1), .B(_450_), .Y(_451_) );
OR2X2 OR2X2_412 ( .gnd(gnd), .vdd(vdd), .A(_255__bF_buf6), .B(_321_), .Y(_452_) );
AND2X2 AND2X2_544 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_212__bF_buf3), .Y(_453_) );
AND2X2 AND2X2_545 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_451_), .Y(_454_) );
OR2X2 OR2X2_413 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf2), .B(_454_), .Y(_455_) );
OR2X2 OR2X2_414 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_445_), .Y(_456_) );
AND2X2 AND2X2_546 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_444_), .Y(_457_) );
AND2X2 AND2X2_547 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_443_), .Y(_459_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[26]), .B(ULA_B[26]), .Y(_460_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf3), .B(_460_), .Y(_461_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(ULA_A[26]), .C(ULA_B[26]), .Y(_462_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_462_), .C(_138__bF_buf1), .Y(_463_) );
OR2X2 OR2X2_415 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_459_), .Y(_464_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_464_), .Y(_0__26_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[27]), .B(ULA_B[27]), .Y(_465_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf0), .B(_465_), .Y(_466_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .B(ULA_A[27]), .C(ULA_B[27]), .Y(_467_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_467_), .C(_138__bF_buf0), .Y(_469_) );
OR2X2 OR2X2_416 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_966_), .Y(_470_) );
OR2X2 OR2X2_417 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf2), .B(_1434_), .Y(_471_) );
OR2X2 OR2X2_418 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[27]), .B(ULA_B[27]), .Y(_472_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf1), .B(ULA_A[27]), .C(ULA_B[27]), .Y(_473_) );
AND2X2 AND2X2_548 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_472_), .Y(_474_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf3), .B(_474_), .C(_106__bF_buf3), .Y(_475_) );
AND2X2 AND2X2_549 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_475_), .Y(_476_) );
AND2X2 AND2X2_550 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_470_), .Y(_477_) );
OR2X2 OR2X2_419 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_1428_), .Y(_478_) );
AND2X2 AND2X2_551 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(ULA_B_3_bF_buf2), .Y(_480_) );
AND2X2 AND2X2_552 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(ULA_B_2_bF_buf7), .Y(_481_) );
AND2X2 AND2X2_553 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(ULA_B_1_bF_buf3), .Y(_482_) );
MUX2X1 MUX2X1_101 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[26]), .B(ULA_A[27]), .S(ULA_B_0_bF_buf2), .Y(_483_) );
AND2X2 AND2X2_554 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_684__bF_buf5), .Y(_484_) );
OR2X2 OR2X2_420 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_484_), .Y(_485_) );
AND2X2 AND2X2_555 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_255__bF_buf4), .Y(_486_) );
OR2X2 OR2X2_421 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_486_), .Y(_487_) );
AND2X2 AND2X2_556 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_212__bF_buf3), .Y(_488_) );
OR2X2 OR2X2_422 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf2), .B(_488_), .Y(_489_) );
OR2X2 OR2X2_423 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_489_), .Y(_491_) );
AND2X2 AND2X2_557 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_491_), .Y(_492_) );
AND2X2 AND2X2_558 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_477_), .Y(_493_) );
OR2X2 OR2X2_424 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_493_), .Y(_494_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_494_), .Y(_0__27_) );
AND2X2 AND2X2_559 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[28]), .B(ULA_B[28]), .Y(_495_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(_495_), .Y(_496_) );
AND2X2 AND2X2_560 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_496_), .Y(_497_) );
OR2X2 OR2X2_425 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_1469_), .Y(_498_) );
OR2X2 OR2X2_426 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf4), .B(_1475_), .Y(_499_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[28]), .B(ULA_B[28]), .Y(_501_) );
AND2X2 AND2X2_561 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(ULA_ctrl_1_bF_buf2), .Y(_502_) );
OR2X2 OR2X2_427 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_501_), .Y(_503_) );
AND2X2 AND2X2_562 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(ULA_ctrl[2]), .Y(_504_) );
OR2X2 OR2X2_428 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl[3]), .B(_504_), .Y(_505_) );
AND2X2 AND2X2_563 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_505_), .Y(_506_) );
AND2X2 AND2X2_564 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_506_), .Y(_507_) );
OR2X2 OR2X2_429 ( .gnd(gnd), .vdd(vdd), .A(_277__bF_buf2), .B(_654_), .Y(_508_) );
OR2X2 OR2X2_430 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_376_), .Y(_509_) );
AND2X2 AND2X2_565 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(ULA_B_2_bF_buf1), .Y(_510_) );
MUX2X1 MUX2X1_102 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[27]), .B(ULA_A[28]), .S(ULA_B_0_bF_buf2), .Y(_512_) );
AND2X2 AND2X2_566 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_684__bF_buf5), .Y(_513_) );
AND2X2 AND2X2_567 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(ULA_B_1_bF_buf3), .Y(_514_) );
OR2X2 OR2X2_431 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_514_), .Y(_515_) );
AND2X2 AND2X2_568 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_255__bF_buf1), .Y(_516_) );
OR2X2 OR2X2_432 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_516_), .Y(_517_) );
OR2X2 OR2X2_433 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf2), .B(_517_), .Y(_518_) );
OR2X2 OR2X2_434 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf5), .B(_257_), .Y(_519_) );
AND2X2 AND2X2_569 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_519_), .Y(_520_) );
OR2X2 OR2X2_435 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf2), .B(_520_), .Y(_521_) );
AND2X2 AND2X2_570 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_509_), .Y(_523_) );
AND2X2 AND2X2_571 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_507_), .Y(_524_) );
OR2X2 OR2X2_436 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_524_), .Y(_525_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_525_), .Y(_0__28_) );
AND2X2 AND2X2_572 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(ULA_B_4_bF_buf0), .Y(_526_) );
AND2X2 AND2X2_573 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(ULA_B_3_bF_buf1), .Y(_527_) );
AND2X2 AND2X2_574 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(ULA_B_1_bF_buf5), .Y(_528_) );
MUX2X1 MUX2X1_103 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[28]), .B(ULA_A[29]), .S(ULA_B_0_bF_buf2), .Y(_529_) );
AND2X2 AND2X2_575 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_684__bF_buf5), .Y(_530_) );
OR2X2 OR2X2_437 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_530_), .Y(_531_) );
AND2X2 AND2X2_576 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_255__bF_buf4), .Y(_533_) );
AND2X2 AND2X2_577 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(ULA_B_2_bF_buf7), .Y(_534_) );
OR2X2 OR2X2_438 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_534_), .Y(_535_) );
AND2X2 AND2X2_578 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_212__bF_buf5), .Y(_536_) );
OR2X2 OR2X2_439 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_536_), .Y(_537_) );
AND2X2 AND2X2_579 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_728_), .Y(_538_) );
OR2X2 OR2X2_440 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_538_), .Y(_539_) );
OR2X2 OR2X2_441 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_539_), .Y(_540_) );
OR2X2 OR2X2_442 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_376_), .Y(_541_) );
OR2X2 OR2X2_443 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf2), .B(_38_), .Y(_542_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[29]), .B(ULA_B[29]), .Y(_544_) );
AND2X2 AND2X2_580 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[29]), .B(ULA_B[29]), .Y(_545_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf0), .B(_545_), .C(_544_), .Y(_546_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf4), .B(_546_), .C(_106__bF_buf1), .Y(_547_) );
AND2X2 AND2X2_581 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_542_), .Y(_548_) );
AND2X2 AND2X2_582 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_541_), .Y(_549_) );
AND2X2 AND2X2_583 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_549_), .Y(_550_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(_545_), .Y(_551_) );
AND2X2 AND2X2_584 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_551_), .Y(_552_) );
OR2X2 OR2X2_444 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_550_), .Y(_553_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_553_), .Y(_0__29_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[30]), .B(ULA_B[30]), .Y(_555_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf3), .B(_555_), .Y(_556_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf5), .B(ULA_A[30]), .C(ULA_B[30]), .Y(_557_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_557_), .C(_138__bF_buf1), .Y(_558_) );
OR2X2 OR2X2_445 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_78_), .Y(_559_) );
OR2X2 OR2X2_446 ( .gnd(gnd), .vdd(vdd), .A(_705__bF_buf4), .B(_80_), .Y(_560_) );
OR2X2 OR2X2_447 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[30]), .B(ULA_B[30]), .Y(_561_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf2), .B(ULA_A[30]), .C(ULA_B[30]), .Y(_562_) );
AND2X2 AND2X2_585 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_561_), .Y(_563_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf1), .B(_563_), .C(_106__bF_buf2), .Y(_565_) );
AND2X2 AND2X2_586 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_565_), .Y(_566_) );
AND2X2 AND2X2_587 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_566_), .Y(_567_) );
OR2X2 OR2X2_448 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_376_), .Y(_568_) );
MUX2X1 MUX2X1_104 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[29]), .B(ULA_A[30]), .S(ULA_B_0_bF_buf2), .Y(_569_) );
AND2X2 AND2X2_588 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_684__bF_buf5), .Y(_570_) );
AND2X2 AND2X2_589 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(ULA_B_1_bF_buf5), .Y(_571_) );
OR2X2 OR2X2_449 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_2_bF_buf7), .B(_571_), .Y(_572_) );
OR2X2 OR2X2_450 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_572_), .Y(_573_) );
OR2X2 OR2X2_451 ( .gnd(gnd), .vdd(vdd), .A(_255__bF_buf4), .B(_450_), .Y(_574_) );
AND2X2 AND2X2_590 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_573_), .Y(_576_) );
OR2X2 OR2X2_452 ( .gnd(gnd), .vdd(vdd), .A(ULA_B_3_bF_buf2), .B(_576_), .Y(_577_) );
OR2X2 OR2X2_453 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_326_), .Y(_578_) );
OR2X2 OR2X2_454 ( .gnd(gnd), .vdd(vdd), .A(_212__bF_buf0), .B(_578_), .Y(_579_) );
AND2X2 AND2X2_591 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_579_), .Y(_580_) );
OR2X2 OR2X2_455 ( .gnd(gnd), .vdd(vdd), .A(_842__bF_buf3), .B(_580_), .Y(_581_) );
AND2X2 AND2X2_592 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_568_), .Y(_582_) );
AND2X2 AND2X2_593 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_567_), .Y(_583_) );
OR2X2 OR2X2_456 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_583_), .Y(_584_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_584_), .Y(_0__30_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .B(ULA_B[31]), .Y(_586_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_149__bF_buf4), .B(_586_), .Y(_587_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_586_), .Y(_588_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_0_bF_buf4), .B(_588_), .Y(_589_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_589_), .C(_138__bF_buf2), .Y(_590_) );
AND2X2 AND2X2_594 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(ULA_B_3_bF_buf1), .Y(_591_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .B(_960_), .Y(_592_) );
OR2X2 OR2X2_457 ( .gnd(gnd), .vdd(vdd), .A(_684__bF_buf1), .B(_529_), .Y(_593_) );
AND2X2 AND2X2_595 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_593_), .Y(_594_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_684__bF_buf5), .B(ULA_B_0_bF_buf2), .C(ULA_A[30]), .Y(_595_) );
AND2X2 AND2X2_596 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_255__bF_buf6), .Y(_597_) );
AND2X2 AND2X2_597 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_597_), .Y(_598_) );
AND2X2 AND2X2_598 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(ULA_B_2_bF_buf1), .Y(_599_) );
OR2X2 OR2X2_458 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_598_), .Y(_600_) );
AND2X2 AND2X2_599 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_212__bF_buf5), .Y(_601_) );
OR2X2 OR2X2_459 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_601_), .Y(_602_) );
AND2X2 AND2X2_600 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_728_), .Y(_603_) );
AND2X2 AND2X2_601 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(ULA_B_4_bF_buf2), .Y(_604_) );
OR2X2 OR2X2_460 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_604_), .Y(_605_) );
OR2X2 OR2X2_461 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_603_), .Y(_606_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_447__bF_buf2), .C(_705__bF_buf2), .Y(_608_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(ULA_A[31]), .C(_731_), .Y(_609_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(ULA_A[31]), .B(ULA_B[31]), .Y(_610_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(ULA_ctrl_1_bF_buf1), .B(_588_), .C(_610_), .Y(_611_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_74__bF_buf3), .B(_611_), .C(_106__bF_buf3), .Y(_612_) );
AND2X2 AND2X2_602 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_612_), .Y(_613_) );
AND2X2 AND2X2_603 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_613_), .Y(_614_) );
OR2X2 OR2X2_462 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_614_), .Y(_615_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_615_), .Y(_0__31_) );
AND2X2 AND2X2_604 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(_10_), .Y(_616_) );
AND2X2 AND2X2_605 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1410_), .Y(_618_) );
AND2X2 AND2X2_606 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_618_), .Y(_619_) );
AND2X2 AND2X2_607 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_90_), .Y(_620_) );
AND2X2 AND2X2_608 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_130_), .Y(_621_) );
AND2X2 AND2X2_609 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_621_), .Y(_622_) );
AND2X2 AND2X2_610 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1032_), .Y(_623_) );
AND2X2 AND2X2_611 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_955_), .Y(_624_) );
AND2X2 AND2X2_612 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_624_), .Y(_625_) );
AND2X2 AND2X2_613 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1331_), .Y(_626_) );
AND2X2 AND2X2_614 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1213_), .Y(_627_) );
AND2X2 AND2X2_615 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_626_), .Y(_628_) );
AND2X2 AND2X2_616 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_628_), .Y(_629_) );
AND2X2 AND2X2_617 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_622_), .Y(_630_) );
AND2X2 AND2X2_618 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_402_), .Y(_631_) );
AND2X2 AND2X2_619 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_494_), .Y(_632_) );
AND2X2 AND2X2_620 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_632_), .Y(_633_) );
AND2X2 AND2X2_621 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_370_), .Y(_634_) );
AND2X2 AND2X2_622 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_307_), .Y(_635_) );
AND2X2 AND2X2_623 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_635_), .Y(_636_) );
AND2X2 AND2X2_624 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_633_), .Y(_637_) );
AND2X2 AND2X2_625 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_214_), .Y(_640_) );
AND2X2 AND2X2_626 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_243_), .Y(_641_) );
AND2X2 AND2X2_627 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_641_), .Y(_642_) );
AND2X2 AND2X2_628 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_584_), .Y(_643_) );
AND2X2 AND2X2_629 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_525_), .Y(_644_) );
AND2X2 AND2X2_630 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_644_), .Y(_645_) );
AND2X2 AND2X2_631 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_747_), .Y(_646_) );
AND2X2 AND2X2_632 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_646_), .Y(_647_) );
AND2X2 AND2X2_633 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_637_), .Y(_648_) );
AND2X2 AND2X2_634 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_648_), .Y(zero) );
BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(_1476__0_), .Y(ULA_OUT[0]) );
BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(_1476__1_), .Y(ULA_OUT[1]) );
BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(_1476__2_), .Y(ULA_OUT[2]) );
BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(_1476__3_), .Y(ULA_OUT[3]) );
BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(_1476__4_), .Y(ULA_OUT[4]) );
BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(_1476__5_), .Y(ULA_OUT[5]) );
BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(_1476__6_), .Y(ULA_OUT[6]) );
BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(_1476__7_), .Y(ULA_OUT[7]) );
BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(_1476__8_), .Y(ULA_OUT[8]) );
BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(_1476__9_), .Y(ULA_OUT[9]) );
BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(_1476__10_), .Y(ULA_OUT[10]) );
BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(_1476__11_), .Y(ULA_OUT[11]) );
BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(_1476__12_), .Y(ULA_OUT[12]) );
BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(_1476__13_), .Y(ULA_OUT[13]) );
BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(_1476__14_), .Y(ULA_OUT[14]) );
BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(_1476__15_), .Y(ULA_OUT[15]) );
BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(_1476__16_), .Y(ULA_OUT[16]) );
BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(_1476__17_), .Y(ULA_OUT[17]) );
BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(_1476__18_), .Y(ULA_OUT[18]) );
BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(_1476__19_), .Y(ULA_OUT[19]) );
BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(_1476__20_), .Y(ULA_OUT[20]) );
BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(_1476__21_), .Y(ULA_OUT[21]) );
BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(_1476__22_), .Y(ULA_OUT[22]) );
BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(_1476__23_), .Y(ULA_OUT[23]) );
BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(_1476__24_), .Y(ULA_OUT[24]) );
BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(_1476__25_), .Y(ULA_OUT[25]) );
BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(_1476__26_), .Y(ULA_OUT[26]) );
BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(_1476__27_), .Y(ULA_OUT[27]) );
BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(_1476__28_), .Y(ULA_OUT[28]) );
BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(_1476__29_), .Y(ULA_OUT[29]) );
BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(_1476__30_), .Y(ULA_OUT[30]) );
BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(_1476__31_), .Y(ULA_OUT[31]) );
BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(ULA_flags[0]) );
BUFX2 BUFX2_173 ( .gnd(gnd), .vdd(vdd), .A(_1477__1_), .Y(ULA_flags[1]) );
BUFX2 BUFX2_174 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(ULA_flags[2]) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(zero), .Q(_1477__1_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__0_), .Q(_1476__0_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__1_), .Q(_1476__1_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__2_), .Q(_1476__2_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__3_), .Q(_1476__3_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__4_), .Q(_1476__4_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__5_), .Q(_1476__5_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__6_), .Q(_1476__6_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__7_), .Q(_1476__7_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__8_), .Q(_1476__8_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__9_), .Q(_1476__9_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__10_), .Q(_1476__10_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__11_), .Q(_1476__11_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__12_), .Q(_1476__12_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__13_), .Q(_1476__13_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__14_), .Q(_1476__14_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__15_), .Q(_1476__15_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__16_), .Q(_1476__16_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__17_), .Q(_1476__17_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__18_), .Q(_1476__18_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__19_), .Q(_1476__19_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__20_), .Q(_1476__20_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__21_), .Q(_1476__21_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__22_), .Q(_1476__22_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__23_), .Q(_1476__23_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__24_), .Q(_1476__24_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__25_), .Q(_1476__25_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__26_), .Q(_1476__26_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__27_), .Q(_1476__27_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__28_), .Q(_1476__28_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__29_), .Q(_1476__29_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__30_), .Q(_1476__30_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__31_), .Q(_1476__31_) );
endmodule
