`include "const.v"

module NRISC_UP(
IDATA_CORE_addr,
IDATA_CORE_out,
IDATA_CORE_clk,
DDATA_CORE_addr,
DDATA_CORE_out,
DDATA_CORE_in,
DDATA_CORE_load,
DDATA_CORE_write,
DDATA_CORE_ctrl,
CORE_ctrl,
clk,											//Main clk source
rst
);

//Parameter numero de bits
parameter TAM = `TAM;
//D-Data defs
parameter N_DData =  `N_DData;
//I-Data Defs
parameter N_IData = `N_IData;
//PC Defs
parameter STACK_TAM =`STACK_TAM;
parameter ADDR_TAM  =`ADDR_TAM;


input wire clk;
input wire rst;
//-------------portas de entrada------------------------------------------------------------------
 wire [TAM-1:0] ULA_A;
 wire [TAM-1:0] ULA_B;
// wire incdec;
  wire [3:0] ULA_ctrl;// 3fios operacao 1 fio complemento

//-------------portas de saida--------------------------------------------------------------------
 wire [TAM-1:0] ULA_OUT;
 wire [2:0] ULA_flags;
//CORE

 input wire [2:0] CORE_ctrl;
 wire [4:0] CORE_Status_ctrl;
//Instruction
 wire [15:0] CORE_InstructionIN;
 wire [1:0]CORE_InstructionToULAMux;
 //REG
 wire [TAM-1:0] STACK_R1;
 wire [TAM-1:0] REG_A;
 wire [TAM-1:0] REG_B;
 wire CORE_REG_write;
 wire [3:0] CORE_REG_RFD;

//ULA
 wire [2:0] CORE_ULA_flags;
 wire [3:0] CORE_ULA_ctrl;
 wire CORE_ULAMux_inc_dec;
 wire CORE_ULA_REGA_Stall;
 wire CORE_ULA_REGB_Stall;
//wire ctrl
 wire [3:0] CORE_wire_RD;
 wire [3:0] CORE_wire_RF1;
 wire [3:0] CORE_wire_RF2;
 wire CORE_wire_write;

//STACK
 wire [1:0] CORE_STACK_ctrl;
//PC
 wire [1:0] CORE_PC_ctrl;
 wire CORE_PC_clk;
//Interrupt Vector
 wire [7:0] CORE_INT_CHA ;
 wire [1:0] CORE_INT_ctrl ;

 //I-Data

  output wire [N_IData-1:0] IDATA_CORE_addr;
  input wire [TAM-1:0] IDATA_CORE_out;
  output wire IDATA_CORE_clk;

  //D-Data
  output wire [N_DData-1:0] DDATA_CORE_addr;
  input wire [TAM-1:0] DDATA_CORE_out;
  output wire [N_DData-1:0] DDATA_CORE_in;
  output wire DDATA_CORE_load;
  output wire DDATA_CORE_write;
  output wire [2:0] DDATA_CORE_ctrl;


  wire CORE_DATA_ADDR_mux;				//DATA clk
  wire CORE_DATA_REGMux;					//DATA to REGs MUX


// pc ctrl
  wire [TAM-1:0] REG_R1;
  wire [7:0] INTERRUPT_ch;
  wire INTERRUPT_flag;

// Pipeline ID
  reg [7:0] InstructionIN;
  always @ ( posedge clk ) begin
    InstructionIN= CORE_InstructionIN[7:0];
  end

// Pipeline EXEC
    //REGS
    reg [3:0] REG_RFD_exec_pipe;
    reg REG_Write_exec_pipe;
    //D-Data
    reg CORE_DATA_write_exec_pipe;
    reg CORE_DATA_load_exec_pipe;
    reg [2:0]CORE_DATA_ctrl_exec_pipe;
    reg CORE_DATA_ADDR_mux_exec_pipe;
    reg CORE_DATA_REGMux_exec_pipe;
    reg [TAM-1:0] ULA_out_exec_pipe;

    always @ ( posedge clk ) begin
      REG_RFD_exec_pipe= CORE_REG_RFD;
      REG_Write_exec_pipe=CORE_REG_write;
      CORE_DATA_write_exec_pipe = DDATA_CORE_write;
      CORE_DATA_load_exec_pipe =DDATA_CORE_load;
      CORE_DATA_ctrl_exec_pipe =DDATA_CORE_ctrl;
      CORE_DATA_ADDR_mux_exec_pipe =	ULA_A;
      CORE_DATA_REGMux_exec_pipe =CORE_DATA_REGMux;
      ULA_out_exec_pipe=ULA_OUT;
    end

    assign ULA_B= CORE_InstructionToULAMux[0] | CORE_InstructionToULAMux[1] ?
                  (CORE_InstructionToULAMux[1] ?
                      {{(TAM-9){CORE_InstructionToULAMux[0]&InstructionIN[7]}},InstructionIN[7:0]} :
                      {{(TAM-5){1'b0}},InstructionIN[3:0]} ) :
                  CORE_ULA_REGB_Stall ? ULA_out_exec_pipe : REG_B;
    assign ULA_A= CORE_ULA_REGA_Stall ? ULA_out_exec_pipe : REG_A;


    //WB Pipeline
    reg [3:0] REG_RFD_wb_pipe;
    reg REG_Write_wb_pipe;
    reg [TAM-1:0] REG_RD_wb_pipe;
    always @ ( posedge clk ) begin
      REG_RFD_wb_pipe= REG_RFD_exec_pipe;
      REG_Write_wb_pipe=REG_Write_exec_pipe;
      REG_RD_wb_pipe= CORE_DATA_REGMux_exec_pipe ? DDATA_CORE_out : ULA_out_exec_pipe;
    end

NRISC_PC_ctrl PC(
                .IDATA_CORE_out(IDATA_CORE_out),
                .IDATA_CORE_addr(IDATA_CORE_addr),
                .IDATA_clk(IDATA_CORE_clk),
                .CORE_InstructionIN(CORE_InstructionIN),
                .CORE_PC_ctrl(CORE_PC_ctrl),
                .CORE_STACK_ctrl(CORE_STACK_ctrl),
                .ULA_OUT(ULA_OUT),
                .REG_R1(REG_R1),
                .INTERRUPT_ch(INTERRUPT_ch),
                .INTERRUPT_flag(INTERRUPT_flag),
                .clk(clk),
                .rst(rst)
                );

NRISC_InstructionDecoder ID(
								.CORE_InstructionIN(CORE_InstructionIN),				//instruction input
								.CORE_InstructionToULAMux(CORE_InstructionToULAMux),	//MUX ctrl of instruction in to REGs
								.CORE_ctrl(CORE_ctrl),								//CORE external  ctrl BUS
								.CORE_Status_ctrl(CORE_Status_ctrl),					//CORE status output
								.CORE_ULA_ctrl(CORE_ULA_ctrl),						//ULA  ctrl BUS
								.CORE_ULA_flags(CORE_ULA_flags),						//ULA flags  {M,Z,C}
                .CORE_ULA_REGA_Stall(CORE_ULA_REGA_Stall),
								.CORE_ULA_REGB_Stall(CORE_ULA_REGB_Stall),
								.CORE_REG_RF1(CORE_REG_RF1),							//REGs to ULA ctrl 1
								.CORE_REG_RF2(CORE_REG_RF2),							//REGs to ULA ctrl 2
								.CORE_REG_RFD(CORE_REG_RFD),							//REGs inputs ctrl
								.CORE_REG_write(CORE_REG_write),						//REGs write ctrl
								.CORE_DATA_write(DDATA_CORE_write),					//DATA write ctrl
								.CORE_DATA_load(DDATA_CORE_load),						//DATA load ctrl
								.CORE_DATA_ctrl(DDATA_CORE_ctrl),						//DATA size load/store ctrl
								.CORE_DATA_ADDR_mux(CORE_DATA_ADDR_mux),				//DATA clk
								.CORE_DATA_REGMux(CORE_DATA_REGMux),					//DATA to REGs MUX
								.CORE_STACK_ctrl(CORE_STACK_ctrl),					//CORE to STACK ctrl
								.CORE_PC_ctrl(CORE_PC_ctrl),							//CORE to PC ctrl MUX
								.CORE_PC_clk(CORE_PC_clk),							//PC clk
								.CORE_INT_CHA(CORE_INT_CHA),							//CORE to interrupt vector channel
								.CORE_INT_ctrl(CORE_INT_ctrl),						//CORE to interrupt vector control
								.clk(clk),											//Main clk source
								.rst(rst)												//general rst
								);

NRISC_REGs REGs(
                    .REG_A(REG_A),
                    .REG_B(REG_B),
                    .REG_D(REG_RD_wb_pipe),
                    .REG_RF1(CORE_REG_RF1),
                    .REG_RF2(CORE_REG_RF2),
                    .REG_RFD(REG_RFD_wb_pipe),
                    .REG_R1(STACK_R1),
                    .REG_Write(REG_Write_exec_pipe),
                    .REG_Interrupt_flag(INTERRUPT_flag),
                    .clk(clk),
                    .rst(rst)
                    );

NRISC_ULA ULA(
                    .ULA_A(ULA_A),      //ULA  A
                    .ULA_B(ULA_B),      //ULA  B
                    .ULA_OUT(ULA_OUT),    //  output
                    .ULA_ctrl(CORE_ULA_ctrl),   // comando
                    .ULA_flags(CORE_ULA_flags)  // minus, carry, zero
                    );

endmodule
