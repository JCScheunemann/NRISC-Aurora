magic
tech scmos
magscale 1 4
timestamp 1516325494
use BUFX2  BUFX2_885
timestamp 1516325494
transform 1 0 2 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_526
timestamp 1516325494
transform -1 0 70 0 1 2620
box 0 0 53 49
use BUFX2  BUFX2_898
timestamp 1516325494
transform -1 0 85 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_526
timestamp 1516325494
transform 1 0 86 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_526
timestamp 1516325494
transform -1 0 131 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_520
timestamp 1516325494
transform -1 0 184 0 1 2620
box 0 0 53 49
use MUX2X1  MUX2X1_520
timestamp 1516325494
transform 1 0 184 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_520
timestamp 1516325494
transform -1 0 230 0 1 2620
box 0 0 15 49
use INVX1  INVX1_194
timestamp 1516325494
transform 1 0 230 0 1 2620
box 0 0 11 49
use BUFX2  BUFX2_900
timestamp 1516325494
transform -1 0 256 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_78
timestamp 1516325494
transform -1 0 272 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_494
timestamp 1516325494
transform 1 0 272 0 1 2620
box 0 0 53 49
use BUFX2  BUFX2_902
timestamp 1516325494
transform 1 0 325 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_558
timestamp 1516325494
transform 1 0 340 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_558
timestamp 1516325494
transform -1 0 385 0 1 2620
box 0 0 30 49
use BUFX2  BUFX2_899
timestamp 1516325494
transform 1 0 386 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_488
timestamp 1516325494
transform 1 0 401 0 1 2620
box 0 0 53 49
use MUX2X1  MUX2X1_552
timestamp 1516325494
transform 1 0 454 0 1 2620
box 0 0 30 49
use BUFX2  BUFX2_891
timestamp 1516325494
transform 1 0 485 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_904
timestamp 1516325494
transform -1 0 515 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_890
timestamp 1516325494
transform -1 0 530 0 1 2620
box 0 0 15 49
use INVX1  INVX1_191
timestamp 1516325494
transform 1 0 530 0 1 2620
box 0 0 11 49
use BUFX2  BUFX2_897
timestamp 1516325494
transform -1 0 557 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_124
timestamp 1516325494
transform -1 0 610 0 1 2620
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_508
timestamp 1516325494
transform 1 0 610 0 1 2620
box 0 0 53 49
use BUFX2  BUFX2_894
timestamp 1516325494
transform -1 0 678 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_27
timestamp 1516325494
transform 1 0 678 0 1 2620
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_539
timestamp 1516325494
transform 1 0 732 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_539
timestamp 1516325494
transform 1 0 785 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_880
timestamp 1516325494
transform -1 0 815 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_571
timestamp 1516325494
transform 1 0 815 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_571
timestamp 1516325494
transform -1 0 861 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_507
timestamp 1516325494
transform -1 0 914 0 1 2620
box 0 0 53 49
use BUFX2  BUFX2_893
timestamp 1516325494
transform -1 0 929 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_103
timestamp 1516325494
transform 1 0 929 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_71
timestamp 1516325494
transform 1 0 982 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_71
timestamp 1516325494
transform -1 0 1028 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_519
timestamp 1516325494
transform 1 0 1028 0 1 2620
box 0 0 53 49
use MUX2X1  MUX2X1_519
timestamp 1516325494
transform 1 0 1081 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_519
timestamp 1516325494
transform -1 0 1127 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_461
timestamp 1516325494
transform 1 0 1127 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_333
timestamp 1516325494
transform 1 0 1180 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_333
timestamp 1516325494
transform 1 0 1195 0 1 2620
box 0 0 30 49
use MUX2X1  MUX2X1_119
timestamp 1516325494
transform 1 0 1226 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_119
timestamp 1516325494
transform -1 0 1271 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_23
timestamp 1516325494
transform -1 0 1324 0 1 2620
box 0 0 53 49
use OR2X2  OR2X2_1698
timestamp 1516325494
transform 1 0 1324 0 1 2620
box 0 0 19 49
use MUX2X1  MUX2X1_535
timestamp 1516325494
transform 1 0 1343 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_535
timestamp 1516325494
transform -1 0 1427 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_535
timestamp 1516325494
transform -1 0 1442 0 1 2620
box 0 0 15 49
use OR2X2  OR2X2_1697
timestamp 1516325494
transform 1 0 1442 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1831
timestamp 1516325494
transform 1 0 1461 0 1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_504
timestamp 1516325494
transform -1 0 1488 0 1 2620
box 0 0 8 49
use BUFX2  BUFX2_504
timestamp 1516325494
transform -1 0 1503 0 1 2620
box 0 0 15 49
use OR2X2  OR2X2_1694
timestamp 1516325494
transform 1 0 1503 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1829
timestamp 1516325494
transform -1 0 1541 0 1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_343
timestamp 1516325494
transform 1 0 1541 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_343
timestamp 1516325494
transform 1 0 1556 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_471
timestamp 1516325494
transform 1 0 1587 0 1 2620
box 0 0 53 49
use OR2X2  OR2X2_1695
timestamp 1516325494
transform -1 0 1659 0 1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_87
timestamp 1516325494
transform 1 0 1659 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_151
timestamp 1516325494
transform 1 0 1712 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_151
timestamp 1516325494
transform 1 0 1727 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_740
timestamp 1516325494
transform -1 0 1773 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_742
timestamp 1516325494
transform -1 0 1788 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_375
timestamp 1516325494
transform 1 0 1788 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_933
timestamp 1516325494
transform 1 0 1841 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_878
timestamp 1516325494
transform 1 0 1856 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_736
timestamp 1516325494
transform 1 0 1887 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_407
timestamp 1516325494
transform 1 0 1902 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_183
timestamp 1516325494
transform -1 0 1970 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_183
timestamp 1516325494
transform 1 0 1970 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_357
timestamp 1516325494
transform 1 0 2001 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_915
timestamp 1516325494
transform 1 0 2054 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_860
timestamp 1516325494
transform 1 0 2069 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_165
timestamp 1516325494
transform 1 0 2100 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_165
timestamp 1516325494
transform 1 0 2115 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_746
timestamp 1516325494
transform 1 0 2145 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_744
timestamp 1516325494
transform 1 0 2160 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_389
timestamp 1516325494
transform -1 0 2229 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_741
timestamp 1516325494
transform -1 0 2244 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_165
timestamp 1516325494
transform 1 0 2244 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_716
timestamp 1516325494
transform 1 0 2297 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_229
timestamp 1516325494
transform 1 0 2312 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_229
timestamp 1516325494
transform -1 0 2358 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_722
timestamp 1516325494
transform -1 0 2373 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_721
timestamp 1516325494
transform 1 0 2373 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_745
timestamp 1516325494
transform 1 0 2388 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_613
timestamp 1516325494
transform 1 0 2404 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_197
timestamp 1516325494
transform -1 0 2487 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_737
timestamp 1516325494
transform 1 0 2487 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_719
timestamp 1516325494
transform 1 0 2502 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_613
timestamp 1516325494
transform -1 0 2533 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_732
timestamp 1516325494
transform -1 0 2548 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_232
timestamp 1516325494
transform 1 0 2548 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_232
timestamp 1516325494
transform -1 0 2593 0 1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_616
timestamp 1516325494
transform 1 0 2594 0 1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_616
timestamp 1516325494
transform -1 0 2639 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_200
timestamp 1516325494
transform -1 0 2692 0 1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_717
timestamp 1516325494
transform 1 0 2692 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_796
timestamp 1516325494
transform 1 0 2708 0 1 2620
box 0 0 53 49
use AND2X2  AND2X2_1188
timestamp 1516325494
transform -1 0 2780 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1193
timestamp 1516325494
transform -1 0 2799 0 1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_828
timestamp 1516325494
transform 1 0 2799 0 1 2620
box 0 0 53 49
use OR2X2  OR2X2_998
timestamp 1516325494
transform -1 0 2871 0 1 2620
box 0 0 19 49
use BUFX2  BUFX2_879
timestamp 1516325494
transform 1 0 2871 0 1 2620
box 0 0 15 49
use AND2X2  AND2X2_1266
timestamp 1516325494
transform -1 0 2905 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1264
timestamp 1516325494
transform -1 0 2924 0 1 2620
box 0 0 19 49
use OR2X2  OR2X2_997
timestamp 1516325494
transform -1 0 2943 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1265
timestamp 1516325494
transform -1 0 2962 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1280
timestamp 1516325494
transform -1 0 2981 0 1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_859
timestamp 1516325494
transform 1 0 2981 0 1 2620
box 0 0 15 49
use OAI21X1  OAI21X1_149
timestamp 1516325494
transform -1 0 3015 0 1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_169
timestamp 1516325494
transform -1 0 3034 0 1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_170
timestamp 1516325494
transform -1 0 3053 0 1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_877
timestamp 1516325494
transform -1 0 3068 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_873
timestamp 1516325494
transform 1 0 3069 0 1 2620
box 0 0 15 49
use OAI21X1  OAI21X1_164
timestamp 1516325494
transform -1 0 3103 0 1 2620
box 0 0 19 49
use BUFX2  BUFX2_914
timestamp 1516325494
transform -1 0 3118 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_872
timestamp 1516325494
transform -1 0 3133 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_818
timestamp 1516325494
transform 1 0 3133 0 1 2620
box 0 0 53 49
use OR2X2  OR2X2_1006
timestamp 1516325494
transform -1 0 3205 0 1 2620
box 0 0 19 49
use AND2X2  AND2X2_1273
timestamp 1516325494
transform -1 0 3224 0 1 2620
box 0 0 19 49
use INVX1  INVX1_296
timestamp 1516325494
transform -1 0 3235 0 1 2620
box 0 0 11 49
use INVX1  INVX1_285
timestamp 1516325494
transform -1 0 3247 0 1 2620
box 0 0 11 49
use BUFX2  BUFX2_913
timestamp 1516325494
transform -1 0 3262 0 1 2620
box 0 0 15 49
use NOR2X1  NOR2X1_148
timestamp 1516325494
transform 1 0 3262 0 1 2620
box 0 0 15 49
use OR2X2  OR2X2_992
timestamp 1516325494
transform 1 0 3278 0 1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_825
timestamp 1516325494
transform -1 0 3350 0 1 2620
box 0 0 53 49
use INVX1  INVX1_297
timestamp 1516325494
transform 1 0 3350 0 1 2620
box 0 0 11 49
use NAND2X1  NAND2X1_851
timestamp 1516325494
transform 1 0 3361 0 1 2620
box 0 0 15 49
use NOR2X1  NOR2X1_143
timestamp 1516325494
transform 1 0 3376 0 1 2620
box 0 0 15 49
use OR2X2  OR2X2_980
timestamp 1516325494
transform 1 0 3392 0 1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_833
timestamp 1516325494
transform -1 0 3464 0 1 2620
box 0 0 53 49
use BUFX2  BUFX2_911
timestamp 1516325494
transform 1 0 3464 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_867
timestamp 1516325494
transform -1 0 3494 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_862
timestamp 1516325494
transform -1 0 3509 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_865
timestamp 1516325494
transform -1 0 3524 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_868
timestamp 1516325494
transform -1 0 3540 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_910
timestamp 1516325494
transform -1 0 3555 0 1 2620
box 0 0 15 49
use NOR2X1  NOR2X1_153
timestamp 1516325494
transform 1 0 3555 0 1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_340
timestamp 1516325494
transform -1 0 3623 0 1 2620
box 0 0 53 49
use FILL  FILL_BUFX2_192
timestamp 1516325494
transform 1 0 3623 0 1 2620
box 0 0 8 49
use BUFX2  BUFX2_192
timestamp 1516325494
transform 1 0 3631 0 1 2620
box 0 0 15 49
use AND2X2  AND2X2_2083
timestamp 1516325494
transform -1 0 3665 0 1 2620
box 0 0 19 49
use INVX1  INVX1_312
timestamp 1516325494
transform -1 0 3676 0 1 2620
box 0 0 11 49
use MUX2X1  MUX2X1_275
timestamp 1516325494
transform -1 0 3707 0 1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_819
timestamp 1516325494
transform 1 0 3707 0 1 2620
box 0 0 53 49
use FILL  FILL_BUFX2_188
timestamp 1516325494
transform 1 0 3760 0 1 2620
box 0 0 8 49
use BUFX2  BUFX2_188
timestamp 1516325494
transform 1 0 3768 0 1 2620
box 0 0 15 49
use INVX1  INVX1_170
timestamp 1516325494
transform 1 0 3783 0 1 2620
box 0 0 11 49
use NOR2X1  NOR2X1_160
timestamp 1516325494
transform -1 0 3809 0 1 2620
box 0 0 15 49
use BUFX2  BUFX2_906
timestamp 1516325494
transform -1 0 3825 0 1 2620
box 0 0 15 49
use INVX1  INVX1_318
timestamp 1516325494
transform -1 0 3836 0 1 2620
box 0 0 11 49
use BUFX2  BUFX2_876
timestamp 1516325494
transform -1 0 3851 0 1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_281
timestamp 1516325494
transform -1 0 3866 0 1 2620
box 0 0 15 49
use INVX1  INVX1_179
timestamp 1516325494
transform -1 0 13 0 -1 2620
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_14
timestamp 1516325494
transform 1 0 13 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_110
timestamp 1516325494
transform 1 0 67 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_110
timestamp 1516325494
transform -1 0 112 0 -1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_8
timestamp 1516325494
transform 1 0 112 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_104
timestamp 1516325494
transform 1 0 165 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_104
timestamp 1516325494
transform -1 0 211 0 -1 2620
box 0 0 30 49
use MUX2X1  MUX2X1_78
timestamp 1516325494
transform 1 0 211 0 -1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_110
timestamp 1516325494
transform -1 0 294 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1430
timestamp 1516325494
transform 1 0 295 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1626
timestamp 1516325494
transform 1 0 314 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1429
timestamp 1516325494
transform -1 0 352 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_104
timestamp 1516325494
transform 1 0 352 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1250
timestamp 1516325494
transform 1 0 405 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1488
timestamp 1516325494
transform 1 0 424 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1249
timestamp 1516325494
transform -1 0 462 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_552
timestamp 1516325494
transform 1 0 462 0 -1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_456
timestamp 1516325494
transform 1 0 477 0 -1 2620
box 0 0 53 49
use MUX2X1  MUX2X1_92
timestamp 1516325494
transform 1 0 530 0 -1 2620
box 0 0 30 49
use OR2X2  OR2X2_1849
timestamp 1516325494
transform 1 0 561 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1948
timestamp 1516325494
transform -1 0 599 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1850
timestamp 1516325494
transform -1 0 618 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_92
timestamp 1516325494
transform 1 0 618 0 -1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_572
timestamp 1516325494
transform 1 0 633 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_572
timestamp 1516325494
transform -1 0 678 0 -1 2620
box 0 0 30 49
use FILL  FILL_BUFX2_223
timestamp 1516325494
transform -1 0 686 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_223
timestamp 1516325494
transform -1 0 701 0 -1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_360
timestamp 1516325494
transform 1 0 701 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1817
timestamp 1516325494
transform 1 0 754 0 -1 2620
box 0 0 19 49
use MUX2X1  MUX2X1_539
timestamp 1516325494
transform 1 0 773 0 -1 2620
box 0 0 30 49
use BUFX2  BUFX2_884
timestamp 1516325494
transform -1 0 819 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_1818
timestamp 1516325494
transform 1 0 819 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1923
timestamp 1516325494
transform 1 0 838 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_123
timestamp 1516325494
transform 1 0 857 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_123
timestamp 1516325494
transform -1 0 902 0 -1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_487
timestamp 1516325494
transform 1 0 903 0 -1 2620
box 0 0 53 49
use FILL  FILL_BUFX2_511
timestamp 1516325494
transform 1 0 956 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_511
timestamp 1516325494
transform 1 0 963 0 -1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_551
timestamp 1516325494
transform 1 0 979 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_551
timestamp 1516325494
transform -1 0 1024 0 -1 2620
box 0 0 30 49
use OR2X2  OR2X2_1220
timestamp 1516325494
transform 1 0 1024 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1219
timestamp 1516325494
transform 1 0 1043 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1465
timestamp 1516325494
transform 1 0 1062 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1819
timestamp 1516325494
transform 1 0 1081 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_485
timestamp 1516325494
transform 1 0 1100 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_549
timestamp 1516325494
transform 1 0 1153 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_549
timestamp 1516325494
transform -1 0 1199 0 -1 2620
box 0 0 30 49
use OR2X2  OR2X2_1159
timestamp 1516325494
transform 1 0 1199 0 -1 2620
box 0 0 19 49
use MUX2X1  MUX2X1_69
timestamp 1516325494
transform 1 0 1218 0 -1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_69
timestamp 1516325494
transform -1 0 1263 0 -1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_101
timestamp 1516325494
transform -1 0 1317 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1160
timestamp 1516325494
transform 1 0 1317 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1419
timestamp 1516325494
transform 1 0 1336 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_507
timestamp 1516325494
transform -1 0 1363 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_507
timestamp 1516325494
transform -1 0 1377 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_1217
timestamp 1516325494
transform 1 0 1378 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_31
timestamp 1516325494
transform -1 0 1405 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_31
timestamp 1516325494
transform -1 0 1419 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_1394
timestamp 1516325494
transform 1 0 1419 0 -1 2620
box 0 0 19 49
use MUX2X1  MUX2X1_517
timestamp 1516325494
transform 1 0 1438 0 -1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_517
timestamp 1516325494
transform -1 0 1484 0 -1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_517
timestamp 1516325494
transform -1 0 1537 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1157
timestamp 1516325494
transform 1 0 1537 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1599
timestamp 1516325494
transform -1 0 1575 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1395
timestamp 1516325494
transform -1 0 1594 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_77
timestamp 1516325494
transform 1 0 1594 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_141
timestamp 1516325494
transform 1 0 1647 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_141
timestamp 1516325494
transform 1 0 1663 0 -1 2620
box 0 0 30 49
use MUX2X1  MUX2X1_327
timestamp 1516325494
transform 1 0 1693 0 -1 2620
box 0 0 30 49
use NAND2X1  NAND2X1_327
timestamp 1516325494
transform -1 0 1738 0 -1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_455
timestamp 1516325494
transform -1 0 1792 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1214
timestamp 1516325494
transform 1 0 1792 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1461
timestamp 1516325494
transform -1 0 1830 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1215
timestamp 1516325494
transform -1 0 1849 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_71
timestamp 1516325494
transform 1 0 1849 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_135
timestamp 1516325494
transform 1 0 1902 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_135
timestamp 1516325494
transform 1 0 1917 0 -1 2620
box 0 0 30 49
use OR2X2  OR2X2_1692
timestamp 1516325494
transform 1 0 1948 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1827
timestamp 1516325494
transform -1 0 1986 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1693
timestamp 1516325494
transform -1 0 2005 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_517
timestamp 1516325494
transform -1 0 2013 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_517
timestamp 1516325494
transform -1 0 2027 0 -1 2620
box 0 0 15 49
use FILL  FILL_BUFX2_477
timestamp 1516325494
transform 1 0 2027 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_477
timestamp 1516325494
transform 1 0 2035 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_1152
timestamp 1516325494
transform 1 0 2050 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1413
timestamp 1516325494
transform -1 0 2088 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1153
timestamp 1516325494
transform -1 0 2107 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_551
timestamp 1516325494
transform 1 0 2107 0 -1 2620
box 0 0 53 49
use AND2X2  AND2X2_1459
timestamp 1516325494
transform -1 0 2179 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1212
timestamp 1516325494
transform -1 0 2198 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1213
timestamp 1516325494
transform -1 0 2217 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_359
timestamp 1516325494
transform 1 0 2217 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_917
timestamp 1516325494
transform 1 0 2271 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_862
timestamp 1516325494
transform -1 0 2316 0 -1 2620
box 0 0 30 49
use FILL  FILL_BUFX2_485
timestamp 1516325494
transform -1 0 2324 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_485
timestamp 1516325494
transform -1 0 2339 0 -1 2620
box 0 0 15 49
use NAND2X1  NAND2X1_167
timestamp 1516325494
transform 1 0 2339 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_167
timestamp 1516325494
transform 1 0 2354 0 -1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_391
timestamp 1516325494
transform -1 0 2438 0 -1 2620
box 0 0 53 49
use FILL  FILL_BUFX2_422
timestamp 1516325494
transform -1 0 2446 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_422
timestamp 1516325494
transform -1 0 2460 0 -1 2620
box 0 0 15 49
use FILL  FILL_AND2X2_10
timestamp 1516325494
transform -1 0 2469 0 -1 2620
box 0 0 8 49
use AND2X2  AND2X2_10
timestamp 1516325494
transform -1 0 2487 0 -1 2620
box 0 0 19 49
use FILL  FILL_OR2X2_12
timestamp 1516325494
transform 1 0 2487 0 -1 2620
box 0 0 8 49
use OR2X2  OR2X2_12
timestamp 1516325494
transform 1 0 2495 0 -1 2620
box 0 0 19 49
use FILL  FILL_AND2X2_11
timestamp 1516325494
transform -1 0 2522 0 -1 2620
box 0 0 8 49
use AND2X2  AND2X2_11
timestamp 1516325494
transform -1 0 2540 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1398
timestamp 1516325494
transform -1 0 2559 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1135
timestamp 1516325494
transform 1 0 2559 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1399
timestamp 1516325494
transform -1 0 2597 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_727
timestamp 1516325494
transform -1 0 2612 0 -1 2620
box 0 0 15 49
use AND2X2  AND2X2_1467
timestamp 1516325494
transform 1 0 2613 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1468
timestamp 1516325494
transform 1 0 2632 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1225
timestamp 1516325494
transform 1 0 2651 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_168
timestamp 1516325494
transform -1 0 2723 0 -1 2620
box 0 0 53 49
use FILL  FILL_AND2X2_55
timestamp 1516325494
transform 1 0 2723 0 -1 2620
box 0 0 8 49
use AND2X2  AND2X2_55
timestamp 1516325494
transform 1 0 2730 0 -1 2620
box 0 0 19 49
use FILL  FILL_AND2X2_56
timestamp 1516325494
transform 1 0 2749 0 -1 2620
box 0 0 8 49
use AND2X2  AND2X2_56
timestamp 1516325494
transform 1 0 2757 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_804
timestamp 1516325494
transform -1 0 2829 0 -1 2620
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_199
timestamp 1516325494
transform 1 0 2829 0 -1 2620
box 0 0 53 49
use INVX1  INVX1_173
timestamp 1516325494
transform -1 0 2893 0 -1 2620
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_797
timestamp 1516325494
transform 1 0 2894 0 -1 2620
box 0 0 53 49
use AND2X2  AND2X2_1194
timestamp 1516325494
transform -1 0 2966 0 -1 2620
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_820
timestamp 1516325494
transform 1 0 2966 0 -1 2620
box 0 0 53 49
use NAND2X1  NAND2X1_876
timestamp 1516325494
transform -1 0 3034 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_1010
timestamp 1516325494
transform -1 0 3053 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1279
timestamp 1516325494
transform -1 0 3072 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1281
timestamp 1516325494
transform -1 0 3091 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1009
timestamp 1516325494
transform -1 0 3110 0 -1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_150
timestamp 1516325494
transform -1 0 3129 0 -1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_171
timestamp 1516325494
transform -1 0 3148 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_860
timestamp 1516325494
transform 1 0 3148 0 -1 2620
box 0 0 15 49
use OAI21X1  OAI21X1_151
timestamp 1516325494
transform -1 0 3183 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1250
timestamp 1516325494
transform -1 0 3202 0 -1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_129
timestamp 1516325494
transform -1 0 3221 0 -1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_130
timestamp 1516325494
transform 1 0 3221 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_843
timestamp 1516325494
transform 1 0 3240 0 -1 2620
box 0 0 15 49
use OAI21X1  OAI21X1_165
timestamp 1516325494
transform -1 0 3274 0 -1 2620
box 0 0 19 49
use OAI21X1  OAI21X1_163
timestamp 1516325494
transform -1 0 3293 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1274
timestamp 1516325494
transform 1 0 3293 0 -1 2620
box 0 0 19 49
use OR2X2  OR2X2_1005
timestamp 1516325494
transform 1 0 3312 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1275
timestamp 1516325494
transform -1 0 3350 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_86
timestamp 1516325494
transform 1 0 3350 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_86
timestamp 1516325494
transform 1 0 3357 0 -1 2620
box 0 0 15 49
use MUX2X1  MUX2X1_815
timestamp 1516325494
transform 1 0 3373 0 -1 2620
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_812
timestamp 1516325494
transform 1 0 3403 0 -1 2620
box 0 0 53 49
use AND2X2  AND2X2_1236
timestamp 1516325494
transform -1 0 3475 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_84
timestamp 1516325494
transform 1 0 3475 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_84
timestamp 1516325494
transform 1 0 3483 0 -1 2620
box 0 0 15 49
use AND2X2  AND2X2_1257
timestamp 1516325494
transform -1 0 3517 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_254
timestamp 1516325494
transform 1 0 3517 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_254
timestamp 1516325494
transform 1 0 3525 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_991
timestamp 1516325494
transform 1 0 3540 0 -1 2620
box 0 0 19 49
use NAND3X1  NAND3X1_96
timestamp 1516325494
transform 1 0 3559 0 -1 2620
box 0 0 19 49
use FILL  FILL_BUFX2_256
timestamp 1516325494
transform -1 0 3586 0 -1 2620
box 0 0 8 49
use BUFX2  BUFX2_256
timestamp 1516325494
transform -1 0 3600 0 -1 2620
box 0 0 15 49
use OR2X2  OR2X2_979
timestamp 1516325494
transform 1 0 3601 0 -1 2620
box 0 0 19 49
use NAND3X1  NAND3X1_94
timestamp 1516325494
transform 1 0 3620 0 -1 2620
box 0 0 19 49
use NAND2X1  NAND2X1_834
timestamp 1516325494
transform -1 0 3654 0 -1 2620
box 0 0 15 49
use INVX1  INVX1_294
timestamp 1516325494
transform 1 0 3654 0 -1 2620
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_817
timestamp 1516325494
transform 1 0 3665 0 -1 2620
box 0 0 53 49
use OR2X2  OR2X2_1004
timestamp 1516325494
transform -1 0 3737 0 -1 2620
box 0 0 19 49
use AND2X2  AND2X2_1272
timestamp 1516325494
transform -1 0 3756 0 -1 2620
box 0 0 19 49
use INVX1  INVX1_300
timestamp 1516325494
transform 1 0 3756 0 -1 2620
box 0 0 11 49
use BUFX2  BUFX2_864
timestamp 1516325494
transform 1 0 3768 0 -1 2620
box 0 0 15 49
use BUFX2  BUFX2_863
timestamp 1516325494
transform -1 0 3798 0 -1 2620
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_345
timestamp 1516325494
transform 1 0 3798 0 -1 2620
box 0 0 53 49
use NOR2X1  NOR2X1_172
timestamp 1516325494
transform -1 0 3866 0 -1 2620
box 0 0 15 49
use NOR2X1  NOR2X1_103
timestamp 1516325494
transform -1 0 17 0 1 2521
box 0 0 15 49
use INVX1  INVX1_128
timestamp 1516325494
transform 1 0 17 0 1 2521
box 0 0 11 49
use INVX1  INVX1_125
timestamp 1516325494
transform 1 0 29 0 1 2521
box 0 0 11 49
use AND2X2  AND2X2_1112
timestamp 1516325494
transform -1 0 59 0 1 2521
box 0 0 19 49
use OR2X2  OR2X2_907
timestamp 1516325494
transform -1 0 78 0 1 2521
box 0 0 19 49
use XOR2X1  XOR2X1_57
timestamp 1516325494
transform -1 0 112 0 1 2521
box 0 0 34 49
use AND2X2  AND2X2_1111
timestamp 1516325494
transform -1 0 131 0 1 2521
box 0 0 19 49
use NOR2X1  NOR2X1_98
timestamp 1516325494
transform 1 0 131 0 1 2521
box 0 0 15 49
use INVX1  INVX1_113
timestamp 1516325494
transform 1 0 146 0 1 2521
box 0 0 11 49
use INVX1  INVX1_112
timestamp 1516325494
transform -1 0 169 0 1 2521
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_26
timestamp 1516325494
transform 1 0 169 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_122
timestamp 1516325494
transform 1 0 222 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_122
timestamp 1516325494
transform -1 0 268 0 1 2521
box 0 0 30 49
use OR2X2  OR2X2_1428
timestamp 1516325494
transform 1 0 268 0 1 2521
box 0 0 19 49
use OR2X2  OR2X2_1248
timestamp 1516325494
transform 1 0 287 0 1 2521
box 0 0 19 49
use XOR2X1  XOR2X1_53
timestamp 1516325494
transform -1 0 340 0 1 2521
box 0 0 34 49
use OR2X2  OR2X2_1427
timestamp 1516325494
transform 1 0 340 0 1 2521
box 0 0 19 49
use OR2X2  OR2X2_1247
timestamp 1516325494
transform 1 0 359 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1486
timestamp 1516325494
transform 1 0 378 0 1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_34
timestamp 1516325494
transform 1 0 397 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_34
timestamp 1516325494
transform 1 0 405 0 1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_72
timestamp 1516325494
transform 1 0 420 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_72
timestamp 1516325494
transform -1 0 465 0 1 2521
box 0 0 30 49
use MUX2X1  MUX2X1_90
timestamp 1516325494
transform 1 0 466 0 1 2521
box 0 0 30 49
use BUFX2  BUFX2_895
timestamp 1516325494
transform 1 0 496 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_122
timestamp 1516325494
transform -1 0 564 0 1 2521
box 0 0 53 49
use FILL  FILL_BUFX2_453
timestamp 1516325494
transform 1 0 564 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_453
timestamp 1516325494
transform 1 0 572 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_328
timestamp 1516325494
transform -1 0 617 0 1 2521
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_114
timestamp 1516325494
transform 1 0 618 0 1 2521
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_506
timestamp 1516325494
transform -1 0 724 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_570
timestamp 1516325494
transform 1 0 724 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_570
timestamp 1516325494
transform -1 0 769 0 1 2521
box 0 0 30 49
use FILL  FILL_BUFX2_471
timestamp 1516325494
transform -1 0 778 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_471
timestamp 1516325494
transform -1 0 792 0 1 2521
box 0 0 15 49
use INVX1  INVX1_174
timestamp 1516325494
transform 1 0 792 0 1 2521
box 0 0 11 49
use FILL  FILL_BUFX2_651
timestamp 1516325494
transform 1 0 804 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_651
timestamp 1516325494
transform 1 0 811 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_348
timestamp 1516325494
transform 1 0 827 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_348
timestamp 1516325494
transform -1 0 872 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_650
timestamp 1516325494
transform -1 0 880 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_650
timestamp 1516325494
transform -1 0 895 0 1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_918
timestamp 1516325494
transform 1 0 895 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_863
timestamp 1516325494
transform 1 0 910 0 1 2521
box 0 0 30 49
use INVX1  INVX1_127
timestamp 1516325494
transform -1 0 13 0 -1 2521
box 0 0 11 49
use AND2X2  AND2X2_1113
timestamp 1516325494
transform 1 0 13 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_908
timestamp 1516325494
transform -1 0 51 0 -1 2521
box 0 0 19 49
use XNOR2X1  XNOR2X1_51
timestamp 1516325494
transform -1 0 85 0 -1 2521
box 0 0 34 49
use INVX1  INVX1_126
timestamp 1516325494
transform 1 0 86 0 -1 2521
box 0 0 11 49
use XOR2X1  XOR2X1_58
timestamp 1516325494
transform 1 0 97 0 -1 2521
box 0 0 34 49
use INVX1  INVX1_123
timestamp 1516325494
transform -1 0 142 0 -1 2521
box 0 0 11 49
use XNOR2X1  XNOR2X1_49
timestamp 1516325494
transform -1 0 177 0 -1 2521
box 0 0 34 49
use NOR2X1  NOR2X1_102
timestamp 1516325494
transform -1 0 192 0 -1 2521
box 0 0 15 49
use INVX1  INVX1_124
timestamp 1516325494
transform -1 0 203 0 -1 2521
box 0 0 11 49
use INVX1  INVX1_122
timestamp 1516325494
transform -1 0 214 0 -1 2521
box 0 0 11 49
use XNOR2X1  XNOR2X1_41
timestamp 1516325494
transform 1 0 215 0 -1 2521
box 0 0 34 49
use INVX1  INVX1_120
timestamp 1516325494
transform -1 0 260 0 -1 2521
box 0 0 11 49
use OR2X2  OR2X2_906
timestamp 1516325494
transform -1 0 279 0 -1 2521
box 0 0 19 49
use XOR2X1  XOR2X1_56
timestamp 1516325494
transform -1 0 313 0 -1 2521
box 0 0 34 49
use INVX1  INVX1_111
timestamp 1516325494
transform 1 0 314 0 -1 2521
box 0 0 11 49
use OR2X2  OR2X2_903
timestamp 1516325494
transform 1 0 325 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1108
timestamp 1516325494
transform 1 0 344 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1624
timestamp 1516325494
transform 1 0 363 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1788
timestamp 1516325494
transform 1 0 382 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1900
timestamp 1516325494
transform 1 0 401 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1787
timestamp 1516325494
transform -1 0 439 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_538
timestamp 1516325494
transform 1 0 439 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_538
timestamp 1516325494
transform -1 0 484 0 -1 2521
box 0 0 30 49
use INVX1  INVX1_196
timestamp 1516325494
transform -1 0 496 0 -1 2521
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_28
timestamp 1516325494
transform 1 0 496 0 -1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_90
timestamp 1516325494
transform -1 0 564 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_124
timestamp 1516325494
transform 1 0 564 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_124
timestamp 1516325494
transform -1 0 610 0 -1 2521
box 0 0 30 49
use OR2X2  OR2X2_1790
timestamp 1516325494
transform 1 0 610 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_251
timestamp 1516325494
transform -1 0 637 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_251
timestamp 1516325494
transform -1 0 652 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_530
timestamp 1516325494
transform 1 0 652 0 -1 2521
box 0 0 53 49
use OR2X2  OR2X2_1550
timestamp 1516325494
transform 1 0 705 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1902
timestamp 1516325494
transform 1 0 724 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1789
timestamp 1516325494
transform -1 0 762 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_328
timestamp 1516325494
transform -1 0 777 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_46
timestamp 1516325494
transform 1 0 777 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_46
timestamp 1516325494
transform 1 0 785 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_82
timestamp 1516325494
transform 1 0 800 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_82
timestamp 1516325494
transform -1 0 845 0 -1 2521
box 0 0 30 49
use OR2X2  OR2X2_1244
timestamp 1516325494
transform -1 0 865 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_56
timestamp 1516325494
transform -1 0 873 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_56
timestamp 1516325494
transform -1 0 887 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_474
timestamp 1516325494
transform 1 0 887 0 -1 2521
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_392
timestamp 1516325494
transform 1 0 941 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_168
timestamp 1516325494
transform 1 0 994 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_168
timestamp 1516325494
transform 1 0 1009 0 1 2521
box 0 0 30 49
use MUX2X1  MUX2X1_882
timestamp 1516325494
transform 1 0 1039 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_937
timestamp 1516325494
transform -1 0 1085 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_379
timestamp 1516325494
transform -1 0 1138 0 1 2521
box 0 0 53 49
use OR2X2  OR2X2_1812
timestamp 1516325494
transform 1 0 1138 0 1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_123
timestamp 1516325494
transform 1 0 1157 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_91
timestamp 1516325494
transform 1 0 1210 0 1 2521
box 0 0 15 49
use OR2X2  OR2X2_1784
timestamp 1516325494
transform -1 0 960 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_346
timestamp 1516325494
transform 1 0 960 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_346
timestamp 1516325494
transform -1 0 1005 0 -1 2521
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_476
timestamp 1516325494
transform -1 0 1058 0 -1 2521
box 0 0 53 49
use OR2X2  OR2X2_1844
timestamp 1516325494
transform 1 0 1058 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1242
timestamp 1516325494
transform 1 0 1077 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1482
timestamp 1516325494
transform -1 0 1115 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1243
timestamp 1516325494
transform 1 0 1115 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_11
timestamp 1516325494
transform 1 0 1134 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_11
timestamp 1516325494
transform 1 0 1142 0 -1 2521
box 0 0 15 49
use BUFX2  BUFX2_892
timestamp 1516325494
transform -1 0 1172 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_402
timestamp 1516325494
transform 1 0 1172 0 -1 2521
box 0 0 53 49
use MUX2X1  MUX2X1_91
timestamp 1516325494
transform -1 0 1256 0 1 2521
box 0 0 30 49
use OR2X2  OR2X2_1820
timestamp 1516325494
transform 1 0 1256 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1925
timestamp 1516325494
transform 1 0 1275 0 1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_726
timestamp 1516325494
transform 1 0 1294 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_726
timestamp 1516325494
transform 1 0 1302 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_207
timestamp 1516325494
transform 1 0 1317 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_207
timestamp 1516325494
transform 1 0 1324 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_451
timestamp 1516325494
transform -1 0 1348 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_451
timestamp 1516325494
transform -1 0 1362 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_567
timestamp 1516325494
transform 1 0 1362 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_567
timestamp 1516325494
transform -1 0 1408 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_503
timestamp 1516325494
transform -1 0 1461 0 1 2521
box 0 0 53 49
use OR2X2  OR2X2_1699
timestamp 1516325494
transform 1 0 1461 0 1 2521
box 0 0 19 49
use MUX2X1  MUX2X1_103
timestamp 1516325494
transform 1 0 1480 0 1 2521
box 0 0 30 49
use MUX2X1  MUX2X1_187
timestamp 1516325494
transform -1 0 1256 0 -1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_187
timestamp 1516325494
transform -1 0 1271 0 -1 2521
box 0 0 15 49
use OR2X2  OR2X2_1813
timestamp 1516325494
transform 1 0 1271 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1919
timestamp 1516325494
transform 1 0 1290 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_419
timestamp 1516325494
transform 1 0 1309 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_419
timestamp 1516325494
transform 1 0 1317 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_229
timestamp 1516325494
transform -1 0 1340 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_229
timestamp 1516325494
transform -1 0 1355 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_525
timestamp 1516325494
transform 1 0 1355 0 -1 2521
box 0 0 53 49
use MUX2X1  MUX2X1_525
timestamp 1516325494
transform 1 0 1408 0 -1 2521
box 0 0 30 49
use OR2X2  OR2X2_1400
timestamp 1516325494
transform -1 0 1457 0 -1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_109
timestamp 1516325494
transform 1 0 1457 0 -1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_103
timestamp 1516325494
transform -1 0 1526 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_7
timestamp 1516325494
transform -1 0 1579 0 1 2521
box 0 0 53 49
use OR2X2  OR2X2_1218
timestamp 1516325494
transform 1 0 1579 0 1 2521
box 0 0 19 49
use OR2X2  OR2X2_1814
timestamp 1516325494
transform 1 0 1598 0 1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_475
timestamp 1516325494
transform 1 0 1617 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_347
timestamp 1516325494
transform 1 0 1670 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_347
timestamp 1516325494
transform 1 0 1685 0 1 2521
box 0 0 30 49
use FILL  FILL_BUFX2_649
timestamp 1516325494
transform -1 0 1724 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_649
timestamp 1516325494
transform -1 0 1738 0 1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_101
timestamp 1516325494
transform -1 0 1754 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_101
timestamp 1516325494
transform -1 0 1784 0 1 2521
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_5
timestamp 1516325494
transform -1 0 1837 0 1 2521
box 0 0 53 49
use FILL  FILL_BUFX2_342
timestamp 1516325494
transform 1 0 1837 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_342
timestamp 1516325494
transform 1 0 1845 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_554
timestamp 1516325494
transform 1 0 1860 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_554
timestamp 1516325494
transform 1 0 1868 0 1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_25
timestamp 1516325494
transform 1 0 1883 0 1 2521
box 0 0 19 49
use INVX2  INVX2_14
timestamp 1516325494
transform 1 0 1902 0 1 2521
box 0 0 11 49
use NAND2X1  NAND2X1_723
timestamp 1516325494
transform 1 0 1913 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_325
timestamp 1516325494
transform 1 0 1929 0 1 2521
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_453
timestamp 1516325494
transform -1 0 2012 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_325
timestamp 1516325494
transform -1 0 2027 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_677
timestamp 1516325494
transform 1 0 2027 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_677
timestamp 1516325494
transform 1 0 2035 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_577
timestamp 1516325494
transform 1 0 2050 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_577
timestamp 1516325494
transform 1 0 2058 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_552
timestamp 1516325494
transform -1 0 2081 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_552
timestamp 1516325494
transform -1 0 2096 0 1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_44
timestamp 1516325494
transform 1 0 2096 0 1 2521
box 0 0 19 49
use INVX2  INVX2_33
timestamp 1516325494
transform 1 0 2115 0 1 2521
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_679
timestamp 1516325494
transform 1 0 2126 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_295
timestamp 1516325494
transform 1 0 2179 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_295
timestamp 1516325494
transform -1 0 2225 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_455
timestamp 1516325494
transform 1 0 2225 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_455
timestamp 1516325494
transform -1 0 2270 0 1 2521
box 0 0 30 49
use FILL  FILL_BUFX2_648
timestamp 1516325494
transform -1 0 2279 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_648
timestamp 1516325494
transform -1 0 2293 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_365
timestamp 1516325494
transform -1 0 2346 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_77
timestamp 1516325494
transform 1 0 1511 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_77
timestamp 1516325494
transform -1 0 1556 0 -1 2521
box 0 0 30 49
use AND2X2  AND2X2_1463
timestamp 1516325494
transform -1 0 1575 0 -1 2521
box 0 0 19 49
use MUX2X1  MUX2X1_87
timestamp 1516325494
transform 1 0 1575 0 -1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_87
timestamp 1516325494
transform -1 0 1621 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_119
timestamp 1516325494
transform -1 0 1674 0 -1 2521
box 0 0 53 49
use OR2X2  OR2X2_1700
timestamp 1516325494
transform 1 0 1674 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1833
timestamp 1516325494
transform 1 0 1693 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1921
timestamp 1516325494
transform -1 0 1731 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1417
timestamp 1516325494
transform -1 0 1750 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1158
timestamp 1516325494
transform -1 0 1769 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1815
timestamp 1516325494
transform -1 0 1788 0 -1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_91
timestamp 1516325494
transform 1 0 1788 0 -1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_155
timestamp 1516325494
transform 1 0 1841 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_155
timestamp 1516325494
transform -1 0 1886 0 -1 2521
box 0 0 30 49
use FILL  FILL_AND2X2_52
timestamp 1516325494
transform 1 0 1887 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_52
timestamp 1516325494
transform 1 0 1894 0 -1 2521
box 0 0 19 49
use FILL  FILL_OR2X2_49
timestamp 1516325494
transform -1 0 1921 0 -1 2521
box 0 0 8 49
use OR2X2  OR2X2_49
timestamp 1516325494
transform -1 0 1940 0 -1 2521
box 0 0 19 49
use FILL  FILL_AND2X2_51
timestamp 1516325494
transform -1 0 1948 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_51
timestamp 1516325494
transform -1 0 1967 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1462
timestamp 1516325494
transform 1 0 1967 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1460
timestamp 1516325494
transform 1 0 1986 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1216
timestamp 1516325494
transform 1 0 2005 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1415
timestamp 1516325494
transform 1 0 2024 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1154
timestamp 1516325494
transform -1 0 2062 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1414
timestamp 1516325494
transform -1 0 2081 0 -1 2521
box 0 0 19 49
use FILL  FILL_AND2X2_21
timestamp 1516325494
transform -1 0 2089 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_21
timestamp 1516325494
transform -1 0 2107 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1821
timestamp 1516325494
transform -1 0 2126 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1683
timestamp 1516325494
transform -1 0 2145 0 -1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_567
timestamp 1516325494
transform 1 0 2145 0 -1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_471
timestamp 1516325494
transform 1 0 2198 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_471
timestamp 1516325494
transform -1 0 2244 0 -1 2521
box 0 0 30 49
use OR2X2  OR2X2_1204
timestamp 1516325494
transform 1 0 2244 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1453
timestamp 1516325494
transform 1 0 2263 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1203
timestamp 1516325494
transform -1 0 2301 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_450
timestamp 1516325494
transform 1 0 2301 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_450
timestamp 1516325494
transform 1 0 2309 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_343
timestamp 1516325494
transform 1 0 2324 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_343
timestamp 1516325494
transform 1 0 2331 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_868
timestamp 1516325494
transform -1 0 2377 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_923
timestamp 1516325494
transform 1 0 2377 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_344
timestamp 1516325494
transform 1 0 2392 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_344
timestamp 1516325494
transform 1 0 2400 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_676
timestamp 1516325494
transform 1 0 2415 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_676
timestamp 1516325494
transform 1 0 2423 0 1 2521
box 0 0 15 49
use INVX2  INVX2_11
timestamp 1516325494
transform -1 0 2449 0 1 2521
box 0 0 11 49
use OAI21X1  OAI21X1_22
timestamp 1516325494
transform 1 0 2449 0 1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_40
timestamp 1516325494
transform 1 0 2468 0 1 2521
box 0 0 19 49
use INVX2  INVX2_29
timestamp 1516325494
transform 1 0 2487 0 1 2521
box 0 0 11 49
use OAI21X1  OAI21X1_30
timestamp 1516325494
transform 1 0 2499 0 1 2521
box 0 0 19 49
use INVX2  INVX2_19
timestamp 1516325494
transform 1 0 2518 0 1 2521
box 0 0 11 49
use MUX2X1  MUX2X1_293
timestamp 1516325494
transform 1 0 2529 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_293
timestamp 1516325494
transform -1 0 2574 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_677
timestamp 1516325494
transform -1 0 2628 0 1 2521
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_173
timestamp 1516325494
transform -1 0 2681 0 1 2521
box 0 0 53 49
use FILL  FILL_BUFX2_576
timestamp 1516325494
transform 1 0 2681 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_576
timestamp 1516325494
transform 1 0 2689 0 1 2521
box 0 0 15 49
use AND2X2  AND2X2_1582
timestamp 1516325494
transform -1 0 2723 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1583
timestamp 1516325494
transform -1 0 2742 0 1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_621
timestamp 1516325494
transform 1 0 2742 0 1 2521
box 0 0 15 49
use FILL  FILL_OR2X2_54
timestamp 1516325494
transform 1 0 2757 0 1 2521
box 0 0 8 49
use OR2X2  OR2X2_54
timestamp 1516325494
transform 1 0 2765 0 1 2521
box 0 0 19 49
use MUX2X1  MUX2X1_621
timestamp 1516325494
transform -1 0 2814 0 1 2521
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_205
timestamp 1516325494
transform -1 0 2867 0 1 2521
box 0 0 53 49
use MUX2X1  MUX2X1_231
timestamp 1516325494
transform 1 0 2867 0 1 2521
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_167
timestamp 1516325494
transform -1 0 2951 0 1 2521
box 0 0 53 49
use NAND2X1  NAND2X1_615
timestamp 1516325494
transform 1 0 2951 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_615
timestamp 1516325494
transform -1 0 2996 0 1 2521
box 0 0 30 49
use AND2X2  AND2X2_1189
timestamp 1516325494
transform 1 0 2996 0 1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_836
timestamp 1516325494
transform 1 0 3015 0 1 2521
box 0 0 53 49
use OR2X2  OR2X2_986
timestamp 1516325494
transform -1 0 3088 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1249
timestamp 1516325494
transform -1 0 3107 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1251
timestamp 1516325494
transform -1 0 3126 0 1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_103
timestamp 1516325494
transform 1 0 3126 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_103
timestamp 1516325494
transform 1 0 3133 0 1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_821
timestamp 1516325494
transform -1 0 3201 0 1 2521
box 0 0 53 49
use MUX2X1  MUX2X1_823
timestamp 1516325494
transform 1 0 3202 0 1 2521
box 0 0 30 49
use INVX1  INVX1_301
timestamp 1516325494
transform -1 0 3243 0 1 2521
box 0 0 11 49
use OR2X2  OR2X2_985
timestamp 1516325494
transform -1 0 3262 0 1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_131
timestamp 1516325494
transform -1 0 3281 0 1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_842
timestamp 1516325494
transform 1 0 3281 0 1 2521
box 0 0 15 49
use NAND3X1  NAND3X1_84
timestamp 1516325494
transform 1 0 3297 0 1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_784
timestamp 1516325494
transform -1 0 3331 0 1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_820
timestamp 1516325494
transform -1 0 3361 0 1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_783
timestamp 1516325494
transform -1 0 3376 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_857
timestamp 1516325494
transform 1 0 3376 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_857
timestamp 1516325494
transform 1 0 3384 0 1 2521
box 0 0 15 49
use AND2X2  AND2X2_1235
timestamp 1516325494
transform -1 0 3418 0 1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_107
timestamp 1516325494
transform -1 0 3437 0 1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_817
timestamp 1516325494
transform -1 0 3452 0 1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_108
timestamp 1516325494
transform 1 0 3452 0 1 2521
box 0 0 19 49
use OR2X2  OR2X2_975
timestamp 1516325494
transform 1 0 3471 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1246
timestamp 1516325494
transform -1 0 3509 0 1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_122
timestamp 1516325494
transform 1 0 3509 0 1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_838
timestamp 1516325494
transform 1 0 3528 0 1 2521
box 0 0 15 49
use OR2X2  OR2X2_981
timestamp 1516325494
transform 1 0 3544 0 1 2521
box 0 0 19 49
use AND2X2  AND2X2_1247
timestamp 1516325494
transform 1 0 3563 0 1 2521
box 0 0 19 49
use OR2X2  OR2X2_982
timestamp 1516325494
transform 1 0 3582 0 1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_834
timestamp 1516325494
transform -1 0 3654 0 1 2521
box 0 0 53 49
use NAND3X1  NAND3X1_97
timestamp 1516325494
transform -1 0 3673 0 1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_852
timestamp 1516325494
transform -1 0 3688 0 1 2521
box 0 0 15 49
use AND2X2  AND2X2_1244
timestamp 1516325494
transform -1 0 3707 0 1 2521
box 0 0 19 49
use NAND3X1  NAND3X1_95
timestamp 1516325494
transform -1 0 3726 0 1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_106
timestamp 1516325494
transform 1 0 3726 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_106
timestamp 1516325494
transform 1 0 3734 0 1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_87
timestamp 1516325494
transform -1 0 3757 0 1 2521
box 0 0 8 49
use BUFX2  BUFX2_87
timestamp 1516325494
transform -1 0 3771 0 1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_869
timestamp 1516325494
transform 1 0 3772 0 1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_868
timestamp 1516325494
transform 1 0 3787 0 1 2521
box 0 0 15 49
use OR2X2  OR2X2_1003
timestamp 1516325494
transform 1 0 3802 0 1 2521
box 0 0 19 49
use NAND3X1  NAND3X1_98
timestamp 1516325494
transform 1 0 3821 0 1 2521
box 0 0 19 49
use NAND3X1  NAND3X1_99
timestamp 1516325494
transform 1 0 3840 0 1 2521
box 0 0 19 49
use FILL  FILL_52_1
timestamp 1516325494
transform 1 0 3859 0 1 2521
box 0 0 8 49
use OR2X2  OR2X2_1144
timestamp 1516325494
transform -1 0 2366 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1392
timestamp 1516325494
transform -1 0 2385 0 -1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_24
timestamp 1516325494
transform 1 0 2385 0 -1 2521
box 0 0 19 49
use INVX2  INVX2_13
timestamp 1516325494
transform 1 0 2404 0 -1 2521
box 0 0 11 49
use OR2X2  OR2X2_1684
timestamp 1516325494
transform -1 0 2434 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_262
timestamp 1516325494
transform 1 0 2434 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_262
timestamp 1516325494
transform 1 0 2442 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_311
timestamp 1516325494
transform 1 0 2457 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_695
timestamp 1516325494
transform 1 0 2472 0 -1 2521
box 0 0 53 49
use MUX2X1  MUX2X1_311
timestamp 1516325494
transform -1 0 2555 0 -1 2521
box 0 0 30 49
use FILL  FILL_BUFX2_555
timestamp 1516325494
transform -1 0 2564 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_555
timestamp 1516325494
transform -1 0 2578 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_553
timestamp 1516325494
transform -1 0 2586 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_553
timestamp 1516325494
transform -1 0 2601 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_341
timestamp 1516325494
transform -1 0 2609 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_341
timestamp 1516325494
transform -1 0 2624 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_237
timestamp 1516325494
transform 1 0 2624 0 -1 2521
box 0 0 30 49
use NAND2X1  NAND2X1_237
timestamp 1516325494
transform -1 0 2669 0 -1 2521
box 0 0 15 49
use FILL  FILL_AND2X2_130
timestamp 1516325494
transform -1 0 2678 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_130
timestamp 1516325494
transform -1 0 2696 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1375
timestamp 1516325494
transform -1 0 2715 0 -1 2521
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_237
timestamp 1516325494
transform -1 0 2768 0 -1 2521
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_232
timestamp 1516325494
transform -1 0 2821 0 -1 2521
box 0 0 53 49
use FILL  FILL_AND2X2_131
timestamp 1516325494
transform -1 0 2830 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_131
timestamp 1516325494
transform -1 0 2848 0 -1 2521
box 0 0 19 49
use FILL  FILL_AND2X2_41
timestamp 1516325494
transform -1 0 2856 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_41
timestamp 1516325494
transform -1 0 2875 0 -1 2521
box 0 0 19 49
use FILL  FILL_AND2X2_40
timestamp 1516325494
transform -1 0 2883 0 -1 2521
box 0 0 8 49
use AND2X2  AND2X2_40
timestamp 1516325494
transform -1 0 2901 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_231
timestamp 1516325494
transform -1 0 2916 0 -1 2521
box 0 0 15 49
use AND2X2  AND2X2_1445
timestamp 1516325494
transform -1 0 2936 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1444
timestamp 1516325494
transform -1 0 2955 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_421
timestamp 1516325494
transform -1 0 2963 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_421
timestamp 1516325494
transform -1 0 2977 0 -1 2521
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_215
timestamp 1516325494
transform 1 0 2977 0 -1 2521
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_826
timestamp 1516325494
transform 1 0 3031 0 -1 2521
box 0 0 53 49
use OR2X2  OR2X2_994
timestamp 1516325494
transform -1 0 3103 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1258
timestamp 1516325494
transform -1 0 3122 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1260
timestamp 1516325494
transform -1 0 3141 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1284
timestamp 1516325494
transform -1 0 3160 0 -1 2521
box 0 0 19 49
use OR2X2  OR2X2_1013
timestamp 1516325494
transform -1 0 3179 0 -1 2521
box 0 0 19 49
use NOR2X1  NOR2X1_154
timestamp 1516325494
transform -1 0 3194 0 -1 2521
box 0 0 15 49
use OR2X2  OR2X2_993
timestamp 1516325494
transform -1 0 3213 0 -1 2521
box 0 0 19 49
use AND2X2  AND2X2_1259
timestamp 1516325494
transform -1 0 3232 0 -1 2521
box 0 0 19 49
use NOR2X1  NOR2X1_155
timestamp 1516325494
transform -1 0 3247 0 -1 2521
box 0 0 15 49
use MUX2X1  MUX2X1_817
timestamp 1516325494
transform 1 0 3247 0 -1 2521
box 0 0 30 49
use AOI22X1  AOI22X1_15
timestamp 1516325494
transform -1 0 3301 0 -1 2521
box 0 0 23 49
use OAI21X1  OAI21X1_145
timestamp 1516325494
transform -1 0 3319 0 -1 2521
box 0 0 19 49
use AOI22X1  AOI22X1_25
timestamp 1516325494
transform -1 0 3342 0 -1 2521
box 0 0 23 49
use NAND2X1  NAND2X1_819
timestamp 1516325494
transform 1 0 3342 0 -1 2521
box 0 0 15 49
use NAND3X1  NAND3X1_93
timestamp 1516325494
transform 1 0 3357 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_818
timestamp 1516325494
transform -1 0 3391 0 -1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_143
timestamp 1516325494
transform 1 0 3392 0 -1 2521
box 0 0 19 49
use FILL  FILL_BUFX2_711
timestamp 1516325494
transform 1 0 3411 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_711
timestamp 1516325494
transform 1 0 3418 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_820
timestamp 1516325494
transform 1 0 3433 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_821
timestamp 1516325494
transform 1 0 3449 0 -1 2521
box 0 0 15 49
use AOI22X1  AOI22X1_26
timestamp 1516325494
transform 1 0 3464 0 -1 2521
box 0 0 23 49
use NAND2X1  NAND2X1_856
timestamp 1516325494
transform 1 0 3487 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_855
timestamp 1516325494
transform 1 0 3502 0 -1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_144
timestamp 1516325494
transform -1 0 3536 0 -1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_123
timestamp 1516325494
transform 1 0 3536 0 -1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_124
timestamp 1516325494
transform 1 0 3555 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_839
timestamp 1516325494
transform -1 0 3589 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_710
timestamp 1516325494
transform -1 0 3597 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_710
timestamp 1516325494
transform -1 0 3612 0 -1 2521
box 0 0 15 49
use FILL  FILL_BUFX2_856
timestamp 1516325494
transform -1 0 3620 0 -1 2521
box 0 0 8 49
use BUFX2  BUFX2_856
timestamp 1516325494
transform -1 0 3635 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_854
timestamp 1516325494
transform 1 0 3635 0 -1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_142
timestamp 1516325494
transform 1 0 3650 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_853
timestamp 1516325494
transform -1 0 3684 0 -1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_141
timestamp 1516325494
transform -1 0 3703 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_837
timestamp 1516325494
transform 1 0 3703 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_835
timestamp 1516325494
transform 1 0 3718 0 -1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_121
timestamp 1516325494
transform 1 0 3734 0 -1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_120
timestamp 1516325494
transform 1 0 3753 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_836
timestamp 1516325494
transform -1 0 3787 0 -1 2521
box 0 0 15 49
use OAI21X1  OAI21X1_162
timestamp 1516325494
transform 1 0 3787 0 -1 2521
box 0 0 19 49
use OAI21X1  OAI21X1_161
timestamp 1516325494
transform 1 0 3806 0 -1 2521
box 0 0 19 49
use NAND2X1  NAND2X1_870
timestamp 1516325494
transform 1 0 3825 0 -1 2521
box 0 0 15 49
use NAND2X1  NAND2X1_871
timestamp 1516325494
transform 1 0 3840 0 -1 2521
box 0 0 15 49
use BUFX2  BUFX2_869
timestamp 1516325494
transform -1 0 3870 0 -1 2521
box 0 0 15 49
use XOR2X1  XOR2X1_59
timestamp 1516325494
transform -1 0 36 0 1 2422
box 0 0 34 49
use OR2X2  OR2X2_909
timestamp 1516325494
transform 1 0 36 0 1 2422
box 0 0 19 49
use XNOR2X1  XNOR2X1_50
timestamp 1516325494
transform -1 0 89 0 1 2422
box 0 0 34 49
use INVX1  INVX1_100
timestamp 1516325494
transform 1 0 89 0 1 2422
box 0 0 11 49
use AND2X2  AND2X2_1114
timestamp 1516325494
transform 1 0 101 0 1 2422
box 0 0 19 49
use INVX1  INVX1_131
timestamp 1516325494
transform -1 0 131 0 1 2422
box 0 0 11 49
use XNOR2X1  XNOR2X1_40
timestamp 1516325494
transform -1 0 165 0 1 2422
box 0 0 34 49
use XOR2X1  XOR2X1_60
timestamp 1516325494
transform 1 0 165 0 1 2422
box 0 0 34 49
use INVX1  INVX1_134
timestamp 1516325494
transform -1 0 211 0 1 2422
box 0 0 11 49
use NOR2X1  NOR2X1_105
timestamp 1516325494
transform -1 0 226 0 1 2422
box 0 0 15 49
use INVX1  INVX1_133
timestamp 1516325494
transform -1 0 237 0 1 2422
box 0 0 11 49
use XNOR2X1  XNOR2X1_47
timestamp 1516325494
transform -1 0 272 0 1 2422
box 0 0 34 49
use NOR2X1  NOR2X1_101
timestamp 1516325494
transform -1 0 287 0 1 2422
box 0 0 15 49
use INVX1  INVX1_121
timestamp 1516325494
transform -1 0 298 0 1 2422
box 0 0 11 49
use AND2X2  AND2X2_1110
timestamp 1516325494
transform -1 0 317 0 1 2422
box 0 0 19 49
use INVX1  INVX1_119
timestamp 1516325494
transform -1 0 328 0 1 2422
box 0 0 11 49
use XOR2X1  XOR2X1_54
timestamp 1516325494
transform -1 0 363 0 1 2422
box 0 0 34 49
use OR2X2  OR2X2_904
timestamp 1516325494
transform 1 0 363 0 1 2422
box 0 0 19 49
use INVX1  INVX1_114
timestamp 1516325494
transform -1 0 393 0 1 2422
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_538
timestamp 1516325494
transform 1 0 393 0 1 2422
box 0 0 53 49
use AND2X2  AND2X2_1107
timestamp 1516325494
transform -1 0 466 0 1 2422
box 0 0 19 49
use INVX1  INVX1_110
timestamp 1516325494
transform -1 0 477 0 1 2422
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_540
timestamp 1516325494
transform 1 0 477 0 1 2422
box 0 0 53 49
use INVX1  INVX1_189
timestamp 1516325494
transform -1 0 541 0 1 2422
box 0 0 11 49
use NAND2X1  NAND2X1_540
timestamp 1516325494
transform 1 0 542 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_540
timestamp 1516325494
transform -1 0 587 0 1 2422
box 0 0 30 49
use BUFX2  BUFX2_901
timestamp 1516325494
transform -1 0 602 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_114
timestamp 1516325494
transform 1 0 602 0 1 2422
box 0 0 30 49
use FILL  FILL_BUFX2_50
timestamp 1516325494
transform 1 0 633 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_50
timestamp 1516325494
transform 1 0 640 0 1 2422
box 0 0 15 49
use OR2X2  OR2X2_1547
timestamp 1516325494
transform 1 0 656 0 1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_530
timestamp 1516325494
transform 1 0 675 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_530
timestamp 1516325494
transform -1 0 720 0 1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_466
timestamp 1516325494
transform 1 0 720 0 1 2422
box 0 0 53 49
use MUX2X1  MUX2X1_338
timestamp 1516325494
transform -1 0 803 0 1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_338
timestamp 1516325494
transform -1 0 819 0 1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_476
timestamp 1516325494
transform 1 0 819 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_476
timestamp 1516325494
transform 1 0 827 0 1 2422
box 0 0 15 49
use AND2X2  AND2X2_1484
timestamp 1516325494
transform -1 0 861 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1245
timestamp 1516325494
transform -1 0 880 0 1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_72
timestamp 1516325494
transform 1 0 880 0 1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_136
timestamp 1516325494
transform 1 0 933 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_136
timestamp 1516325494
transform 1 0 948 0 1 2422
box 0 0 30 49
use OR2X2  OR2X2_1544
timestamp 1516325494
transform 1 0 979 0 1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_156
timestamp 1516325494
transform -1 0 1013 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_156
timestamp 1516325494
transform 1 0 1013 0 1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_92
timestamp 1516325494
transform -1 0 1096 0 1 2422
box 0 0 53 49
use OR2X2  OR2X2_1845
timestamp 1516325494
transform 1 0 1096 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1543
timestamp 1516325494
transform -1 0 1134 0 1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_827
timestamp 1516325494
transform 1 0 1134 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_827
timestamp 1516325494
transform 1 0 1142 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_873
timestamp 1516325494
transform -1 0 1187 0 1 2422
box 0 0 30 49
use XOR2X1  XOR2X1_49
timestamp 1516325494
transform -1 0 36 0 -1 2422
box 0 0 34 49
use OR2X2  OR2X2_899
timestamp 1516325494
transform 1 0 36 0 -1 2422
box 0 0 19 49
use INVX1  INVX1_99
timestamp 1516325494
transform -1 0 66 0 -1 2422
box 0 0 11 49
use XNOR2X1  XNOR2X1_33
timestamp 1516325494
transform 1 0 67 0 -1 2422
box 0 0 34 49
use NOR2X1  NOR2X1_94
timestamp 1516325494
transform 1 0 101 0 -1 2422
box 0 0 15 49
use INVX1  INVX1_101
timestamp 1516325494
transform 1 0 116 0 -1 2422
box 0 0 11 49
use AND2X2  AND2X2_1104
timestamp 1516325494
transform 1 0 127 0 -1 2422
box 0 0 19 49
use INVX1  INVX1_129
timestamp 1516325494
transform -1 0 157 0 -1 2422
box 0 0 11 49
use NOR2X1  NOR2X1_104
timestamp 1516325494
transform -1 0 173 0 -1 2422
box 0 0 15 49
use XNOR2X1  XNOR2X1_53
timestamp 1516325494
transform 1 0 173 0 -1 2422
box 0 0 34 49
use INVX1  INVX1_130
timestamp 1516325494
transform 1 0 207 0 -1 2422
box 0 0 11 49
use AND2X2  AND2X2_1115
timestamp 1516325494
transform -1 0 238 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_910
timestamp 1516325494
transform -1 0 257 0 -1 2422
box 0 0 19 49
use INVX1  INVX1_132
timestamp 1516325494
transform -1 0 268 0 -1 2422
box 0 0 11 49
use XNOR2X1  XNOR2X1_55
timestamp 1516325494
transform 1 0 268 0 -1 2422
box 0 0 34 49
use XNOR2X1  XNOR2X1_46
timestamp 1516325494
transform 1 0 302 0 -1 2422
box 0 0 34 49
use OR2X2  OR2X2_905
timestamp 1516325494
transform -1 0 355 0 -1 2422
box 0 0 19 49
use XOR2X1  XOR2X1_55
timestamp 1516325494
transform -1 0 389 0 -1 2422
box 0 0 34 49
use AND2X2  AND2X2_1109
timestamp 1516325494
transform 1 0 390 0 -1 2422
box 0 0 19 49
use INVX1  INVX1_116
timestamp 1516325494
transform 1 0 409 0 -1 2422
box 0 0 11 49
use INVX1  INVX1_192
timestamp 1516325494
transform -1 0 431 0 -1 2422
box 0 0 11 49
use XNOR2X1  XNOR2X1_38
timestamp 1516325494
transform -1 0 465 0 -1 2422
box 0 0 34 49
use NOR2X1  NOR2X1_97
timestamp 1516325494
transform 1 0 466 0 -1 2422
box 0 0 15 49
use INVX1  INVX1_109
timestamp 1516325494
transform -1 0 492 0 -1 2422
box 0 0 11 49
use XNOR2X1  XNOR2X1_39
timestamp 1516325494
transform 1 0 492 0 -1 2422
box 0 0 34 49
use INVX1  INVX1_193
timestamp 1516325494
transform -1 0 537 0 -1 2422
box 0 0 11 49
use OR2X2  OR2X2_1847
timestamp 1516325494
transform 1 0 538 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1848
timestamp 1516325494
transform 1 0 557 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1946
timestamp 1516325494
transform 1 0 576 0 -1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_222
timestamp 1516325494
transform 1 0 595 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_222
timestamp 1516325494
transform 1 0 602 0 -1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_18
timestamp 1516325494
transform -1 0 671 0 -1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_114
timestamp 1516325494
transform -1 0 686 0 -1 2422
box 0 0 15 49
use OR2X2  OR2X2_1548
timestamp 1516325494
transform 1 0 686 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1716
timestamp 1516325494
transform -1 0 724 0 -1 2422
box 0 0 19 49
use INVX1  INVX1_184
timestamp 1516325494
transform -1 0 735 0 -1 2422
box 0 0 11 49
use AND2X2  AND2X2_1718
timestamp 1516325494
transform 1 0 735 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1549
timestamp 1516325494
transform -1 0 773 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_562
timestamp 1516325494
transform 1 0 773 0 -1 2422
box 0 0 15 49
use INVX1  INVX1_178
timestamp 1516325494
transform 1 0 789 0 -1 2422
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_498
timestamp 1516325494
transform 1 0 800 0 -1 2422
box 0 0 53 49
use MUX2X1  MUX2X1_562
timestamp 1516325494
transform -1 0 883 0 -1 2422
box 0 0 30 49
use FILL  FILL_OR2X2_63
timestamp 1516325494
transform -1 0 892 0 -1 2422
box 0 0 8 49
use OR2X2  OR2X2_63
timestamp 1516325494
transform -1 0 910 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_67
timestamp 1516325494
transform -1 0 918 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_67
timestamp 1516325494
transform -1 0 937 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_66
timestamp 1516325494
transform -1 0 945 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_66
timestamp 1516325494
transform -1 0 963 0 -1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_172
timestamp 1516325494
transform -1 0 971 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_172
timestamp 1516325494
transform -1 0 986 0 -1 2422
box 0 0 15 49
use INVX1  INVX1_186
timestamp 1516325494
transform 1 0 986 0 -1 2422
box 0 0 11 49
use FILL  FILL_AND2X2_217
timestamp 1516325494
transform 1 0 998 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_217
timestamp 1516325494
transform 1 0 1005 0 -1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_203
timestamp 1516325494
transform -1 0 1032 0 -1 2422
box 0 0 8 49
use OR2X2  OR2X2_203
timestamp 1516325494
transform -1 0 1051 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_216
timestamp 1516325494
transform -1 0 1059 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_216
timestamp 1516325494
transform -1 0 1077 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1944
timestamp 1516325494
transform -1 0 1096 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1712
timestamp 1516325494
transform -1 0 1115 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1542
timestamp 1516325494
transform -1 0 1134 0 -1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_370
timestamp 1516325494
transform 1 0 1134 0 -1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_178
timestamp 1516325494
transform 1 0 1188 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_178
timestamp 1516325494
transform 1 0 1203 0 1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_411
timestamp 1516325494
transform -1 0 1286 0 1 2422
box 0 0 53 49
use FILL  FILL_BUFX2_431
timestamp 1516325494
transform 1 0 1286 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_431
timestamp 1516325494
transform 1 0 1294 0 1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_214
timestamp 1516325494
transform -1 0 1317 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_214
timestamp 1516325494
transform -1 0 1332 0 1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_493
timestamp 1516325494
transform 1 0 1332 0 1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_557
timestamp 1516325494
transform 1 0 1385 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_557
timestamp 1516325494
transform -1 0 1430 0 1 2422
box 0 0 30 49
use MUX2X1  MUX2X1_830
timestamp 1516325494
transform 1 0 1431 0 1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_885
timestamp 1516325494
transform -1 0 1476 0 1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_615
timestamp 1516325494
transform -1 0 1529 0 1 2422
box 0 0 53 49
use AND2X2  AND2X2_1924
timestamp 1516325494
transform 1 0 1530 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1821
timestamp 1516325494
transform -1 0 1568 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_1926
timestamp 1516325494
transform -1 0 1587 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_354
timestamp 1516325494
transform -1 0 1606 0 1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_54
timestamp 1516325494
transform 1 0 1606 0 1 2422
box 0 0 8 49
use AND2X2  AND2X2_54
timestamp 1516325494
transform 1 0 1613 0 1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_53
timestamp 1516325494
transform 1 0 1632 0 1 2422
box 0 0 8 49
use AND2X2  AND2X2_53
timestamp 1516325494
transform 1 0 1640 0 1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_50
timestamp 1516325494
transform 1 0 1659 0 1 2422
box 0 0 8 49
use OR2X2  OR2X2_50
timestamp 1516325494
transform 1 0 1666 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_293
timestamp 1516325494
transform 1 0 1685 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_294
timestamp 1516325494
transform -1 0 1723 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_1834
timestamp 1516325494
transform 1 0 1723 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_1832
timestamp 1516325494
transform 1 0 1742 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1701
timestamp 1516325494
transform 1 0 1761 0 1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_23
timestamp 1516325494
transform 1 0 1780 0 1 2422
box 0 0 8 49
use AND2X2  AND2X2_23
timestamp 1516325494
transform 1 0 1788 0 1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_51
timestamp 1516325494
transform -1 0 1815 0 1 2422
box 0 0 8 49
use OR2X2  OR2X2_51
timestamp 1516325494
transform -1 0 1834 0 1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_21
timestamp 1516325494
transform -1 0 1842 0 1 2422
box 0 0 8 49
use OR2X2  OR2X2_21
timestamp 1516325494
transform -1 0 1860 0 1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_22
timestamp 1516325494
transform -1 0 1868 0 1 2422
box 0 0 8 49
use AND2X2  AND2X2_22
timestamp 1516325494
transform -1 0 1887 0 1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_203
timestamp 1516325494
transform 1 0 1887 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_203
timestamp 1516325494
transform 1 0 1894 0 1 2422
box 0 0 15 49
use AND2X2  AND2X2_1416
timestamp 1516325494
transform 1 0 1910 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1156
timestamp 1516325494
transform 1 0 1929 0 1 2422
box 0 0 19 49
use INVX1  INVX1_139
timestamp 1516325494
transform 1 0 1948 0 1 2422
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_39
timestamp 1516325494
transform -1 0 2012 0 1 2422
box 0 0 53 49
use OR2X2  OR2X2_1155
timestamp 1516325494
transform -1 0 2031 0 1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_55
timestamp 1516325494
transform 1 0 2031 0 1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_133
timestamp 1516325494
transform 1 0 2084 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_133
timestamp 1516325494
transform 1 0 2100 0 1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_69
timestamp 1516325494
transform -1 0 2183 0 1 2422
box 0 0 53 49
use FILL  FILL_BUFX2_461
timestamp 1516325494
transform -1 0 2191 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_461
timestamp 1516325494
transform -1 0 2206 0 1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_164
timestamp 1516325494
transform 1 0 2206 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_164
timestamp 1516325494
transform 1 0 2214 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_453
timestamp 1516325494
transform -1 0 2259 0 1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_557
timestamp 1516325494
transform 1 0 2259 0 1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_461
timestamp 1516325494
transform 1 0 2312 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_461
timestamp 1516325494
transform -1 0 2358 0 1 2422
box 0 0 30 49
use AND2X2  AND2X2_1597
timestamp 1516325494
transform -1 0 2377 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1393
timestamp 1516325494
transform -1 0 2396 0 1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_397
timestamp 1516325494
transform 1 0 2396 0 1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_173
timestamp 1516325494
transform 1 0 2449 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_173
timestamp 1516325494
transform -1 0 2494 0 1 2422
box 0 0 30 49
use OAI21X1  OAI21X1_35
timestamp 1516325494
transform 1 0 2495 0 1 2422
box 0 0 19 49
use INVX2  INVX2_24
timestamp 1516325494
transform 1 0 2514 0 1 2422
box 0 0 11 49
use FILL  FILL_BUFX2_583
timestamp 1516325494
transform 1 0 2525 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_583
timestamp 1516325494
transform 1 0 2533 0 1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_264
timestamp 1516325494
transform -1 0 2556 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_264
timestamp 1516325494
transform -1 0 2571 0 1 2422
box 0 0 15 49
use NAND2X1  NAND2X1_720
timestamp 1516325494
transform 1 0 2571 0 1 2422
box 0 0 15 49
use FILL  FILL_OR2X2_125
timestamp 1516325494
transform 1 0 2586 0 1 2422
box 0 0 8 49
use OR2X2  OR2X2_125
timestamp 1516325494
transform 1 0 2594 0 1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_132
timestamp 1516325494
transform -1 0 2621 0 1 2422
box 0 0 8 49
use AND2X2  AND2X2_132
timestamp 1516325494
transform -1 0 2639 0 1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_124
timestamp 1516325494
transform -1 0 2647 0 1 2422
box 0 0 8 49
use OR2X2  OR2X2_124
timestamp 1516325494
transform -1 0 2666 0 1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_230
timestamp 1516325494
transform 1 0 2666 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_230
timestamp 1516325494
transform 1 0 2673 0 1 2422
box 0 0 15 49
use NAND2X1  NAND2X1_205
timestamp 1516325494
transform 1 0 2689 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_205
timestamp 1516325494
transform -1 0 2734 0 1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_200
timestamp 1516325494
transform -1 0 2749 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_200
timestamp 1516325494
transform -1 0 2779 0 1 2422
box 0 0 30 49
use FILL  FILL_OR2X2_40
timestamp 1516325494
transform -1 0 2788 0 1 2422
box 0 0 8 49
use OR2X2  OR2X2_40
timestamp 1516325494
transform -1 0 2806 0 1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_215
timestamp 1516325494
transform 1 0 2806 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_215
timestamp 1516325494
transform -1 0 2852 0 1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_247
timestamp 1516325494
transform -1 0 2905 0 1 2422
box 0 0 53 49
use OR2X2  OR2X2_1195
timestamp 1516325494
transform -1 0 2924 0 1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_631
timestamp 1516325494
transform 1 0 2924 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_631
timestamp 1516325494
transform -1 0 2969 0 1 2422
box 0 0 30 49
use MUX2X1  MUX2X1_247
timestamp 1516325494
transform 1 0 2970 0 1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_247
timestamp 1516325494
transform -1 0 3015 0 1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_183
timestamp 1516325494
transform -1 0 3068 0 1 2422
box 0 0 53 49
use FILL  FILL_BUFX2_216
timestamp 1516325494
transform 1 0 3069 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_216
timestamp 1516325494
transform 1 0 3076 0 1 2422
box 0 0 15 49
use AND2X2  AND2X2_1186
timestamp 1516325494
transform 1 0 3091 0 1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_794
timestamp 1516325494
transform 1 0 3110 0 1 2422
box 0 0 53 49
use OR2X2  OR2X2_1012
timestamp 1516325494
transform -1 0 3183 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_1283
timestamp 1516325494
transform -1 0 3202 0 1 2422
box 0 0 19 49
use OR2X2  OR2X2_1011
timestamp 1516325494
transform -1 0 3221 0 1 2422
box 0 0 19 49
use AND2X2  AND2X2_1282
timestamp 1516325494
transform -1 0 3240 0 1 2422
box 0 0 19 49
use OAI21X1  OAI21X1_173
timestamp 1516325494
transform -1 0 3259 0 1 2422
box 0 0 19 49
use AOI21X1  AOI21X1_66
timestamp 1516325494
transform -1 0 3278 0 1 2422
box 0 0 19 49
use OAI21X1  OAI21X1_172
timestamp 1516325494
transform 1 0 3278 0 1 2422
box 0 0 19 49
use NOR2X1  NOR2X1_156
timestamp 1516325494
transform -1 0 3312 0 1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_818
timestamp 1516325494
transform -1 0 3342 0 1 2422
box 0 0 30 49
use MUX2X1  MUX2X1_821
timestamp 1516325494
transform -1 0 3372 0 1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_928
timestamp 1516325494
transform 1 0 1188 0 -1 2422
box 0 0 15 49
use OR2X2  OR2X2_1843
timestamp 1516325494
transform -1 0 1222 0 -1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_412
timestamp 1516325494
transform 1 0 1222 0 -1 2422
box 0 0 53 49
use NAND2X1  NAND2X1_188
timestamp 1516325494
transform 1 0 1275 0 -1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_188
timestamp 1516325494
transform 1 0 1290 0 -1 2422
box 0 0 30 49
use FILL  FILL_BUFX2_828
timestamp 1516325494
transform 1 0 1321 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_828
timestamp 1516325494
transform 1 0 1328 0 -1 2422
box 0 0 15 49
use AND2X2  AND2X2_1920
timestamp 1516325494
transform -1 0 1362 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_351
timestamp 1516325494
transform 1 0 1362 0 -1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_32
timestamp 1516325494
transform -1 0 1389 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_32
timestamp 1516325494
transform -1 0 1404 0 -1 2422
box 0 0 15 49
use OR2X2  OR2X2_1399
timestamp 1516325494
transform 1 0 1404 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_525
timestamp 1516325494
transform 1 0 1423 0 -1 2422
box 0 0 15 49
use AND2X2  AND2X2_1603
timestamp 1516325494
transform 1 0 1438 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1397
timestamp 1516325494
transform 1 0 1457 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1206
timestamp 1516325494
transform 1 0 1476 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_330
timestamp 1516325494
transform -1 0 1514 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_353
timestamp 1516325494
transform -1 0 1533 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1466
timestamp 1516325494
transform 1 0 1533 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1464
timestamp 1516325494
transform 1 0 1552 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1221
timestamp 1516325494
transform 1 0 1571 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_142
timestamp 1516325494
transform 1 0 1590 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_142
timestamp 1516325494
transform 1 0 1598 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1600
timestamp 1516325494
transform -1 0 1636 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1420
timestamp 1516325494
transform 1 0 1636 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_141
timestamp 1516325494
transform -1 0 1663 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_141
timestamp 1516325494
transform -1 0 1682 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_275
timestamp 1516325494
transform -1 0 1701 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_274
timestamp 1516325494
transform 1 0 1701 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_24
timestamp 1516325494
transform 1 0 1720 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_24
timestamp 1516325494
transform 1 0 1727 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1418
timestamp 1516325494
transform 1 0 1746 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1161
timestamp 1516325494
transform 1 0 1765 0 -1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_22
timestamp 1516325494
transform 1 0 1784 0 -1 2422
box 0 0 8 49
use OR2X2  OR2X2_22
timestamp 1516325494
transform 1 0 1792 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1702
timestamp 1516325494
transform 1 0 1811 0 -1 2422
box 0 0 19 49
use FILL  FILL_OR2X2_23
timestamp 1516325494
transform 1 0 1830 0 -1 2422
box 0 0 8 49
use OR2X2  OR2X2_23
timestamp 1516325494
transform 1 0 1837 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1696
timestamp 1516325494
transform -1 0 1875 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1830
timestamp 1516325494
transform -1 0 1894 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_292
timestamp 1516325494
transform 1 0 1894 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_273
timestamp 1516325494
transform -1 0 1932 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_291
timestamp 1516325494
transform -1 0 1951 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1828
timestamp 1516325494
transform -1 0 1970 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1162
timestamp 1516325494
transform 1 0 1970 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1455
timestamp 1516325494
transform -1 0 2008 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1207
timestamp 1516325494
transform -1 0 2027 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1222
timestamp 1516325494
transform 1 0 2027 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1687
timestamp 1516325494
transform -1 0 2065 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_423
timestamp 1516325494
transform 1 0 2065 0 -1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_423
timestamp 1516325494
transform -1 0 2111 0 -1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_439
timestamp 1516325494
transform 1 0 2111 0 -1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_439
timestamp 1516325494
transform -1 0 2156 0 -1 2422
box 0 0 30 49
use FILL  FILL_BUFX2_166
timestamp 1516325494
transform 1 0 2157 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_166
timestamp 1516325494
transform 1 0 2164 0 -1 2422
box 0 0 15 49
use AND2X2  AND2X2_1407
timestamp 1516325494
transform -1 0 2198 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1143
timestamp 1516325494
transform -1 0 2217 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_453
timestamp 1516325494
transform 1 0 2217 0 -1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_549
timestamp 1516325494
transform 1 0 2233 0 -1 2422
box 0 0 53 49
use AND2X2  AND2X2_1591
timestamp 1516325494
transform -1 0 2305 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1383
timestamp 1516325494
transform -1 0 2324 0 -1 2422
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_429
timestamp 1516325494
transform -1 0 2377 0 -1 2422
box 0 0 53 49
use INVX1  INVX1_141
timestamp 1516325494
transform -1 0 2388 0 -1 2422
box 0 0 11 49
use OR2X2  OR2X2_1384
timestamp 1516325494
transform -1 0 2407 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_301
timestamp 1516325494
transform 1 0 2407 0 -1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_685
timestamp 1516325494
transform 1 0 2423 0 -1 2422
box 0 0 53 49
use MUX2X1  MUX2X1_301
timestamp 1516325494
transform -1 0 2506 0 -1 2422
box 0 0 30 49
use FILL  FILL_BUFX2_263
timestamp 1516325494
transform 1 0 2506 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_263
timestamp 1516325494
transform 1 0 2514 0 -1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_589
timestamp 1516325494
transform 1 0 2529 0 -1 2422
box 0 0 30 49
use NAND2X1  NAND2X1_589
timestamp 1516325494
transform -1 0 2574 0 -1 2422
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_269
timestamp 1516325494
transform -1 0 2628 0 -1 2422
box 0 0 53 49
use FILL  FILL_OR2X2_126
timestamp 1516325494
transform -1 0 2636 0 -1 2422
box 0 0 8 49
use OR2X2  OR2X2_126
timestamp 1516325494
transform -1 0 2654 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1376
timestamp 1516325494
transform 1 0 2654 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1584
timestamp 1516325494
transform -1 0 2692 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1377
timestamp 1516325494
transform 1 0 2692 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1227
timestamp 1516325494
transform 1 0 2711 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1226
timestamp 1516325494
transform -1 0 2749 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1469
timestamp 1516325494
transform -1 0 2768 0 -1 2422
box 0 0 19 49
use FILL  FILL_AND2X2_57
timestamp 1516325494
transform 1 0 2768 0 -1 2422
box 0 0 8 49
use AND2X2  AND2X2_57
timestamp 1516325494
transform 1 0 2776 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_282
timestamp 1516325494
transform 1 0 2795 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_265
timestamp 1516325494
transform 1 0 2814 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_266
timestamp 1516325494
transform -1 0 2852 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1814
timestamp 1516325494
transform 1 0 2852 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_264
timestamp 1516325494
transform -1 0 2890 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_280
timestamp 1516325494
transform -1 0 2909 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_281
timestamp 1516325494
transform -1 0 2928 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_599
timestamp 1516325494
transform 1 0 2928 0 -1 2422
box 0 0 15 49
use MUX2X1  MUX2X1_599
timestamp 1516325494
transform -1 0 2973 0 -1 2422
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_279
timestamp 1516325494
transform 1 0 2974 0 -1 2422
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_805
timestamp 1516325494
transform -1 0 3080 0 -1 2422
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_802
timestamp 1516325494
transform 1 0 3080 0 -1 2422
box 0 0 53 49
use INVX1  INVX1_283
timestamp 1516325494
transform 1 0 3133 0 -1 2422
box 0 0 11 49
use OR2X2  OR2X2_1001
timestamp 1516325494
transform -1 0 3164 0 -1 2422
box 0 0 19 49
use NOR2X1  NOR2X1_149
timestamp 1516325494
transform 1 0 3164 0 -1 2422
box 0 0 15 49
use INVX1  INVX1_298
timestamp 1516325494
transform -1 0 3190 0 -1 2422
box 0 0 11 49
use AND2X2  AND2X2_1269
timestamp 1516325494
transform -1 0 3209 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_1000
timestamp 1516325494
transform -1 0 3228 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1268
timestamp 1516325494
transform -1 0 3247 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_999
timestamp 1516325494
transform -1 0 3266 0 -1 2422
box 0 0 19 49
use NOR2X1  NOR2X1_150
timestamp 1516325494
transform -1 0 3281 0 -1 2422
box 0 0 15 49
use AND2X2  AND2X2_1267
timestamp 1516325494
transform -1 0 3300 0 -1 2422
box 0 0 19 49
use AOI21X1  AOI21X1_63
timestamp 1516325494
transform 1 0 3300 0 -1 2422
box 0 0 19 49
use OAI21X1  OAI21X1_153
timestamp 1516325494
transform 1 0 3319 0 -1 2422
box 0 0 19 49
use OAI21X1  OAI21X1_152
timestamp 1516325494
transform -1 0 3357 0 -1 2422
box 0 0 19 49
use NOR2X1  NOR2X1_151
timestamp 1516325494
transform -1 0 3372 0 -1 2422
box 0 0 15 49
use XNOR2X1  XNOR2X1_61
timestamp 1516325494
transform -1 0 3407 0 1 2422
box 0 0 34 49
use AOI22X1  AOI22X1_12
timestamp 1516325494
transform -1 0 3430 0 1 2422
box 0 0 23 49
use AOI21X1  AOI21X1_51
timestamp 1516325494
transform -1 0 3449 0 1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_780
timestamp 1516325494
transform -1 0 3464 0 1 2422
box 0 0 15 49
use NAND2X1  NAND2X1_809
timestamp 1516325494
transform 1 0 3464 0 1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_408
timestamp 1516325494
transform 1 0 3479 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_408
timestamp 1516325494
transform 1 0 3487 0 1 2422
box 0 0 15 49
use AOI22X1  AOI22X1_20
timestamp 1516325494
transform 1 0 3502 0 1 2422
box 0 0 23 49
use INVX1  INVX1_280
timestamp 1516325494
transform 1 0 3525 0 1 2422
box 0 0 11 49
use MUX2X1  MUX2X1_816
timestamp 1516325494
transform 1 0 3536 0 1 2422
box 0 0 30 49
use FILL  FILL_BUFX2_409
timestamp 1516325494
transform -1 0 3574 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_409
timestamp 1516325494
transform -1 0 3589 0 1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_709
timestamp 1516325494
transform -1 0 3597 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_709
timestamp 1516325494
transform -1 0 3612 0 1 2422
box 0 0 15 49
use AND2X2  AND2X2_1245
timestamp 1516325494
transform -1 0 3631 0 1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_235
timestamp 1516325494
transform -1 0 3639 0 1 2422
box 0 0 8 49
use BUFX2  BUFX2_235
timestamp 1516325494
transform -1 0 3654 0 1 2422
box 0 0 15 49
use INVX1  INVX1_281
timestamp 1516325494
transform -1 0 3665 0 1 2422
box 0 0 11 49
use AND2X2  AND2X2_1227
timestamp 1516325494
transform 1 0 3665 0 1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_779
timestamp 1516325494
transform 1 0 3684 0 1 2422
box 0 0 15 49
use NAND3X1  NAND3X1_82
timestamp 1516325494
transform -1 0 3718 0 1 2422
box 0 0 19 49
use AOI22X1  AOI22X1_11
timestamp 1516325494
transform 1 0 3718 0 1 2422
box 0 0 23 49
use NAND2X1  NAND2X1_778
timestamp 1516325494
transform -1 0 3756 0 1 2422
box 0 0 15 49
use OAI21X1  OAI21X1_102
timestamp 1516325494
transform 1 0 3756 0 1 2422
box 0 0 19 49
use OAI21X1  OAI21X1_101
timestamp 1516325494
transform 1 0 3775 0 1 2422
box 0 0 19 49
use AOI22X1  AOI22X1_19
timestamp 1516325494
transform -1 0 3817 0 1 2422
box 0 0 23 49
use NAND2X1  NAND2X1_805
timestamp 1516325494
transform 1 0 3817 0 1 2422
box 0 0 15 49
use NAND2X1  NAND2X1_806
timestamp 1516325494
transform 1 0 3832 0 1 2422
box 0 0 15 49
use INVX1  INVX1_284
timestamp 1516325494
transform 1 0 3848 0 1 2422
box 0 0 11 49
use FILL  FILL_50_1
timestamp 1516325494
transform 1 0 3859 0 1 2422
box 0 0 8 49
use AND2X2  AND2X2_1237
timestamp 1516325494
transform -1 0 3392 0 -1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_491
timestamp 1516325494
transform 1 0 3392 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_491
timestamp 1516325494
transform 1 0 3399 0 -1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_855
timestamp 1516325494
transform 1 0 3414 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_855
timestamp 1516325494
transform 1 0 3422 0 -1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_609
timestamp 1516325494
transform 1 0 3437 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_609
timestamp 1516325494
transform 1 0 3445 0 -1 2422
box 0 0 15 49
use FILL  FILL_BUFX2_492
timestamp 1516325494
transform 1 0 3460 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_492
timestamp 1516325494
transform 1 0 3468 0 -1 2422
box 0 0 15 49
use INVX1  INVX1_290
timestamp 1516325494
transform -1 0 3494 0 -1 2422
box 0 0 11 49
use NAND2X1  NAND2X1_808
timestamp 1516325494
transform 1 0 3494 0 -1 2422
box 0 0 15 49
use NAND3X1  NAND3X1_91
timestamp 1516325494
transform 1 0 3509 0 -1 2422
box 0 0 19 49
use AOI22X1  AOI22X1_13
timestamp 1516325494
transform -1 0 3551 0 -1 2422
box 0 0 23 49
use XNOR2X1  XNOR2X1_60
timestamp 1516325494
transform -1 0 3585 0 -1 2422
box 0 0 34 49
use AND2X2  AND2X2_1232
timestamp 1516325494
transform -1 0 3604 0 -1 2422
box 0 0 19 49
use INVX1  INVX1_293
timestamp 1516325494
transform -1 0 3615 0 -1 2422
box 0 0 11 49
use AND2X2  AND2X2_1230
timestamp 1516325494
transform -1 0 3635 0 -1 2422
box 0 0 19 49
use XOR2X1  XOR2X1_74
timestamp 1516325494
transform 1 0 3635 0 -1 2422
box 0 0 34 49
use OR2X2  OR2X2_972
timestamp 1516325494
transform -1 0 3688 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_971
timestamp 1516325494
transform -1 0 3707 0 -1 2422
box 0 0 19 49
use AND2X2  AND2X2_1228
timestamp 1516325494
transform 1 0 3707 0 -1 2422
box 0 0 19 49
use FILL  FILL_BUFX2_490
timestamp 1516325494
transform -1 0 3734 0 -1 2422
box 0 0 8 49
use BUFX2  BUFX2_490
timestamp 1516325494
transform -1 0 3749 0 -1 2422
box 0 0 15 49
use AND2X2  AND2X2_1226
timestamp 1516325494
transform 1 0 3749 0 -1 2422
box 0 0 19 49
use OR2X2  OR2X2_970
timestamp 1516325494
transform -1 0 3787 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_803
timestamp 1516325494
transform -1 0 3802 0 -1 2422
box 0 0 15 49
use AND2X2  AND2X2_1225
timestamp 1516325494
transform -1 0 3821 0 -1 2422
box 0 0 19 49
use NAND2X1  NAND2X1_804
timestamp 1516325494
transform 1 0 3821 0 -1 2422
box 0 0 15 49
use AOI21X1  AOI21X1_56
timestamp 1516325494
transform 1 0 3836 0 -1 2422
box 0 0 19 49
use FILL  FILL_49_1
timestamp 1516325494
transform -1 0 3863 0 -1 2422
box 0 0 8 49
use FILL  FILL_49_2
timestamp 1516325494
transform -1 0 3871 0 -1 2422
box 0 0 8 49
use OR2X2  OR2X2_769
timestamp 1516325494
transform -1 0 21 0 1 2324
box 0 0 19 49
use XOR2X1  XOR2X1_16
timestamp 1516325494
transform -1 0 55 0 1 2324
box 0 0 34 49
use XNOR2X1  XNOR2X1_32
timestamp 1516325494
transform -1 0 89 0 1 2324
box 0 0 34 49
use NOR2X1  NOR2X1_59
timestamp 1516325494
transform -1 0 104 0 1 2324
box 0 0 15 49
use NAND2X1  NAND2X1_682
timestamp 1516325494
transform 1 0 105 0 1 2324
box 0 0 15 49
use AOI21X1  AOI21X1_17
timestamp 1516325494
transform 1 0 120 0 1 2324
box 0 0 19 49
use XNOR2X1  XNOR2X1_52
timestamp 1516325494
transform -1 0 173 0 1 2324
box 0 0 34 49
use XOR2X1  XOR2X1_22
timestamp 1516325494
transform -1 0 207 0 1 2324
box 0 0 34 49
use AND2X2  AND2X2_984
timestamp 1516325494
transform 1 0 207 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_990
timestamp 1516325494
transform 1 0 226 0 1 2324
box 0 0 19 49
use OAI21X1  OAI21X1_16
timestamp 1516325494
transform 1 0 245 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_826
timestamp 1516325494
transform -1 0 283 0 1 2324
box 0 0 19 49
use NAND2X1  NAND2X1_695
timestamp 1516325494
transform 1 0 283 0 1 2324
box 0 0 15 49
use XNOR2X1  XNOR2X1_54
timestamp 1516325494
transform 1 0 298 0 1 2324
box 0 0 34 49
use NAND2X1  NAND2X1_694
timestamp 1516325494
transform -1 0 348 0 1 2324
box 0 0 15 49
use INVX1  INVX1_117
timestamp 1516325494
transform -1 0 359 0 1 2324
box 0 0 11 49
use XNOR2X1  XNOR2X1_45
timestamp 1516325494
transform -1 0 393 0 1 2324
box 0 0 34 49
use NOR2X1  NOR2X1_100
timestamp 1516325494
transform 1 0 393 0 1 2324
box 0 0 15 49
use NOR2X1  NOR2X1_99
timestamp 1516325494
transform -1 0 424 0 1 2324
box 0 0 15 49
use INVX1  INVX1_115
timestamp 1516325494
transform -1 0 435 0 1 2324
box 0 0 11 49
use XNOR2X1  XNOR2X1_43
timestamp 1516325494
transform 1 0 435 0 1 2324
box 0 0 34 49
use XNOR2X1  XNOR2X1_42
timestamp 1516325494
transform 1 0 469 0 1 2324
box 0 0 34 49
use INVX1  INVX1_108
timestamp 1516325494
transform 1 0 504 0 1 2324
box 0 0 11 49
use OAI21X1  OAI21X1_80
timestamp 1516325494
transform -1 0 534 0 1 2324
box 0 0 19 49
use OAI21X1  OAI21X1_73
timestamp 1516325494
transform -1 0 553 0 1 2324
box 0 0 19 49
use OAI21X1  OAI21X1_76
timestamp 1516325494
transform -1 0 572 0 1 2324
box 0 0 19 49
use INVX1  INVX1_195
timestamp 1516325494
transform 1 0 572 0 1 2324
box 0 0 11 49
use MUX2X1  MUX2X1_769
timestamp 1516325494
transform 1 0 583 0 1 2324
box 0 0 30 49
use INVX1  INVX1_157
timestamp 1516325494
transform -1 0 625 0 1 2324
box 0 0 11 49
use BUFX2  BUFX2_889
timestamp 1516325494
transform -1 0 640 0 1 2324
box 0 0 15 49
use FILL  FILL_AND2X2_68
timestamp 1516325494
transform 1 0 640 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_68
timestamp 1516325494
transform 1 0 648 0 1 2324
box 0 0 19 49
use BUFX2  BUFX2_903
timestamp 1516325494
transform -1 0 682 0 1 2324
box 0 0 15 49
use AND2X2  AND2X2_1717
timestamp 1516325494
transform -1 0 701 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_218
timestamp 1516325494
transform 1 0 701 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_218
timestamp 1516325494
transform 1 0 709 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1551
timestamp 1516325494
transform 1 0 728 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1719
timestamp 1516325494
transform -1 0 766 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_219
timestamp 1516325494
transform 1 0 766 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_219
timestamp 1516325494
transform 1 0 773 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_204
timestamp 1516325494
transform 1 0 792 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_204
timestamp 1516325494
transform 1 0 800 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_69
timestamp 1516325494
transform 1 0 819 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_69
timestamp 1516325494
transform 1 0 827 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_64
timestamp 1516325494
transform 1 0 846 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_64
timestamp 1516325494
transform 1 0 853 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1246
timestamp 1516325494
transform -1 0 891 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1485
timestamp 1516325494
transform -1 0 910 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1483
timestamp 1516325494
transform -1 0 929 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1898
timestamp 1516325494
transform -1 0 948 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1546
timestamp 1516325494
transform -1 0 967 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1715
timestamp 1516325494
transform -1 0 986 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1714
timestamp 1516325494
transform -1 0 1005 0 1 2324
box 0 0 19 49
use FILL  FILL_BUFX2_539
timestamp 1516325494
transform 1 0 1005 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_539
timestamp 1516325494
transform 1 0 1013 0 1 2324
box 0 0 15 49
use FILL  FILL_OR2X2_205
timestamp 1516325494
transform 1 0 1028 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_205
timestamp 1516325494
transform 1 0 1036 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1713
timestamp 1516325494
transform -1 0 1074 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1782
timestamp 1516325494
transform 1 0 1074 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1942
timestamp 1516325494
transform -1 0 1112 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1842
timestamp 1516325494
transform -1 0 1131 0 1 2324
box 0 0 19 49
use NAND2X1  NAND2X1_936
timestamp 1516325494
transform 1 0 1131 0 1 2324
box 0 0 15 49
use MUX2X1  MUX2X1_881
timestamp 1516325494
transform 1 0 1146 0 1 2324
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_378
timestamp 1516325494
transform -1 0 1229 0 1 2324
box 0 0 53 49
use FILL  FILL_BUFX2_144
timestamp 1516325494
transform 1 0 1229 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_144
timestamp 1516325494
transform 1 0 1237 0 1 2324
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_380
timestamp 1516325494
transform 1 0 1252 0 1 2324
box 0 0 53 49
use AND2X2  AND2X2_1922
timestamp 1516325494
transform 1 0 1305 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1816
timestamp 1516325494
transform 1 0 1324 0 1 2324
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_13
timestamp 1516325494
transform 1 0 1343 0 1 2324
box 0 0 53 49
use MUX2X1  MUX2X1_109
timestamp 1516325494
transform 1 0 1397 0 1 2324
box 0 0 30 49
use NAND2X1  NAND2X1_109
timestamp 1516325494
transform -1 0 1442 0 1 2324
box 0 0 15 49
use OR2X2  OR2X2_1398
timestamp 1516325494
transform 1 0 1442 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1601
timestamp 1516325494
transform 1 0 1461 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_329
timestamp 1516325494
transform 1 0 1480 0 1 2324
box 0 0 19 49
use BUFX2  BUFX2_883
timestamp 1516325494
transform -1 0 1514 0 1 2324
box 0 0 15 49
use AND2X2  AND2X2_352
timestamp 1516325494
transform -1 0 1533 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_143
timestamp 1516325494
transform 1 0 1533 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_143
timestamp 1516325494
transform 1 0 1541 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_134
timestamp 1516325494
transform 1 0 1560 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_134
timestamp 1516325494
transform 1 0 1568 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_144
timestamp 1516325494
transform -1 0 1595 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_144
timestamp 1516325494
transform -1 0 1613 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_135
timestamp 1516325494
transform -1 0 1621 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_135
timestamp 1516325494
transform -1 0 1640 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_133
timestamp 1516325494
transform -1 0 1648 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_133
timestamp 1516325494
transform -1 0 1666 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1396
timestamp 1516325494
transform -1 0 1685 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1598
timestamp 1516325494
transform -1 0 1704 0 1 2324
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_571
timestamp 1516325494
transform 1 0 1704 0 1 2324
box 0 0 53 49
use NAND2X1  NAND2X1_475
timestamp 1516325494
transform 1 0 1758 0 1 2324
box 0 0 15 49
use MUX2X1  MUX2X1_475
timestamp 1516325494
transform -1 0 1803 0 1 2324
box 0 0 30 49
use OR2X2  OR2X2_1704
timestamp 1516325494
transform -1 0 1822 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1703
timestamp 1516325494
transform -1 0 1841 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1691
timestamp 1516325494
transform -1 0 1860 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_138
timestamp 1516325494
transform -1 0 1868 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_138
timestamp 1516325494
transform -1 0 1887 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1592
timestamp 1516325494
transform -1 0 1906 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1685
timestamp 1516325494
transform -1 0 1925 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1822
timestamp 1516325494
transform -1 0 1944 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_46
timestamp 1516325494
transform -1 0 1952 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_46
timestamp 1516325494
transform -1 0 1970 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_47
timestamp 1516325494
transform -1 0 1978 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_47
timestamp 1516325494
transform -1 0 1997 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1454
timestamp 1516325494
transform -1 0 2016 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_48
timestamp 1516325494
transform -1 0 2024 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_48
timestamp 1516325494
transform -1 0 2043 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1223
timestamp 1516325494
transform 1 0 2043 0 1 2324
box 0 0 19 49
use FILL  FILL_BUFX2_675
timestamp 1516325494
transform 1 0 2062 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_675
timestamp 1516325494
transform 1 0 2069 0 1 2324
box 0 0 15 49
use AND2X2  AND2X2_1451
timestamp 1516325494
transform -1 0 2103 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1201
timestamp 1516325494
transform -1 0 2122 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1202
timestamp 1516325494
transform -1 0 2141 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1148
timestamp 1516325494
transform -1 0 2160 0 1 2324
box 0 0 19 49
use NAND2X1  NAND2X1_37
timestamp 1516325494
transform 1 0 2160 0 1 2324
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_645
timestamp 1516325494
transform 1 0 2176 0 1 2324
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_423
timestamp 1516325494
transform 1 0 2229 0 1 2324
box 0 0 53 49
use NAND2X1  NAND2X1_391
timestamp 1516325494
transform 1 0 2282 0 1 2324
box 0 0 15 49
use MUX2X1  MUX2X1_391
timestamp 1516325494
transform -1 0 2327 0 1 2324
box 0 0 30 49
use MUX2X1  MUX2X1_397
timestamp 1516325494
transform -1 0 2358 0 1 2324
box 0 0 30 49
use MUX2X1  MUX2X1_493
timestamp 1516325494
transform 1 0 2358 0 1 2324
box 0 0 30 49
use NAND2X1  NAND2X1_493
timestamp 1516325494
transform -1 0 2403 0 1 2324
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_301
timestamp 1516325494
transform 1 0 2404 0 1 2324
box 0 0 53 49
use NAND2X1  NAND2X1_45
timestamp 1516325494
transform 1 0 2457 0 1 2324
box 0 0 15 49
use MUX2X1  MUX2X1_45
timestamp 1516325494
transform -1 0 2502 0 1 2324
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_653
timestamp 1516325494
transform -1 0 2555 0 1 2324
box 0 0 53 49
use FILL  FILL_BUFX2_261
timestamp 1516325494
transform -1 0 2564 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_261
timestamp 1516325494
transform -1 0 2578 0 1 2324
box 0 0 15 49
use FILL  FILL_AND2X2_133
timestamp 1516325494
transform 1 0 2578 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_133
timestamp 1516325494
transform 1 0 2586 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1585
timestamp 1516325494
transform 1 0 2605 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1401
timestamp 1516325494
transform 1 0 2624 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1136
timestamp 1516325494
transform 1 0 2643 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1137
timestamp 1516325494
transform 1 0 2662 0 1 2324
box 0 0 19 49
use MUX2X1  MUX2X1_584
timestamp 1516325494
transform 1 0 2681 0 1 2324
box 0 0 30 49
use NAND2X1  NAND2X1_584
timestamp 1516325494
transform -1 0 2726 0 1 2324
box 0 0 15 49
use AND2X2  AND2X2_1470
timestamp 1516325494
transform 1 0 2727 0 1 2324
box 0 0 19 49
use FILL  FILL_AND2X2_58
timestamp 1516325494
transform 1 0 2746 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_58
timestamp 1516325494
transform 1 0 2753 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_55
timestamp 1516325494
transform 1 0 2772 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_55
timestamp 1516325494
transform 1 0 2780 0 1 2324
box 0 0 19 49
use FILL  FILL_OR2X2_56
timestamp 1516325494
transform 1 0 2799 0 1 2324
box 0 0 8 49
use OR2X2  OR2X2_56
timestamp 1516325494
transform 1 0 2806 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_283
timestamp 1516325494
transform -1 0 2844 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1815
timestamp 1516325494
transform 1 0 2844 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1676
timestamp 1516325494
transform 1 0 2863 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1680
timestamp 1516325494
transform -1 0 2901 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1677
timestamp 1516325494
transform -1 0 2920 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1813
timestamp 1516325494
transform 1 0 2920 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_1675
timestamp 1516325494
transform -1 0 2958 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1812
timestamp 1516325494
transform -1 0 2977 0 1 2324
box 0 0 19 49
use FILL  FILL_BUFX2_184
timestamp 1516325494
transform 1 0 2977 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_184
timestamp 1516325494
transform 1 0 2985 0 1 2324
box 0 0 15 49
use MUX2X1  MUX2X1_360
timestamp 1516325494
transform -1 0 3030 0 1 2324
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_328
timestamp 1516325494
transform -1 0 3084 0 1 2324
box 0 0 53 49
use FILL  FILL_BUFX2_195
timestamp 1516325494
transform -1 0 3092 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_195
timestamp 1516325494
transform -1 0 3106 0 1 2324
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_829
timestamp 1516325494
transform -1 0 3160 0 1 2324
box 0 0 53 49
use OR2X2  OR2X2_988
timestamp 1516325494
transform -1 0 3179 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1253
timestamp 1516325494
transform -1 0 3198 0 1 2324
box 0 0 19 49
use OR2X2  OR2X2_987
timestamp 1516325494
transform -1 0 3217 0 1 2324
box 0 0 19 49
use AOI21X1  AOI21X1_60
timestamp 1516325494
transform -1 0 3236 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1252
timestamp 1516325494
transform -1 0 3255 0 1 2324
box 0 0 19 49
use AOI22X1  AOI22X1_16
timestamp 1516325494
transform 1 0 3255 0 1 2324
box 0 0 23 49
use NAND3X1  NAND3X1_85
timestamp 1516325494
transform 1 0 3278 0 1 2324
box 0 0 19 49
use XOR2X1  XOR2X1_76
timestamp 1516325494
transform -1 0 3331 0 1 2324
box 0 0 34 49
use FILL  FILL_BUFX2_403
timestamp 1516325494
transform 1 0 3331 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_403
timestamp 1516325494
transform 1 0 3338 0 1 2324
box 0 0 15 49
use FILL  FILL_BUFX2_104
timestamp 1516325494
transform 1 0 3354 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_104
timestamp 1516325494
transform 1 0 3361 0 1 2324
box 0 0 15 49
use NAND2X1  NAND2X1_824
timestamp 1516325494
transform 1 0 3376 0 1 2324
box 0 0 15 49
use FILL  FILL_BUFX2_693
timestamp 1516325494
transform -1 0 3400 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_693
timestamp 1516325494
transform -1 0 3414 0 1 2324
box 0 0 15 49
use OAI21X1  OAI21X1_103
timestamp 1516325494
transform 1 0 3414 0 1 2324
box 0 0 19 49
use FILL  FILL_BUFX2_268
timestamp 1516325494
transform 1 0 3433 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_268
timestamp 1516325494
transform 1 0 3441 0 1 2324
box 0 0 15 49
use OAI21X1  OAI21X1_104
timestamp 1516325494
transform 1 0 3456 0 1 2324
box 0 0 19 49
use AOI22X1  AOI22X1_21
timestamp 1516325494
transform -1 0 3498 0 1 2324
box 0 0 23 49
use NAND2X1  NAND2X1_813
timestamp 1516325494
transform -1 0 3513 0 1 2324
box 0 0 15 49
use NAND2X1  NAND2X1_812
timestamp 1516325494
transform -1 0 3528 0 1 2324
box 0 0 15 49
use FILL  FILL_BUFX2_266
timestamp 1516325494
transform 1 0 3528 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_266
timestamp 1516325494
transform 1 0 3536 0 1 2324
box 0 0 15 49
use AND2X2  AND2X2_1234
timestamp 1516325494
transform -1 0 3570 0 1 2324
box 0 0 19 49
use XNOR2X1  XNOR2X1_62
timestamp 1516325494
transform 1 0 3570 0 1 2324
box 0 0 34 49
use DFFPOSX1  DFFPOSX1_835
timestamp 1516325494
transform 1 0 3604 0 1 2324
box 0 0 53 49
use NAND2X1  NAND2X1_840
timestamp 1516325494
transform -1 0 3673 0 1 2324
box 0 0 15 49
use OAI21X1  OAI21X1_166
timestamp 1516325494
transform 1 0 3673 0 1 2324
box 0 0 19 49
use FILL  FILL_BUFX2_404
timestamp 1516325494
transform 1 0 3692 0 1 2324
box 0 0 8 49
use BUFX2  BUFX2_404
timestamp 1516325494
transform 1 0 3699 0 1 2324
box 0 0 15 49
use OAI21X1  OAI21X1_147
timestamp 1516325494
transform 1 0 3715 0 1 2324
box 0 0 19 49
use OAI21X1  OAI21X1_146
timestamp 1516325494
transform 1 0 3734 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1262
timestamp 1516325494
transform 1 0 3753 0 1 2324
box 0 0 19 49
use AND2X2  AND2X2_1277
timestamp 1516325494
transform 1 0 3772 0 1 2324
box 0 0 19 49
use INVX1  INVX1_295
timestamp 1516325494
transform -1 0 3802 0 1 2324
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_809
timestamp 1516325494
transform 1 0 3802 0 1 2324
box 0 0 53 49
use FILL  FILL_48_1
timestamp 1516325494
transform 1 0 3855 0 1 2324
box 0 0 8 49
use FILL  FILL_48_2
timestamp 1516325494
transform 1 0 3863 0 1 2324
box 0 0 8 49
use AND2X2  AND2X2_922
timestamp 1516325494
transform 1 0 2 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_921
timestamp 1516325494
transform -1 0 40 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_770
timestamp 1516325494
transform -1 0 59 0 -1 2323
box 0 0 19 49
use XNOR2X1  XNOR2X1_56
timestamp 1516325494
transform -1 0 93 0 -1 2323
box 0 0 34 49
use OR2X2  OR2X2_866
timestamp 1516325494
transform -1 0 112 0 -1 2323
box 0 0 19 49
use NOR2X1  NOR2X1_80
timestamp 1516325494
transform -1 0 127 0 -1 2323
box 0 0 15 49
use AOI21X1  AOI21X1_26
timestamp 1516325494
transform -1 0 146 0 -1 2323
box 0 0 19 49
use NAND2X1  NAND2X1_704
timestamp 1516325494
transform -1 0 161 0 -1 2323
box 0 0 15 49
use XOR2X1  XOR2X1_61
timestamp 1516325494
transform 1 0 162 0 -1 2323
box 0 0 34 49
use XOR2X1  XOR2X1_62
timestamp 1516325494
transform -1 0 230 0 -1 2323
box 0 0 34 49
use OR2X2  OR2X2_822
timestamp 1516325494
transform 1 0 230 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_15
timestamp 1516325494
transform 1 0 249 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_986
timestamp 1516325494
transform -1 0 287 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_992
timestamp 1516325494
transform 1 0 287 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_827
timestamp 1516325494
transform -1 0 325 0 -1 2323
box 0 0 19 49
use XOR2X1  XOR2X1_23
timestamp 1516325494
transform 1 0 325 0 -1 2323
box 0 0 34 49
use OR2X2  OR2X2_821
timestamp 1516325494
transform -1 0 378 0 -1 2323
box 0 0 19 49
use XNOR2X1  XNOR2X1_44
timestamp 1516325494
transform -1 0 412 0 -1 2323
box 0 0 34 49
use INVX1  INVX1_118
timestamp 1516325494
transform -1 0 423 0 -1 2323
box 0 0 11 49
use OAI21X1  OAI21X1_79
timestamp 1516325494
transform -1 0 443 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_66
timestamp 1516325494
transform -1 0 462 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_83
timestamp 1516325494
transform -1 0 481 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1117
timestamp 1516325494
transform -1 0 500 0 -1 2323
box 0 0 19 49
use INVX1  INVX1_199
timestamp 1516325494
transform -1 0 511 0 -1 2323
box 0 0 11 49
use OR2X2  OR2X2_902
timestamp 1516325494
transform -1 0 530 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_78
timestamp 1516325494
transform -1 0 549 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_82
timestamp 1516325494
transform -1 0 568 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_84
timestamp 1516325494
transform -1 0 587 0 -1 2323
box 0 0 19 49
use MUX2X1  MUX2X1_800
timestamp 1516325494
transform 1 0 587 0 -1 2323
box 0 0 30 49
use INVX1  INVX1_222
timestamp 1516325494
transform -1 0 629 0 -1 2323
box 0 0 11 49
use AND2X2  AND2X2_338
timestamp 1516325494
transform 1 0 629 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1901
timestamp 1516325494
transform 1 0 648 0 -1 2323
box 0 0 19 49
use INVX1  INVX1_197
timestamp 1516325494
transform -1 0 678 0 -1 2323
box 0 0 11 49
use AND2X2  AND2X2_1487
timestamp 1516325494
transform 1 0 678 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_316
timestamp 1516325494
transform 1 0 697 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_339
timestamp 1516325494
transform -1 0 735 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1791
timestamp 1516325494
transform 1 0 735 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1903
timestamp 1516325494
transform -1 0 773 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1489
timestamp 1516325494
transform 1 0 773 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1251
timestamp 1516325494
transform 1 0 792 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1552
timestamp 1516325494
transform 1 0 811 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1792
timestamp 1516325494
transform 1 0 830 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1252
timestamp 1516325494
transform 1 0 849 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_65
timestamp 1516325494
transform 1 0 868 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_65
timestamp 1516325494
transform 1 0 876 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1786
timestamp 1516325494
transform -1 0 914 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1899
timestamp 1516325494
transform -1 0 933 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_337
timestamp 1516325494
transform -1 0 952 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1785
timestamp 1516325494
transform -1 0 971 0 -1 2323
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_90
timestamp 1516325494
transform 1 0 971 0 -1 2323
box 0 0 53 49
use MUX2X1  MUX2X1_154
timestamp 1516325494
transform -1 0 1054 0 -1 2323
box 0 0 30 49
use NAND2X1  NAND2X1_154
timestamp 1516325494
transform 1 0 1055 0 -1 2323
box 0 0 15 49
use AND2X2  AND2X2_367
timestamp 1516325494
transform -1 0 1089 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1943
timestamp 1516325494
transform 1 0 1089 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1846
timestamp 1516325494
transform 1 0 1108 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1945
timestamp 1516325494
transform -1 0 1146 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1896
timestamp 1516325494
transform -1 0 1165 0 -1 2323
box 0 0 19 49
use FILL  FILL_BUFX2_412
timestamp 1516325494
transform -1 0 1173 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_412
timestamp 1516325494
transform -1 0 1187 0 -1 2323
box 0 0 15 49
use OR2X2  OR2X2_1783
timestamp 1516325494
transform -1 0 1207 0 -1 2323
box 0 0 19 49
use NAND2X1  NAND2X1_186
timestamp 1516325494
transform 1 0 1207 0 -1 2323
box 0 0 15 49
use MUX2X1  MUX2X1_186
timestamp 1516325494
transform 1 0 1222 0 -1 2323
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_410
timestamp 1516325494
transform -1 0 1305 0 -1 2323
box 0 0 53 49
use NAND2X1  NAND2X1_938
timestamp 1516325494
transform 1 0 1305 0 -1 2323
box 0 0 15 49
use MUX2X1  MUX2X1_883
timestamp 1516325494
transform -1 0 1351 0 -1 2323
box 0 0 30 49
use FILL  FILL_BUFX2_143
timestamp 1516325494
transform 1 0 1351 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_143
timestamp 1516325494
transform 1 0 1359 0 -1 2323
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_621
timestamp 1516325494
transform -1 0 1427 0 -1 2323
box 0 0 53 49
use NAND2X1  NAND2X1_891
timestamp 1516325494
transform 1 0 1427 0 -1 2323
box 0 0 15 49
use MUX2X1  MUX2X1_836
timestamp 1516325494
transform -1 0 1472 0 -1 2323
box 0 0 30 49
use OR2X2  OR2X2_1822
timestamp 1516325494
transform 1 0 1473 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_331
timestamp 1516325494
transform 1 0 1492 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1604
timestamp 1516325494
transform -1 0 1530 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1602
timestamp 1516325494
transform 1 0 1530 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1401
timestamp 1516325494
transform 1 0 1549 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1402
timestamp 1516325494
transform 1 0 1568 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1403
timestamp 1516325494
transform -1 0 1606 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1391
timestamp 1516325494
transform -1 0 1625 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_277
timestamp 1516325494
transform -1 0 1644 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_276
timestamp 1516325494
transform -1 0 1663 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_130
timestamp 1516325494
transform -1 0 1671 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_130
timestamp 1516325494
transform -1 0 1689 0 -1 2323
box 0 0 19 49
use FILL  FILL_AND2X2_137
timestamp 1516325494
transform -1 0 1697 0 -1 2323
box 0 0 8 49
use AND2X2  AND2X2_137
timestamp 1516325494
transform -1 0 1716 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_272
timestamp 1516325494
transform -1 0 1735 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_271
timestamp 1516325494
transform -1 0 1754 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1385
timestamp 1516325494
transform -1 0 1773 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1590
timestamp 1516325494
transform -1 0 1792 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_52
timestamp 1516325494
transform -1 0 1800 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_52
timestamp 1516325494
transform -1 0 1818 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_48
timestamp 1516325494
transform -1 0 1826 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_48
timestamp 1516325494
transform -1 0 1845 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_270
timestamp 1516325494
transform -1 0 1864 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_287
timestamp 1516325494
transform -1 0 1883 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_288
timestamp 1516325494
transform -1 0 1902 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1820
timestamp 1516325494
transform 1 0 1902 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1452
timestamp 1516325494
transform -1 0 1940 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1205
timestamp 1516325494
transform 1 0 1940 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1211
timestamp 1516325494
transform 1 0 1959 0 -1 2323
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_37
timestamp 1516325494
transform 1 0 1978 0 -1 2323
box 0 0 53 49
use MUX2X1  MUX2X1_421
timestamp 1516325494
transform 1 0 2031 0 -1 2323
box 0 0 30 49
use OR2X2  OR2X2_1147
timestamp 1516325494
transform -1 0 2081 0 -1 2323
box 0 0 19 49
use NAND2X1  NAND2X1_421
timestamp 1516325494
transform 1 0 2081 0 -1 2323
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_583
timestamp 1516325494
transform 1 0 2096 0 -1 2323
box 0 0 53 49
use NAND2X1  NAND2X1_7
timestamp 1516325494
transform 1 0 2149 0 -1 2323
box 0 0 15 49
use MUX2X1  MUX2X1_7
timestamp 1516325494
transform -1 0 2194 0 -1 2323
box 0 0 30 49
use MUX2X1  MUX2X1_37
timestamp 1516325494
transform -1 0 2225 0 -1 2323
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_647
timestamp 1516325494
transform 1 0 2225 0 -1 2323
box 0 0 53 49
use AND2X2  AND2X2_1589
timestamp 1516325494
transform -1 0 2297 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1382
timestamp 1516325494
transform -1 0 2316 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1381
timestamp 1516325494
transform -1 0 2335 0 -1 2323
box 0 0 19 49
use NAND2X1  NAND2X1_397
timestamp 1516325494
transform -1 0 2350 0 -1 2323
box 0 0 15 49
use AND2X2  AND2X2_1595
timestamp 1516325494
transform -1 0 2369 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1388
timestamp 1516325494
transform -1 0 2388 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1389
timestamp 1516325494
transform -1 0 2407 0 -1 2323
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_589
timestamp 1516325494
transform 1 0 2407 0 -1 2323
box 0 0 53 49
use NAND2X1  NAND2X1_13
timestamp 1516325494
transform 1 0 2461 0 -1 2323
box 0 0 15 49
use MUX2X1  MUX2X1_13
timestamp 1516325494
transform -1 0 2506 0 -1 2323
box 0 0 30 49
use FILL  FILL_AND2X2_13
timestamp 1516325494
transform 1 0 2506 0 -1 2323
box 0 0 8 49
use AND2X2  AND2X2_13
timestamp 1516325494
transform 1 0 2514 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_13
timestamp 1516325494
transform 1 0 2533 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_13
timestamp 1516325494
transform 1 0 2540 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_14
timestamp 1516325494
transform 1 0 2559 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_14
timestamp 1516325494
transform 1 0 2567 0 -1 2323
box 0 0 19 49
use FILL  FILL_OR2X2_129
timestamp 1516325494
transform -1 0 2594 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_129
timestamp 1516325494
transform -1 0 2613 0 -1 2323
box 0 0 19 49
use FILL  FILL_AND2X2_12
timestamp 1516325494
transform -1 0 2621 0 -1 2323
box 0 0 8 49
use AND2X2  AND2X2_12
timestamp 1516325494
transform -1 0 2639 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1400
timestamp 1516325494
transform -1 0 2658 0 -1 2323
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_264
timestamp 1516325494
transform -1 0 2711 0 -1 2323
box 0 0 53 49
use OR2X2  OR2X2_1230
timestamp 1516325494
transform -1 0 2730 0 -1 2323
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_263
timestamp 1516325494
transform 1 0 2730 0 -1 2323
box 0 0 53 49
use FILL  FILL_OR2X2_42
timestamp 1516325494
transform 1 0 2784 0 -1 2323
box 0 0 8 49
use OR2X2  OR2X2_42
timestamp 1516325494
transform 1 0 2791 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_269
timestamp 1516325494
transform -1 0 2829 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1224
timestamp 1516325494
transform 1 0 2829 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1196
timestamp 1516325494
transform 1 0 2848 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1197
timestamp 1516325494
transform 1 0 2867 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1200
timestamp 1516325494
transform -1 0 2905 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_1199
timestamp 1516325494
transform -1 0 2924 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1448
timestamp 1516325494
transform -1 0 2943 0 -1 2323
box 0 0 19 49
use FILL  FILL_AND2X2_44
timestamp 1516325494
transform -1 0 2951 0 -1 2323
box 0 0 8 49
use AND2X2  AND2X2_44
timestamp 1516325494
transform -1 0 2970 0 -1 2323
box 0 0 19 49
use FILL  FILL_BUFX2_488
timestamp 1516325494
transform -1 0 2978 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_488
timestamp 1516325494
transform -1 0 2992 0 -1 2323
box 0 0 15 49
use NAND2X1  NAND2X1_360
timestamp 1516325494
transform -1 0 3008 0 -1 2323
box 0 0 15 49
use MUX2X1  MUX2X1_264
timestamp 1516325494
transform 1 0 3008 0 -1 2323
box 0 0 30 49
use NAND2X1  NAND2X1_264
timestamp 1516325494
transform -1 0 3053 0 -1 2323
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_136
timestamp 1516325494
transform -1 0 3106 0 -1 2323
box 0 0 53 49
use AND2X2  AND2X2_1254
timestamp 1516325494
transform -1 0 3126 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_989
timestamp 1516325494
transform 1 0 3126 0 -1 2323
box 0 0 19 49
use NOR2X1  NOR2X1_144
timestamp 1516325494
transform -1 0 3160 0 -1 2323
box 0 0 15 49
use OAI21X1  OAI21X1_133
timestamp 1516325494
transform 1 0 3160 0 -1 2323
box 0 0 19 49
use OAI21X1  OAI21X1_132
timestamp 1516325494
transform -1 0 3198 0 -1 2323
box 0 0 19 49
use NOR2X1  NOR2X1_145
timestamp 1516325494
transform -1 0 3213 0 -1 2323
box 0 0 15 49
use NAND2X1  NAND2X1_823
timestamp 1516325494
transform 1 0 3213 0 -1 2323
box 0 0 15 49
use OAI21X1  OAI21X1_110
timestamp 1516325494
transform 1 0 3228 0 -1 2323
box 0 0 19 49
use AOI22X1  AOI22X1_27
timestamp 1516325494
transform 1 0 3247 0 -1 2323
box 0 0 23 49
use INVX1  INVX1_289
timestamp 1516325494
transform -1 0 3281 0 -1 2323
box 0 0 11 49
use NAND2X1  NAND2X1_785
timestamp 1516325494
transform -1 0 3296 0 -1 2323
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_813
timestamp 1516325494
transform -1 0 3350 0 -1 2323
box 0 0 53 49
use FILL  FILL_BUFX2_694
timestamp 1516325494
transform -1 0 3358 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_694
timestamp 1516325494
transform -1 0 3372 0 -1 2323
box 0 0 15 49
use NAND2X1  NAND2X1_822
timestamp 1516325494
transform 1 0 3373 0 -1 2323
box 0 0 15 49
use FILL  FILL_BUFX2_708
timestamp 1516325494
transform 1 0 3388 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_708
timestamp 1516325494
transform 1 0 3395 0 -1 2323
box 0 0 15 49
use NAND2X1  NAND2X1_810
timestamp 1516325494
transform 1 0 3411 0 -1 2323
box 0 0 15 49
use AOI21X1  AOI21X1_57
timestamp 1516325494
transform -1 0 3445 0 -1 2323
box 0 0 19 49
use NAND2X1  NAND2X1_807
timestamp 1516325494
transform -1 0 3460 0 -1 2323
box 0 0 15 49
use NAND2X1  NAND2X1_811
timestamp 1516325494
transform 1 0 3460 0 -1 2323
box 0 0 15 49
use AND2X2  AND2X2_1231
timestamp 1516325494
transform -1 0 3494 0 -1 2323
box 0 0 19 49
use FILL  FILL_BUFX2_692
timestamp 1516325494
transform -1 0 3502 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_692
timestamp 1516325494
transform -1 0 3517 0 -1 2323
box 0 0 15 49
use INVX1  INVX1_277
timestamp 1516325494
transform 1 0 3517 0 -1 2323
box 0 0 11 49
use FILL  FILL_BUFX2_253
timestamp 1516325494
transform 1 0 3528 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_253
timestamp 1516325494
transform 1 0 3536 0 -1 2323
box 0 0 15 49
use FILL  FILL_BUFX2_255
timestamp 1516325494
transform -1 0 3559 0 -1 2323
box 0 0 8 49
use BUFX2  BUFX2_255
timestamp 1516325494
transform -1 0 3574 0 -1 2323
box 0 0 15 49
use XOR2X1  XOR2X1_75
timestamp 1516325494
transform 1 0 3574 0 -1 2323
box 0 0 34 49
use NAND2X1  NAND2X1_814
timestamp 1516325494
transform -1 0 3623 0 -1 2323
box 0 0 15 49
use OAI21X1  OAI21X1_128
timestamp 1516325494
transform 1 0 3623 0 -1 2323
box 0 0 19 49
use AOI22X1  AOI22X1_22
timestamp 1516325494
transform -1 0 3665 0 -1 2323
box 0 0 23 49
use NAND2X1  NAND2X1_874
timestamp 1516325494
transform 1 0 3665 0 -1 2323
box 0 0 15 49
use OAI21X1  OAI21X1_167
timestamp 1516325494
transform 1 0 3680 0 -1 2323
box 0 0 19 49
use NAND2X1  NAND2X1_857
timestamp 1516325494
transform 1 0 3699 0 -1 2323
box 0 0 15 49
use NAND2X1  NAND2X1_858
timestamp 1516325494
transform 1 0 3715 0 -1 2323
box 0 0 15 49
use OAI21X1  OAI21X1_148
timestamp 1516325494
transform -1 0 3749 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_995
timestamp 1516325494
transform 1 0 3749 0 -1 2323
box 0 0 19 49
use AND2X2  AND2X2_1263
timestamp 1516325494
transform 1 0 3768 0 -1 2323
box 0 0 19 49
use OR2X2  OR2X2_996
timestamp 1516325494
transform 1 0 3787 0 -1 2323
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_827
timestamp 1516325494
transform -1 0 3859 0 -1 2323
box 0 0 53 49
use INVX1  INVX1_287
timestamp 1516325494
transform -1 0 3870 0 -1 2323
box 0 0 11 49
use BUFX2  BUFX2_896
timestamp 1516325494
transform 1 0 2 0 1 2225
box 0 0 15 49
use AND2X2  AND2X2_1103
timestamp 1516325494
transform -1 0 36 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_898
timestamp 1516325494
transform -1 0 55 0 1 2225
box 0 0 19 49
use INVX1  INVX1_98
timestamp 1516325494
transform -1 0 66 0 1 2225
box 0 0 11 49
use AND2X2  AND2X2_1044
timestamp 1516325494
transform -1 0 86 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1045
timestamp 1516325494
transform 1 0 86 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_867
timestamp 1516325494
transform -1 0 124 0 1 2225
box 0 0 19 49
use XOR2X1  XOR2X1_27
timestamp 1516325494
transform -1 0 158 0 1 2225
box 0 0 34 49
use FILL  FILL_BUFX2_789
timestamp 1516325494
transform 1 0 158 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_789
timestamp 1516325494
transform 1 0 165 0 1 2225
box 0 0 15 49
use NAND2X1  NAND2X1_700
timestamp 1516325494
transform -1 0 196 0 1 2225
box 0 0 15 49
use AOI21X1  AOI21X1_25
timestamp 1516325494
transform 1 0 196 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_853
timestamp 1516325494
transform -1 0 234 0 1 2225
box 0 0 19 49
use NOR2X1  NOR2X1_77
timestamp 1516325494
transform -1 0 249 0 1 2225
box 0 0 15 49
use AND2X2  AND2X2_985
timestamp 1516325494
transform 1 0 249 0 1 2225
box 0 0 19 49
use XNOR2X1  XNOR2X1_48
timestamp 1516325494
transform -1 0 302 0 1 2225
box 0 0 34 49
use AND2X2  AND2X2_991
timestamp 1516325494
transform -1 0 321 0 1 2225
box 0 0 19 49
use FILL  FILL_BUFX2_565
timestamp 1516325494
transform 1 0 321 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_565
timestamp 1516325494
transform 1 0 329 0 1 2225
box 0 0 15 49
use INVX1  INVX1_190
timestamp 1516325494
transform -1 0 355 0 1 2225
box 0 0 11 49
use NAND3X1  NAND3X1_59
timestamp 1516325494
transform 1 0 355 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_974
timestamp 1516325494
transform 1 0 374 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_973
timestamp 1516325494
transform -1 0 412 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_812
timestamp 1516325494
transform -1 0 431 0 1 2225
box 0 0 19 49
use OAI21X1  OAI21X1_81
timestamp 1516325494
transform -1 0 450 0 1 2225
box 0 0 19 49
use OAI21X1  OAI21X1_77
timestamp 1516325494
transform -1 0 469 0 1 2225
box 0 0 19 49
use NOR2X1  NOR2X1_69
timestamp 1516325494
transform -1 0 484 0 1 2225
box 0 0 15 49
use NOR2X1  NOR2X1_66
timestamp 1516325494
transform 1 0 485 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_784
timestamp 1516325494
transform 1 0 500 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_784
timestamp 1516325494
transform 1 0 507 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_782
timestamp 1516325494
transform -1 0 531 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_782
timestamp 1516325494
transform -1 0 545 0 1 2225
box 0 0 15 49
use XOR2X1  XOR2X1_52
timestamp 1516325494
transform -1 0 579 0 1 2225
box 0 0 34 49
use FILL  FILL_BUFX2_852
timestamp 1516325494
transform 1 0 580 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_852
timestamp 1516325494
transform 1 0 587 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_741
timestamp 1516325494
transform -1 0 655 0 1 2225
box 0 0 53 49
use FILL  FILL_BUFX2_180
timestamp 1516325494
transform 1 0 656 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_180
timestamp 1516325494
transform 1 0 663 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_759
timestamp 1516325494
transform 1 0 678 0 1 2225
box 0 0 30 49
use MUX2X1  MUX2X1_773
timestamp 1516325494
transform 1 0 709 0 1 2225
box 0 0 30 49
use MUX2X1  MUX2X1_804
timestamp 1516325494
transform -1 0 769 0 1 2225
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_533
timestamp 1516325494
transform 1 0 770 0 1 2225
box 0 0 53 49
use OR2X2  OR2X2_317
timestamp 1516325494
transform 1 0 823 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_533
timestamp 1516325494
transform 1 0 842 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_533
timestamp 1516325494
transform -1 0 887 0 1 2225
box 0 0 30 49
use AND2X2  AND2X2_368
timestamp 1516325494
transform 1 0 887 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1947
timestamp 1516325494
transform 1 0 906 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_315
timestamp 1516325494
transform -1 0 944 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_336
timestamp 1516325494
transform -1 0 963 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1897
timestamp 1516325494
transform -1 0 982 0 1 2225
box 0 0 19 49
use FILL  FILL_BUFX2_500
timestamp 1516325494
transform 1 0 982 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_500
timestamp 1516325494
transform 1 0 990 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_483
timestamp 1516325494
transform 1 0 1005 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_483
timestamp 1516325494
transform 1 0 1013 0 1 2225
box 0 0 15 49
use AND2X2  AND2X2_1949
timestamp 1516325494
transform 1 0 1028 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1851
timestamp 1516325494
transform 1 0 1047 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_343
timestamp 1516325494
transform 1 0 1066 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_366
timestamp 1516325494
transform -1 0 1104 0 1 2225
box 0 0 19 49
use INVX1  INVX1_212
timestamp 1516325494
transform -1 0 1115 0 1 2225
box 0 0 11 49
use OR2X2  OR2X2_1852
timestamp 1516325494
transform 1 0 1115 0 1 2225
box 0 0 19 49
use FILL  FILL_BUFX2_112
timestamp 1516325494
transform 1 0 1134 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_112
timestamp 1516325494
transform 1 0 1142 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_1
timestamp 1516325494
transform 1 0 1157 0 1 2225
box 0 0 53 49
use OR2X2  OR2X2_1037
timestamp 1516325494
transform 1 0 1210 0 1 2225
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_513
timestamp 1516325494
transform 1 0 1229 0 1 2225
box 0 0 53 49
use NAND2X1  NAND2X1_513
timestamp 1516325494
transform 1 0 1283 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_513
timestamp 1516325494
transform -1 0 1328 0 1 2225
box 0 0 30 49
use FILL  FILL_BUFX2_202
timestamp 1516325494
transform -1 0 1336 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_202
timestamp 1516325494
transform -1 0 1351 0 1 2225
box 0 0 15 49
use NAND2X1  NAND2X1_735
timestamp 1516325494
transform -1 0 1366 0 1 2225
box 0 0 15 49
use OAI21X1  OAI21X1_43
timestamp 1516325494
transform 1 0 1366 0 1 2225
box 0 0 19 49
use INVX2  INVX2_32
timestamp 1516325494
transform -1 0 1396 0 1 2225
box 0 0 11 49
use FILL  FILL_BUFX2_499
timestamp 1516325494
transform 1 0 1397 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_499
timestamp 1516325494
transform 1 0 1404 0 1 2225
box 0 0 15 49
use OR2X2  OR2X2_1386
timestamp 1516325494
transform 1 0 1419 0 1 2225
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_469
timestamp 1516325494
transform 1 0 1438 0 1 2225
box 0 0 53 49
use NAND2X1  NAND2X1_733
timestamp 1516325494
transform 1 0 1492 0 1 2225
box 0 0 15 49
use OR2X2  OR2X2_1824
timestamp 1516325494
transform -1 0 1526 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1823
timestamp 1516325494
transform -1 0 1545 0 1 2225
box 0 0 19 49
use FILL  FILL_OR2X2_137
timestamp 1516325494
transform -1 0 1553 0 1 2225
box 0 0 8 49
use OR2X2  OR2X2_137
timestamp 1516325494
transform -1 0 1571 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1404
timestamp 1516325494
transform -1 0 1590 0 1 2225
box 0 0 19 49
use FILL  FILL_OR2X2_136
timestamp 1516325494
transform -1 0 1598 0 1 2225
box 0 0 8 49
use OR2X2  OR2X2_136
timestamp 1516325494
transform -1 0 1617 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_332
timestamp 1516325494
transform 1 0 1617 0 1 2225
box 0 0 19 49
use FILL  FILL_OR2X2_132
timestamp 1516325494
transform -1 0 1644 0 1 2225
box 0 0 8 49
use OR2X2  OR2X2_132
timestamp 1516325494
transform -1 0 1663 0 1 2225
box 0 0 19 49
use FILL  FILL_OR2X2_131
timestamp 1516325494
transform -1 0 1671 0 1 2225
box 0 0 8 49
use OR2X2  OR2X2_131
timestamp 1516325494
transform -1 0 1689 0 1 2225
box 0 0 19 49
use FILL  FILL_AND2X2_140
timestamp 1516325494
transform -1 0 1697 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_140
timestamp 1516325494
transform -1 0 1716 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1390
timestamp 1516325494
transform -1 0 1735 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1596
timestamp 1516325494
transform -1 0 1754 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_289
timestamp 1516325494
transform -1 0 1773 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_290
timestamp 1516325494
transform -1 0 1792 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1826
timestamp 1516325494
transform 1 0 1792 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1824
timestamp 1516325494
transform 1 0 1811 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1690
timestamp 1516325494
transform 1 0 1830 0 1 2225
box 0 0 19 49
use FILL  FILL_OR2X2_47
timestamp 1516325494
transform -1 0 1857 0 1 2225
box 0 0 8 49
use OR2X2  OR2X2_47
timestamp 1516325494
transform -1 0 1875 0 1 2225
box 0 0 19 49
use FILL  FILL_AND2X2_49
timestamp 1516325494
transform -1 0 1883 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_49
timestamp 1516325494
transform -1 0 1902 0 1 2225
box 0 0 19 49
use FILL  FILL_AND2X2_50
timestamp 1516325494
transform -1 0 1910 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_50
timestamp 1516325494
transform -1 0 1929 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1456
timestamp 1516325494
transform 1 0 1929 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1210
timestamp 1516325494
transform 1 0 1948 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1458
timestamp 1516325494
transform -1 0 1986 0 1 2225
box 0 0 19 49
use FILL  FILL_AND2X2_18
timestamp 1516325494
transform -1 0 1994 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_18
timestamp 1516325494
transform -1 0 2012 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1823
timestamp 1516325494
transform -1 0 2031 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1686
timestamp 1516325494
transform -1 0 2050 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1409
timestamp 1516325494
transform -1 0 2069 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1408
timestamp 1516325494
transform -1 0 2088 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1146
timestamp 1516325494
transform -1 0 2107 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_883
timestamp 1516325494
transform 1 0 2107 0 1 2225
box 0 0 15 49
use NAND2X1  NAND2X1_901
timestamp 1516325494
transform 1 0 2122 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_421
timestamp 1516325494
transform 1 0 2138 0 1 2225
box 0 0 53 49
use NAND2X1  NAND2X1_389
timestamp 1516325494
transform 1 0 2191 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_389
timestamp 1516325494
transform -1 0 2236 0 1 2225
box 0 0 30 49
use AND2X2  AND2X2_1457
timestamp 1516325494
transform -1 0 2255 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1208
timestamp 1516325494
transform -1 0 2274 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_39
timestamp 1516325494
transform 1 0 2274 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_39
timestamp 1516325494
transform -1 0 2320 0 1 2225
box 0 0 30 49
use OR2X2  OR2X2_1209
timestamp 1516325494
transform -1 0 2339 0 1 2225
box 0 0 19 49
use FILL  FILL_BUFX2_674
timestamp 1516325494
transform -1 0 2347 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_674
timestamp 1516325494
transform -1 0 2362 0 1 2225
box 0 0 15 49
use AND2X2  AND2X2_1819
timestamp 1516325494
transform -1 0 2381 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1681
timestamp 1516325494
transform -1 0 2400 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_23
timestamp 1516325494
transform 1 0 2400 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_599
timestamp 1516325494
transform 1 0 2415 0 1 2225
box 0 0 53 49
use MUX2X1  MUX2X1_23
timestamp 1516325494
transform -1 0 2498 0 1 2225
box 0 0 30 49
use FILL  FILL_BUFX2_416
timestamp 1516325494
transform 1 0 2499 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_416
timestamp 1516325494
transform 1 0 2506 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_168
timestamp 1516325494
transform 1 0 2521 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_168
timestamp 1516325494
transform 1 0 2529 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_261
timestamp 1516325494
transform 1 0 2544 0 1 2225
box 0 0 53 49
use MUX2X1  MUX2X1_581
timestamp 1516325494
transform 1 0 2597 0 1 2225
box 0 0 30 49
use NAND2X1  NAND2X1_581
timestamp 1516325494
transform 1 0 2628 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_229
timestamp 1516325494
transform 1 0 2643 0 1 2225
box 0 0 53 49
use OR2X2  OR2X2_1380
timestamp 1516325494
transform -1 0 2715 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_197
timestamp 1516325494
transform 1 0 2715 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_197
timestamp 1516325494
transform -1 0 2760 0 1 2225
box 0 0 30 49
use FILL  FILL_AND2X2_43
timestamp 1516325494
transform 1 0 2761 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_43
timestamp 1516325494
transform 1 0 2768 0 1 2225
box 0 0 19 49
use FILL  FILL_OR2X2_41
timestamp 1516325494
transform -1 0 2795 0 1 2225
box 0 0 8 49
use OR2X2  OR2X2_41
timestamp 1516325494
transform -1 0 2814 0 1 2225
box 0 0 19 49
use FILL  FILL_AND2X2_42
timestamp 1516325494
transform -1 0 2822 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_42
timestamp 1516325494
transform -1 0 2841 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1446
timestamp 1516325494
transform 1 0 2841 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1447
timestamp 1516325494
transform -1 0 2879 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_583
timestamp 1516325494
transform 1 0 2879 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_583
timestamp 1516325494
transform -1 0 2924 0 1 2225
box 0 0 30 49
use MUX2X1  MUX2X1_753
timestamp 1516325494
transform -1 0 2954 0 1 2225
box 0 0 30 49
use OR2X2  OR2X2_1229
timestamp 1516325494
transform -1 0 2974 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1471
timestamp 1516325494
transform -1 0 2993 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1228
timestamp 1516325494
transform -1 0 3012 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1473
timestamp 1516325494
transform -1 0 3031 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1472
timestamp 1516325494
transform -1 0 3050 0 1 2225
box 0 0 19 49
use FILL  FILL_AND2X2_59
timestamp 1516325494
transform 1 0 3050 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_59
timestamp 1516325494
transform 1 0 3057 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1450
timestamp 1516325494
transform 1 0 3076 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1198
timestamp 1516325494
transform -1 0 3114 0 1 2225
box 0 0 19 49
use MUX2X1  MUX2X1_359
timestamp 1516325494
transform 1 0 3114 0 1 2225
box 0 0 30 49
use NAND2X1  NAND2X1_359
timestamp 1516325494
transform -1 0 3160 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_327
timestamp 1516325494
transform -1 0 3213 0 1 2225
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_837
timestamp 1516325494
transform -1 0 3266 0 1 2225
box 0 0 53 49
use FILL  FILL_BUFX2_257
timestamp 1516325494
transform 1 0 3266 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_257
timestamp 1516325494
transform 1 0 3274 0 1 2225
box 0 0 15 49
use NOR2X1  NOR2X1_146
timestamp 1516325494
transform -1 0 3304 0 1 2225
box 0 0 15 49
use AND2X2  AND2X2_1240
timestamp 1516325494
transform -1 0 3323 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_977
timestamp 1516325494
transform -1 0 3342 0 1 2225
box 0 0 19 49
use OAI21X1  OAI21X1_112
timestamp 1516325494
transform 1 0 3342 0 1 2225
box 0 0 19 49
use NAND2X1  NAND2X1_826
timestamp 1516325494
transform 1 0 3361 0 1 2225
box 0 0 15 49
use INVX1  INVX1_288
timestamp 1516325494
transform -1 0 3387 0 1 2225
box 0 0 11 49
use NAND2X1  NAND2X1_825
timestamp 1516325494
transform 1 0 3388 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_305
timestamp 1516325494
transform 1 0 3403 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_305
timestamp 1516325494
transform 1 0 3411 0 1 2225
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_810
timestamp 1516325494
transform -1 0 3479 0 1 2225
box 0 0 53 49
use FILL  FILL_BUFX2_854
timestamp 1516325494
transform 1 0 3479 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_854
timestamp 1516325494
transform 1 0 3487 0 1 2225
box 0 0 15 49
use INVX1  INVX1_273
timestamp 1516325494
transform -1 0 3513 0 1 2225
box 0 0 11 49
use FILL  FILL_BUFX2_407
timestamp 1516325494
transform -1 0 3521 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_407
timestamp 1516325494
transform -1 0 3536 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_612
timestamp 1516325494
transform -1 0 3544 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_612
timestamp 1516325494
transform -1 0 3559 0 1 2225
box 0 0 15 49
use FILL  FILL_BUFX2_259
timestamp 1516325494
transform 1 0 3559 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_259
timestamp 1516325494
transform 1 0 3566 0 1 2225
box 0 0 15 49
use OAI21X1  OAI21X1_125
timestamp 1516325494
transform 1 0 3582 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_984
timestamp 1516325494
transform 1 0 3601 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1248
timestamp 1516325494
transform 1 0 3620 0 1 2225
box 0 0 19 49
use AOI22X1  AOI22X1_32
timestamp 1516325494
transform 1 0 3639 0 1 2225
box 0 0 23 49
use OAI21X1  OAI21X1_126
timestamp 1516325494
transform -1 0 3680 0 1 2225
box 0 0 19 49
use FILL  FILL_BUFX2_304
timestamp 1516325494
transform -1 0 3688 0 1 2225
box 0 0 8 49
use BUFX2  BUFX2_304
timestamp 1516325494
transform -1 0 3703 0 1 2225
box 0 0 15 49
use NAND2X1  NAND2X1_875
timestamp 1516325494
transform 1 0 3703 0 1 2225
box 0 0 15 49
use NAND2X1  NAND2X1_782
timestamp 1516325494
transform 1 0 3718 0 1 2225
box 0 0 15 49
use MUX2X1  MUX2X1_819
timestamp 1516325494
transform -1 0 3764 0 1 2225
box 0 0 30 49
use OAI21X1  OAI21X1_168
timestamp 1516325494
transform 1 0 3764 0 1 2225
box 0 0 19 49
use OR2X2  OR2X2_1007
timestamp 1516325494
transform 1 0 3783 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1261
timestamp 1516325494
transform -1 0 3821 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1276
timestamp 1516325494
transform 1 0 3821 0 1 2225
box 0 0 19 49
use AND2X2  AND2X2_1278
timestamp 1516325494
transform 1 0 3840 0 1 2225
box 0 0 19 49
use FILL  FILL_46_1
timestamp 1516325494
transform 1 0 3859 0 1 2225
box 0 0 8 49
use AND2X2  AND2X2_1102
timestamp 1516325494
transform 1 0 2 0 -1 2224
box 0 0 19 49
use INVX1  INVX1_95
timestamp 1516325494
transform -1 0 32 0 -1 2224
box 0 0 11 49
use XOR2X1  XOR2X1_48
timestamp 1516325494
transform 1 0 32 0 -1 2224
box 0 0 34 49
use INVX1  INVX1_96
timestamp 1516325494
transform -1 0 78 0 -1 2224
box 0 0 11 49
use NOR2X1  NOR2X1_93
timestamp 1516325494
transform -1 0 93 0 -1 2224
box 0 0 15 49
use INVX1  INVX1_97
timestamp 1516325494
transform -1 0 104 0 -1 2224
box 0 0 11 49
use INVX1  INVX1_92
timestamp 1516325494
transform -1 0 13 0 1 2126
box 0 0 11 49
use OR2X2  OR2X2_897
timestamp 1516325494
transform -1 0 32 0 1 2126
box 0 0 19 49
use INVX1  INVX1_93
timestamp 1516325494
transform -1 0 43 0 1 2126
box 0 0 11 49
use XNOR2X1  XNOR2X1_29
timestamp 1516325494
transform -1 0 78 0 1 2126
box 0 0 34 49
use NOR2X1  NOR2X1_92
timestamp 1516325494
transform -1 0 93 0 1 2126
box 0 0 15 49
use INVX1  INVX1_94
timestamp 1516325494
transform -1 0 104 0 1 2126
box 0 0 11 49
use XNOR2X1  XNOR2X1_31
timestamp 1516325494
transform 1 0 105 0 -1 2224
box 0 0 34 49
use XOR2X1  XOR2X1_26
timestamp 1516325494
transform -1 0 173 0 -1 2224
box 0 0 34 49
use NAND2X1  NAND2X1_701
timestamp 1516325494
transform 1 0 173 0 -1 2224
box 0 0 15 49
use AND2X2  AND2X2_1023
timestamp 1516325494
transform 1 0 188 0 -1 2224
box 0 0 19 49
use FILL  FILL_BUFX2_786
timestamp 1516325494
transform -1 0 215 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_786
timestamp 1516325494
transform -1 0 230 0 -1 2224
box 0 0 15 49
use AND2X2  AND2X2_1024
timestamp 1516325494
transform 1 0 230 0 -1 2224
box 0 0 19 49
use NOR2X1  NOR2X1_79
timestamp 1516325494
transform 1 0 249 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_848
timestamp 1516325494
transform -1 0 283 0 -1 2224
box 0 0 19 49
use NOR2X1  NOR2X1_75
timestamp 1516325494
transform -1 0 298 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_862
timestamp 1516325494
transform 1 0 298 0 -1 2224
box 0 0 19 49
use OAI21X1  OAI21X1_17
timestamp 1516325494
transform -1 0 336 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1039
timestamp 1516325494
transform -1 0 355 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1038
timestamp 1516325494
transform -1 0 374 0 -1 2224
box 0 0 19 49
use NAND3X1  NAND3X1_60
timestamp 1516325494
transform -1 0 393 0 -1 2224
box 0 0 19 49
use NOR2X1  NOR2X1_70
timestamp 1516325494
transform -1 0 408 0 -1 2224
box 0 0 15 49
use NAND2X1  NAND2X1_691
timestamp 1516325494
transform -1 0 424 0 -1 2224
box 0 0 15 49
use AOI21X1  AOI21X1_22
timestamp 1516325494
transform -1 0 443 0 -1 2224
box 0 0 19 49
use XOR2X1  XOR2X1_21
timestamp 1516325494
transform 1 0 443 0 -1 2224
box 0 0 34 49
use NAND2X1  NAND2X1_690
timestamp 1516325494
transform -1 0 492 0 -1 2224
box 0 0 15 49
use NOR2X1  NOR2X1_71
timestamp 1516325494
transform 1 0 492 0 -1 2224
box 0 0 15 49
use NAND2X1  NAND2X1_686
timestamp 1516325494
transform 1 0 507 0 -1 2224
box 0 0 15 49
use AOI21X1  AOI21X1_19
timestamp 1516325494
transform 1 0 523 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_795
timestamp 1516325494
transform 1 0 542 0 -1 2224
box 0 0 19 49
use NOR2X1  NOR2X1_65
timestamp 1516325494
transform -1 0 576 0 -1 2224
box 0 0 15 49
use NOR2X1  NOR2X1_64
timestamp 1516325494
transform -1 0 591 0 -1 2224
box 0 0 15 49
use INVX1  INVX1_43
timestamp 1516325494
transform 1 0 591 0 -1 2224
box 0 0 11 49
use FILL  FILL_BUFX2_849
timestamp 1516325494
transform -1 0 610 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_849
timestamp 1516325494
transform -1 0 625 0 -1 2224
box 0 0 15 49
use INVX1  INVX1_183
timestamp 1516325494
transform -1 0 636 0 -1 2224
box 0 0 11 49
use XNOR2X1  XNOR2X1_28
timestamp 1516325494
transform -1 0 139 0 1 2126
box 0 0 34 49
use XNOR2X1  XNOR2X1_30
timestamp 1516325494
transform -1 0 173 0 1 2126
box 0 0 34 49
use NAND3X1  NAND3X1_47
timestamp 1516325494
transform 1 0 173 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_680
timestamp 1516325494
transform 1 0 192 0 1 2126
box 0 0 15 49
use NAND2X1  NAND2X1_679
timestamp 1516325494
transform -1 0 222 0 1 2126
box 0 0 15 49
use NOR2X1  NOR2X1_76
timestamp 1516325494
transform 1 0 222 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_150
timestamp 1516325494
transform 1 0 238 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_150
timestamp 1516325494
transform 1 0 245 0 1 2126
box 0 0 15 49
use NAND3X1  NAND3X1_55
timestamp 1516325494
transform 1 0 260 0 1 2126
box 0 0 19 49
use AOI21X1  AOI21X1_24
timestamp 1516325494
transform -1 0 298 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_699
timestamp 1516325494
transform -1 0 313 0 1 2126
box 0 0 15 49
use NAND2X1  NAND2X1_698
timestamp 1516325494
transform -1 0 329 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_622
timestamp 1516325494
transform 1 0 329 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_622
timestamp 1516325494
transform 1 0 336 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_625
timestamp 1516325494
transform -1 0 360 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_625
timestamp 1516325494
transform -1 0 374 0 1 2126
box 0 0 15 49
use AOI21X1  AOI21X1_10
timestamp 1516325494
transform -1 0 393 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1037
timestamp 1516325494
transform -1 0 412 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_703
timestamp 1516325494
transform -1 0 427 0 1 2126
box 0 0 15 49
use NAND2X1  NAND2X1_702
timestamp 1516325494
transform -1 0 443 0 1 2126
box 0 0 15 49
use NOR2X1  NOR2X1_72
timestamp 1516325494
transform 1 0 443 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_562
timestamp 1516325494
transform -1 0 466 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_562
timestamp 1516325494
transform -1 0 481 0 1 2126
box 0 0 15 49
use AND2X2  AND2X2_952
timestamp 1516325494
transform -1 0 500 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_687
timestamp 1516325494
transform -1 0 515 0 1 2126
box 0 0 15 49
use XOR2X1  XOR2X1_19
timestamp 1516325494
transform -1 0 549 0 1 2126
box 0 0 34 49
use NOR2X1  NOR2X1_68
timestamp 1516325494
transform 1 0 549 0 1 2126
box 0 0 15 49
use OR2X2  OR2X2_901
timestamp 1516325494
transform 1 0 564 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1106
timestamp 1516325494
transform 1 0 583 0 1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_148
timestamp 1516325494
transform 1 0 602 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_148
timestamp 1516325494
transform 1 0 610 0 1 2126
box 0 0 15 49
use INVX1  INVX1_107
timestamp 1516325494
transform -1 0 636 0 1 2126
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_731
timestamp 1516325494
transform -1 0 690 0 -1 2224
box 0 0 53 49
use INVX1  INVX1_147
timestamp 1516325494
transform 1 0 690 0 -1 2224
box 0 0 11 49
use AND2X2  AND2X2_1625
timestamp 1516325494
transform 1 0 701 0 -1 2224
box 0 0 19 49
use INVX1  INVX1_161
timestamp 1516325494
transform 1 0 720 0 -1 2224
box 0 0 11 49
use FILL  FILL_AND2X2_158
timestamp 1516325494
transform 1 0 732 0 -1 2224
box 0 0 8 49
use AND2X2  AND2X2_158
timestamp 1516325494
transform 1 0 739 0 -1 2224
box 0 0 19 49
use INVX1  INVX1_226
timestamp 1516325494
transform -1 0 769 0 -1 2224
box 0 0 11 49
use MUX2X1  MUX2X1_790
timestamp 1516325494
transform -1 0 800 0 -1 2224
box 0 0 30 49
use INVX1  INVX1_177
timestamp 1516325494
transform 1 0 800 0 -1 2224
box 0 0 11 49
use MUX2X1  MUX2X1_85
timestamp 1516325494
transform 1 0 811 0 -1 2224
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_117
timestamp 1516325494
transform -1 0 895 0 -1 2224
box 0 0 53 49
use NAND2X1  NAND2X1_85
timestamp 1516325494
transform -1 0 910 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_754
timestamp 1516325494
transform 1 0 910 0 -1 2224
box 0 0 30 49
use OR2X2  OR2X2_1640
timestamp 1516325494
transform 1 0 941 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_66
timestamp 1516325494
transform 1 0 960 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_66
timestamp 1516325494
transform 1 0 967 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1787
timestamp 1516325494
transform 1 0 986 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1253
timestamp 1516325494
transform 1 0 1005 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1254
timestamp 1516325494
transform -1 0 1043 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_67
timestamp 1516325494
transform -1 0 1051 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_67
timestamp 1516325494
transform -1 0 1070 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_369
timestamp 1516325494
transform 1 0 1070 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_344
timestamp 1516325494
transform 1 0 1089 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_345
timestamp 1516325494
transform 1 0 1108 0 -1 2224
box 0 0 19 49
use MUX2X1  MUX2X1_321
timestamp 1516325494
transform 1 0 1127 0 -1 2224
box 0 0 30 49
use NAND2X1  NAND2X1_321
timestamp 1516325494
transform -1 0 1172 0 -1 2224
box 0 0 15 49
use NAND2X1  NAND2X1_97
timestamp 1516325494
transform 1 0 1172 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_97
timestamp 1516325494
transform -1 0 1218 0 -1 2224
box 0 0 30 49
use OR2X2  OR2X2_1038
timestamp 1516325494
transform 1 0 1218 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1324
timestamp 1516325494
transform 1 0 1237 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1783
timestamp 1516325494
transform -1 0 1275 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1635
timestamp 1516325494
transform -1 0 1294 0 -1 2224
box 0 0 19 49
use NAND2X1  NAND2X1_149
timestamp 1516325494
transform 1 0 1294 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_149
timestamp 1516325494
transform 1 0 1309 0 -1 2224
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_85
timestamp 1516325494
transform -1 0 1393 0 -1 2224
box 0 0 53 49
use OR2X2  OR2X2_1634
timestamp 1516325494
transform -1 0 1412 0 -1 2224
box 0 0 19 49
use FILL  FILL_BUFX2_579
timestamp 1516325494
transform 1 0 1412 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_579
timestamp 1516325494
transform 1 0 1419 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_1639
timestamp 1516325494
transform -1 0 1454 0 -1 2224
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_501
timestamp 1516325494
transform 1 0 1454 0 -1 2224
box 0 0 53 49
use NAND2X1  NAND2X1_565
timestamp 1516325494
transform 1 0 1507 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_565
timestamp 1516325494
transform -1 0 1552 0 -1 2224
box 0 0 30 49
use NAND2X1  NAND2X1_341
timestamp 1516325494
transform 1 0 1552 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_341
timestamp 1516325494
transform -1 0 1598 0 -1 2224
box 0 0 30 49
use FILL  FILL_BUFX2_466
timestamp 1516325494
transform -1 0 1606 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_466
timestamp 1516325494
transform -1 0 1621 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_333
timestamp 1516325494
transform -1 0 1640 0 -1 2224
box 0 0 19 49
use FILL  FILL_BUFX2_113
timestamp 1516325494
transform 1 0 1640 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_113
timestamp 1516325494
transform 1 0 1647 0 -1 2224
box 0 0 15 49
use OAI21X1  OAI21X1_71
timestamp 1516325494
transform 1 0 637 0 1 2126
box 0 0 19 49
use INVX1  INVX1_48
timestamp 1516325494
transform 1 0 656 0 1 2126
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_745
timestamp 1516325494
transform -1 0 720 0 1 2126
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_746
timestamp 1516325494
transform -1 0 773 0 1 2126
box 0 0 53 49
use MUX2X1  MUX2X1_774
timestamp 1516325494
transform 1 0 773 0 1 2126
box 0 0 30 49
use FILL  FILL_OR2X2_148
timestamp 1516325494
transform 1 0 804 0 1 2126
box 0 0 8 49
use OR2X2  OR2X2_148
timestamp 1516325494
transform 1 0 811 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_159
timestamp 1516325494
transform -1 0 838 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_159
timestamp 1516325494
transform -1 0 857 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_117
timestamp 1516325494
transform 1 0 857 0 1 2126
box 0 0 15 49
use OR2X2  OR2X2_1637
timestamp 1516325494
transform 1 0 872 0 1 2126
box 0 0 19 49
use INVX1  INVX1_162
timestamp 1516325494
transform 1 0 891 0 1 2126
box 0 0 11 49
use AND2X2  AND2X2_1101
timestamp 1516325494
transform 1 0 2 0 -1 2126
box 0 0 19 49
use NOR2X1  NOR2X1_91
timestamp 1516325494
transform -1 0 36 0 -1 2126
box 0 0 15 49
use INVX1  INVX1_91
timestamp 1516325494
transform -1 0 47 0 -1 2126
box 0 0 11 49
use XNOR2X1  XNOR2X1_27
timestamp 1516325494
transform 1 0 48 0 -1 2126
box 0 0 34 49
use XOR2X1  XOR2X1_47
timestamp 1516325494
transform -1 0 116 0 -1 2126
box 0 0 34 49
use AND2X2  AND2X2_897
timestamp 1516325494
transform -1 0 135 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_751
timestamp 1516325494
transform -1 0 154 0 -1 2126
box 0 0 19 49
use NOR2X1  NOR2X1_55
timestamp 1516325494
transform -1 0 169 0 -1 2126
box 0 0 15 49
use AND2X2  AND2X2_896
timestamp 1516325494
transform -1 0 188 0 -1 2126
box 0 0 19 49
use NAND3X1  NAND3X1_48
timestamp 1516325494
transform -1 0 207 0 -1 2126
box 0 0 19 49
use AOI21X1  AOI21X1_16
timestamp 1516325494
transform 1 0 207 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_966
timestamp 1516325494
transform -1 0 245 0 -1 2126
box 0 0 19 49
use INVX1  INVX1_44
timestamp 1516325494
transform 1 0 245 0 -1 2126
box 0 0 11 49
use AOI21X1  AOI21X1_21
timestamp 1516325494
transform -1 0 276 0 -1 2126
box 0 0 19 49
use NAND3X1  NAND3X1_56
timestamp 1516325494
transform -1 0 295 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1017
timestamp 1516325494
transform 1 0 295 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1018
timestamp 1516325494
transform 1 0 314 0 -1 2126
box 0 0 19 49
use XOR2X1  XOR2X1_20
timestamp 1516325494
transform -1 0 367 0 -1 2126
box 0 0 34 49
use OR2X2  OR2X2_697
timestamp 1516325494
transform -1 0 386 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_688
timestamp 1516325494
transform 1 0 386 0 -1 2126
box 0 0 15 49
use AOI21X1  AOI21X1_20
timestamp 1516325494
transform 1 0 401 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_805
timestamp 1516325494
transform -1 0 439 0 -1 2126
box 0 0 19 49
use NOR2X1  NOR2X1_67
timestamp 1516325494
transform -1 0 454 0 -1 2126
box 0 0 15 49
use OR2X2  OR2X2_844
timestamp 1516325494
transform 1 0 454 0 -1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_564
timestamp 1516325494
transform 1 0 473 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_564
timestamp 1516325494
transform 1 0 481 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_147
timestamp 1516325494
transform 1 0 496 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_147
timestamp 1516325494
transform 1 0 504 0 -1 2126
box 0 0 15 49
use XOR2X1  XOR2X1_51
timestamp 1516325494
transform 1 0 519 0 -1 2126
box 0 0 34 49
use AND2X2  AND2X2_953
timestamp 1516325494
transform 1 0 553 0 -1 2126
box 0 0 19 49
use INVX1  INVX1_105
timestamp 1516325494
transform -1 0 583 0 -1 2126
box 0 0 11 49
use XNOR2X1  XNOR2X1_37
timestamp 1516325494
transform 1 0 583 0 -1 2126
box 0 0 34 49
use NOR2X1  NOR2X1_96
timestamp 1516325494
transform 1 0 618 0 -1 2126
box 0 0 15 49
use INVX1  INVX1_106
timestamp 1516325494
transform -1 0 644 0 -1 2126
box 0 0 11 49
use AND2X2  AND2X2_1070
timestamp 1516325494
transform -1 0 663 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_833
timestamp 1516325494
transform -1 0 682 0 -1 2126
box 0 0 19 49
use INVX1  INVX1_49
timestamp 1516325494
transform 1 0 682 0 -1 2126
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_744
timestamp 1516325494
transform -1 0 747 0 -1 2126
box 0 0 53 49
use FILL  FILL_BUFX2_221
timestamp 1516325494
transform -1 0 755 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_221
timestamp 1516325494
transform -1 0 769 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_726
timestamp 1516325494
transform -1 0 823 0 -1 2126
box 0 0 53 49
use OR2X2  OR2X2_1431
timestamp 1516325494
transform 1 0 823 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1627
timestamp 1516325494
transform -1 0 861 0 -1 2126
box 0 0 19 49
use INVX1  INVX1_185
timestamp 1516325494
transform -1 0 872 0 -1 2126
box 0 0 11 49
use MUX2X1  MUX2X1_117
timestamp 1516325494
transform -1 0 902 0 -1 2126
box 0 0 30 49
use INVX1  INVX1_187
timestamp 1516325494
transform 1 0 903 0 1 2126
box 0 0 11 49
use OR2X2  OR2X2_1638
timestamp 1516325494
transform 1 0 914 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1785
timestamp 1516325494
transform 1 0 933 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1786
timestamp 1516325494
transform 1 0 952 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1641
timestamp 1516325494
transform -1 0 990 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1788
timestamp 1516325494
transform -1 0 1009 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_264
timestamp 1516325494
transform -1 0 1017 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_264
timestamp 1516325494
transform -1 0 1036 0 1 2126
box 0 0 19 49
use INVX1  INVX1_207
timestamp 1516325494
transform -1 0 1047 0 1 2126
box 0 0 11 49
use FILL  FILL_BUFX2_129
timestamp 1516325494
transform 1 0 1047 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_129
timestamp 1516325494
transform 1 0 1055 0 1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_78
timestamp 1516325494
transform 1 0 1070 0 1 2126
box 0 0 53 49
use MUX2X1  MUX2X1_142
timestamp 1516325494
transform -1 0 1153 0 1 2126
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_449
timestamp 1516325494
transform -1 0 1206 0 1 2126
box 0 0 53 49
use OR2X2  OR2X2_1034
timestamp 1516325494
transform 1 0 1207 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1545
timestamp 1516325494
transform -1 0 1245 0 1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_65
timestamp 1516325494
transform 1 0 1245 0 1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_129
timestamp 1516325494
transform 1 0 1298 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_129
timestamp 1516325494
transform -1 0 1343 0 1 2126
box 0 0 30 49
use FILL  FILL_BUFX2_550
timestamp 1516325494
transform 1 0 1343 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_550
timestamp 1516325494
transform 1 0 1351 0 1 2126
box 0 0 15 49
use OAI21X1  OAI21X1_45
timestamp 1516325494
transform 1 0 1366 0 1 2126
box 0 0 19 49
use INVX2  INVX2_34
timestamp 1516325494
transform 1 0 1385 0 1 2126
box 0 0 11 49
use OAI21X1  OAI21X1_38
timestamp 1516325494
transform 1 0 1397 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_728
timestamp 1516325494
transform -1 0 1431 0 1 2126
box 0 0 15 49
use INVX2  INVX2_27
timestamp 1516325494
transform 1 0 1431 0 1 2126
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_63
timestamp 1516325494
transform 1 0 1442 0 1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_447
timestamp 1516325494
transform 1 0 1495 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_447
timestamp 1516325494
transform -1 0 1541 0 1 2126
box 0 0 30 49
use FILL  FILL_BUFX2_122
timestamp 1516325494
transform 1 0 1541 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_122
timestamp 1516325494
transform 1 0 1549 0 1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_45
timestamp 1516325494
transform -1 0 1617 0 1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_715
timestamp 1516325494
transform -1 0 1632 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_429
timestamp 1516325494
transform 1 0 1632 0 1 2126
box 0 0 30 49
use FILL  FILL_BUFX2_120
timestamp 1516325494
transform 1 0 1663 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_120
timestamp 1516325494
transform 1 0 1670 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_328
timestamp 1516325494
transform -1 0 1704 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1593
timestamp 1516325494
transform 1 0 1704 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1594
timestamp 1516325494
transform -1 0 1742 0 -1 2224
box 0 0 19 49
use FILL  FILL_AND2X2_139
timestamp 1516325494
transform 1 0 1742 0 -1 2224
box 0 0 8 49
use AND2X2  AND2X2_139
timestamp 1516325494
transform 1 0 1750 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_326
timestamp 1516325494
transform -1 0 1788 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_347
timestamp 1516325494
transform -1 0 1807 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1803
timestamp 1516325494
transform 1 0 1807 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_53
timestamp 1516325494
transform 1 0 1826 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_53
timestamp 1516325494
transform 1 0 1834 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_24
timestamp 1516325494
transform 1 0 1853 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_24
timestamp 1516325494
transform 1 0 1860 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_20
timestamp 1516325494
transform -1 0 1887 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_20
timestamp 1516325494
transform -1 0 1906 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_19
timestamp 1516325494
transform -1 0 1914 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_19
timestamp 1516325494
transform -1 0 1932 0 -1 2224
box 0 0 19 49
use FILL  FILL_AND2X2_19
timestamp 1516325494
transform -1 0 1940 0 -1 2224
box 0 0 8 49
use AND2X2  AND2X2_19
timestamp 1516325494
transform -1 0 1959 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_18
timestamp 1516325494
transform -1 0 1967 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_18
timestamp 1516325494
transform -1 0 1986 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1410
timestamp 1516325494
transform 1 0 1986 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1150
timestamp 1516325494
transform 1 0 2005 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1151
timestamp 1516325494
transform 1 0 2024 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1163
timestamp 1516325494
transform 1 0 2043 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1145
timestamp 1516325494
transform -1 0 2081 0 -1 2224
box 0 0 19 49
use FILL  FILL_BUFX2_117
timestamp 1516325494
transform -1 0 2089 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_117
timestamp 1516325494
transform -1 0 2103 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_828
timestamp 1516325494
transform 1 0 2103 0 -1 2224
box 0 0 30 49
use AND2X2  AND2X2_1411
timestamp 1516325494
transform -1 0 2153 0 -1 2224
box 0 0 19 49
use MUX2X1  MUX2X1_846
timestamp 1516325494
transform -1 0 2183 0 -1 2224
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_631
timestamp 1516325494
transform -1 0 2236 0 -1 2224
box 0 0 53 49
use OR2X2  OR2X2_1142
timestamp 1516325494
transform 1 0 2236 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1405
timestamp 1516325494
transform 1 0 2255 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1149
timestamp 1516325494
transform -1 0 2293 0 -1 2224
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_293
timestamp 1516325494
transform 1 0 2293 0 -1 2224
box 0 0 53 49
use NAND2X1  NAND2X1_485
timestamp 1516325494
transform 1 0 2347 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_485
timestamp 1516325494
transform -1 0 2392 0 -1 2224
box 0 0 30 49
use MUX2X1  MUX2X1_487
timestamp 1516325494
transform 1 0 2392 0 -1 2224
box 0 0 30 49
use NAND2X1  NAND2X1_487
timestamp 1516325494
transform -1 0 2438 0 -1 2224
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_295
timestamp 1516325494
transform -1 0 2491 0 -1 2224
box 0 0 53 49
use OR2X2  OR2X2_1141
timestamp 1516325494
transform -1 0 2510 0 -1 2224
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_581
timestamp 1516325494
transform 1 0 2510 0 -1 2224
box 0 0 53 49
use NAND2X1  NAND2X1_5
timestamp 1516325494
transform 1 0 2563 0 -1 2224
box 0 0 15 49
use MUX2X1  MUX2X1_5
timestamp 1516325494
transform -1 0 2608 0 -1 2224
box 0 0 30 49
use MUX2X1  MUX2X1_251
timestamp 1516325494
transform 1 0 2609 0 -1 2224
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_187
timestamp 1516325494
transform -1 0 2692 0 -1 2224
box 0 0 53 49
use NAND2X1  NAND2X1_251
timestamp 1516325494
transform -1 0 2707 0 -1 2224
box 0 0 15 49
use AND2X2  AND2X2_1904
timestamp 1516325494
transform -1 0 2727 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_340
timestamp 1516325494
transform 1 0 2727 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1140
timestamp 1516325494
transform 1 0 2746 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_1164
timestamp 1516325494
transform 1 0 2765 0 -1 2224
box 0 0 19 49
use MUX2X1  MUX2X1_199
timestamp 1516325494
transform 1 0 2784 0 -1 2224
box 0 0 30 49
use NAND2X1  NAND2X1_199
timestamp 1516325494
transform -1 0 2829 0 -1 2224
box 0 0 15 49
use FILL  FILL_OR2X2_45
timestamp 1516325494
transform -1 0 2837 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_45
timestamp 1516325494
transform -1 0 2856 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_59
timestamp 1516325494
transform -1 0 2864 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_59
timestamp 1516325494
transform -1 0 2882 0 -1 2224
box 0 0 19 49
use FILL  FILL_BUFX2_473
timestamp 1516325494
transform 1 0 2882 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_473
timestamp 1516325494
transform 1 0 2890 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_1679
timestamp 1516325494
transform -1 0 2924 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_44
timestamp 1516325494
transform -1 0 2932 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_44
timestamp 1516325494
transform -1 0 2951 0 -1 2224
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_155
timestamp 1516325494
transform 1 0 2951 0 -1 2224
box 0 0 53 49
use OR2X2  OR2X2_1139
timestamp 1516325494
transform -1 0 3023 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1402
timestamp 1516325494
transform 1 0 3023 0 -1 2224
box 0 0 19 49
use FILL  FILL_AND2X2_14
timestamp 1516325494
transform -1 0 3050 0 -1 2224
box 0 0 8 49
use AND2X2  AND2X2_14
timestamp 1516325494
transform -1 0 3069 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_58
timestamp 1516325494
transform -1 0 3077 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_58
timestamp 1516325494
transform -1 0 3095 0 -1 2224
box 0 0 19 49
use FILL  FILL_OR2X2_57
timestamp 1516325494
transform -1 0 3103 0 -1 2224
box 0 0 8 49
use OR2X2  OR2X2_57
timestamp 1516325494
transform -1 0 3122 0 -1 2224
box 0 0 19 49
use FILL  FILL_AND2X2_60
timestamp 1516325494
transform -1 0 3130 0 -1 2224
box 0 0 8 49
use AND2X2  AND2X2_60
timestamp 1516325494
transform -1 0 3148 0 -1 2224
box 0 0 19 49
use MUX2X1  MUX2X1_263
timestamp 1516325494
transform 1 0 3148 0 -1 2224
box 0 0 30 49
use NAND2X1  NAND2X1_263
timestamp 1516325494
transform -1 0 3194 0 -1 2224
box 0 0 15 49
use AND2X2  AND2X2_1449
timestamp 1516325494
transform -1 0 3213 0 -1 2224
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_135
timestamp 1516325494
transform -1 0 3266 0 -1 2224
box 0 0 53 49
use OAI21X1  OAI21X1_109
timestamp 1516325494
transform -1 0 3285 0 -1 2224
box 0 0 19 49
use INVX1  INVX1_291
timestamp 1516325494
transform -1 0 3296 0 -1 2224
box 0 0 11 49
use NAND2X1  NAND2X1_786
timestamp 1516325494
transform 1 0 3297 0 -1 2224
box 0 0 15 49
use INVX1  INVX1_292
timestamp 1516325494
transform 1 0 3312 0 -1 2224
box 0 0 11 49
use AND2X2  AND2X2_1238
timestamp 1516325494
transform 1 0 3323 0 -1 2224
box 0 0 19 49
use OR2X2  OR2X2_976
timestamp 1516325494
transform 1 0 3342 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1239
timestamp 1516325494
transform 1 0 3361 0 -1 2224
box 0 0 19 49
use OAI21X1  OAI21X1_111
timestamp 1516325494
transform 1 0 3380 0 -1 2224
box 0 0 19 49
use AOI22X1  AOI22X1_28
timestamp 1516325494
transform 1 0 3399 0 -1 2224
box 0 0 23 49
use FILL  FILL_BUFX2_105
timestamp 1516325494
transform 1 0 3422 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_105
timestamp 1516325494
transform 1 0 3430 0 -1 2224
box 0 0 15 49
use FILL  FILL_BUFX2_265
timestamp 1516325494
transform -1 0 3453 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_265
timestamp 1516325494
transform -1 0 3467 0 -1 2224
box 0 0 15 49
use NAND2X1  NAND2X1_429
timestamp 1516325494
transform -1 0 1678 0 1 2126
box 0 0 15 49
use OR2X2  OR2X2_1387
timestamp 1516325494
transform 1 0 1678 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_327
timestamp 1516325494
transform -1 0 1716 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1810
timestamp 1516325494
transform 1 0 1716 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1811
timestamp 1516325494
transform -1 0 1754 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_349
timestamp 1516325494
transform -1 0 1773 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1916
timestamp 1516325494
transform -1 0 1792 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1915
timestamp 1516325494
transform -1 0 1811 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1806
timestamp 1516325494
transform -1 0 1830 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1913
timestamp 1516325494
transform 1 0 1830 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_348
timestamp 1516325494
transform -1 0 1868 0 1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_727
timestamp 1516325494
transform 1 0 1868 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_727
timestamp 1516325494
transform 1 0 1875 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_805
timestamp 1516325494
transform 1 0 903 0 -1 2126
box 0 0 30 49
use INVX1  INVX1_227
timestamp 1516325494
transform -1 0 944 0 -1 2126
box 0 0 11 49
use FILL  FILL_AND2X2_263
timestamp 1516325494
transform 1 0 944 0 -1 2126
box 0 0 8 49
use AND2X2  AND2X2_263
timestamp 1516325494
transform 1 0 952 0 -1 2126
box 0 0 19 49
use FILL  FILL_OR2X2_246
timestamp 1516325494
transform 1 0 971 0 -1 2126
box 0 0 8 49
use OR2X2  OR2X2_246
timestamp 1516325494
transform 1 0 979 0 -1 2126
box 0 0 19 49
use FILL  FILL_OR2X2_247
timestamp 1516325494
transform 1 0 998 0 -1 2126
box 0 0 8 49
use OR2X2  OR2X2_247
timestamp 1516325494
transform 1 0 1005 0 -1 2126
box 0 0 19 49
use MUX2X1  MUX2X1_785
timestamp 1516325494
transform 1 0 1024 0 -1 2126
box 0 0 30 49
use AND2X2  AND2X2_1784
timestamp 1516325494
transform -1 0 1074 0 -1 2126
box 0 0 19 49
use FILL  FILL_OR2X2_245
timestamp 1516325494
transform -1 0 1082 0 -1 2126
box 0 0 8 49
use OR2X2  OR2X2_245
timestamp 1516325494
transform -1 0 1100 0 -1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_261
timestamp 1516325494
transform -1 0 1108 0 -1 2126
box 0 0 8 49
use AND2X2  AND2X2_261
timestamp 1516325494
transform -1 0 1127 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_142
timestamp 1516325494
transform 1 0 1127 0 -1 2126
box 0 0 15 49
use FILL  FILL_AND2X2_262
timestamp 1516325494
transform 1 0 1142 0 -1 2126
box 0 0 8 49
use AND2X2  AND2X2_262
timestamp 1516325494
transform 1 0 1150 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1425
timestamp 1516325494
transform 1 0 1169 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1853
timestamp 1516325494
transform 1 0 1188 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1854
timestamp 1516325494
transform -1 0 1226 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1321
timestamp 1516325494
transform -1 0 1245 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1035
timestamp 1516325494
transform -1 0 1264 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_346
timestamp 1516325494
transform 1 0 1264 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_347
timestamp 1516325494
transform -1 0 1302 0 -1 2126
box 0 0 19 49
use INVX1  INVX1_142
timestamp 1516325494
transform 1 0 1302 0 -1 2126
box 0 0 11 49
use AND2X2  AND2X2_412
timestamp 1516325494
transform 1 0 1313 0 -1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_323
timestamp 1516325494
transform 1 0 1332 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_323
timestamp 1516325494
transform 1 0 1340 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_385
timestamp 1516325494
transform 1 0 1355 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_385
timestamp 1516325494
transform 1 0 1362 0 -1 2126
box 0 0 15 49
use OAI21X1  OAI21X1_31
timestamp 1516325494
transform 1 0 1378 0 -1 2126
box 0 0 19 49
use INVX2  INVX2_20
timestamp 1516325494
transform 1 0 1397 0 -1 2126
box 0 0 11 49
use AND2X2  AND2X2_2007
timestamp 1516325494
transform -1 0 1427 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1927
timestamp 1516325494
transform -1 0 1446 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1926
timestamp 1516325494
transform -1 0 1465 0 -1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_384
timestamp 1516325494
transform -1 0 1473 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_384
timestamp 1516325494
transform -1 0 1488 0 -1 2126
box 0 0 15 49
use OR2X2  OR2X2_1939
timestamp 1516325494
transform -1 0 1507 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_511
timestamp 1516325494
transform 1 0 1507 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_575
timestamp 1516325494
transform 1 0 1560 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_575
timestamp 1516325494
transform -1 0 1605 0 -1 2126
box 0 0 30 49
use FILL  FILL_BUFX2_433
timestamp 1516325494
transform -1 0 1614 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_433
timestamp 1516325494
transform -1 0 1628 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_639
timestamp 1516325494
transform 1 0 1628 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_909
timestamp 1516325494
transform 1 0 1682 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_854
timestamp 1516325494
transform -1 0 1727 0 -1 2126
box 0 0 30 49
use FILL  FILL_BUFX2_325
timestamp 1516325494
transform -1 0 1735 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_325
timestamp 1516325494
transform -1 0 1750 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_41
timestamp 1516325494
transform 1 0 1750 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_41
timestamp 1516325494
transform 1 0 1758 0 -1 2126
box 0 0 15 49
use OR2X2  OR2X2_1804
timestamp 1516325494
transform 1 0 1773 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_635
timestamp 1516325494
transform 1 0 1792 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_905
timestamp 1516325494
transform 1 0 1845 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_850
timestamp 1516325494
transform -1 0 1890 0 -1 2126
box 0 0 30 49
use INVX1  INVX1_206
timestamp 1516325494
transform 1 0 1891 0 1 2126
box 0 0 11 49
use FILL  FILL_OR2X2_25
timestamp 1516325494
transform 1 0 1902 0 1 2126
box 0 0 8 49
use OR2X2  OR2X2_25
timestamp 1516325494
transform 1 0 1910 0 1 2126
box 0 0 19 49
use INVX1  INVX1_204
timestamp 1516325494
transform -1 0 1940 0 1 2126
box 0 0 11 49
use AND2X2  AND2X2_1914
timestamp 1516325494
transform 1 0 1940 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1805
timestamp 1516325494
transform -1 0 1978 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1912
timestamp 1516325494
transform -1 0 1997 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_20
timestamp 1516325494
transform -1 0 2005 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_20
timestamp 1516325494
transform -1 0 2024 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1412
timestamp 1516325494
transform -1 0 2043 0 1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_60
timestamp 1516325494
transform 1 0 2043 0 1 2126
box 0 0 53 49
use MUX2X1  MUX2X1_444
timestamp 1516325494
transform -1 0 2126 0 1 2126
box 0 0 30 49
use AND2X2  AND2X2_1406
timestamp 1516325494
transform -1 0 2145 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_17
timestamp 1516325494
transform -1 0 2153 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_17
timestamp 1516325494
transform -1 0 2172 0 1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_613
timestamp 1516325494
transform -1 0 2225 0 1 2126
box 0 0 53 49
use FILL  FILL_BUFX2_729
timestamp 1516325494
transform 1 0 2225 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_729
timestamp 1516325494
transform 1 0 2233 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_234
timestamp 1516325494
transform 1 0 2248 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_234
timestamp 1516325494
transform 1 0 2255 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_178
timestamp 1516325494
transform -1 0 2279 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_178
timestamp 1516325494
transform -1 0 2293 0 1 2126
box 0 0 15 49
use AND2X2  AND2X2_1911
timestamp 1516325494
transform -1 0 2312 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1801
timestamp 1516325494
transform -1 0 2331 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1825
timestamp 1516325494
transform -1 0 2350 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1688
timestamp 1516325494
transform -1 0 2369 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1689
timestamp 1516325494
transform -1 0 2388 0 1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_311
timestamp 1516325494
transform 1 0 2388 0 1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_503
timestamp 1516325494
transform 1 0 2442 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_503
timestamp 1516325494
transform -1 0 2487 0 1 2126
box 0 0 30 49
use OR2X2  OR2X2_1682
timestamp 1516325494
transform -1 0 2506 0 1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_663
timestamp 1516325494
transform 1 0 2506 0 1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_55
timestamp 1516325494
transform 1 0 2559 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_55
timestamp 1516325494
transform -1 0 2605 0 1 2126
box 0 0 30 49
use FILL  FILL_OR2X2_17
timestamp 1516325494
transform -1 0 2613 0 1 2126
box 0 0 8 49
use OR2X2  OR2X2_17
timestamp 1516325494
transform -1 0 2632 0 1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_442
timestamp 1516325494
transform 1 0 2632 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_442
timestamp 1516325494
transform 1 0 2639 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_728
timestamp 1516325494
transform -1 0 2662 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_728
timestamp 1516325494
transform -1 0 2677 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_42
timestamp 1516325494
transform -1 0 2685 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_42
timestamp 1516325494
transform -1 0 2700 0 1 2126
box 0 0 15 49
use OR2X2  OR2X2_325
timestamp 1516325494
transform -1 0 2719 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_322
timestamp 1516325494
transform -1 0 2738 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_320
timestamp 1516325494
transform -1 0 2757 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_341
timestamp 1516325494
transform -1 0 2776 0 1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_231
timestamp 1516325494
transform -1 0 2829 0 1 2126
box 0 0 53 49
use OR2X2  OR2X2_324
timestamp 1516325494
transform -1 0 2848 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_344
timestamp 1516325494
transform -1 0 2867 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_323
timestamp 1516325494
transform -1 0 2886 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_345
timestamp 1516325494
transform -1 0 2905 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1816
timestamp 1516325494
transform 1 0 2905 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_1678
timestamp 1516325494
transform -1 0 2943 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1817
timestamp 1516325494
transform -1 0 2962 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1818
timestamp 1516325494
transform -1 0 2981 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_283
timestamp 1516325494
transform 1 0 2981 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_283
timestamp 1516325494
transform -1 0 3026 0 1 2126
box 0 0 30 49
use FILL  FILL_OR2X2_16
timestamp 1516325494
transform -1 0 3035 0 1 2126
box 0 0 8 49
use OR2X2  OR2X2_16
timestamp 1516325494
transform -1 0 3053 0 1 2126
box 0 0 19 49
use FILL  FILL_OR2X2_15
timestamp 1516325494
transform -1 0 3061 0 1 2126
box 0 0 8 49
use OR2X2  OR2X2_15
timestamp 1516325494
transform -1 0 3080 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_61
timestamp 1516325494
transform 1 0 3080 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_61
timestamp 1516325494
transform 1 0 3088 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_15
timestamp 1516325494
transform -1 0 3115 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_15
timestamp 1516325494
transform -1 0 3133 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_46
timestamp 1516325494
transform 1 0 3133 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_46
timestamp 1516325494
transform 1 0 3141 0 1 2126
box 0 0 19 49
use FILL  FILL_OR2X2_43
timestamp 1516325494
transform -1 0 3168 0 1 2126
box 0 0 8 49
use OR2X2  OR2X2_43
timestamp 1516325494
transform -1 0 3186 0 1 2126
box 0 0 19 49
use FILL  FILL_AND2X2_45
timestamp 1516325494
transform -1 0 3194 0 1 2126
box 0 0 8 49
use AND2X2  AND2X2_45
timestamp 1516325494
transform -1 0 3213 0 1 2126
box 0 0 19 49
use OR2X2  OR2X2_960
timestamp 1516325494
transform 1 0 3213 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1209
timestamp 1516325494
transform 1 0 3232 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1199
timestamp 1516325494
transform 1 0 3251 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1202
timestamp 1516325494
transform 1 0 3270 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1211
timestamp 1516325494
transform 1 0 3289 0 1 2126
box 0 0 19 49
use AOI22X1  AOI22X1_30
timestamp 1516325494
transform -1 0 3331 0 1 2126
box 0 0 23 49
use OAI21X1  OAI21X1_116
timestamp 1516325494
transform 1 0 3331 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_831
timestamp 1516325494
transform -1 0 3365 0 1 2126
box 0 0 15 49
use AND2X2  AND2X2_1242
timestamp 1516325494
transform 1 0 3365 0 1 2126
box 0 0 19 49
use INVX1  INVX1_274
timestamp 1516325494
transform 1 0 3384 0 1 2126
box 0 0 11 49
use OR2X2  OR2X2_978
timestamp 1516325494
transform -1 0 3414 0 1 2126
box 0 0 19 49
use AND2X2  AND2X2_1223
timestamp 1516325494
transform -1 0 3433 0 1 2126
box 0 0 19 49
use NAND3X1  NAND3X1_90
timestamp 1516325494
transform -1 0 3452 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_799
timestamp 1516325494
transform -1 0 3467 0 1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_406
timestamp 1516325494
transform 1 0 3468 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_406
timestamp 1516325494
transform 1 0 3475 0 -1 2224
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_793
timestamp 1516325494
transform 1 0 3490 0 -1 2224
box 0 0 53 49
use AND2X2  AND2X2_1191
timestamp 1516325494
transform -1 0 3563 0 -1 2224
box 0 0 19 49
use FILL  FILL_BUFX2_267
timestamp 1516325494
transform -1 0 3571 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_267
timestamp 1516325494
transform -1 0 3585 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_983
timestamp 1516325494
transform -1 0 3604 0 -1 2224
box 0 0 19 49
use AOI22X1  AOI22X1_23
timestamp 1516325494
transform -1 0 3627 0 -1 2224
box 0 0 23 49
use FILL  FILL_BUFX2_402
timestamp 1516325494
transform 1 0 3627 0 -1 2224
box 0 0 8 49
use BUFX2  BUFX2_402
timestamp 1516325494
transform 1 0 3635 0 -1 2224
box 0 0 15 49
use NAND2X1  NAND2X1_841
timestamp 1516325494
transform 1 0 3650 0 -1 2224
box 0 0 15 49
use OAI21X1  OAI21X1_127
timestamp 1516325494
transform -1 0 3684 0 -1 2224
box 0 0 19 49
use OAI21X1  OAI21X1_105
timestamp 1516325494
transform 1 0 3684 0 -1 2224
box 0 0 19 49
use NAND2X1  NAND2X1_816
timestamp 1516325494
transform 1 0 3703 0 -1 2224
box 0 0 15 49
use OAI21X1  OAI21X1_106
timestamp 1516325494
transform 1 0 3718 0 -1 2224
box 0 0 19 49
use AOI22X1  AOI22X1_24
timestamp 1516325494
transform -1 0 3760 0 -1 2224
box 0 0 23 49
use MUX2X1  MUX2X1_814
timestamp 1516325494
transform 1 0 3760 0 -1 2224
box 0 0 30 49
use NAND2X1  NAND2X1_815
timestamp 1516325494
transform 1 0 3791 0 -1 2224
box 0 0 15 49
use OR2X2  OR2X2_974
timestamp 1516325494
transform 1 0 3806 0 -1 2224
box 0 0 19 49
use NAND3X1  NAND3X1_92
timestamp 1516325494
transform 1 0 3825 0 -1 2224
box 0 0 19 49
use AND2X2  AND2X2_1334
timestamp 1516325494
transform 1 0 3844 0 -1 2224
box 0 0 19 49
use FILL  FILL_45_1
timestamp 1516325494
transform -1 0 3871 0 -1 2224
box 0 0 8 49
use OAI21X1  OAI21X1_99
timestamp 1516325494
transform -1 0 3487 0 1 2126
box 0 0 19 49
use AOI22X1  AOI22X1_18
timestamp 1516325494
transform 1 0 3487 0 1 2126
box 0 0 23 49
use NAND2X1  NAND2X1_802
timestamp 1516325494
transform -1 0 3524 0 1 2126
box 0 0 15 49
use AND2X2  AND2X2_1917
timestamp 1516325494
transform -1 0 1910 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1807
timestamp 1516325494
transform -1 0 1929 0 -1 2126
box 0 0 19 49
use MUX2X1  MUX2X1_782
timestamp 1516325494
transform 1 0 1929 0 -1 2126
box 0 0 30 49
use MUX2X1  MUX2X1_784
timestamp 1516325494
transform 1 0 1959 0 -1 2126
box 0 0 30 49
use OR2X2  OR2X2_1837
timestamp 1516325494
transform -1 0 2008 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_424
timestamp 1516325494
transform 1 0 2008 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_40
timestamp 1516325494
transform 1 0 2024 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_444
timestamp 1516325494
transform 1 0 2077 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_424
timestamp 1516325494
transform -1 0 2122 0 -1 2126
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_59
timestamp 1516325494
transform 1 0 2122 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_443
timestamp 1516325494
transform 1 0 2176 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_443
timestamp 1516325494
transform -1 0 2221 0 -1 2126
box 0 0 30 49
use OR2X2  OR2X2_1808
timestamp 1516325494
transform -1 0 2240 0 -1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_516
timestamp 1516325494
transform -1 0 2248 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_516
timestamp 1516325494
transform -1 0 2263 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_27
timestamp 1516325494
transform 1 0 2263 0 -1 2126
box 0 0 30 49
use NAND2X1  NAND2X1_27
timestamp 1516325494
transform -1 0 2308 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_603
timestamp 1516325494
transform -1 0 2362 0 -1 2126
box 0 0 53 49
use OR2X2  OR2X2_1802
timestamp 1516325494
transform -1 0 2381 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_443
timestamp 1516325494
transform 1 0 2381 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_411
timestamp 1516325494
transform 1 0 2434 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_411
timestamp 1516325494
transform -1 0 2479 0 -1 2126
box 0 0 30 49
use MUX2X1  MUX2X1_407
timestamp 1516325494
transform 1 0 2480 0 -1 2126
box 0 0 30 49
use NAND2X1  NAND2X1_407
timestamp 1516325494
transform -1 0 2525 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_667
timestamp 1516325494
transform 1 0 2525 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_59
timestamp 1516325494
transform 1 0 2578 0 -1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_59
timestamp 1516325494
transform -1 0 2624 0 -1 2126
box 0 0 30 49
use OR2X2  OR2X2_1800
timestamp 1516325494
transform -1 0 2643 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1797
timestamp 1516325494
transform -1 0 2662 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1795
timestamp 1516325494
transform -1 0 2681 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_251
timestamp 1516325494
transform 1 0 2681 0 -1 2126
box 0 0 53 49
use AND2X2  AND2X2_1905
timestamp 1516325494
transform -1 0 2753 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_219
timestamp 1516325494
transform 1 0 2753 0 -1 2126
box 0 0 53 49
use MUX2X1  MUX2X1_751
timestamp 1516325494
transform -1 0 2836 0 -1 2126
box 0 0 30 49
use OR2X2  OR2X2_268
timestamp 1516325494
transform -1 0 2856 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_284
timestamp 1516325494
transform -1 0 2875 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1799
timestamp 1516325494
transform -1 0 2894 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1908
timestamp 1516325494
transform -1 0 2913 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1798
timestamp 1516325494
transform -1 0 2932 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1909
timestamp 1516325494
transform -1 0 2951 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_267
timestamp 1516325494
transform -1 0 2970 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_286
timestamp 1516325494
transform -1 0 2989 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_151
timestamp 1516325494
transform 1 0 2989 0 -1 2126
box 0 0 53 49
use FILL  FILL_AND2X2_16
timestamp 1516325494
transform 1 0 3042 0 -1 2126
box 0 0 8 49
use AND2X2  AND2X2_16
timestamp 1516325494
transform 1 0 3050 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1404
timestamp 1516325494
transform 1 0 3069 0 -1 2126
box 0 0 19 49
use OR2X2  OR2X2_1138
timestamp 1516325494
transform -1 0 3107 0 -1 2126
box 0 0 19 49
use AND2X2  AND2X2_1403
timestamp 1516325494
transform -1 0 3126 0 -1 2126
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_133
timestamp 1516325494
transform -1 0 3179 0 -1 2126
box 0 0 53 49
use INVX2  INVX2_6
timestamp 1516325494
transform -1 0 3190 0 -1 2126
box 0 0 11 49
use AND2X2  AND2X2_1204
timestamp 1516325494
transform -1 0 3209 0 -1 2126
box 0 0 19 49
use XOR2X1  XOR2X1_70
timestamp 1516325494
transform -1 0 3243 0 -1 2126
box 0 0 34 49
use XOR2X1  XOR2X1_72
timestamp 1516325494
transform 1 0 3243 0 -1 2126
box 0 0 34 49
use DFFPOSX1  DFFPOSX1_831
timestamp 1516325494
transform 1 0 3278 0 -1 2126
box 0 0 53 49
use OAI21X1  OAI21X1_117
timestamp 1516325494
transform -1 0 3350 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_830
timestamp 1516325494
transform -1 0 3365 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_307
timestamp 1516325494
transform -1 0 3373 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_307
timestamp 1516325494
transform -1 0 3388 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_808
timestamp 1516325494
transform -1 0 3441 0 -1 2126
box 0 0 53 49
use NAND2X1  NAND2X1_800
timestamp 1516325494
transform -1 0 3456 0 -1 2126
box 0 0 15 49
use AND2X2  AND2X2_1214
timestamp 1516325494
transform -1 0 3475 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_798
timestamp 1516325494
transform -1 0 3490 0 -1 2126
box 0 0 15 49
use AOI21X1  AOI21X1_59
timestamp 1516325494
transform 1 0 3490 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_801
timestamp 1516325494
transform 1 0 3509 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_691
timestamp 1516325494
transform -1 0 3533 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_691
timestamp 1516325494
transform -1 0 3547 0 1 2126
box 0 0 15 49
use NOR3X1  NOR3X1_30
timestamp 1516325494
transform -1 0 3566 0 1 2126
box 0 0 19 49
use OAI21X1  OAI21X1_100
timestamp 1516325494
transform -1 0 3585 0 1 2126
box 0 0 19 49
use NOR2X1  NOR2X1_142
timestamp 1516325494
transform 1 0 3585 0 1 2126
box 0 0 15 49
use XNOR2X1  XNOR2X1_59
timestamp 1516325494
transform 1 0 3601 0 1 2126
box 0 0 34 49
use AND2X2  AND2X2_1224
timestamp 1516325494
transform 1 0 3635 0 1 2126
box 0 0 19 49
use FILL  FILL_BUFX2_489
timestamp 1516325494
transform -1 0 3662 0 1 2126
box 0 0 8 49
use BUFX2  BUFX2_489
timestamp 1516325494
transform -1 0 3676 0 1 2126
box 0 0 15 49
use INVX1  INVX1_286
timestamp 1516325494
transform 1 0 3677 0 1 2126
box 0 0 11 49
use AOI22X1  AOI22X1_14
timestamp 1516325494
transform 1 0 3688 0 1 2126
box 0 0 23 49
use INVX1  INVX1_282
timestamp 1516325494
transform -1 0 3722 0 1 2126
box 0 0 11 49
use NAND3X1  NAND3X1_83
timestamp 1516325494
transform 1 0 3722 0 1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_781
timestamp 1516325494
transform -1 0 3756 0 1 2126
box 0 0 15 49
use MUX2X1  MUX2X1_822
timestamp 1516325494
transform 1 0 3756 0 1 2126
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_811
timestamp 1516325494
transform 1 0 3787 0 1 2126
box 0 0 53 49
use AND2X2  AND2X2_1233
timestamp 1516325494
transform 1 0 3840 0 1 2126
box 0 0 19 49
use FILL  FILL_44_1
timestamp 1516325494
transform 1 0 3859 0 1 2126
box 0 0 8 49
use OAI21X1  OAI21X1_118
timestamp 1516325494
transform 1 0 3525 0 -1 2126
box 0 0 19 49
use OAI21X1  OAI21X1_119
timestamp 1516325494
transform 1 0 3544 0 -1 2126
box 0 0 19 49
use AOI22X1  AOI22X1_31
timestamp 1516325494
transform 1 0 3563 0 -1 2126
box 0 0 23 49
use AND2X2  AND2X2_1243
timestamp 1516325494
transform -1 0 3604 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_832
timestamp 1516325494
transform 1 0 3604 0 -1 2126
box 0 0 15 49
use NAND2X1  NAND2X1_833
timestamp 1516325494
transform 1 0 3620 0 -1 2126
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_832
timestamp 1516325494
transform -1 0 3688 0 -1 2126
box 0 0 53 49
use FILL  FILL_BUFX2_258
timestamp 1516325494
transform 1 0 3688 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_258
timestamp 1516325494
transform 1 0 3696 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_260
timestamp 1516325494
transform -1 0 3719 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_260
timestamp 1516325494
transform -1 0 3733 0 -1 2126
box 0 0 15 49
use FILL  FILL_BUFX2_306
timestamp 1516325494
transform -1 0 3742 0 -1 2126
box 0 0 8 49
use BUFX2  BUFX2_306
timestamp 1516325494
transform -1 0 3756 0 -1 2126
box 0 0 15 49
use AND2X2  AND2X2_1210
timestamp 1516325494
transform -1 0 3775 0 -1 2126
box 0 0 19 49
use OAI21X1  OAI21X1_134
timestamp 1516325494
transform 1 0 3775 0 -1 2126
box 0 0 19 49
use OAI21X1  OAI21X1_135
timestamp 1516325494
transform 1 0 3794 0 -1 2126
box 0 0 19 49
use NAND2X1  NAND2X1_844
timestamp 1516325494
transform -1 0 3828 0 -1 2126
box 0 0 15 49
use INVX1  INVX1_317
timestamp 1516325494
transform -1 0 3840 0 -1 2126
box 0 0 11 49
use NOR2X1  NOR2X1_157
timestamp 1516325494
transform -1 0 3855 0 -1 2126
box 0 0 15 49
use FILL  FILL_43_1
timestamp 1516325494
transform -1 0 3863 0 -1 2126
box 0 0 8 49
use FILL  FILL_43_2
timestamp 1516325494
transform -1 0 3871 0 -1 2126
box 0 0 8 49
use OR2X2  OR2X2_896
timestamp 1516325494
transform -1 0 21 0 1 2027
box 0 0 19 49
use XNOR2X1  XNOR2X1_26
timestamp 1516325494
transform -1 0 55 0 1 2027
box 0 0 34 49
use INVX1  INVX1_90
timestamp 1516325494
transform -1 0 66 0 1 2027
box 0 0 11 49
use AND2X2  AND2X2_1100
timestamp 1516325494
transform 1 0 2 0 -1 2027
box 0 0 19 49
use INVX1  INVX1_89
timestamp 1516325494
transform -1 0 32 0 -1 2027
box 0 0 11 49
use XOR2X1  XOR2X1_46
timestamp 1516325494
transform 1 0 32 0 -1 2027
box 0 0 34 49
use XNOR2X1  XNOR2X1_18
timestamp 1516325494
transform -1 0 101 0 1 2027
box 0 0 34 49
use NOR2X1  NOR2X1_52
timestamp 1516325494
transform 1 0 101 0 1 2027
box 0 0 15 49
use OR2X2  OR2X2_745
timestamp 1516325494
transform 1 0 116 0 1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_642
timestamp 1516325494
transform 1 0 135 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_642
timestamp 1516325494
transform 1 0 143 0 1 2027
box 0 0 15 49
use AOI21X1  AOI21X1_15
timestamp 1516325494
transform -1 0 177 0 1 2027
box 0 0 19 49
use XOR2X1  XOR2X1_50
timestamp 1516325494
transform 1 0 177 0 1 2027
box 0 0 34 49
use OR2X2  OR2X2_900
timestamp 1516325494
transform 1 0 211 0 1 2027
box 0 0 19 49
use INVX1  INVX1_102
timestamp 1516325494
transform -1 0 241 0 1 2027
box 0 0 11 49
use OR2X2  OR2X2_696
timestamp 1516325494
transform 1 0 241 0 1 2027
box 0 0 19 49
use OAI21X1  OAI21X1_11
timestamp 1516325494
transform -1 0 279 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1105
timestamp 1516325494
transform 1 0 279 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_827
timestamp 1516325494
transform -1 0 317 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_698
timestamp 1516325494
transform -1 0 336 0 1 2027
box 0 0 19 49
use NOR2X1  NOR2X1_42
timestamp 1516325494
transform -1 0 351 0 1 2027
box 0 0 15 49
use AND2X2  AND2X2_826
timestamp 1516325494
transform -1 0 371 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_668
timestamp 1516325494
transform -1 0 386 0 1 2027
box 0 0 15 49
use OR2X2  OR2X2_823
timestamp 1516325494
transform 1 0 386 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_941
timestamp 1516325494
transform -1 0 424 0 1 2027
box 0 0 19 49
use NAND3X1  NAND3X1_52
timestamp 1516325494
transform -1 0 443 0 1 2027
box 0 0 19 49
use NAND3X1  NAND3X1_51
timestamp 1516325494
transform -1 0 462 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_684
timestamp 1516325494
transform 1 0 462 0 1 2027
box 0 0 15 49
use XNOR2X1  XNOR2X1_36
timestamp 1516325494
transform -1 0 511 0 1 2027
box 0 0 34 49
use INVX1  INVX1_47
timestamp 1516325494
transform 1 0 511 0 1 2027
box 0 0 11 49
use AND2X2  AND2X2_1069
timestamp 1516325494
transform -1 0 542 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1071
timestamp 1516325494
transform 1 0 542 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_797
timestamp 1516325494
transform -1 0 580 0 1 2027
box 0 0 19 49
use MUX2X1  MUX2X1_772
timestamp 1516325494
transform 1 0 580 0 1 2027
box 0 0 30 49
use FILL  FILL_BUFX2_781
timestamp 1516325494
transform -1 0 618 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_781
timestamp 1516325494
transform -1 0 633 0 1 2027
box 0 0 15 49
use INVX1  INVX1_31
timestamp 1516325494
transform 1 0 633 0 1 2027
box 0 0 11 49
use INVX1  INVX1_160
timestamp 1516325494
transform 1 0 644 0 1 2027
box 0 0 11 49
use MUX2X1  MUX2X1_803
timestamp 1516325494
transform -1 0 686 0 1 2027
box 0 0 30 49
use INVX1  INVX1_225
timestamp 1516325494
transform -1 0 697 0 1 2027
box 0 0 11 49
use FILL  FILL_BUFX2_317
timestamp 1516325494
transform 1 0 697 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_317
timestamp 1516325494
transform 1 0 705 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_21
timestamp 1516325494
transform 1 0 720 0 1 2027
box 0 0 53 49
use INVX1  INVX1_165
timestamp 1516325494
transform 1 0 773 0 1 2027
box 0 0 11 49
use MUX2X1  MUX2X1_795
timestamp 1516325494
transform 1 0 785 0 1 2027
box 0 0 30 49
use MUX2X1  MUX2X1_309
timestamp 1516325494
transform 1 0 815 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_309
timestamp 1516325494
transform -1 0 861 0 1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_335
timestamp 1516325494
transform 1 0 861 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_335
timestamp 1516325494
transform 1 0 868 0 1 2027
box 0 0 15 49
use INVX1  INVX1_155
timestamp 1516325494
transform 1 0 884 0 1 2027
box 0 0 11 49
use OR2X2  OR2X2_1642
timestamp 1516325494
transform -1 0 914 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1636
timestamp 1516325494
transform -1 0 933 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1782
timestamp 1516325494
transform -1 0 952 0 1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_589
timestamp 1516325494
transform 1 0 952 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_589
timestamp 1516325494
transform 1 0 960 0 1 2027
box 0 0 15 49
use FILL  FILL_OR2X2_62
timestamp 1516325494
transform -1 0 983 0 1 2027
box 0 0 8 49
use OR2X2  OR2X2_62
timestamp 1516325494
transform -1 0 1001 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_248
timestamp 1516325494
transform -1 0 1020 0 1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_605
timestamp 1516325494
transform 1 0 1020 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_605
timestamp 1516325494
transform 1 0 1028 0 1 2027
box 0 0 15 49
use OR2X2  OR2X2_1241
timestamp 1516325494
transform -1 0 1062 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1240
timestamp 1516325494
transform -1 0 1081 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_414
timestamp 1516325494
transform 1 0 1081 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1479
timestamp 1516325494
transform -1 0 1119 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_2018
timestamp 1516325494
transform 1 0 1119 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_2012
timestamp 1516325494
transform 1 0 1138 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1936
timestamp 1516325494
transform 1 0 1157 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_2014
timestamp 1516325494
transform -1 0 1195 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1841
timestamp 1516325494
transform -1 0 1214 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1840
timestamp 1516325494
transform -1 0 1233 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1939
timestamp 1516325494
transform -1 0 1252 0 1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_7
timestamp 1516325494
transform 1 0 1252 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_7
timestamp 1516325494
transform 1 0 1260 0 1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_362
timestamp 1516325494
transform 1 0 1275 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_362
timestamp 1516325494
transform 1 0 1283 0 1 2027
box 0 0 15 49
use OR2X2  OR2X2_342
timestamp 1516325494
transform -1 0 1317 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_2013
timestamp 1516325494
transform -1 0 1336 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1935
timestamp 1516325494
transform -1 0 1355 0 1 2027
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_95
timestamp 1516325494
transform 1 0 1355 0 1 2027
box 0 0 53 49
use AND2X2  AND2X2_2017
timestamp 1516325494
transform -1 0 1427 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_159
timestamp 1516325494
transform 1 0 1427 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_159
timestamp 1516325494
transform 1 0 1442 0 1 2027
box 0 0 30 49
use FILL  FILL_BUFX2_794
timestamp 1516325494
transform 1 0 1473 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_794
timestamp 1516325494
transform 1 0 1480 0 1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_65
timestamp 1516325494
transform 1 0 1495 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_65
timestamp 1516325494
transform 1 0 1503 0 1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_607
timestamp 1516325494
transform -1 0 1526 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_607
timestamp 1516325494
transform -1 0 1541 0 1 2027
box 0 0 15 49
use AND2X2  AND2X2_1918
timestamp 1516325494
transform -1 0 1560 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_350
timestamp 1516325494
transform 1 0 1560 0 1 2027
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_31
timestamp 1516325494
transform 1 0 1579 0 1 2027
box 0 0 53 49
use NAND2X1  NAND2X1_127
timestamp 1516325494
transform 1 0 1632 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_127
timestamp 1516325494
transform -1 0 1677 0 1 2027
box 0 0 30 49
use FILL  FILL_BUFX2_100
timestamp 1516325494
transform 1 0 1678 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_100
timestamp 1516325494
transform 1 0 1685 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_315
timestamp 1516325494
transform 1 0 1701 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_315
timestamp 1516325494
transform -1 0 1746 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_699
timestamp 1516325494
transform -1 0 1799 0 1 2027
box 0 0 53 49
use MUX2X1  MUX2X1_507
timestamp 1516325494
transform 1 0 1799 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_507
timestamp 1516325494
transform -1 0 1845 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_315
timestamp 1516325494
transform -1 0 1898 0 1 2027
box 0 0 53 49
use OR2X2  OR2X2_1809
timestamp 1516325494
transform 1 0 1898 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1478
timestamp 1516325494
transform -1 0 1936 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1237
timestamp 1516325494
transform -1 0 1955 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1236
timestamp 1516325494
transform -1 0 1974 0 1 2027
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_616
timestamp 1516325494
transform 1 0 1974 0 1 2027
box 0 0 53 49
use NAND2X1  NAND2X1_886
timestamp 1516325494
transform 1 0 2027 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_831
timestamp 1516325494
transform -1 0 2073 0 1 2027
box 0 0 30 49
use FILL  FILL_BUFX2_798
timestamp 1516325494
transform 1 0 2073 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_798
timestamp 1516325494
transform 1 0 2081 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_68
timestamp 1516325494
transform 1 0 2096 0 1 2027
box 0 0 53 49
use MUX2X1  MUX2X1_132
timestamp 1516325494
transform 1 0 2149 0 1 2027
box 0 0 30 49
use AND2X2  AND2X2_1781
timestamp 1516325494
transform -1 0 2198 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1632
timestamp 1516325494
transform -1 0 2217 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1633
timestamp 1516325494
transform -1 0 2236 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_931
timestamp 1516325494
transform 1 0 2236 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_373
timestamp 1516325494
transform 1 0 2252 0 1 2027
box 0 0 53 49
use MUX2X1  MUX2X1_876
timestamp 1516325494
transform -1 0 2335 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_181
timestamp 1516325494
transform 1 0 2335 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_405
timestamp 1516325494
transform 1 0 2350 0 1 2027
box 0 0 53 49
use MUX2X1  MUX2X1_181
timestamp 1516325494
transform -1 0 2434 0 1 2027
box 0 0 30 49
use OAI21X1  OAI21X1_48
timestamp 1516325494
transform 1 0 2434 0 1 2027
box 0 0 19 49
use INVX2  INVX2_37
timestamp 1516325494
transform 1 0 2453 0 1 2027
box 0 0 11 49
use FILL  FILL_BUFX2_5
timestamp 1516325494
transform -1 0 2472 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_5
timestamp 1516325494
transform -1 0 2487 0 1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_439
timestamp 1516325494
transform -1 0 2540 0 1 2027
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_444
timestamp 1516325494
transform 1 0 2540 0 1 2027
box 0 0 53 49
use AND2X2  AND2X2_343
timestamp 1516325494
transform 1 0 2594 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1907
timestamp 1516325494
transform 1 0 2613 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1796
timestamp 1516325494
transform 1 0 2632 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1906
timestamp 1516325494
transform -1 0 2670 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_321
timestamp 1516325494
transform 1 0 2670 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_342
timestamp 1516325494
transform -1 0 2708 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_219
timestamp 1516325494
transform 1 0 2708 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_219
timestamp 1516325494
transform -1 0 2753 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_635
timestamp 1516325494
transform 1 0 2753 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_635
timestamp 1516325494
transform -1 0 2798 0 1 2027
box 0 0 30 49
use INVX1  INVX1_79
timestamp 1516325494
transform -1 0 78 0 -1 2027
box 0 0 11 49
use NOR2X1  NOR2X1_87
timestamp 1516325494
transform -1 0 93 0 -1 2027
box 0 0 15 49
use XNOR2X1  XNOR2X1_19
timestamp 1516325494
transform 1 0 93 0 -1 2027
box 0 0 34 49
use NOR2X1  NOR2X1_54
timestamp 1516325494
transform -1 0 142 0 -1 2027
box 0 0 15 49
use NOR2X1  NOR2X1_58
timestamp 1516325494
transform 1 0 143 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_676
timestamp 1516325494
transform 1 0 158 0 -1 2027
box 0 0 15 49
use XOR2X1  XOR2X1_13
timestamp 1516325494
transform 1 0 173 0 -1 2027
box 0 0 34 49
use NAND2X1  NAND2X1_677
timestamp 1516325494
transform 1 0 207 0 -1 2027
box 0 0 15 49
use AND2X2  AND2X2_887
timestamp 1516325494
transform 1 0 222 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_888
timestamp 1516325494
transform 1 0 241 0 -1 2027
box 0 0 19 49
use XNOR2X1  XNOR2X1_35
timestamp 1516325494
transform -1 0 294 0 -1 2027
box 0 0 34 49
use INVX1  INVX1_103
timestamp 1516325494
transform 1 0 295 0 -1 2027
box 0 0 11 49
use NOR2X1  NOR2X1_95
timestamp 1516325494
transform 1 0 306 0 -1 2027
box 0 0 15 49
use INVX1  INVX1_104
timestamp 1516325494
transform 1 0 321 0 -1 2027
box 0 0 11 49
use AND2X2  AND2X2_828
timestamp 1516325494
transform 1 0 333 0 -1 2027
box 0 0 19 49
use NOR2X1  NOR2X1_74
timestamp 1516325494
transform 1 0 352 0 -1 2027
box 0 0 15 49
use NOR2X1  NOR2X1_60
timestamp 1516325494
transform 1 0 367 0 -1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_788
timestamp 1516325494
transform -1 0 390 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_788
timestamp 1516325494
transform -1 0 405 0 -1 2027
box 0 0 15 49
use AND2X2  AND2X2_942
timestamp 1516325494
transform -1 0 424 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_782
timestamp 1516325494
transform 1 0 424 0 -1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_641
timestamp 1516325494
transform -1 0 451 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_641
timestamp 1516325494
transform -1 0 465 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_685
timestamp 1516325494
transform -1 0 481 0 -1 2027
box 0 0 15 49
use NOR2X1  NOR2X1_78
timestamp 1516325494
transform 1 0 481 0 -1 2027
box 0 0 15 49
use AOI21X1  AOI21X1_18
timestamp 1516325494
transform 1 0 496 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_787
timestamp 1516325494
transform -1 0 534 0 -1 2027
box 0 0 19 49
use NOR2X1  NOR2X1_63
timestamp 1516325494
transform -1 0 549 0 -1 2027
box 0 0 15 49
use OR2X2  OR2X2_813
timestamp 1516325494
transform -1 0 568 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1072
timestamp 1516325494
transform 1 0 568 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1074
timestamp 1516325494
transform 1 0 587 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1075
timestamp 1516325494
transform 1 0 606 0 -1 2027
box 0 0 19 49
use OAI21X1  OAI21X1_70
timestamp 1516325494
transform -1 0 644 0 -1 2027
box 0 0 19 49
use OAI21X1  OAI21X1_75
timestamp 1516325494
transform -1 0 663 0 -1 2027
box 0 0 19 49
use INVX1  INVX1_188
timestamp 1516325494
transform -1 0 674 0 -1 2027
box 0 0 11 49
use OAI21X1  OAI21X1_72
timestamp 1516325494
transform -1 0 694 0 -1 2027
box 0 0 19 49
use INVX1  INVX1_41
timestamp 1516325494
transform 1 0 694 0 -1 2027
box 0 0 11 49
use FILL  FILL_BUFX2_851
timestamp 1516325494
transform -1 0 713 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_851
timestamp 1516325494
transform -1 0 728 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_739
timestamp 1516325494
transform -1 0 781 0 -1 2027
box 0 0 53 49
use MUX2X1  MUX2X1_808
timestamp 1516325494
transform -1 0 811 0 -1 2027
box 0 0 30 49
use INVX1  INVX1_230
timestamp 1516325494
transform -1 0 822 0 -1 2027
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_693
timestamp 1516325494
transform -1 0 876 0 -1 2027
box 0 0 53 49
use INVX1  INVX1_152
timestamp 1516325494
transform -1 0 887 0 -1 2027
box 0 0 11 49
use MUX2X1  MUX2X1_767
timestamp 1516325494
transform 1 0 887 0 -1 2027
box 0 0 30 49
use INVX1  INVX1_217
timestamp 1516325494
transform -1 0 929 0 -1 2027
box 0 0 11 49
use OR2X2  OR2X2_1624
timestamp 1516325494
transform 1 0 929 0 -1 2027
box 0 0 19 49
use MUX2X1  MUX2X1_798
timestamp 1516325494
transform -1 0 978 0 -1 2027
box 0 0 30 49
use INVX1  INVX1_220
timestamp 1516325494
transform -1 0 990 0 -1 2027
box 0 0 11 49
use OR2X2  OR2X2_249
timestamp 1516325494
transform -1 0 1009 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1644
timestamp 1516325494
transform -1 0 1028 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1643
timestamp 1516325494
transform -1 0 1047 0 -1 2027
box 0 0 19 49
use FILL  FILL_OR2X2_60
timestamp 1516325494
transform -1 0 1055 0 -1 2027
box 0 0 8 49
use OR2X2  OR2X2_60
timestamp 1516325494
transform -1 0 1074 0 -1 2027
box 0 0 19 49
use FILL  FILL_OR2X2_61
timestamp 1516325494
transform -1 0 1082 0 -1 2027
box 0 0 8 49
use OR2X2  OR2X2_61
timestamp 1516325494
transform -1 0 1100 0 -1 2027
box 0 0 19 49
use FILL  FILL_AND2X2_64
timestamp 1516325494
transform -1 0 1108 0 -1 2027
box 0 0 8 49
use AND2X2  AND2X2_64
timestamp 1516325494
transform -1 0 1127 0 -1 2027
box 0 0 19 49
use FILL  FILL_AND2X2_65
timestamp 1516325494
transform -1 0 1135 0 -1 2027
box 0 0 8 49
use AND2X2  AND2X2_65
timestamp 1516325494
transform -1 0 1153 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1481
timestamp 1516325494
transform -1 0 1172 0 -1 2027
box 0 0 19 49
use FILL  FILL_OR2X2_206
timestamp 1516325494
transform 1 0 1172 0 -1 2027
box 0 0 8 49
use OR2X2  OR2X2_206
timestamp 1516325494
transform 1 0 1180 0 -1 2027
box 0 0 19 49
use FILL  FILL_OR2X2_207
timestamp 1516325494
transform -1 0 1207 0 -1 2027
box 0 0 8 49
use OR2X2  OR2X2_207
timestamp 1516325494
transform -1 0 1226 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_386
timestamp 1516325494
transform 1 0 1226 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_413
timestamp 1516325494
transform -1 0 1264 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1941
timestamp 1516325494
transform 1 0 1264 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1942
timestamp 1516325494
transform 1 0 1283 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_387
timestamp 1516325494
transform 1 0 1302 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_385
timestamp 1516325494
transform -1 0 1340 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_411
timestamp 1516325494
transform -1 0 1359 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_341
timestamp 1516325494
transform -1 0 1378 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_364
timestamp 1516325494
transform -1 0 1397 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_365
timestamp 1516325494
transform -1 0 1416 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1941
timestamp 1516325494
transform -1 0 1435 0 -1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_804
timestamp 1516325494
transform 1 0 1435 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_804
timestamp 1516325494
transform 1 0 1442 0 -1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_816
timestamp 1516325494
transform 1 0 1457 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_816
timestamp 1516325494
transform 1 0 1465 0 -1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_64
timestamp 1516325494
transform 1 0 1480 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_64
timestamp 1516325494
transform 1 0 1488 0 -1 2027
box 0 0 15 49
use OR2X2  OR2X2_1099
timestamp 1516325494
transform 1 0 1503 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_547
timestamp 1516325494
transform 1 0 1522 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_547
timestamp 1516325494
transform -1 0 1567 0 -1 2027
box 0 0 30 49
use AND2X2  AND2X2_1373
timestamp 1516325494
transform -1 0 1587 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1100
timestamp 1516325494
transform -1 0 1606 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_67
timestamp 1516325494
transform 1 0 1606 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_67
timestamp 1516325494
transform -1 0 1651 0 -1 2027
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_99
timestamp 1516325494
transform -1 0 1704 0 -1 2027
box 0 0 53 49
use OR2X2  OR2X2_1938
timestamp 1516325494
transform 1 0 1704 0 -1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_593
timestamp 1516325494
transform -1 0 1731 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_593
timestamp 1516325494
transform -1 0 1746 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_99
timestamp 1516325494
transform 1 0 1746 0 -1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_99
timestamp 1516325494
transform -1 0 1792 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_3
timestamp 1516325494
transform -1 0 1845 0 -1 2027
box 0 0 53 49
use FILL  FILL_BUFX2_805
timestamp 1516325494
transform -1 0 1853 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_805
timestamp 1516325494
transform -1 0 1868 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_723
timestamp 1516325494
transform -1 0 1921 0 -1 2027
box 0 0 53 49
use AND2X2  AND2X2_1938
timestamp 1516325494
transform -1 0 1940 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1836
timestamp 1516325494
transform -1 0 1959 0 -1 2027
box 0 0 19 49
use FILL  FILL_AND2X2_7
timestamp 1516325494
transform 1 0 1959 0 -1 2027
box 0 0 8 49
use AND2X2  AND2X2_7
timestamp 1516325494
transform 1 0 1967 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1393
timestamp 1516325494
transform 1 0 1986 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_906
timestamp 1516325494
transform 1 0 2005 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_636
timestamp 1516325494
transform 1 0 2020 0 -1 2027
box 0 0 53 49
use MUX2X1  MUX2X1_851
timestamp 1516325494
transform -1 0 2103 0 -1 2027
box 0 0 30 49
use AND2X2  AND2X2_1392
timestamp 1516325494
transform -1 0 2122 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1125
timestamp 1516325494
transform -1 0 2141 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_132
timestamp 1516325494
transform 1 0 2141 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_324
timestamp 1516325494
transform 1 0 2157 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_324
timestamp 1516325494
transform -1 0 2202 0 -1 2027
box 0 0 30 49
use MUX2X1  MUX2X1_8
timestamp 1516325494
transform 1 0 2202 0 -1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_8
timestamp 1516325494
transform -1 0 2248 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_584
timestamp 1516325494
transform -1 0 2301 0 -1 2027
box 0 0 53 49
use FILL  FILL_BUFX2_131
timestamp 1516325494
transform 1 0 2301 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_131
timestamp 1516325494
transform 1 0 2309 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_700
timestamp 1516325494
transform 1 0 2324 0 -1 2027
box 0 0 53 49
use OR2X2  OR2X2_1832
timestamp 1516325494
transform -1 0 2396 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1940
timestamp 1516325494
transform -1 0 2415 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1839
timestamp 1516325494
transform -1 0 2434 0 -1 2027
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_316
timestamp 1516325494
transform 1 0 2434 0 -1 2027
box 0 0 53 49
use NAND2X1  NAND2X1_508
timestamp 1516325494
transform 1 0 2487 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_508
timestamp 1516325494
transform -1 0 2532 0 -1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_412
timestamp 1516325494
transform 1 0 2533 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_412
timestamp 1516325494
transform -1 0 2578 0 -1 2027
box 0 0 30 49
use FILL  FILL_BUFX2_114
timestamp 1516325494
transform -1 0 2586 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_114
timestamp 1516325494
transform -1 0 2601 0 -1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_215
timestamp 1516325494
transform 1 0 2601 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_215
timestamp 1516325494
transform 1 0 2609 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_603
timestamp 1516325494
transform 1 0 2624 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_603
timestamp 1516325494
transform -1 0 2669 0 -1 2027
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_283
timestamp 1516325494
transform -1 0 2723 0 -1 2027
box 0 0 53 49
use NAND2X1  NAND2X1_597
timestamp 1516325494
transform 1 0 2723 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_597
timestamp 1516325494
transform -1 0 2768 0 -1 2027
box 0 0 30 49
use MUX2X1  MUX2X1_213
timestamp 1516325494
transform 1 0 2768 0 -1 2027
box 0 0 30 49
use FILL  FILL_OR2X2_128
timestamp 1516325494
transform -1 0 2807 0 1 2027
box 0 0 8 49
use OR2X2  OR2X2_128
timestamp 1516325494
transform -1 0 2825 0 1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_382
timestamp 1516325494
transform 1 0 2825 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_382
timestamp 1516325494
transform 1 0 2833 0 1 2027
box 0 0 15 49
use FILL  FILL_AND2X2_134
timestamp 1516325494
transform -1 0 2856 0 1 2027
box 0 0 8 49
use AND2X2  AND2X2_134
timestamp 1516325494
transform -1 0 2875 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_1379
timestamp 1516325494
transform -1 0 2894 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1586
timestamp 1516325494
transform -1 0 2913 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_346
timestamp 1516325494
transform -1 0 2932 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1910
timestamp 1516325494
transform -1 0 2951 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_285
timestamp 1516325494
transform 1 0 2951 0 1 2027
box 0 0 19 49
use MUX2X1  MUX2X1_375
timestamp 1516325494
transform -1 0 3000 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_279
timestamp 1516325494
transform 1 0 3000 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_279
timestamp 1516325494
transform -1 0 3045 0 1 2027
box 0 0 30 49
use MUX2X1  MUX2X1_357
timestamp 1516325494
transform 1 0 3046 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_357
timestamp 1516325494
transform -1 0 3091 0 1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_261
timestamp 1516325494
transform 1 0 3091 0 1 2027
box 0 0 30 49
use NAND2X1  NAND2X1_261
timestamp 1516325494
transform -1 0 3137 0 1 2027
box 0 0 15 49
use OR2X2  OR2X2_959
timestamp 1516325494
transform 1 0 3137 0 1 2027
box 0 0 19 49
use XOR2X1  XOR2X1_71
timestamp 1516325494
transform 1 0 3156 0 1 2027
box 0 0 34 49
use AND2X2  AND2X2_1195
timestamp 1516325494
transform 1 0 3190 0 1 2027
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_788
timestamp 1516325494
transform 1 0 3209 0 1 2027
box 0 0 53 49
use NOR2X1  NOR2X1_139
timestamp 1516325494
transform -1 0 3277 0 1 2027
box 0 0 15 49
use NOR2X1  NOR2X1_136
timestamp 1516325494
transform 1 0 3278 0 1 2027
box 0 0 15 49
use INVX1  INVX1_269
timestamp 1516325494
transform -1 0 3304 0 1 2027
box 0 0 11 49
use NOR2X1  NOR2X1_137
timestamp 1516325494
transform 1 0 3304 0 1 2027
box 0 0 15 49
use AND2X2  AND2X2_1241
timestamp 1516325494
transform -1 0 3338 0 1 2027
box 0 0 19 49
use AOI21X1  AOI21X1_55
timestamp 1516325494
transform -1 0 3357 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1217
timestamp 1516325494
transform -1 0 3376 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_792
timestamp 1516325494
transform -1 0 3391 0 1 2027
box 0 0 15 49
use AOI22X1  AOI22X1_17
timestamp 1516325494
transform -1 0 3415 0 1 2027
box 0 0 23 49
use OAI21X1  OAI21X1_98
timestamp 1516325494
transform 1 0 3414 0 1 2027
box 0 0 19 49
use NAND3X1  NAND3X1_89
timestamp 1516325494
transform -1 0 3452 0 1 2027
box 0 0 19 49
use AOI22X1  AOI22X1_8
timestamp 1516325494
transform -1 0 3475 0 1 2027
box 0 0 23 49
use INVX1  INVX1_276
timestamp 1516325494
transform 1 0 3475 0 1 2027
box 0 0 11 49
use OAI21X1  OAI21X1_113
timestamp 1516325494
transform 1 0 3487 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_828
timestamp 1516325494
transform -1 0 3521 0 1 2027
box 0 0 15 49
use AOI21X1  AOI21X1_53
timestamp 1516325494
transform 1 0 3521 0 1 2027
box 0 0 19 49
use AOI21X1  AOI21X1_52
timestamp 1516325494
transform 1 0 3540 0 1 2027
box 0 0 19 49
use OAI21X1  OAI21X1_97
timestamp 1516325494
transform 1 0 3559 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_789
timestamp 1516325494
transform -1 0 3593 0 1 2027
box 0 0 15 49
use OR2X2  OR2X2_958
timestamp 1516325494
transform -1 0 3612 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1221
timestamp 1516325494
transform -1 0 3631 0 1 2027
box 0 0 19 49
use OR2X2  OR2X2_969
timestamp 1516325494
transform -1 0 3650 0 1 2027
box 0 0 19 49
use AOI22X1  AOI22X1_10
timestamp 1516325494
transform -1 0 3673 0 1 2027
box 0 0 23 49
use OR2X2  OR2X2_967
timestamp 1516325494
transform -1 0 3692 0 1 2027
box 0 0 19 49
use AND2X2  AND2X2_1220
timestamp 1516325494
transform -1 0 3711 0 1 2027
box 0 0 19 49
use FILL  FILL_BUFX2_405
timestamp 1516325494
transform -1 0 3719 0 1 2027
box 0 0 8 49
use BUFX2  BUFX2_405
timestamp 1516325494
transform -1 0 3733 0 1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_774
timestamp 1516325494
transform 1 0 3734 0 1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_845
timestamp 1516325494
transform 1 0 3749 0 1 2027
box 0 0 15 49
use NOR2X1  NOR2X1_147
timestamp 1516325494
transform 1 0 3764 0 1 2027
box 0 0 15 49
use AOI21X1  AOI21X1_61
timestamp 1516325494
transform 1 0 3779 0 1 2027
box 0 0 19 49
use AOI22X1  AOI22X1_6
timestamp 1516325494
transform -1 0 3821 0 1 2027
box 0 0 23 49
use NAND3X1  NAND3X1_81
timestamp 1516325494
transform 1 0 3821 0 1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_775
timestamp 1516325494
transform -1 0 3855 0 1 2027
box 0 0 15 49
use INVX1  INVX1_275
timestamp 1516325494
transform -1 0 3866 0 1 2027
box 0 0 11 49
use NAND2X1  NAND2X1_213
timestamp 1516325494
transform -1 0 2814 0 -1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_9
timestamp 1516325494
transform -1 0 2822 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_9
timestamp 1516325494
transform -1 0 2837 0 -1 2027
box 0 0 15 49
use FILL  FILL_BUFX2_115
timestamp 1516325494
transform -1 0 2845 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_115
timestamp 1516325494
transform -1 0 2859 0 -1 2027
box 0 0 15 49
use FILL  FILL_OR2X2_127
timestamp 1516325494
transform -1 0 2868 0 -1 2027
box 0 0 8 49
use OR2X2  OR2X2_127
timestamp 1516325494
transform -1 0 2886 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_1378
timestamp 1516325494
transform -1 0 2905 0 -1 2027
box 0 0 19 49
use FILL  FILL_AND2X2_136
timestamp 1516325494
transform -1 0 2913 0 -1 2027
box 0 0 8 49
use AND2X2  AND2X2_136
timestamp 1516325494
transform -1 0 2932 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1588
timestamp 1516325494
transform -1 0 2951 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_379
timestamp 1516325494
transform 1 0 2951 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_375
timestamp 1516325494
transform -1 0 2981 0 -1 2027
box 0 0 15 49
use MUX2X1  MUX2X1_379
timestamp 1516325494
transform -1 0 3011 0 -1 2027
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_343
timestamp 1516325494
transform -1 0 3065 0 -1 2027
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_325
timestamp 1516325494
transform -1 0 3118 0 -1 2027
box 0 0 53 49
use AND2X2  AND2X2_1206
timestamp 1516325494
transform 1 0 3118 0 -1 2027
box 0 0 19 49
use XNOR2X1  XNOR2X1_58
timestamp 1516325494
transform -1 0 3171 0 -1 2027
box 0 0 34 49
use AND2X2  AND2X2_1197
timestamp 1516325494
transform 1 0 3171 0 -1 2027
box 0 0 19 49
use NAND3X1  NAND3X1_86
timestamp 1516325494
transform 1 0 3190 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_957
timestamp 1516325494
transform 1 0 3209 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1198
timestamp 1516325494
transform 1 0 3228 0 -1 2027
box 0 0 19 49
use INVX1  INVX1_268
timestamp 1516325494
transform 1 0 3247 0 -1 2027
box 0 0 11 49
use NOR2X1  NOR2X1_135
timestamp 1516325494
transform 1 0 3259 0 -1 2027
box 0 0 15 49
use NOR2X1  NOR2X1_138
timestamp 1516325494
transform -1 0 3289 0 -1 2027
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_807
timestamp 1516325494
transform 1 0 3289 0 -1 2027
box 0 0 53 49
use NAND2X1  NAND2X1_795
timestamp 1516325494
transform -1 0 3357 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_794
timestamp 1516325494
transform -1 0 3372 0 -1 2027
box 0 0 15 49
use NAND2X1  NAND2X1_793
timestamp 1516325494
transform -1 0 3388 0 -1 2027
box 0 0 15 49
use AND2X2  AND2X2_1215
timestamp 1516325494
transform 1 0 3388 0 -1 2027
box 0 0 19 49
use AOI22X1  AOI22X1_29
timestamp 1516325494
transform 1 0 3407 0 -1 2027
box 0 0 23 49
use NAND2X1  NAND2X1_797
timestamp 1516325494
transform -1 0 3445 0 -1 2027
box 0 0 15 49
use OR2X2  OR2X2_964
timestamp 1516325494
transform 1 0 3445 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_965
timestamp 1516325494
transform 1 0 3464 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_966
timestamp 1516325494
transform 1 0 3483 0 -1 2027
box 0 0 19 49
use XOR2X1  XOR2X1_73
timestamp 1516325494
transform 1 0 3502 0 -1 2027
box 0 0 34 49
use AND2X2  AND2X2_1201
timestamp 1516325494
transform -1 0 3555 0 -1 2027
box 0 0 19 49
use NAND3X1  NAND3X1_88
timestamp 1516325494
transform -1 0 3574 0 -1 2027
box 0 0 19 49
use NAND3X1  NAND3X1_87
timestamp 1516325494
transform -1 0 3593 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1218
timestamp 1516325494
transform 1 0 3593 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_968
timestamp 1516325494
transform 1 0 3612 0 -1 2027
box 0 0 19 49
use AND2X2  AND2X2_1200
timestamp 1516325494
transform 1 0 3631 0 -1 2027
box 0 0 19 49
use INVX1  INVX1_271
timestamp 1516325494
transform -1 0 3661 0 -1 2027
box 0 0 11 49
use FILL  FILL_BUFX2_85
timestamp 1516325494
transform 1 0 3661 0 -1 2027
box 0 0 8 49
use BUFX2  BUFX2_85
timestamp 1516325494
transform 1 0 3669 0 -1 2027
box 0 0 15 49
use INVX1  INVX1_299
timestamp 1516325494
transform -1 0 3695 0 -1 2027
box 0 0 11 49
use OR2X2  OR2X2_962
timestamp 1516325494
transform 1 0 3696 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_963
timestamp 1516325494
transform -1 0 3734 0 -1 2027
box 0 0 19 49
use OR2X2  OR2X2_961
timestamp 1516325494
transform -1 0 3753 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_829
timestamp 1516325494
transform 1 0 3753 0 -1 2027
box 0 0 15 49
use AOI21X1  AOI21X1_58
timestamp 1516325494
transform 1 0 3768 0 -1 2027
box 0 0 19 49
use NOR2X1  NOR2X1_141
timestamp 1516325494
transform -1 0 3802 0 -1 2027
box 0 0 15 49
use AND2X2  AND2X2_1212
timestamp 1516325494
transform -1 0 3821 0 -1 2027
box 0 0 19 49
use NAND2X1  NAND2X1_827
timestamp 1516325494
transform 1 0 3821 0 -1 2027
box 0 0 15 49
use OAI21X1  OAI21X1_114
timestamp 1516325494
transform 1 0 3836 0 -1 2027
box 0 0 19 49
use FILL  FILL_41_1
timestamp 1516325494
transform -1 0 3863 0 -1 2027
box 0 0 8 49
use FILL  FILL_41_2
timestamp 1516325494
transform -1 0 3871 0 -1 2027
box 0 0 8 49
use OR2X2  OR2X2_895
timestamp 1516325494
transform -1 0 21 0 1 1928
box 0 0 19 49
use INVX1  INVX1_87
timestamp 1516325494
transform -1 0 32 0 1 1928
box 0 0 11 49
use NOR2X1  NOR2X1_90
timestamp 1516325494
transform -1 0 47 0 1 1928
box 0 0 15 49
use XOR2X1  XOR2X1_45
timestamp 1516325494
transform 1 0 2 0 -1 1928
box 0 0 34 49
use INVX1  INVX1_88
timestamp 1516325494
transform -1 0 47 0 -1 1928
box 0 0 11 49
use BUFX2  BUFX2_886
timestamp 1516325494
transform 1 0 2 0 1 1830
box 0 0 15 49
use AND2X2  AND2X2_1099
timestamp 1516325494
transform -1 0 36 0 1 1830
box 0 0 19 49
use INVX1  INVX1_83
timestamp 1516325494
transform -1 0 47 0 1 1830
box 0 0 11 49
use XNOR2X1  XNOR2X1_25
timestamp 1516325494
transform 1 0 48 0 1 1928
box 0 0 34 49
use INVX1  INVX1_80
timestamp 1516325494
transform -1 0 93 0 1 1928
box 0 0 11 49
use XNOR2X1  XNOR2X1_24
timestamp 1516325494
transform -1 0 127 0 1 1928
box 0 0 34 49
use AND2X2  AND2X2_876
timestamp 1516325494
transform -1 0 146 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_875
timestamp 1516325494
transform -1 0 165 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_737
timestamp 1516325494
transform -1 0 184 0 1 1928
box 0 0 19 49
use NOR2X1  NOR2X1_50
timestamp 1516325494
transform -1 0 199 0 1 1928
box 0 0 15 49
use AOI21X1  AOI21X1_14
timestamp 1516325494
transform -1 0 219 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_674
timestamp 1516325494
transform 1 0 219 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_151
timestamp 1516325494
transform 1 0 234 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_151
timestamp 1516325494
transform 1 0 241 0 1 1928
box 0 0 15 49
use INVX2  INVX2_2
timestamp 1516325494
transform 1 0 257 0 1 1928
box 0 0 11 49
use FILL  FILL_BUFX2_743
timestamp 1516325494
transform 1 0 268 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_743
timestamp 1516325494
transform 1 0 276 0 1 1928
box 0 0 15 49
use XNOR2X1  XNOR2X1_34
timestamp 1516325494
transform -1 0 325 0 1 1928
box 0 0 34 49
use FILL  FILL_BUFX2_628
timestamp 1516325494
transform 1 0 325 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_628
timestamp 1516325494
transform 1 0 333 0 1 1928
box 0 0 15 49
use NOR2X1  NOR2X1_57
timestamp 1516325494
transform 1 0 348 0 1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_681
timestamp 1516325494
transform 1 0 363 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_744
timestamp 1516325494
transform -1 0 386 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_744
timestamp 1516325494
transform -1 0 401 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_154
timestamp 1516325494
transform -1 0 409 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_154
timestamp 1516325494
transform -1 0 424 0 1 1928
box 0 0 15 49
use OAI21X1  OAI21X1_4
timestamp 1516325494
transform -1 0 443 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_729
timestamp 1516325494
transform -1 0 462 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_613
timestamp 1516325494
transform -1 0 481 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_661
timestamp 1516325494
transform -1 0 496 0 1 1928
box 0 0 15 49
use OR2X2  OR2X2_806
timestamp 1516325494
transform 1 0 496 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_629
timestamp 1516325494
transform -1 0 523 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_629
timestamp 1516325494
transform -1 0 538 0 1 1928
box 0 0 15 49
use NOR2X1  NOR2X1_62
timestamp 1516325494
transform 1 0 538 0 1 1928
box 0 0 15 49
use OR2X2  OR2X2_788
timestamp 1516325494
transform 1 0 553 0 1 1928
box 0 0 19 49
use AOI21X1  AOI21X1_8
timestamp 1516325494
transform -1 0 591 0 1 1928
box 0 0 19 49
use XOR2X1  XOR2X1_10
timestamp 1516325494
transform -1 0 625 0 1 1928
box 0 0 34 49
use AND2X2  AND2X2_1073
timestamp 1516325494
transform -1 0 644 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_665
timestamp 1516325494
transform -1 0 659 0 1 1928
box 0 0 15 49
use OAI21X1  OAI21X1_74
timestamp 1516325494
transform -1 0 678 0 1 1928
box 0 0 19 49
use OAI21X1  OAI21X1_64
timestamp 1516325494
transform -1 0 697 0 1 1928
box 0 0 19 49
use INVX1  INVX1_42
timestamp 1516325494
transform 1 0 697 0 1 1928
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_749
timestamp 1516325494
transform -1 0 762 0 1 1928
box 0 0 53 49
use INVX1  INVX1_46
timestamp 1516325494
transform 1 0 762 0 1 1928
box 0 0 11 49
use OAI21X1  OAI21X1_61
timestamp 1516325494
transform 1 0 773 0 1 1928
box 0 0 19 49
use MUX2X1  MUX2X1_777
timestamp 1516325494
transform 1 0 792 0 1 1928
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_736
timestamp 1516325494
transform -1 0 876 0 1 1928
box 0 0 53 49
use MUX2X1  MUX2X1_764
timestamp 1516325494
transform 1 0 876 0 1 1928
box 0 0 30 49
use OR2X2  OR2X2_319
timestamp 1516325494
transform -1 0 925 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_318
timestamp 1516325494
transform -1 0 944 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1794
timestamp 1516325494
transform -1 0 963 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1793
timestamp 1516325494
transform -1 0 982 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1775
timestamp 1516325494
transform 1 0 982 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1623
timestamp 1516325494
transform -1 0 1020 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_469
timestamp 1516325494
transform 1 0 1020 0 1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_469
timestamp 1516325494
transform -1 0 1066 0 1 1928
box 0 0 30 49
use FILL  FILL_AND2X2_63
timestamp 1516325494
transform -1 0 1074 0 1 1928
box 0 0 8 49
use AND2X2  AND2X2_63
timestamp 1516325494
transform -1 0 1093 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1477
timestamp 1516325494
transform 1 0 1093 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1235
timestamp 1516325494
transform -1 0 1131 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1239
timestamp 1516325494
transform 1 0 1131 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1480
timestamp 1516325494
transform 1 0 1150 0 1 1928
box 0 0 19 49
use FILL  FILL_OR2X2_244
timestamp 1516325494
transform -1 0 1177 0 1 1928
box 0 0 8 49
use OR2X2  OR2X2_244
timestamp 1516325494
transform -1 0 1195 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1475
timestamp 1516325494
transform -1 0 1214 0 1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_62
timestamp 1516325494
transform -1 0 1222 0 1 1928
box 0 0 8 49
use AND2X2  AND2X2_62
timestamp 1516325494
transform -1 0 1241 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_537
timestamp 1516325494
transform 1 0 1241 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_537
timestamp 1516325494
transform 1 0 1248 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_283
timestamp 1516325494
transform 1 0 1264 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_283
timestamp 1516325494
transform 1 0 1271 0 1 1928
box 0 0 15 49
use FILL  FILL_OR2X2_243
timestamp 1516325494
transform -1 0 1294 0 1 1928
box 0 0 8 49
use OR2X2  OR2X2_243
timestamp 1516325494
transform -1 0 1313 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_2016
timestamp 1516325494
transform -1 0 1332 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_389
timestamp 1516325494
transform -1 0 1351 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_388
timestamp 1516325494
transform -1 0 1370 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1835
timestamp 1516325494
transform -1 0 1389 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1935
timestamp 1516325494
transform -1 0 1408 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1937
timestamp 1516325494
transform -1 0 1427 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_340
timestamp 1516325494
transform -1 0 1446 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_362
timestamp 1516325494
transform -1 0 1465 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_363
timestamp 1516325494
transform -1 0 1484 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_483
timestamp 1516325494
transform 1 0 1484 0 1 1928
box 0 0 53 49
use OR2X2  OR2X2_1934
timestamp 1516325494
transform -1 0 1556 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_479
timestamp 1516325494
transform 1 0 1556 0 1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_351
timestamp 1516325494
transform 1 0 1609 0 1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_351
timestamp 1516325494
transform 1 0 1625 0 1 1928
box 0 0 30 49
use FILL  FILL_BUFX2_740
timestamp 1516325494
transform 1 0 1655 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_740
timestamp 1516325494
transform 1 0 1663 0 1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_476
timestamp 1516325494
transform 1 0 1678 0 1 1928
box 0 0 30 49
use NAND2X1  NAND2X1_476
timestamp 1516325494
transform -1 0 1723 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_2015
timestamp 1516325494
transform 1 0 1723 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_572
timestamp 1516325494
transform -1 0 1795 0 1 1928
box 0 0 53 49
use OR2X2  OR2X2_1833
timestamp 1516325494
transform 1 0 1796 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1936
timestamp 1516325494
transform -1 0 1834 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1098
timestamp 1516325494
transform -1 0 1853 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_332
timestamp 1516325494
transform 1 0 1853 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_332
timestamp 1516325494
transform 1 0 1860 0 1 1928
box 0 0 15 49
use OR2X2  OR2X2_1834
timestamp 1516325494
transform -1 0 1894 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1397
timestamp 1516325494
transform 1 0 1894 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1131
timestamp 1516325494
transform 1 0 1913 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_284
timestamp 1516325494
transform 1 0 1932 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_284
timestamp 1516325494
transform 1 0 1940 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_196
timestamp 1516325494
transform 1 0 1955 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_196
timestamp 1516325494
transform 1 0 1963 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_737
timestamp 1516325494
transform 1 0 1978 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_737
timestamp 1516325494
transform 1 0 1986 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_134
timestamp 1516325494
transform -1 0 2009 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_134
timestamp 1516325494
transform -1 0 2023 0 1 1928
box 0 0 15 49
use OR2X2  OR2X2_1132
timestamp 1516325494
transform 1 0 2024 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1126
timestamp 1516325494
transform -1 0 2062 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_452
timestamp 1516325494
transform 1 0 2062 0 1 1928
box 0 0 53 49
use OR2X2  OR2X2_1124
timestamp 1516325494
transform -1 0 2134 0 1 1928
box 0 0 19 49
use MUX2X1  MUX2X1_28
timestamp 1516325494
transform 1 0 2134 0 1 1928
box 0 0 30 49
use NAND2X1  NAND2X1_28
timestamp 1516325494
transform -1 0 2179 0 1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_604
timestamp 1516325494
transform -1 0 2232 0 1 1928
box 0 0 53 49
use AND2X2  AND2X2_2011
timestamp 1516325494
transform 1 0 2233 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1231
timestamp 1516325494
transform -1 0 2271 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1831
timestamp 1516325494
transform 1 0 2271 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1934
timestamp 1516325494
transform -1 0 2309 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_1932
timestamp 1516325494
transform -1 0 2328 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_316
timestamp 1516325494
transform 1 0 2328 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_19
timestamp 1516325494
transform -1 0 2351 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_19
timestamp 1516325494
transform -1 0 2365 0 1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_316
timestamp 1516325494
transform -1 0 2396 0 1 1928
box 0 0 30 49
use FILL  FILL_BUFX2_25
timestamp 1516325494
transform 1 0 2396 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_25
timestamp 1516325494
transform 1 0 2404 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_578
timestamp 1516325494
transform 1 0 2419 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_578
timestamp 1516325494
transform 1 0 2426 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_1097
timestamp 1516325494
transform -1 0 67 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_892
timestamp 1516325494
transform -1 0 86 0 -1 1928
box 0 0 19 49
use INVX1  INVX1_78
timestamp 1516325494
transform -1 0 97 0 -1 1928
box 0 0 11 49
use XOR2X1  XOR2X1_42
timestamp 1516325494
transform -1 0 131 0 -1 1928
box 0 0 34 49
use NOR2X1  NOR2X1_56
timestamp 1516325494
transform -1 0 146 0 -1 1928
box 0 0 15 49
use NOR2X1  NOR2X1_51
timestamp 1516325494
transform 1 0 146 0 -1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_675
timestamp 1516325494
transform -1 0 177 0 -1 1928
box 0 0 15 49
use OR2X2  OR2X2_752
timestamp 1516325494
transform 1 0 177 0 -1 1928
box 0 0 19 49
use XOR2X1  XOR2X1_12
timestamp 1516325494
transform 1 0 196 0 -1 1928
box 0 0 34 49
use FILL  FILL_BUFX2_640
timestamp 1516325494
transform -1 0 238 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_640
timestamp 1516325494
transform -1 0 253 0 -1 1928
box 0 0 15 49
use XOR2X1  XOR2X1_25
timestamp 1516325494
transform -1 0 287 0 -1 1928
box 0 0 34 49
use NAND2X1  NAND2X1_696
timestamp 1516325494
transform -1 0 302 0 -1 1928
box 0 0 15 49
use OR2X2  OR2X2_875
timestamp 1516325494
transform 1 0 302 0 -1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_787
timestamp 1516325494
transform 1 0 321 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_787
timestamp 1516325494
transform 1 0 329 0 -1 1928
box 0 0 15 49
use XOR2X1  XOR2X1_15
timestamp 1516325494
transform -1 0 378 0 -1 1928
box 0 0 34 49
use OR2X2  OR2X2_760
timestamp 1516325494
transform 1 0 378 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_908
timestamp 1516325494
transform 1 0 397 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_730
timestamp 1516325494
transform -1 0 435 0 -1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_741
timestamp 1516325494
transform -1 0 443 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_741
timestamp 1516325494
transform -1 0 458 0 -1 1928
box 0 0 15 49
use NAND3X1  NAND3X1_37
timestamp 1516325494
transform -1 0 477 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_662
timestamp 1516325494
transform -1 0 492 0 -1 1928
box 0 0 15 49
use NAND3X1  NAND3X1_36
timestamp 1516325494
transform -1 0 511 0 -1 1928
box 0 0 19 49
use XNOR2X1  XNOR2X1_9
timestamp 1516325494
transform -1 0 545 0 -1 1928
box 0 0 34 49
use INVX1  INVX1_37
timestamp 1516325494
transform 1 0 545 0 -1 1928
box 0 0 11 49
use OR2X2  OR2X2_671
timestamp 1516325494
transform -1 0 576 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_670
timestamp 1516325494
transform 1 0 576 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_865
timestamp 1516325494
transform 1 0 595 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1076
timestamp 1516325494
transform 1 0 614 0 -1 1928
box 0 0 19 49
use INVX1  INVX1_53
timestamp 1516325494
transform 1 0 633 0 -1 1928
box 0 0 11 49
use NOR2X1  NOR2X1_39
timestamp 1516325494
transform -1 0 659 0 -1 1928
box 0 0 15 49
use AND2X2  AND2X2_1084
timestamp 1516325494
transform 1 0 659 0 -1 1928
box 0 0 19 49
use XNOR2X1  XNOR2X1_14
timestamp 1516325494
transform 1 0 678 0 -1 1928
box 0 0 34 49
use DFFPOSX1  DFFPOSX1_740
timestamp 1516325494
transform -1 0 766 0 -1 1928
box 0 0 53 49
use INVX1  INVX1_45
timestamp 1516325494
transform 1 0 766 0 -1 1928
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_743
timestamp 1516325494
transform -1 0 830 0 -1 1928
box 0 0 53 49
use INVX1  INVX1_56
timestamp 1516325494
transform 1 0 830 0 -1 1928
box 0 0 11 49
use FILL  FILL_BUFX2_320
timestamp 1516325494
transform 1 0 842 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_320
timestamp 1516325494
transform 1 0 849 0 -1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_750
timestamp 1516325494
transform -1 0 918 0 -1 1928
box 0 0 53 49
use OR2X2  OR2X2_1554
timestamp 1516325494
transform -1 0 937 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1553
timestamp 1516325494
transform -1 0 956 0 -1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_680
timestamp 1516325494
transform 1 0 956 0 -1 1928
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_565
timestamp 1516325494
transform 1 0 1009 0 -1 1928
box 0 0 53 49
use OR2X2  OR2X2_1631
timestamp 1516325494
transform -1 0 1081 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1625
timestamp 1516325494
transform -1 0 1100 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1776
timestamp 1516325494
transform -1 0 1119 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_258
timestamp 1516325494
transform 1 0 1119 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_258
timestamp 1516325494
transform 1 0 1127 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1774
timestamp 1516325494
transform -1 0 1165 0 -1 1928
box 0 0 19 49
use FILL  FILL_OR2X2_242
timestamp 1516325494
transform 1 0 1165 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_242
timestamp 1516325494
transform 1 0 1172 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_257
timestamp 1516325494
transform -1 0 1199 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_257
timestamp 1516325494
transform -1 0 1218 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1630
timestamp 1516325494
transform -1 0 1237 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1778
timestamp 1516325494
transform -1 0 1256 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1780
timestamp 1516325494
transform -1 0 1275 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_259
timestamp 1516325494
transform 1 0 1275 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_259
timestamp 1516325494
transform 1 0 1283 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_260
timestamp 1516325494
transform -1 0 1310 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_260
timestamp 1516325494
transform -1 0 1328 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1944
timestamp 1516325494
transform -1 0 1347 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1943
timestamp 1516325494
transform -1 0 1366 0 -1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_540
timestamp 1516325494
transform 1 0 1366 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_540
timestamp 1516325494
transform 1 0 1374 0 -1 1928
box 0 0 15 49
use AND2X2  AND2X2_2008
timestamp 1516325494
transform -1 0 1408 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_409
timestamp 1516325494
transform 1 0 1408 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1931
timestamp 1516325494
transform -1 0 1446 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1930
timestamp 1516325494
transform -1 0 1465 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_384
timestamp 1516325494
transform -1 0 1484 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_383
timestamp 1516325494
transform -1 0 1503 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_410
timestamp 1516325494
transform -1 0 1522 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_2010
timestamp 1516325494
transform 1 0 1522 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1929
timestamp 1516325494
transform -1 0 1560 0 -1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_296
timestamp 1516325494
transform 1 0 1560 0 -1 1928
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_575
timestamp 1516325494
transform 1 0 1613 0 -1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_488
timestamp 1516325494
transform 1 0 1666 0 -1 1928
box 0 0 15 49
use NOR2X1  NOR2X1_88
timestamp 1516325494
transform -1 0 63 0 1 1830
box 0 0 15 49
use INVX1  INVX1_82
timestamp 1516325494
transform -1 0 74 0 1 1830
box 0 0 11 49
use XNOR2X1  XNOR2X1_21
timestamp 1516325494
transform 1 0 74 0 1 1830
box 0 0 34 49
use AND2X2  AND2X2_1096
timestamp 1516325494
transform -1 0 127 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_891
timestamp 1516325494
transform -1 0 146 0 1 1830
box 0 0 19 49
use XNOR2X1  XNOR2X1_20
timestamp 1516325494
transform -1 0 180 0 1 1830
box 0 0 34 49
use AND2X2  AND2X2_1054
timestamp 1516325494
transform 1 0 181 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1046
timestamp 1516325494
transform -1 0 219 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_669
timestamp 1516325494
transform 1 0 219 0 1 1830
box 0 0 15 49
use NAND2X1  NAND2X1_670
timestamp 1516325494
transform -1 0 249 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_841
timestamp 1516325494
transform -1 0 268 0 1 1830
box 0 0 19 49
use XOR2X1  XOR2X1_11
timestamp 1516325494
transform 1 0 268 0 1 1830
box 0 0 34 49
use XOR2X1  XOR2X1_24
timestamp 1516325494
transform -1 0 336 0 1 1830
box 0 0 34 49
use OR2X2  OR2X2_859
timestamp 1516325494
transform 1 0 336 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_759
timestamp 1516325494
transform 1 0 355 0 1 1830
box 0 0 19 49
use XOR2X1  XOR2X1_14
timestamp 1516325494
transform 1 0 374 0 1 1830
box 0 0 34 49
use OR2X2  OR2X2_779
timestamp 1516325494
transform -1 0 428 0 1 1830
box 0 0 19 49
use NOR2X1  NOR2X1_61
timestamp 1516325494
transform -1 0 443 0 1 1830
box 0 0 15 49
use NOR2X1  NOR2X1_43
timestamp 1516325494
transform 1 0 443 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_746
timestamp 1516325494
transform 1 0 458 0 1 1830
box 0 0 19 49
use XOR2X1  XOR2X1_17
timestamp 1516325494
transform 1 0 477 0 1 1830
box 0 0 34 49
use NAND2X1  NAND2X1_683
timestamp 1516325494
transform -1 0 526 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_851
timestamp 1516325494
transform 1 0 526 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1081
timestamp 1516325494
transform 1 0 545 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1082
timestamp 1516325494
transform 1 0 564 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_624
timestamp 1516325494
transform -1 0 591 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_624
timestamp 1516325494
transform -1 0 606 0 1 1830
box 0 0 15 49
use AND2X2  AND2X2_1077
timestamp 1516325494
transform 1 0 606 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1078
timestamp 1516325494
transform 1 0 625 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1083
timestamp 1516325494
transform 1 0 644 0 1 1830
box 0 0 19 49
use INVX1  INVX1_74
timestamp 1516325494
transform -1 0 674 0 1 1830
box 0 0 11 49
use XNOR2X1  XNOR2X1_15
timestamp 1516325494
transform -1 0 709 0 1 1830
box 0 0 34 49
use INVX1  INVX1_72
timestamp 1516325494
transform 1 0 709 0 1 1830
box 0 0 11 49
use NOR2X1  NOR2X1_85
timestamp 1516325494
transform 1 0 720 0 1 1830
box 0 0 15 49
use INVX1  INVX1_52
timestamp 1516325494
transform 1 0 735 0 1 1830
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_748
timestamp 1516325494
transform -1 0 800 0 1 1830
box 0 0 53 49
use MUX2X1  MUX2X1_776
timestamp 1516325494
transform 1 0 800 0 1 1830
box 0 0 30 49
use MUX2X1  MUX2X1_771
timestamp 1516325494
transform 1 0 830 0 1 1830
box 0 0 30 49
use INVX1  INVX1_164
timestamp 1516325494
transform 1 0 861 0 1 1830
box 0 0 11 49
use MUX2X1  MUX2X1_768
timestamp 1516325494
transform 1 0 872 0 1 1830
box 0 0 30 49
use INVX1  INVX1_51
timestamp 1516325494
transform 1 0 903 0 1 1830
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_121
timestamp 1516325494
transform 1 0 914 0 1 1830
box 0 0 53 49
use OR2X2  OR2X2_1234
timestamp 1516325494
transform 1 0 967 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1476
timestamp 1516325494
transform 1 0 986 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_296
timestamp 1516325494
transform 1 0 1005 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_296
timestamp 1516325494
transform -1 0 1050 0 1 1830
box 0 0 30 49
use OR2X2  OR2X2_1781
timestamp 1516325494
transform -1 0 1070 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_314
timestamp 1516325494
transform -1 0 1089 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1780
timestamp 1516325494
transform -1 0 1108 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1893
timestamp 1516325494
transform -1 0 1127 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_313
timestamp 1516325494
transform -1 0 1146 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_334
timestamp 1516325494
transform -1 0 1165 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1895
timestamp 1516325494
transform -1 0 1184 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_335
timestamp 1516325494
transform -1 0 1203 0 1 1830
box 0 0 19 49
use FILL  FILL_OR2X2_202
timestamp 1516325494
transform -1 0 1211 0 1 1830
box 0 0 8 49
use OR2X2  OR2X2_202
timestamp 1516325494
transform -1 0 1229 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1541
timestamp 1516325494
transform -1 0 1248 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_138
timestamp 1516325494
transform 1 0 1248 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_138
timestamp 1516325494
transform 1 0 1256 0 1 1830
box 0 0 15 49
use FILL  FILL_OR2X2_201
timestamp 1516325494
transform -1 0 1279 0 1 1830
box 0 0 8 49
use OR2X2  OR2X2_201
timestamp 1516325494
transform -1 0 1298 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1540
timestamp 1516325494
transform -1 0 1317 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1709
timestamp 1516325494
transform -1 0 1336 0 1 1830
box 0 0 19 49
use FILL  FILL_AND2X2_214
timestamp 1516325494
transform -1 0 1344 0 1 1830
box 0 0 8 49
use AND2X2  AND2X2_214
timestamp 1516325494
transform -1 0 1362 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1711
timestamp 1516325494
transform -1 0 1381 0 1 1830
box 0 0 19 49
use FILL  FILL_AND2X2_215
timestamp 1516325494
transform -1 0 1389 0 1 1830
box 0 0 8 49
use AND2X2  AND2X2_215
timestamp 1516325494
transform -1 0 1408 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_2004
timestamp 1516325494
transform -1 0 1427 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1925
timestamp 1516325494
transform 1 0 1427 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_2006
timestamp 1516325494
transform -1 0 1465 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_408
timestamp 1516325494
transform 1 0 1465 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_382
timestamp 1516325494
transform -1 0 1503 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_407
timestamp 1516325494
transform -1 0 1522 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_2009
timestamp 1516325494
transform -1 0 1541 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1928
timestamp 1516325494
transform -1 0 1560 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1777
timestamp 1516325494
transform -1 0 1579 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_2005
timestamp 1516325494
transform -1 0 1598 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1923
timestamp 1516325494
transform -1 0 1617 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1626
timestamp 1516325494
transform -1 0 1636 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_479
timestamp 1516325494
transform 1 0 1636 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_479
timestamp 1516325494
transform -1 0 1681 0 1 1830
box 0 0 30 49
use MUX2X1  MUX2X1_488
timestamp 1516325494
transform -1 0 1712 0 -1 1928
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_319
timestamp 1516325494
transform 1 0 1712 0 -1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_511
timestamp 1516325494
transform 1 0 1765 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_511
timestamp 1516325494
transform -1 0 1810 0 -1 1928
box 0 0 30 49
use FILL  FILL_BUFX2_98
timestamp 1516325494
transform 1 0 1811 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_98
timestamp 1516325494
transform 1 0 1818 0 -1 1928
box 0 0 15 49
use AND2X2  AND2X2_1371
timestamp 1516325494
transform 1 0 1834 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1372
timestamp 1516325494
transform 1 0 1853 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_2106
timestamp 1516325494
transform 1 0 1872 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_9
timestamp 1516325494
transform 1 0 1891 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_9
timestamp 1516325494
transform 1 0 1898 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1395
timestamp 1516325494
transform -1 0 1936 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_8
timestamp 1516325494
transform 1 0 1936 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_8
timestamp 1516325494
transform 1 0 1944 0 -1 1928
box 0 0 19 49
use FILL  FILL_OR2X2_8
timestamp 1516325494
transform 1 0 1963 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_8
timestamp 1516325494
transform 1 0 1970 0 -1 1928
box 0 0 19 49
use FILL  FILL_OR2X2_9
timestamp 1516325494
transform 1 0 1989 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_9
timestamp 1516325494
transform 1 0 1997 0 -1 1928
box 0 0 19 49
use FILL  FILL_OR2X2_7
timestamp 1516325494
transform -1 0 2024 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_7
timestamp 1516325494
transform -1 0 2043 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_6
timestamp 1516325494
transform -1 0 2051 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_6
timestamp 1516325494
transform -1 0 2069 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1391
timestamp 1516325494
transform -1 0 2088 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1474
timestamp 1516325494
transform -1 0 2107 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1232
timestamp 1516325494
transform -1 0 2126 0 -1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_424
timestamp 1516325494
transform 1 0 2126 0 -1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_392
timestamp 1516325494
transform 1 0 2179 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_392
timestamp 1516325494
transform -1 0 2225 0 -1 1928
box 0 0 30 49
use OR2X2  OR2X2_1933
timestamp 1516325494
transform -1 0 2244 0 -1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_415
timestamp 1516325494
transform 1 0 2244 0 -1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_191
timestamp 1516325494
transform 1 0 2297 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_191
timestamp 1516325494
transform 1 0 2312 0 -1 1928
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_383
timestamp 1516325494
transform 1 0 2343 0 -1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_941
timestamp 1516325494
transform 1 0 2396 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_886
timestamp 1516325494
transform -1 0 2441 0 -1 1928
box 0 0 30 49
use MUX2X1  MUX2X1_859
timestamp 1516325494
transform 1 0 2442 0 1 1928
box 0 0 30 49
use INVX1  INVX1_272
timestamp 1516325494
transform 1 0 2472 0 1 1928
box 0 0 11 49
use OR2X2  OR2X2_1838
timestamp 1516325494
transform -1 0 2502 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_718
timestamp 1516325494
transform 1 0 2502 0 1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_388
timestamp 1516325494
transform 1 0 2518 0 1 1928
box 0 0 53 49
use OR2X2  OR2X2_1123
timestamp 1516325494
transform -1 0 2590 0 1 1928
box 0 0 19 49
use MUX2X1  MUX2X1_60
timestamp 1516325494
transform 1 0 2590 0 1 1928
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_668
timestamp 1516325494
transform -1 0 2673 0 1 1928
box 0 0 53 49
use FILL  FILL_BUFX2_773
timestamp 1516325494
transform 1 0 2673 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_773
timestamp 1516325494
transform 1 0 2681 0 1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_277
timestamp 1516325494
transform 1 0 2696 0 1 1928
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_245
timestamp 1516325494
transform -1 0 2802 0 1 1928
box 0 0 53 49
use FILL  FILL_BUFX2_707
timestamp 1516325494
transform 1 0 2803 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_707
timestamp 1516325494
transform 1 0 2810 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_835
timestamp 1516325494
transform 1 0 2825 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_835
timestamp 1516325494
transform 1 0 2833 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_397
timestamp 1516325494
transform 1 0 2848 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_397
timestamp 1516325494
transform 1 0 2856 0 1 1928
box 0 0 15 49
use FILL  FILL_AND2X2_135
timestamp 1516325494
transform -1 0 2879 0 1 1928
box 0 0 8 49
use AND2X2  AND2X2_135
timestamp 1516325494
transform -1 0 2898 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_559
timestamp 1516325494
transform 1 0 2898 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_559
timestamp 1516325494
transform 1 0 2905 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_1587
timestamp 1516325494
transform -1 0 2939 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_347
timestamp 1516325494
transform 1 0 2939 0 1 1928
box 0 0 53 49
use FILL  FILL_BUFX2_534
timestamp 1516325494
transform 1 0 2993 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_534
timestamp 1516325494
transform 1 0 3000 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_768
timestamp 1516325494
transform 1 0 3015 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_768
timestamp 1516325494
transform 1 0 3023 0 1 1928
box 0 0 15 49
use OR2X2  OR2X2_955
timestamp 1516325494
transform 1 0 3038 0 1 1928
box 0 0 19 49
use AOI21X1  AOI21X1_54
timestamp 1516325494
transform 1 0 3057 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1205
timestamp 1516325494
transform 1 0 3076 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_365
timestamp 1516325494
transform 1 0 3095 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_1207
timestamp 1516325494
transform -1 0 3129 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1208
timestamp 1516325494
transform 1 0 3129 0 1 1928
box 0 0 19 49
use INVX1  INVX1_270
timestamp 1516325494
transform 1 0 3148 0 1 1928
box 0 0 11 49
use OR2X2  OR2X2_954
timestamp 1516325494
transform 1 0 3160 0 1 1928
box 0 0 19 49
use OR2X2  OR2X2_956
timestamp 1516325494
transform 1 0 3179 0 1 1928
box 0 0 19 49
use AND2X2  AND2X2_1196
timestamp 1516325494
transform 1 0 3198 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_231
timestamp 1516325494
transform -1 0 3225 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_231
timestamp 1516325494
transform -1 0 3239 0 1 1928
box 0 0 15 49
use NOR2X1  NOR2X1_140
timestamp 1516325494
transform 1 0 3240 0 1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_789
timestamp 1516325494
transform -1 0 3308 0 1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_788
timestamp 1516325494
transform -1 0 3323 0 1 1928
box 0 0 15 49
use OAI21X1  OAI21X1_136
timestamp 1516325494
transform 1 0 3323 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_848
timestamp 1516325494
transform 1 0 3342 0 1 1928
box 0 0 15 49
use OAI21X1  OAI21X1_137
timestamp 1516325494
transform 1 0 3357 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_847
timestamp 1516325494
transform -1 0 3391 0 1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_846
timestamp 1516325494
transform 1 0 3392 0 1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_610
timestamp 1516325494
transform 1 0 3407 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_610
timestamp 1516325494
transform 1 0 3414 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_1213
timestamp 1516325494
transform -1 0 3449 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_863
timestamp 1516325494
transform -1 0 3464 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_1216
timestamp 1516325494
transform -1 0 3483 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_806
timestamp 1516325494
transform 1 0 3483 0 1 1928
box 0 0 53 49
use AND2X2  AND2X2_1256
timestamp 1516325494
transform 1 0 3536 0 1 1928
box 0 0 19 49
use AOI21X1  AOI21X1_62
timestamp 1516325494
transform 1 0 3555 0 1 1928
box 0 0 19 49
use AOI22X1  AOI22X1_33
timestamp 1516325494
transform 1 0 3574 0 1 1928
box 0 0 23 49
use AND2X2  AND2X2_1222
timestamp 1516325494
transform 1 0 3597 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_824
timestamp 1516325494
transform -1 0 3669 0 1 1928
box 0 0 53 49
use AND2X2  AND2X2_1219
timestamp 1516325494
transform 1 0 3669 0 1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_862
timestamp 1516325494
transform -1 0 3703 0 1 1928
box 0 0 15 49
use AOI21X1  AOI21X1_64
timestamp 1516325494
transform 1 0 3703 0 1 1928
box 0 0 19 49
use NOR2X1  NOR2X1_152
timestamp 1516325494
transform -1 0 3737 0 1 1928
box 0 0 15 49
use AND2X2  AND2X2_1203
timestamp 1516325494
transform -1 0 3756 0 1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_101
timestamp 1516325494
transform -1 0 3764 0 1 1928
box 0 0 8 49
use BUFX2  BUFX2_101
timestamp 1516325494
transform -1 0 3779 0 1 1928
box 0 0 15 49
use OAI21X1  OAI21X1_154
timestamp 1516325494
transform 1 0 3779 0 1 1928
box 0 0 19 49
use OAI21X1  OAI21X1_155
timestamp 1516325494
transform 1 0 3798 0 1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_830
timestamp 1516325494
transform 1 0 3817 0 1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_914
timestamp 1516325494
transform -1 0 2457 0 -1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_356
timestamp 1516325494
transform -1 0 2510 0 -1 1928
box 0 0 53 49
use FILL  FILL_BUFX2_185
timestamp 1516325494
transform 1 0 2510 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_185
timestamp 1516325494
transform 1 0 2518 0 -1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_97
timestamp 1516325494
transform 1 0 2533 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_97
timestamp 1516325494
transform 1 0 2540 0 -1 1928
box 0 0 15 49
use AND2X2  AND2X2_1390
timestamp 1516325494
transform -1 0 2575 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1122
timestamp 1516325494
transform -1 0 2594 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_164
timestamp 1516325494
transform 1 0 2594 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_164
timestamp 1516325494
transform -1 0 2639 0 -1 1928
box 0 0 30 49
use NAND2X1  NAND2X1_60
timestamp 1516325494
transform -1 0 2654 0 -1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_219
timestamp 1516325494
transform -1 0 2662 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_219
timestamp 1516325494
transform -1 0 2677 0 -1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_538
timestamp 1516325494
transform -1 0 2685 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_538
timestamp 1516325494
transform -1 0 2700 0 -1 1928
box 0 0 15 49
use FILL  FILL_OR2X2_241
timestamp 1516325494
transform -1 0 2708 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_241
timestamp 1516325494
transform -1 0 2727 0 -1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_775
timestamp 1516325494
transform -1 0 2735 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_775
timestamp 1516325494
transform -1 0 2749 0 -1 1928
box 0 0 15 49
use OR2X2  OR2X2_1616
timestamp 1516325494
transform -1 0 2768 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1769
timestamp 1516325494
transform -1 0 2787 0 -1 1928
box 0 0 19 49
use AND2X2  AND2X2_1768
timestamp 1516325494
transform -1 0 2806 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_602
timestamp 1516325494
transform -1 0 2821 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_602
timestamp 1516325494
transform -1 0 2852 0 -1 1928
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_282
timestamp 1516325494
transform -1 0 2905 0 -1 1928
box 0 0 53 49
use FILL  FILL_OR2X2_240
timestamp 1516325494
transform -1 0 2913 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_240
timestamp 1516325494
transform -1 0 2932 0 -1 1928
box 0 0 19 49
use FILL  FILL_AND2X2_254
timestamp 1516325494
transform -1 0 2940 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_254
timestamp 1516325494
transform -1 0 2958 0 -1 1928
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_250
timestamp 1516325494
transform 1 0 2958 0 -1 1928
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_141
timestamp 1516325494
transform 1 0 3012 0 -1 1928
box 0 0 53 49
use NAND2X1  NAND2X1_269
timestamp 1516325494
transform 1 0 3065 0 -1 1928
box 0 0 15 49
use MUX2X1  MUX2X1_269
timestamp 1516325494
transform -1 0 3110 0 -1 1928
box 0 0 30 49
use MUX2X1  MUX2X1_365
timestamp 1516325494
transform -1 0 3140 0 -1 1928
box 0 0 30 49
use INVX1  INVX1_278
timestamp 1516325494
transform -1 0 3152 0 -1 1928
box 0 0 11 49
use XNOR2X1  XNOR2X1_57
timestamp 1516325494
transform 1 0 3152 0 -1 1928
box 0 0 34 49
use FILL  FILL_BUFX2_209
timestamp 1516325494
transform -1 0 3194 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_209
timestamp 1516325494
transform -1 0 3209 0 -1 1928
box 0 0 15 49
use FILL  FILL_OR2X2_239
timestamp 1516325494
transform -1 0 3217 0 -1 1928
box 0 0 8 49
use OR2X2  OR2X2_239
timestamp 1516325494
transform -1 0 3236 0 -1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_204
timestamp 1516325494
transform 1 0 3236 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_204
timestamp 1516325494
transform 1 0 3243 0 -1 1928
box 0 0 15 49
use FILL  FILL_AND2X2_255
timestamp 1516325494
transform -1 0 3267 0 -1 1928
box 0 0 8 49
use AND2X2  AND2X2_255
timestamp 1516325494
transform -1 0 3285 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_790
timestamp 1516325494
transform 1 0 3285 0 -1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_348
timestamp 1516325494
transform 1 0 3300 0 -1 1928
box 0 0 53 49
use FILL  FILL_BUFX2_521
timestamp 1516325494
transform 1 0 3354 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_521
timestamp 1516325494
transform 1 0 3361 0 -1 1928
box 0 0 15 49
use AND2X2  AND2X2_1255
timestamp 1516325494
transform 1 0 3376 0 -1 1928
box 0 0 19 49
use OAI21X1  OAI21X1_138
timestamp 1516325494
transform 1 0 3395 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_990
timestamp 1516325494
transform -1 0 3433 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_791
timestamp 1516325494
transform -1 0 3448 0 -1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_787
timestamp 1516325494
transform 1 0 3449 0 -1 1928
box 0 0 15 49
use AOI22X1  AOI22X1_7
timestamp 1516325494
transform 1 0 3464 0 -1 1928
box 0 0 23 49
use AND2X2  AND2X2_1185
timestamp 1516325494
transform 1 0 3487 0 -1 1928
box 0 0 19 49
use FILL  FILL_BUFX2_611
timestamp 1516325494
transform -1 0 3514 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_611
timestamp 1516325494
transform -1 0 3528 0 -1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_796
timestamp 1516325494
transform 1 0 3528 0 -1 1928
box 0 0 15 49
use NOR3X1  NOR3X1_31
timestamp 1516325494
transform 1 0 3544 0 -1 1928
box 0 0 19 49
use OAI21X1  OAI21X1_140
timestamp 1516325494
transform -1 0 3582 0 -1 1928
box 0 0 19 49
use OAI21X1  OAI21X1_139
timestamp 1516325494
transform -1 0 3601 0 -1 1928
box 0 0 19 49
use OR2X2  OR2X2_1002
timestamp 1516325494
transform 1 0 3601 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_850
timestamp 1516325494
transform -1 0 3635 0 -1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_776
timestamp 1516325494
transform 1 0 3635 0 -1 1928
box 0 0 15 49
use AOI21X1  AOI21X1_49
timestamp 1516325494
transform 1 0 3650 0 -1 1928
box 0 0 19 49
use NOR3X1  NOR3X1_32
timestamp 1516325494
transform 1 0 3669 0 -1 1928
box 0 0 19 49
use NAND2X1  NAND2X1_849
timestamp 1516325494
transform -1 0 3703 0 -1 1928
box 0 0 15 49
use AOI22X1  AOI22X1_9
timestamp 1516325494
transform 1 0 3703 0 -1 1928
box 0 0 23 49
use NAND2X1  NAND2X1_866
timestamp 1516325494
transform -1 0 3741 0 -1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_244
timestamp 1516325494
transform -1 0 3749 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_244
timestamp 1516325494
transform -1 0 3764 0 -1 1928
box 0 0 15 49
use FILL  FILL_BUFX2_102
timestamp 1516325494
transform -1 0 3772 0 -1 1928
box 0 0 8 49
use BUFX2  BUFX2_102
timestamp 1516325494
transform -1 0 3787 0 -1 1928
box 0 0 15 49
use NAND2X1  NAND2X1_861
timestamp 1516325494
transform 1 0 3787 0 -1 1928
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_814
timestamp 1516325494
transform 1 0 3802 0 -1 1928
box 0 0 53 49
use FILL  FILL_39_1
timestamp 1516325494
transform -1 0 3863 0 -1 1928
box 0 0 8 49
use FILL  FILL_39_2
timestamp 1516325494
transform -1 0 3871 0 -1 1928
box 0 0 8 49
use FILL  FILL_BUFX2_59
timestamp 1516325494
transform 1 0 1682 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_59
timestamp 1516325494
transform 1 0 1689 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_510
timestamp 1516325494
transform 1 0 1704 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_510
timestamp 1516325494
transform 1 0 1712 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_1924
timestamp 1516325494
transform -1 0 1746 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_807
timestamp 1516325494
transform 1 0 1746 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_807
timestamp 1516325494
transform 1 0 1754 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_845
timestamp 1516325494
transform 1 0 1769 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_845
timestamp 1516325494
transform 1 0 1777 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_1937
timestamp 1516325494
transform -1 0 1811 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1368
timestamp 1516325494
transform 1 0 1811 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_130
timestamp 1516325494
transform 1 0 1830 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_130
timestamp 1516325494
transform 1 0 1837 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_133
timestamp 1516325494
transform 1 0 1853 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_133
timestamp 1516325494
transform 1 0 1860 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_1096
timestamp 1516325494
transform 1 0 1875 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1370
timestamp 1516325494
transform -1 0 1913 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_365
timestamp 1516325494
transform 1 0 1913 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_365
timestamp 1516325494
transform 1 0 1921 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_141
timestamp 1516325494
transform 1 0 1936 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_141
timestamp 1516325494
transform 1 0 1944 0 1 1830
box 0 0 15 49
use AND2X2  AND2X2_1773
timestamp 1516325494
transform -1 0 1978 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1621
timestamp 1516325494
transform -1 0 1997 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1622
timestamp 1516325494
transform -1 0 2016 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_60
timestamp 1516325494
transform -1 0 2024 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_60
timestamp 1516325494
transform -1 0 2039 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_806
timestamp 1516325494
transform -1 0 2047 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_806
timestamp 1516325494
transform -1 0 2061 0 1 1830
box 0 0 15 49
use FILL  FILL_AND2X2_4
timestamp 1516325494
transform -1 0 2070 0 1 1830
box 0 0 8 49
use AND2X2  AND2X2_4
timestamp 1516325494
transform -1 0 2088 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1387
timestamp 1516325494
transform 1 0 2088 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1386
timestamp 1516325494
transform -1 0 2126 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1116
timestamp 1516325494
transform -1 0 2145 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_882
timestamp 1516325494
transform 1 0 2145 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_827
timestamp 1516325494
transform -1 0 2190 0 1 1830
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_437
timestamp 1516325494
transform 1 0 2191 0 1 1830
box 0 0 53 49
use NAND2X1  NAND2X1_405
timestamp 1516325494
transform 1 0 2244 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_405
timestamp 1516325494
transform -1 0 2289 0 1 1830
box 0 0 30 49
use FILL  FILL_BUFX2_721
timestamp 1516325494
transform -1 0 2298 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_721
timestamp 1516325494
transform -1 0 2312 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_440
timestamp 1516325494
transform 1 0 2312 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_440
timestamp 1516325494
transform 1 0 2320 0 1 1830
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_703
timestamp 1516325494
transform 1 0 2335 0 1 1830
box 0 0 53 49
use NAND2X1  NAND2X1_319
timestamp 1516325494
transform 1 0 2388 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_319
timestamp 1516325494
transform -1 0 2434 0 1 1830
box 0 0 30 49
use FILL  FILL_BUFX2_432
timestamp 1516325494
transform 1 0 2434 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_432
timestamp 1516325494
transform 1 0 2442 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_844
timestamp 1516325494
transform 1 0 2457 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_844
timestamp 1516325494
transform 1 0 2464 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_644
timestamp 1516325494
transform 1 0 2480 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_644
timestamp 1516325494
transform 1 0 2487 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_57
timestamp 1516325494
transform -1 0 2510 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_57
timestamp 1516325494
transform -1 0 2525 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_291
timestamp 1516325494
transform -1 0 2533 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_291
timestamp 1516325494
transform -1 0 2548 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_16
timestamp 1516325494
transform 1 0 2548 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_16
timestamp 1516325494
transform 1 0 2556 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_26
timestamp 1516325494
transform -1 0 2579 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_26
timestamp 1516325494
transform -1 0 2593 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_99
timestamp 1516325494
transform -1 0 2602 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_99
timestamp 1516325494
transform -1 0 2616 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_319
timestamp 1516325494
transform -1 0 2624 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_319
timestamp 1516325494
transform -1 0 2639 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_311
timestamp 1516325494
transform -1 0 2658 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_308
timestamp 1516325494
transform -1 0 2677 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1620
timestamp 1516325494
transform -1 0 2696 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1617
timestamp 1516325494
transform -1 0 2715 0 1 1830
box 0 0 19 49
use FILL  FILL_OR2X2_238
timestamp 1516325494
transform -1 0 2723 0 1 1830
box 0 0 8 49
use OR2X2  OR2X2_238
timestamp 1516325494
transform -1 0 2742 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_1770
timestamp 1516325494
transform -1 0 2761 0 1 1830
box 0 0 19 49
use FILL  FILL_OR2X2_237
timestamp 1516325494
transform -1 0 2769 0 1 1830
box 0 0 8 49
use OR2X2  OR2X2_237
timestamp 1516325494
transform -1 0 2787 0 1 1830
box 0 0 19 49
use FILL  FILL_AND2X2_253
timestamp 1516325494
transform -1 0 2795 0 1 1830
box 0 0 8 49
use AND2X2  AND2X2_253
timestamp 1516325494
transform -1 0 2814 0 1 1830
box 0 0 19 49
use OR2X2  OR2X2_307
timestamp 1516325494
transform -1 0 2833 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_328
timestamp 1516325494
transform -1 0 2852 0 1 1830
box 0 0 19 49
use FILL  FILL_AND2X2_252
timestamp 1516325494
transform -1 0 2860 0 1 1830
box 0 0 8 49
use AND2X2  AND2X2_252
timestamp 1516325494
transform -1 0 2879 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_600
timestamp 1516325494
transform 1 0 2879 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_600
timestamp 1516325494
transform 1 0 2886 0 1 1830
box 0 0 15 49
use AND2X2  AND2X2_327
timestamp 1516325494
transform -1 0 2920 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_395
timestamp 1516325494
transform 1 0 2920 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_395
timestamp 1516325494
transform 1 0 2928 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_110
timestamp 1516325494
transform 1 0 2943 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_110
timestamp 1516325494
transform 1 0 2951 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_1830
timestamp 1516325494
transform -1 0 2985 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_604
timestamp 1516325494
transform -1 0 3000 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_604
timestamp 1516325494
transform -1 0 3030 0 1 1830
box 0 0 30 49
use MUX2X1  MUX2X1_218
timestamp 1516325494
transform -1 0 3061 0 1 1830
box 0 0 30 49
use FILL  FILL_BUFX2_617
timestamp 1516325494
transform 1 0 3061 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_617
timestamp 1516325494
transform 1 0 3069 0 1 1830
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_333
timestamp 1516325494
transform 1 0 3084 0 1 1830
box 0 0 53 49
use FILL  FILL_BUFX2_280
timestamp 1516325494
transform -1 0 3145 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_280
timestamp 1516325494
transform -1 0 3160 0 1 1830
box 0 0 15 49
use FILL  FILL_BUFX2_656
timestamp 1516325494
transform 1 0 3160 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_656
timestamp 1516325494
transform 1 0 3167 0 1 1830
box 0 0 15 49
use OR2X2  OR2X2_1829
timestamp 1516325494
transform -1 0 3202 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1931
timestamp 1516325494
transform -1 0 3221 0 1 1830
box 0 0 19 49
use FILL  FILL_AND2X2_256
timestamp 1516325494
transform -1 0 3229 0 1 1830
box 0 0 8 49
use AND2X2  AND2X2_256
timestamp 1516325494
transform -1 0 3247 0 1 1830
box 0 0 19 49
use FILL  FILL_BUFX2_326
timestamp 1516325494
transform 1 0 3247 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_326
timestamp 1516325494
transform 1 0 3255 0 1 1830
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_149
timestamp 1516325494
transform 1 0 3270 0 1 1830
box 0 0 53 49
use OR2X2  OR2X2_1828
timestamp 1516325494
transform -1 0 3342 0 1 1830
box 0 0 19 49
use AND2X2  AND2X2_1933
timestamp 1516325494
transform -1 0 3361 0 1 1830
box 0 0 19 49
use MUX2X1  MUX2X1_380
timestamp 1516325494
transform 1 0 3361 0 1 1830
box 0 0 30 49
use NAND2X1  NAND2X1_380
timestamp 1516325494
transform 1 0 3392 0 1 1830
box 0 0 15 49
use AND2X2  AND2X2_361
timestamp 1516325494
transform -1 0 3426 0 1 1830
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_823
timestamp 1516325494
transform -1 0 3479 0 1 1830
box 0 0 53 49
use FILL  FILL_BUFX2_536
timestamp 1516325494
transform 1 0 3479 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_536
timestamp 1516325494
transform 1 0 3487 0 1 1830
box 0 0 15 49
use MUX2X1  MUX2X1_383
timestamp 1516325494
transform 1 0 3502 0 1 1830
box 0 0 30 49
use OAI21X1  OAI21X1_156
timestamp 1516325494
transform 1 0 3532 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_865
timestamp 1516325494
transform 1 0 3551 0 1 1830
box 0 0 15 49
use OAI21X1  OAI21X1_157
timestamp 1516325494
transform -1 0 3585 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_864
timestamp 1516325494
transform -1 0 3600 0 1 1830
box 0 0 15 49
use AND2X2  AND2X2_1270
timestamp 1516325494
transform 1 0 3601 0 1 1830
box 0 0 19 49
use AOI21X1  AOI21X1_65
timestamp 1516325494
transform 1 0 3620 0 1 1830
box 0 0 19 49
use OAI21X1  OAI21X1_159
timestamp 1516325494
transform 1 0 3639 0 1 1830
box 0 0 19 49
use AOI22X1  AOI22X1_34
timestamp 1516325494
transform -1 0 3681 0 1 1830
box 0 0 23 49
use AND2X2  AND2X2_1271
timestamp 1516325494
transform -1 0 3699 0 1 1830
box 0 0 19 49
use OAI21X1  OAI21X1_160
timestamp 1516325494
transform 1 0 3699 0 1 1830
box 0 0 19 49
use NAND2X1  NAND2X1_867
timestamp 1516325494
transform -1 0 3733 0 1 1830
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_816
timestamp 1516325494
transform -1 0 3787 0 1 1830
box 0 0 53 49
use FILL  FILL_BUFX2_522
timestamp 1516325494
transform 1 0 3787 0 1 1830
box 0 0 8 49
use BUFX2  BUFX2_522
timestamp 1516325494
transform 1 0 3794 0 1 1830
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_790
timestamp 1516325494
transform 1 0 3810 0 1 1830
box 0 0 53 49
use FILL  FILL_38_1
timestamp 1516325494
transform 1 0 3863 0 1 1830
box 0 0 8 49
use INVX1  INVX1_180
timestamp 1516325494
transform -1 0 13 0 -1 1829
box 0 0 11 49
use INVX1  INVX1_86
timestamp 1516325494
transform 1 0 13 0 -1 1829
box 0 0 11 49
use AND2X2  AND2X2_1098
timestamp 1516325494
transform 1 0 25 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_893
timestamp 1516325494
transform -1 0 63 0 -1 1829
box 0 0 19 49
use INVX1  INVX1_81
timestamp 1516325494
transform -1 0 74 0 -1 1829
box 0 0 11 49
use XOR2X1  XOR2X1_43
timestamp 1516325494
transform -1 0 108 0 -1 1829
box 0 0 34 49
use INVX1  INVX1_77
timestamp 1516325494
transform -1 0 119 0 -1 1829
box 0 0 11 49
use INVX1  INVX1_75
timestamp 1516325494
transform 1 0 120 0 -1 1829
box 0 0 11 49
use XOR2X1  XOR2X1_41
timestamp 1516325494
transform -1 0 165 0 -1 1829
box 0 0 34 49
use OR2X2  OR2X2_771
timestamp 1516325494
transform 1 0 165 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_844
timestamp 1516325494
transform -1 0 203 0 -1 1829
box 0 0 19 49
use NOR2X1  NOR2X1_45
timestamp 1516325494
transform -1 0 218 0 -1 1829
box 0 0 15 49
use AND2X2  AND2X2_1011
timestamp 1516325494
transform -1 0 238 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1010
timestamp 1516325494
transform -1 0 257 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1009
timestamp 1516325494
transform -1 0 276 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_840
timestamp 1516325494
transform -1 0 295 0 -1 1829
box 0 0 19 49
use NOR2X1  NOR2X1_73
timestamp 1516325494
transform -1 0 310 0 -1 1829
box 0 0 15 49
use NAND3X1  NAND3X1_54
timestamp 1516325494
transform -1 0 329 0 -1 1829
box 0 0 19 49
use NAND3X1  NAND3X1_49
timestamp 1516325494
transform -1 0 348 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_907
timestamp 1516325494
transform -1 0 367 0 -1 1829
box 0 0 19 49
use NAND3X1  NAND3X1_50
timestamp 1516325494
transform -1 0 386 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_931
timestamp 1516325494
transform -1 0 405 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_909
timestamp 1516325494
transform 1 0 405 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_780
timestamp 1516325494
transform -1 0 443 0 -1 1829
box 0 0 19 49
use FILL  FILL_BUFX2_639
timestamp 1516325494
transform -1 0 451 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_639
timestamp 1516325494
transform -1 0 465 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_699
timestamp 1516325494
transform 1 0 466 0 -1 1829
box 0 0 19 49
use XOR2X1  XOR2X1_18
timestamp 1516325494
transform -1 0 519 0 -1 1829
box 0 0 34 49
use OR2X2  OR2X2_762
timestamp 1516325494
transform 1 0 519 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_793
timestamp 1516325494
transform -1 0 557 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1080
timestamp 1516325494
transform 1 0 557 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_794
timestamp 1516325494
transform -1 0 595 0 -1 1829
box 0 0 19 49
use OAI21X1  OAI21X1_69
timestamp 1516325494
transform -1 0 614 0 -1 1829
box 0 0 19 49
use OAI21X1  OAI21X1_67
timestamp 1516325494
transform -1 0 633 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1079
timestamp 1516325494
transform 1 0 633 0 -1 1829
box 0 0 19 49
use INVX1  INVX1_39
timestamp 1516325494
transform 1 0 652 0 -1 1829
box 0 0 11 49
use AND2X2  AND2X2_1095
timestamp 1516325494
transform -1 0 682 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_890
timestamp 1516325494
transform -1 0 701 0 -1 1829
box 0 0 19 49
use XOR2X1  XOR2X1_40
timestamp 1516325494
transform -1 0 735 0 -1 1829
box 0 0 34 49
use INVX1  INVX1_73
timestamp 1516325494
transform -1 0 746 0 -1 1829
box 0 0 11 49
use FILL  FILL_BUFX2_853
timestamp 1516325494
transform 1 0 747 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_853
timestamp 1516325494
transform 1 0 754 0 -1 1829
box 0 0 15 49
use INVX1  INVX1_85
timestamp 1516325494
transform -1 0 13 0 1 1731
box 0 0 11 49
use NOR2X1  NOR2X1_89
timestamp 1516325494
transform -1 0 28 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_894
timestamp 1516325494
transform -1 0 48 0 1 1731
box 0 0 19 49
use XOR2X1  XOR2X1_44
timestamp 1516325494
transform -1 0 82 0 1 1731
box 0 0 34 49
use XNOR2X1  XNOR2X1_17
timestamp 1516325494
transform -1 0 116 0 1 1731
box 0 0 34 49
use NOR2X1  NOR2X1_86
timestamp 1516325494
transform -1 0 131 0 1 1731
box 0 0 15 49
use XNOR2X1  XNOR2X1_16
timestamp 1516325494
transform -1 0 165 0 1 1731
box 0 0 34 49
use AND2X2  AND2X2_845
timestamp 1516325494
transform -1 0 184 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_713
timestamp 1516325494
transform -1 0 203 0 1 1731
box 0 0 19 49
use AOI21X1  AOI21X1_11
timestamp 1516325494
transform -1 0 222 0 1 1731
box 0 0 19 49
use NAND2X1  NAND2X1_667
timestamp 1516325494
transform -1 0 237 0 1 1731
box 0 0 15 49
use NAND2X1  NAND2X1_666
timestamp 1516325494
transform -1 0 253 0 1 1731
box 0 0 15 49
use NAND2X1  NAND2X1_646
timestamp 1516325494
transform -1 0 268 0 1 1731
box 0 0 15 49
use XOR2X1  XOR2X1_6
timestamp 1516325494
transform 1 0 268 0 1 1731
box 0 0 34 49
use AND2X2  AND2X2_649
timestamp 1516325494
transform 1 0 302 0 1 1731
box 0 0 19 49
use OAI21X1  OAI21X1_2
timestamp 1516325494
transform 1 0 321 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_551
timestamp 1516325494
transform -1 0 359 0 1 1731
box 0 0 19 49
use NAND2X1  NAND2X1_654
timestamp 1516325494
transform -1 0 374 0 1 1731
box 0 0 15 49
use AND2X2  AND2X2_472
timestamp 1516325494
transform 1 0 374 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_561
timestamp 1516325494
transform 1 0 393 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_561
timestamp 1516325494
transform 1 0 401 0 1 1731
box 0 0 15 49
use AND2X2  AND2X2_932
timestamp 1516325494
transform -1 0 435 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_742
timestamp 1516325494
transform -1 0 443 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_742
timestamp 1516325494
transform -1 0 458 0 1 1731
box 0 0 15 49
use NAND3X1  NAND3X1_43
timestamp 1516325494
transform 1 0 458 0 1 1731
box 0 0 19 49
use NAND3X1  NAND3X1_44
timestamp 1516325494
transform -1 0 496 0 1 1731
box 0 0 19 49
use NAND2X1  NAND2X1_672
timestamp 1516325494
transform 1 0 496 0 1 1731
box 0 0 15 49
use NAND2X1  NAND2X1_671
timestamp 1516325494
transform -1 0 526 0 1 1731
box 0 0 15 49
use FILL  FILL_BUFX2_563
timestamp 1516325494
transform -1 0 534 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_563
timestamp 1516325494
transform -1 0 549 0 1 1731
box 0 0 15 49
use NOR2X1  NOR2X1_82
timestamp 1516325494
transform 1 0 549 0 1 1731
box 0 0 15 49
use INVX1  INVX1_65
timestamp 1516325494
transform 1 0 564 0 1 1731
box 0 0 11 49
use OR2X2  OR2X2_653
timestamp 1516325494
transform -1 0 595 0 1 1731
box 0 0 19 49
use AOI21X1  AOI21X1_7
timestamp 1516325494
transform -1 0 614 0 1 1731
box 0 0 19 49
use OAI21X1  OAI21X1_65
timestamp 1516325494
transform -1 0 633 0 1 1731
box 0 0 19 49
use INVX1  INVX1_40
timestamp 1516325494
transform 1 0 633 0 1 1731
box 0 0 11 49
use AND2X2  AND2X2_1091
timestamp 1516325494
transform -1 0 663 0 1 1731
box 0 0 19 49
use NAND2X1  NAND2X1_712
timestamp 1516325494
transform -1 0 678 0 1 1731
box 0 0 15 49
use NAND2X1  NAND2X1_711
timestamp 1516325494
transform -1 0 693 0 1 1731
box 0 0 15 49
use NOR2X1  NOR2X1_81
timestamp 1516325494
transform -1 0 709 0 1 1731
box 0 0 15 49
use INVX1  INVX1_62
timestamp 1516325494
transform -1 0 720 0 1 1731
box 0 0 11 49
use XNOR2X1  XNOR2X1_12
timestamp 1516325494
transform 1 0 720 0 1 1731
box 0 0 34 49
use NOR2X1  NOR2X1_84
timestamp 1516325494
transform 1 0 754 0 1 1731
box 0 0 15 49
use INVX1  INVX1_25
timestamp 1516325494
transform -1 0 781 0 -1 1829
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_737
timestamp 1516325494
transform -1 0 834 0 -1 1829
box 0 0 53 49
use INVX1  INVX1_36
timestamp 1516325494
transform 1 0 834 0 -1 1829
box 0 0 11 49
use INVX1  INVX1_159
timestamp 1516325494
transform 1 0 846 0 -1 1829
box 0 0 11 49
use MUX2X1  MUX2X1_760
timestamp 1516325494
transform 1 0 857 0 -1 1829
box 0 0 30 49
use INVX1  INVX1_148
timestamp 1516325494
transform 1 0 887 0 -1 1829
box 0 0 11 49
use INVX1  INVX1_71
timestamp 1516325494
transform 1 0 770 0 1 1731
box 0 0 11 49
use AND2X2  AND2X2_1094
timestamp 1516325494
transform -1 0 800 0 1 1731
box 0 0 19 49
use XNOR2X1  XNOR2X1_13
timestamp 1516325494
transform 1 0 800 0 1 1731
box 0 0 34 49
use DFFPOSX1  DFFPOSX1_732
timestamp 1516325494
transform -1 0 887 0 1 1731
box 0 0 53 49
use INVX1  INVX1_156
timestamp 1516325494
transform 1 0 887 0 1 1731
box 0 0 11 49
use MUX2X1  MUX2X1_791
timestamp 1516325494
transform -1 0 929 0 -1 1829
box 0 0 30 49
use NAND2X1  NAND2X1_89
timestamp 1516325494
transform 1 0 929 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_89
timestamp 1516325494
transform -1 0 974 0 -1 1829
box 0 0 30 49
use OR2X2  OR2X2_1760
timestamp 1516325494
transform 1 0 975 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1233
timestamp 1516325494
transform -1 0 1013 0 -1 1829
box 0 0 19 49
use NAND2X1  NAND2X1_456
timestamp 1516325494
transform 1 0 1013 0 -1 1829
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_552
timestamp 1516325494
transform 1 0 1028 0 -1 1829
box 0 0 53 49
use MUX2X1  MUX2X1_456
timestamp 1516325494
transform -1 0 1111 0 -1 1829
box 0 0 30 49
use MUX2X1  MUX2X1_40
timestamp 1516325494
transform 1 0 1112 0 -1 1829
box 0 0 30 49
use NAND2X1  NAND2X1_40
timestamp 1516325494
transform -1 0 1157 0 -1 1829
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_648
timestamp 1516325494
transform -1 0 1210 0 -1 1829
box 0 0 53 49
use OR2X2  OR2X2_1238
timestamp 1516325494
transform -1 0 1229 0 -1 1829
box 0 0 19 49
use FILL  FILL_BUFX2_686
timestamp 1516325494
transform -1 0 1237 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_686
timestamp 1516325494
transform -1 0 1252 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_1535
timestamp 1516325494
transform -1 0 1271 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1705
timestamp 1516325494
transform -1 0 1290 0 -1 1829
box 0 0 19 49
use FILL  FILL_OR2X2_200
timestamp 1516325494
transform -1 0 1298 0 -1 1829
box 0 0 8 49
use OR2X2  OR2X2_200
timestamp 1516325494
transform -1 0 1317 0 -1 1829
box 0 0 19 49
use FILL  FILL_AND2X2_212
timestamp 1516325494
transform -1 0 1325 0 -1 1829
box 0 0 8 49
use AND2X2  AND2X2_212
timestamp 1516325494
transform -1 0 1343 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_82
timestamp 1516325494
transform 1 0 1343 0 -1 1829
box 0 0 53 49
use MUX2X1  MUX2X1_146
timestamp 1516325494
transform -1 0 1427 0 -1 1829
box 0 0 30 49
use NAND2X1  NAND2X1_146
timestamp 1516325494
transform 1 0 1427 0 -1 1829
box 0 0 15 49
use AND2X2  AND2X2_1708
timestamp 1516325494
transform -1 0 1461 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1536
timestamp 1516325494
transform -1 0 1480 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_626
timestamp 1516325494
transform 1 0 1480 0 -1 1829
box 0 0 53 49
use NAND2X1  NAND2X1_896
timestamp 1516325494
transform 1 0 1533 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_841
timestamp 1516325494
transform -1 0 1579 0 -1 1829
box 0 0 30 49
use NAND2X1  NAND2X1_63
timestamp 1516325494
transform 1 0 1579 0 -1 1829
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_671
timestamp 1516325494
transform 1 0 1594 0 -1 1829
box 0 0 53 49
use MUX2X1  MUX2X1_63
timestamp 1516325494
transform -1 0 1677 0 -1 1829
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_629
timestamp 1516325494
transform 1 0 1678 0 -1 1829
box 0 0 53 49
use NAND2X1  NAND2X1_899
timestamp 1516325494
transform 1 0 1731 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_844
timestamp 1516325494
transform -1 0 1776 0 -1 1829
box 0 0 30 49
use AND2X2  AND2X2_1374
timestamp 1516325494
transform 1 0 1777 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_2107
timestamp 1516325494
transform 1 0 1796 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_67
timestamp 1516325494
transform 1 0 1815 0 -1 1829
box 0 0 53 49
use MUX2X1  MUX2X1_131
timestamp 1516325494
transform -1 0 1898 0 -1 1829
box 0 0 30 49
use NAND2X1  NAND2X1_131
timestamp 1516325494
transform -1 0 1913 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_2013
timestamp 1516325494
transform 1 0 1913 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1101
timestamp 1516325494
transform 1 0 1932 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1102
timestamp 1516325494
transform 1 0 1951 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_2104
timestamp 1516325494
transform 1 0 1970 0 -1 1829
box 0 0 19 49
use FILL  FILL_BUFX2_643
timestamp 1516325494
transform 1 0 1989 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_643
timestamp 1516325494
transform 1 0 1997 0 -1 1829
box 0 0 15 49
use FILL  FILL_BUFX2_683
timestamp 1516325494
transform -1 0 2020 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_683
timestamp 1516325494
transform -1 0 2035 0 -1 1829
box 0 0 15 49
use FILL  FILL_BUFX2_819
timestamp 1516325494
transform -1 0 2043 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_819
timestamp 1516325494
transform -1 0 2058 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_2010
timestamp 1516325494
transform -1 0 2077 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_2102
timestamp 1516325494
transform -1 0 2096 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_2103
timestamp 1516325494
transform -1 0 2115 0 -1 1829
box 0 0 19 49
use FILL  FILL_OR2X2_10
timestamp 1516325494
transform 1 0 2115 0 -1 1829
box 0 0 8 49
use OR2X2  OR2X2_10
timestamp 1516325494
transform 1 0 2122 0 -1 1829
box 0 0 19 49
use FILL  FILL_OR2X2_6
timestamp 1516325494
transform -1 0 2149 0 -1 1829
box 0 0 8 49
use OR2X2  OR2X2_6
timestamp 1516325494
transform -1 0 2168 0 -1 1829
box 0 0 19 49
use FILL  FILL_OR2X2_5
timestamp 1516325494
transform -1 0 2176 0 -1 1829
box 0 0 8 49
use OR2X2  OR2X2_5
timestamp 1516325494
transform -1 0 2195 0 -1 1829
box 0 0 19 49
use FILL  FILL_AND2X2_5
timestamp 1516325494
transform -1 0 2203 0 -1 1829
box 0 0 8 49
use AND2X2  AND2X2_5
timestamp 1516325494
transform -1 0 2221 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1366
timestamp 1516325494
transform 1 0 2221 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1389
timestamp 1516325494
transform 1 0 2240 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1120
timestamp 1516325494
transform 1 0 2259 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1115
timestamp 1516325494
transform 1 0 2278 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1121
timestamp 1516325494
transform 1 0 2297 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1133
timestamp 1516325494
transform 1 0 2316 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_612
timestamp 1516325494
transform -1 0 2388 0 -1 1829
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_419
timestamp 1516325494
transform -1 0 2441 0 -1 1829
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_579
timestamp 1516325494
transform -1 0 2495 0 -1 1829
box 0 0 53 49
use OAI21X1  OAI21X1_21
timestamp 1516325494
transform 1 0 2495 0 -1 1829
box 0 0 19 49
use INVX2  INVX2_10
timestamp 1516325494
transform 1 0 2514 0 -1 1829
box 0 0 11 49
use AND2X2  AND2X2_1710
timestamp 1516325494
transform -1 0 2544 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1539
timestamp 1516325494
transform -1 0 2563 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1388
timestamp 1516325494
transform -1 0 2582 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1119
timestamp 1516325494
transform -1 0 2601 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1118
timestamp 1516325494
transform -1 0 2620 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1538
timestamp 1516325494
transform -1 0 2639 0 -1 1829
box 0 0 19 49
use FILL  FILL_BUFX2_367
timestamp 1516325494
transform -1 0 2647 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_367
timestamp 1516325494
transform -1 0 2662 0 -1 1829
box 0 0 15 49
use NAND2X1  NAND2X1_484
timestamp 1516325494
transform 1 0 2662 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_484
timestamp 1516325494
transform -1 0 2707 0 -1 1829
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_292
timestamp 1516325494
transform -1 0 2761 0 -1 1829
box 0 0 53 49
use MUX2X1  MUX2X1_636
timestamp 1516325494
transform 1 0 2761 0 -1 1829
box 0 0 30 49
use NAND2X1  NAND2X1_636
timestamp 1516325494
transform -1 0 2806 0 -1 1829
box 0 0 15 49
use FILL  FILL_BUFX2_441
timestamp 1516325494
transform 1 0 2806 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_441
timestamp 1516325494
transform 1 0 2814 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_306
timestamp 1516325494
transform -1 0 2848 0 -1 1829
box 0 0 19 49
use FILL  FILL_BUFX2_469
timestamp 1516325494
transform -1 0 2856 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_469
timestamp 1516325494
transform -1 0 2871 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_1767
timestamp 1516325494
transform -1 0 2890 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1766
timestamp 1516325494
transform -1 0 2909 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1884
timestamp 1516325494
transform -1 0 2928 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_339
timestamp 1516325494
transform -1 0 2947 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1883
timestamp 1516325494
transform -1 0 2966 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1827
timestamp 1516325494
transform 1 0 2966 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1826
timestamp 1516325494
transform -1 0 3004 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1930
timestamp 1516325494
transform -1 0 3023 0 -1 1829
box 0 0 19 49
use NAND2X1  NAND2X1_218
timestamp 1516325494
transform 1 0 3023 0 -1 1829
box 0 0 15 49
use AND2X2  AND2X2_1929
timestamp 1516325494
transform -1 0 3057 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_284
timestamp 1516325494
transform -1 0 3110 0 -1 1829
box 0 0 53 49
use FILL  FILL_BUFX2_620
timestamp 1516325494
transform -1 0 3118 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_620
timestamp 1516325494
transform -1 0 3133 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_338
timestamp 1516325494
transform -1 0 3152 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_359
timestamp 1516325494
transform -1 0 3171 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_252
timestamp 1516325494
transform -1 0 3224 0 -1 1829
box 0 0 53 49
use OR2X2  OR2X2_1619
timestamp 1516325494
transform -1 0 3243 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1770
timestamp 1516325494
transform -1 0 3262 0 -1 1829
box 0 0 19 49
use AND2X2  AND2X2_1771
timestamp 1516325494
transform 1 0 3262 0 -1 1829
box 0 0 19 49
use OR2X2  OR2X2_1618
timestamp 1516325494
transform -1 0 3300 0 -1 1829
box 0 0 19 49
use NAND2X1  NAND2X1_277
timestamp 1516325494
transform 1 0 3300 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_277
timestamp 1516325494
transform -1 0 3346 0 -1 1829
box 0 0 30 49
use AND2X2  AND2X2_1772
timestamp 1516325494
transform -1 0 3365 0 -1 1829
box 0 0 19 49
use FILL  FILL_BUFX2_658
timestamp 1516325494
transform -1 0 3373 0 -1 1829
box 0 0 8 49
use BUFX2  BUFX2_658
timestamp 1516325494
transform -1 0 3388 0 -1 1829
box 0 0 15 49
use OR2X2  OR2X2_337
timestamp 1516325494
transform -1 0 3407 0 -1 1829
box 0 0 19 49
use NAND2X1  NAND2X1_284
timestamp 1516325494
transform -1 0 3422 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_284
timestamp 1516325494
transform -1 0 3452 0 -1 1829
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_156
timestamp 1516325494
transform -1 0 3505 0 -1 1829
box 0 0 53 49
use NAND2X1  NAND2X1_287
timestamp 1516325494
transform 1 0 3506 0 -1 1829
box 0 0 15 49
use NAND2X1  NAND2X1_383
timestamp 1516325494
transform -1 0 3536 0 -1 1829
box 0 0 15 49
use MUX2X1  MUX2X1_287
timestamp 1516325494
transform -1 0 3566 0 -1 1829
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_351
timestamp 1516325494
transform -1 0 3619 0 -1 1829
box 0 0 53 49
use OAI21X1  OAI21X1_158
timestamp 1516325494
transform 1 0 3620 0 -1 1829
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_801
timestamp 1516325494
transform 1 0 3639 0 -1 1829
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_815
timestamp 1516325494
transform -1 0 3745 0 -1 1829
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_791
timestamp 1516325494
transform -1 0 3798 0 -1 1829
box 0 0 53 49
use AOI21X1  AOI21X1_50
timestamp 1516325494
transform -1 0 3817 0 -1 1829
box 0 0 19 49
use NAND2X1  NAND2X1_777
timestamp 1516325494
transform 1 0 3817 0 -1 1829
box 0 0 15 49
use AND2X2  AND2X2_1192
timestamp 1516325494
transform 1 0 3832 0 -1 1829
box 0 0 19 49
use BUFX2  BUFX2_870
timestamp 1516325494
transform -1 0 3866 0 -1 1829
box 0 0 15 49
use FILL  FILL_BUFX2_777
timestamp 1516325494
transform 1 0 899 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_777
timestamp 1516325494
transform 1 0 906 0 1 1731
box 0 0 15 49
use INVX1  INVX1_213
timestamp 1516325494
transform -1 0 933 0 1 1731
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_697
timestamp 1516325494
transform 1 0 933 0 1 1731
box 0 0 53 49
use MUX2X1  MUX2X1_313
timestamp 1516325494
transform -1 0 1016 0 1 1731
box 0 0 30 49
use OR2X2  OR2X2_1774
timestamp 1516325494
transform 1 0 1017 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1890
timestamp 1516325494
transform 1 0 1036 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1891
timestamp 1516325494
transform 1 0 1055 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1775
timestamp 1516325494
transform -1 0 1093 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_333
timestamp 1516325494
transform 1 0 1093 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_312
timestamp 1516325494
transform -1 0 1131 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_725
timestamp 1516325494
transform -1 0 1184 0 1 1731
box 0 0 53 49
use FILL  FILL_BUFX2_569
timestamp 1516325494
transform 1 0 1184 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_569
timestamp 1516325494
transform 1 0 1191 0 1 1731
box 0 0 15 49
use AND2X2  AND2X2_1894
timestamp 1516325494
transform -1 0 1226 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_780
timestamp 1516325494
transform 1 0 1226 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_780
timestamp 1516325494
transform 1 0 1233 0 1 1731
box 0 0 15 49
use FILL  FILL_BUFX2_275
timestamp 1516325494
transform -1 0 1256 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_275
timestamp 1516325494
transform -1 0 1271 0 1 1731
box 0 0 15 49
use AND2X2  AND2X2_1707
timestamp 1516325494
transform -1 0 1290 0 1 1731
box 0 0 19 49
use FILL  FILL_AND2X2_213
timestamp 1516325494
transform 1 0 1290 0 1 1731
box 0 0 8 49
use AND2X2  AND2X2_213
timestamp 1516325494
transform 1 0 1298 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1892
timestamp 1516325494
transform -1 0 1336 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1776
timestamp 1516325494
transform -1 0 1355 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_634
timestamp 1516325494
transform 1 0 1355 0 1 1731
box 0 0 53 49
use MUX2X1  MUX2X1_849
timestamp 1516325494
transform 1 0 1408 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_904
timestamp 1516325494
transform 1 0 1438 0 1 1731
box 0 0 15 49
use FILL  FILL_BUFX2_169
timestamp 1516325494
transform -1 0 1462 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_169
timestamp 1516325494
transform -1 0 1476 0 1 1731
box 0 0 15 49
use AND2X2  AND2X2_1706
timestamp 1516325494
transform -1 0 1495 0 1 1731
box 0 0 19 49
use MUX2X1  MUX2X1_466
timestamp 1516325494
transform 1 0 1495 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_466
timestamp 1516325494
transform -1 0 1541 0 1 1731
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_562
timestamp 1516325494
transform -1 0 1594 0 1 1731
box 0 0 53 49
use OR2X2  OR2X2_1533
timestamp 1516325494
transform -1 0 1613 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1779
timestamp 1516325494
transform -1 0 1632 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1628
timestamp 1516325494
transform -1 0 1651 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_661
timestamp 1516325494
transform 1 0 1651 0 1 1731
box 0 0 53 49
use NAND2X1  NAND2X1_53
timestamp 1516325494
transform 1 0 1704 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_53
timestamp 1516325494
transform -1 0 1750 0 1 1731
box 0 0 30 49
use OR2X2  OR2X2_1940
timestamp 1516325494
transform -1 0 1769 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_228
timestamp 1516325494
transform 1 0 1769 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_228
timestamp 1516325494
transform 1 0 1777 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_858
timestamp 1516325494
transform -1 0 1822 0 1 1731
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_355
timestamp 1516325494
transform -1 0 1875 0 1 1731
box 0 0 53 49
use NAND2X1  NAND2X1_913
timestamp 1516325494
transform -1 0 1890 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_1092
timestamp 1516325494
transform 1 0 1891 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1367
timestamp 1516325494
transform 1 0 1910 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1537
timestamp 1516325494
transform -1 0 1948 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_2014
timestamp 1516325494
transform 1 0 1948 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_2012
timestamp 1516325494
transform -1 0 1986 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1097
timestamp 1516325494
transform -1 0 2005 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_2015
timestamp 1516325494
transform -1 0 2024 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_2011
timestamp 1516325494
transform -1 0 2043 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_2009
timestamp 1516325494
transform -1 0 2062 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_2100
timestamp 1516325494
transform -1 0 2081 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_276
timestamp 1516325494
transform 1 0 2081 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_276
timestamp 1516325494
transform 1 0 2088 0 1 1731
box 0 0 15 49
use INVX1  INVX1_203
timestamp 1516325494
transform 1 0 2103 0 1 1731
box 0 0 11 49
use FILL  FILL_OR2X2_11
timestamp 1516325494
transform -1 0 2123 0 1 1731
box 0 0 8 49
use OR2X2  OR2X2_11
timestamp 1516325494
transform -1 0 2141 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1360
timestamp 1516325494
transform 1 0 2141 0 1 1731
box 0 0 19 49
use FILL  FILL_OR2X2_4
timestamp 1516325494
transform -1 0 2168 0 1 1731
box 0 0 8 49
use OR2X2  OR2X2_4
timestamp 1516325494
transform -1 0 2187 0 1 1731
box 0 0 19 49
use FILL  FILL_AND2X2_2
timestamp 1516325494
transform -1 0 2195 0 1 1731
box 0 0 8 49
use AND2X2  AND2X2_2
timestamp 1516325494
transform -1 0 2214 0 1 1731
box 0 0 19 49
use FILL  FILL_AND2X2_3
timestamp 1516325494
transform -1 0 2222 0 1 1731
box 0 0 8 49
use AND2X2  AND2X2_3
timestamp 1516325494
transform -1 0 2240 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1385
timestamp 1516325494
transform 1 0 2240 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1383
timestamp 1516325494
transform 1 0 2259 0 1 1731
box 0 0 19 49
use OAI21X1  OAI21X1_47
timestamp 1516325494
transform -1 0 2297 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1384
timestamp 1516325494
transform -1 0 2316 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1113
timestamp 1516325494
transform -1 0 2335 0 1 1731
box 0 0 19 49
use MUX2X1  MUX2X1_387
timestamp 1516325494
transform 1 0 2335 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_452
timestamp 1516325494
transform 1 0 2366 0 1 1731
box 0 0 15 49
use NAND2X1  NAND2X1_387
timestamp 1516325494
transform -1 0 2396 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_3
timestamp 1516325494
transform 1 0 2396 0 1 1731
box 0 0 30 49
use OR2X2  OR2X2_1082
timestamp 1516325494
transform 1 0 2426 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1359
timestamp 1516325494
transform 1 0 2445 0 1 1731
box 0 0 19 49
use NAND2X1  NAND2X1_3
timestamp 1516325494
transform -1 0 2479 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_1081
timestamp 1516325494
transform -1 0 2499 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_347
timestamp 1516325494
transform -1 0 2507 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_347
timestamp 1516325494
transform -1 0 2521 0 1 1731
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_306
timestamp 1516325494
transform 1 0 2521 0 1 1731
box 0 0 53 49
use NAND2X1  NAND2X1_498
timestamp 1516325494
transform 1 0 2575 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_498
timestamp 1516325494
transform -1 0 2620 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_36
timestamp 1516325494
transform 1 0 2620 0 1 1731
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_218
timestamp 1516325494
transform 1 0 2635 0 1 1731
box 0 0 53 49
use MUX2X1  MUX2X1_634
timestamp 1516325494
transform 1 0 2689 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_634
timestamp 1516325494
transform -1 0 2734 0 1 1731
box 0 0 15 49
use NAND2X1  NAND2X1_50
timestamp 1516325494
transform -1 0 2749 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_1615
timestamp 1516325494
transform -1 0 2768 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_220
timestamp 1516325494
transform -1 0 2821 0 1 1731
box 0 0 53 49
use OR2X2  OR2X2_1920
timestamp 1516325494
transform -1 0 2841 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_326
timestamp 1516325494
transform -1 0 2860 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1882
timestamp 1516325494
transform 1 0 2860 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1765
timestamp 1516325494
transform -1 0 2898 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1928
timestamp 1516325494
transform 1 0 2898 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_356
timestamp 1516325494
transform 1 0 2917 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_336
timestamp 1516325494
transform -1 0 2955 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_1825
timestamp 1516325494
transform -1 0 2974 0 1 1731
box 0 0 19 49
use OR2X2  OR2X2_335
timestamp 1516325494
transform -1 0 2993 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_358
timestamp 1516325494
transform -1 0 3012 0 1 1731
box 0 0 19 49
use INVX1  INVX1_171
timestamp 1516325494
transform 1 0 3012 0 1 1731
box 0 0 11 49
use AND2X2  AND2X2_357
timestamp 1516325494
transform -1 0 3042 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_255
timestamp 1516325494
transform 1 0 3042 0 1 1731
box 0 0 53 49
use NAND2X1  NAND2X1_223
timestamp 1516325494
transform 1 0 3095 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_223
timestamp 1516325494
transform -1 0 3140 0 1 1731
box 0 0 30 49
use FILL  FILL_BUFX2_601
timestamp 1516325494
transform -1 0 3149 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_601
timestamp 1516325494
transform -1 0 3163 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_220
timestamp 1516325494
transform 1 0 3164 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_220
timestamp 1516325494
transform -1 0 3209 0 1 1731
box 0 0 15 49
use FILL  FILL_BUFX2_587
timestamp 1516325494
transform 1 0 3209 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_587
timestamp 1516325494
transform 1 0 3217 0 1 1731
box 0 0 15 49
use FILL  FILL_BUFX2_155
timestamp 1516325494
transform 1 0 3232 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_155
timestamp 1516325494
transform 1 0 3240 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_1769
timestamp 1516325494
transform -1 0 3274 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1885
timestamp 1516325494
transform -1 0 3293 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_341
timestamp 1516325494
transform 1 0 3293 0 1 1731
box 0 0 53 49
use MUX2X1  MUX2X1_373
timestamp 1516325494
transform 1 0 3346 0 1 1731
box 0 0 30 49
use NAND2X1  NAND2X1_373
timestamp 1516325494
transform 1 0 3376 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_1919
timestamp 1516325494
transform -1 0 3411 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_360
timestamp 1516325494
transform -1 0 3430 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_1932
timestamp 1516325494
transform -1 0 3449 0 1 1731
box 0 0 19 49
use FILL  FILL_BUFX2_327
timestamp 1516325494
transform -1 0 3457 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_327
timestamp 1516325494
transform -1 0 3471 0 1 1731
box 0 0 15 49
use OR2X2  OR2X2_1918
timestamp 1516325494
transform -1 0 3490 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_2001
timestamp 1516325494
transform -1 0 3509 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_2002
timestamp 1516325494
transform -1 0 3528 0 1 1731
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_159
timestamp 1516325494
transform 1 0 3528 0 1 1731
box 0 0 53 49
use AND2X2  AND2X2_1380
timestamp 1516325494
transform 1 0 3582 0 1 1731
box 0 0 19 49
use AND2X2  AND2X2_2113
timestamp 1516325494
transform 1 0 3601 0 1 1731
box 0 0 19 49
use NAND2X1  NAND2X1_260
timestamp 1516325494
transform 1 0 3620 0 1 1731
box 0 0 15 49
use MUX2X1  MUX2X1_260
timestamp 1516325494
transform -1 0 3665 0 1 1731
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_132
timestamp 1516325494
transform -1 0 3718 0 1 1731
box 0 0 53 49
use FILL  FILL_BUFX2_584
timestamp 1516325494
transform 1 0 3718 0 1 1731
box 0 0 8 49
use BUFX2  BUFX2_584
timestamp 1516325494
transform 1 0 3726 0 1 1731
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_800
timestamp 1516325494
transform 1 0 3741 0 1 1731
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_792
timestamp 1516325494
transform -1 0 3847 0 1 1731
box 0 0 53 49
use AND2X2  AND2X2_1184
timestamp 1516325494
transform -1 0 3867 0 1 1731
box 0 0 19 49
use XNOR2X1  XNOR2X1_23
timestamp 1516325494
transform -1 0 36 0 -1 1730
box 0 0 34 49
use INVX1  INVX1_84
timestamp 1516325494
transform 1 0 36 0 -1 1730
box 0 0 11 49
use NOR2X1  NOR2X1_48
timestamp 1516325494
transform -1 0 63 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_731
timestamp 1516325494
transform -1 0 82 0 -1 1730
box 0 0 19 49
use NOR2X1  NOR2X1_44
timestamp 1516325494
transform 1 0 82 0 -1 1730
box 0 0 15 49
use INVX1  INVX1_76
timestamp 1516325494
transform 1 0 97 0 -1 1730
box 0 0 11 49
use AND2X2  AND2X2_809
timestamp 1516325494
transform -1 0 127 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_810
timestamp 1516325494
transform 1 0 127 0 -1 1730
box 0 0 19 49
use NAND3X1  NAND3X1_40
timestamp 1516325494
transform 1 0 146 0 -1 1730
box 0 0 19 49
use NAND3X1  NAND3X1_41
timestamp 1516325494
transform -1 0 184 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_683
timestamp 1516325494
transform 1 0 184 0 -1 1730
box 0 0 19 49
use OAI21X1  OAI21X1_9
timestamp 1516325494
transform -1 0 222 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_808
timestamp 1516325494
transform -1 0 241 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_474
timestamp 1516325494
transform -1 0 260 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_552
timestamp 1516325494
transform 1 0 260 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_650
timestamp 1516325494
transform 1 0 279 0 -1 1730
box 0 0 19 49
use XNOR2X1  XNOR2X1_22
timestamp 1516325494
transform -1 0 332 0 -1 1730
box 0 0 34 49
use AND2X2  AND2X2_651
timestamp 1516325494
transform 1 0 333 0 -1 1730
box 0 0 19 49
use FILL  FILL_BUFX2_623
timestamp 1516325494
transform -1 0 360 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_623
timestamp 1516325494
transform -1 0 374 0 -1 1730
box 0 0 15 49
use FILL  FILL_BUFX2_785
timestamp 1516325494
transform -1 0 382 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_785
timestamp 1516325494
transform -1 0 397 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_933
timestamp 1516325494
transform 1 0 397 0 -1 1730
box 0 0 19 49
use NOR2X1  NOR2X1_46
timestamp 1516325494
transform 1 0 416 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_778
timestamp 1516325494
transform -1 0 450 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_654
timestamp 1516325494
transform -1 0 469 0 -1 1730
box 0 0 19 49
use NOR2X1  NOR2X1_38
timestamp 1516325494
transform -1 0 484 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_857
timestamp 1516325494
transform 1 0 485 0 -1 1730
box 0 0 19 49
use AOI21X1  AOI21X1_13
timestamp 1516325494
transform -1 0 523 0 -1 1730
box 0 0 19 49
use INVX1  INVX1_64
timestamp 1516325494
transform 1 0 523 0 -1 1730
box 0 0 11 49
use NAND2X1  NAND2X1_713
timestamp 1516325494
transform 1 0 534 0 -1 1730
box 0 0 15 49
use NAND2X1  NAND2X1_664
timestamp 1516325494
transform -1 0 564 0 -1 1730
box 0 0 15 49
use NAND2X1  NAND2X1_714
timestamp 1516325494
transform 1 0 564 0 -1 1730
box 0 0 15 49
use XOR2X1  XOR2X1_37
timestamp 1516325494
transform -1 0 614 0 -1 1730
box 0 0 34 49
use OR2X2  OR2X2_887
timestamp 1516325494
transform 1 0 614 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1092
timestamp 1516325494
transform 1 0 633 0 -1 1730
box 0 0 19 49
use INVX1  INVX1_63
timestamp 1516325494
transform -1 0 663 0 -1 1730
box 0 0 11 49
use XNOR2X1  XNOR2X1_8
timestamp 1516325494
transform -1 0 697 0 -1 1730
box 0 0 34 49
use XOR2X1  XOR2X1_39
timestamp 1516325494
transform -1 0 731 0 -1 1730
box 0 0 34 49
use INVX1  INVX1_69
timestamp 1516325494
transform -1 0 743 0 -1 1730
box 0 0 11 49
use OR2X2  OR2X2_889
timestamp 1516325494
transform 1 0 743 0 -1 1730
box 0 0 19 49
use INVX1  INVX1_70
timestamp 1516325494
transform -1 0 773 0 -1 1730
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_738
timestamp 1516325494
transform -1 0 826 0 -1 1730
box 0 0 53 49
use INVX1  INVX1_32
timestamp 1516325494
transform 1 0 827 0 -1 1730
box 0 0 11 49
use FILL  FILL_OR2X2_149
timestamp 1516325494
transform 1 0 838 0 -1 1730
box 0 0 8 49
use OR2X2  OR2X2_149
timestamp 1516325494
transform 1 0 846 0 -1 1730
box 0 0 19 49
use INVX1  INVX1_18
timestamp 1516325494
transform 1 0 865 0 -1 1730
box 0 0 11 49
use INVX1  INVX1_23
timestamp 1516325494
transform 1 0 876 0 -1 1730
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_698
timestamp 1516325494
transform 1 0 887 0 -1 1730
box 0 0 53 49
use OR2X2  OR2X2_1744
timestamp 1516325494
transform 1 0 941 0 -1 1730
box 0 0 19 49
use FILL  FILL_BUFX2_247
timestamp 1516325494
transform 1 0 960 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_247
timestamp 1516325494
transform 1 0 967 0 -1 1730
box 0 0 15 49
use NAND2X1  NAND2X1_313
timestamp 1516325494
transform 1 0 982 0 -1 1730
box 0 0 15 49
use NAND2X1  NAND2X1_314
timestamp 1516325494
transform 1 0 998 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_314
timestamp 1516325494
transform -1 0 1043 0 -1 1730
box 0 0 30 49
use OR2X2  OR2X2_1773
timestamp 1516325494
transform -1 0 1062 0 -1 1730
box 0 0 19 49
use NAND2X1  NAND2X1_474
timestamp 1516325494
transform 1 0 1062 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_474
timestamp 1516325494
transform -1 0 1107 0 -1 1730
box 0 0 30 49
use FILL  FILL_BUFX2_239
timestamp 1516325494
transform 1 0 1108 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_239
timestamp 1516325494
transform 1 0 1115 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_58
timestamp 1516325494
transform 1 0 1131 0 -1 1730
box 0 0 30 49
use NAND2X1  NAND2X1_58
timestamp 1516325494
transform -1 0 1176 0 -1 1730
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_666
timestamp 1516325494
transform -1 0 1229 0 -1 1730
box 0 0 53 49
use OR2X2  OR2X2_1778
timestamp 1516325494
transform -1 0 1248 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1622
timestamp 1516325494
transform 1 0 1248 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_473
timestamp 1516325494
transform -1 0 1320 0 -1 1730
box 0 0 53 49
use FILL  FILL_BUFX2_14
timestamp 1516325494
transform 1 0 1321 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_14
timestamp 1516325494
transform 1 0 1328 0 -1 1730
box 0 0 15 49
use OR2X2  OR2X2_1777
timestamp 1516325494
transform -1 0 1362 0 -1 1730
box 0 0 19 49
use NAND2X1  NAND2X1_442
timestamp 1516325494
transform 1 0 1362 0 -1 1730
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_58
timestamp 1516325494
transform 1 0 1378 0 -1 1730
box 0 0 53 49
use MUX2X1  MUX2X1_442
timestamp 1516325494
transform -1 0 1461 0 -1 1730
box 0 0 30 49
use OR2X2  OR2X2_1032
timestamp 1516325494
transform -1 0 1480 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1534
timestamp 1516325494
transform -1 0 1499 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_690
timestamp 1516325494
transform 1 0 1499 0 -1 1730
box 0 0 53 49
use NAND2X1  NAND2X1_306
timestamp 1516325494
transform 1 0 1552 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_306
timestamp 1516325494
transform -1 0 1598 0 -1 1730
box 0 0 30 49
use NAND2X1  NAND2X1_911
timestamp 1516325494
transform 1 0 1598 0 -1 1730
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_353
timestamp 1516325494
transform 1 0 1613 0 -1 1730
box 0 0 53 49
use MUX2X1  MUX2X1_856
timestamp 1516325494
transform -1 0 1696 0 -1 1730
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_462
timestamp 1516325494
transform -1 0 1750 0 -1 1730
box 0 0 53 49
use OR2X2  OR2X2_1424
timestamp 1516325494
transform -1 0 1769 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1629
timestamp 1516325494
transform -1 0 1788 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_309
timestamp 1516325494
transform 1 0 1788 0 -1 1730
box 0 0 53 49
use NAND2X1  NAND2X1_501
timestamp 1516325494
transform 1 0 1841 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_501
timestamp 1516325494
transform -1 0 1886 0 -1 1730
box 0 0 30 49
use FILL  FILL_BUFX2_823
timestamp 1516325494
transform 1 0 1887 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_823
timestamp 1516325494
transform 1 0 1894 0 -1 1730
box 0 0 15 49
use OR2X2  OR2X2_1095
timestamp 1516325494
transform 1 0 1910 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1369
timestamp 1516325494
transform 1 0 1929 0 -1 1730
box 0 0 19 49
use FILL  FILL_BUFX2_2
timestamp 1516325494
transform 1 0 1948 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_2
timestamp 1516325494
transform 1 0 1955 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_2105
timestamp 1516325494
transform -1 0 1989 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_2016
timestamp 1516325494
transform -1 0 2008 0 -1 1730
box 0 0 19 49
use NAND2X1  NAND2X1_21
timestamp 1516325494
transform 1 0 2008 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_21
timestamp 1516325494
transform -1 0 2054 0 -1 1730
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_597
timestamp 1516325494
transform -1 0 2107 0 -1 1730
box 0 0 53 49
use MUX2X1  MUX2X1_781
timestamp 1516325494
transform 1 0 2107 0 -1 1730
box 0 0 30 49
use AND2X2  AND2X2_1364
timestamp 1516325494
transform 1 0 2138 0 -1 1730
box 0 0 19 49
use FILL  FILL_BUFX2_567
timestamp 1516325494
transform -1 0 2165 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_567
timestamp 1516325494
transform -1 0 2179 0 -1 1730
box 0 0 15 49
use OR2X2  OR2X2_1103
timestamp 1516325494
transform 1 0 2179 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1091
timestamp 1516325494
transform -1 0 2217 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1090
timestamp 1516325494
transform -1 0 2236 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1085
timestamp 1516325494
transform -1 0 2255 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_2101
timestamp 1516325494
transform -1 0 2274 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_50
timestamp 1516325494
transform 1 0 2274 0 -1 1730
box 0 0 53 49
use AND2X2  AND2X2_1012
timestamp 1516325494
transform 1 0 2 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1013
timestamp 1516325494
transform 1 0 21 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1015
timestamp 1516325494
transform 1 0 40 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1053
timestamp 1516325494
transform 1 0 59 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_564
timestamp 1516325494
transform -1 0 97 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_490
timestamp 1516325494
transform -1 0 116 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_714
timestamp 1516325494
transform 1 0 116 0 1 1632
box 0 0 19 49
use XOR2X1  XOR2X1_8
timestamp 1516325494
transform -1 0 169 0 1 1632
box 0 0 34 49
use AND2X2  AND2X2_925
timestamp 1516325494
transform 1 0 169 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_475
timestamp 1516325494
transform 1 0 188 0 1 1632
box 0 0 19 49
use OAI21X1  OAI21X1_1
timestamp 1516325494
transform -1 0 226 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_473
timestamp 1516325494
transform -1 0 245 0 1 1632
box 0 0 19 49
use XOR2X1  XOR2X1_9
timestamp 1516325494
transform -1 0 279 0 1 1632
box 0 0 34 49
use NOR3X1  NOR3X1_3
timestamp 1516325494
transform -1 0 298 0 1 1632
box 0 0 19 49
use INVX1  INVX1_8
timestamp 1516325494
transform 1 0 298 0 1 1632
box 0 0 11 49
use XNOR2X1  XNOR2X1_6
timestamp 1516325494
transform -1 0 344 0 1 1632
box 0 0 34 49
use NOR3X1  NOR3X1_2
timestamp 1516325494
transform 1 0 344 0 1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_707
timestamp 1516325494
transform -1 0 378 0 1 1632
box 0 0 15 49
use OR2X2  OR2X2_882
timestamp 1516325494
transform 1 0 378 0 1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_708
timestamp 1516325494
transform 1 0 397 0 1 1632
box 0 0 15 49
use XOR2X1  XOR2X1_34
timestamp 1516325494
transform -1 0 446 0 1 1632
box 0 0 34 49
use OR2X2  OR2X2_883
timestamp 1516325494
transform 1 0 447 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1089
timestamp 1516325494
transform 1 0 466 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_723
timestamp 1516325494
transform -1 0 504 0 1 1632
box 0 0 19 49
use NOR2X1  NOR2X1_47
timestamp 1516325494
transform -1 0 519 0 1 1632
box 0 0 15 49
use OAI21X1  OAI21X1_7
timestamp 1516325494
transform -1 0 538 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_777
timestamp 1516325494
transform -1 0 557 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_652
timestamp 1516325494
transform -1 0 576 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_885
timestamp 1516325494
transform -1 0 595 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1090
timestamp 1516325494
transform 1 0 595 0 1 1632
box 0 0 19 49
use XOR2X1  XOR2X1_36
timestamp 1516325494
transform 1 0 614 0 1 1632
box 0 0 34 49
use OR2X2  OR2X2_886
timestamp 1516325494
transform 1 0 648 0 1 1632
box 0 0 19 49
use OAI21X1  OAI21X1_63
timestamp 1516325494
transform 1 0 667 0 1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_783
timestamp 1516325494
transform 1 0 686 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_783
timestamp 1516325494
transform 1 0 694 0 1 1632
box 0 0 15 49
use XOR2X1  XOR2X1_38
timestamp 1516325494
transform 1 0 709 0 1 1632
box 0 0 34 49
use OR2X2  OR2X2_888
timestamp 1516325494
transform 1 0 743 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1093
timestamp 1516325494
transform 1 0 762 0 1 1632
box 0 0 19 49
use INVX1  INVX1_68
timestamp 1516325494
transform -1 0 792 0 1 1632
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_742
timestamp 1516325494
transform -1 0 845 0 1 1632
box 0 0 53 49
use AND2X2  AND2X2_879
timestamp 1516325494
transform -1 0 21 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_923
timestamp 1516325494
transform -1 0 40 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_878
timestamp 1516325494
transform -1 0 59 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_738
timestamp 1516325494
transform 1 0 59 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_880
timestamp 1516325494
transform -1 0 97 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_877
timestamp 1516325494
transform -1 0 116 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_846
timestamp 1516325494
transform -1 0 135 0 -1 1632
box 0 0 19 49
use NOR2X1  NOR2X1_41
timestamp 1516325494
transform 1 0 135 0 -1 1632
box 0 0 15 49
use AND2X2  AND2X2_924
timestamp 1516325494
transform -1 0 169 0 -1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_650
timestamp 1516325494
transform -1 0 184 0 -1 1632
box 0 0 15 49
use NAND3X1  NAND3X1_21
timestamp 1516325494
transform -1 0 203 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_563
timestamp 1516325494
transform 1 0 203 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_565
timestamp 1516325494
transform 1 0 222 0 -1 1632
box 0 0 19 49
use INVX1  INVX1_14
timestamp 1516325494
transform 1 0 241 0 -1 1632
box 0 0 11 49
use OR2X2  OR2X2_489
timestamp 1516325494
transform -1 0 272 0 -1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_152
timestamp 1516325494
transform 1 0 272 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_152
timestamp 1516325494
transform 1 0 279 0 -1 1632
box 0 0 15 49
use NOR3X1  NOR3X1_1
timestamp 1516325494
transform -1 0 314 0 -1 1632
box 0 0 19 49
use NAND3X1  NAND3X1_20
timestamp 1516325494
transform 1 0 314 0 -1 1632
box 0 0 19 49
use NAND3X1  NAND3X1_12
timestamp 1516325494
transform -1 0 352 0 -1 1632
box 0 0 19 49
use NAND3X1  NAND3X1_22
timestamp 1516325494
transform 1 0 352 0 -1 1632
box 0 0 19 49
use INVX1  INVX1_60
timestamp 1516325494
transform 1 0 371 0 -1 1632
box 0 0 11 49
use INVX1  INVX1_6
timestamp 1516325494
transform -1 0 393 0 -1 1632
box 0 0 11 49
use INVX1  INVX1_7
timestamp 1516325494
transform -1 0 404 0 -1 1632
box 0 0 11 49
use INVX1  INVX1_26
timestamp 1516325494
transform 1 0 405 0 -1 1632
box 0 0 11 49
use OAI21X1  OAI21X1_5
timestamp 1516325494
transform -1 0 435 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_779
timestamp 1516325494
transform -1 0 454 0 -1 1632
box 0 0 19 49
use OAI21X1  OAI21X1_6
timestamp 1516325494
transform -1 0 473 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_756
timestamp 1516325494
transform 1 0 473 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_858
timestamp 1516325494
transform 1 0 492 0 -1 1632
box 0 0 19 49
use XNOR2X1  XNOR2X1_5
timestamp 1516325494
transform -1 0 545 0 -1 1632
box 0 0 34 49
use FILL  FILL_BUFX2_153
timestamp 1516325494
transform -1 0 553 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_153
timestamp 1516325494
transform -1 0 568 0 -1 1632
box 0 0 15 49
use NOR2X1  NOR2X1_27
timestamp 1516325494
transform 1 0 568 0 -1 1632
box 0 0 15 49
use XOR2X1  XOR2X1_35
timestamp 1516325494
transform 1 0 583 0 -1 1632
box 0 0 34 49
use OAI21X1  OAI21X1_68
timestamp 1516325494
transform -1 0 637 0 -1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_710
timestamp 1516325494
transform -1 0 652 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_149
timestamp 1516325494
transform -1 0 660 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_149
timestamp 1516325494
transform -1 0 674 0 -1 1632
box 0 0 15 49
use NOR2X1  NOR2X1_31
timestamp 1516325494
transform 1 0 675 0 -1 1632
box 0 0 15 49
use OAI21X1  OAI21X1_62
timestamp 1516325494
transform -1 0 709 0 -1 1632
box 0 0 19 49
use XNOR2X1  XNOR2X1_10
timestamp 1516325494
transform 1 0 709 0 -1 1632
box 0 0 34 49
use INVX1  INVX1_66
timestamp 1516325494
transform -1 0 754 0 -1 1632
box 0 0 11 49
use XNOR2X1  XNOR2X1_11
timestamp 1516325494
transform 1 0 754 0 -1 1632
box 0 0 34 49
use OR2X2  OR2X2_594
timestamp 1516325494
transform -1 0 808 0 -1 1632
box 0 0 19 49
use NOR2X1  NOR2X1_83
timestamp 1516325494
transform 1 0 808 0 -1 1632
box 0 0 15 49
use INVX1  INVX1_67
timestamp 1516325494
transform -1 0 834 0 -1 1632
box 0 0 11 49
use INVX1  INVX1_10
timestamp 1516325494
transform 1 0 834 0 -1 1632
box 0 0 11 49
use MUX2X1  MUX2X1_807
timestamp 1516325494
transform 1 0 846 0 1 1632
box 0 0 30 49
use OR2X2  OR2X2_1434
timestamp 1516325494
transform -1 0 895 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1433
timestamp 1516325494
transform -1 0 914 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1432
timestamp 1516325494
transform -1 0 933 0 1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_722
timestamp 1516325494
transform -1 0 986 0 1 1632
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_570
timestamp 1516325494
transform 1 0 986 0 1 1632
box 0 0 53 49
use OR2X2  OR2X2_1426
timestamp 1516325494
transform -1 0 1058 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1621
timestamp 1516325494
transform -1 0 1077 0 1 1632
box 0 0 19 49
use FILL  FILL_OR2X2_147
timestamp 1516325494
transform -1 0 1085 0 1 1632
box 0 0 8 49
use OR2X2  OR2X2_147
timestamp 1516325494
transform -1 0 1104 0 1 1632
box 0 0 19 49
use FILL  FILL_AND2X2_157
timestamp 1516325494
transform -1 0 1112 0 1 1632
box 0 0 8 49
use AND2X2  AND2X2_157
timestamp 1516325494
transform -1 0 1131 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1623
timestamp 1516325494
transform -1 0 1150 0 1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_92
timestamp 1516325494
transform 1 0 1150 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_92
timestamp 1516325494
transform 1 0 1157 0 1 1632
box 0 0 15 49
use INVX1  INVX1_202
timestamp 1516325494
transform -1 0 1183 0 1 1632
box 0 0 11 49
use NAND2X1  NAND2X1_345
timestamp 1516325494
transform -1 0 1199 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_345
timestamp 1516325494
transform 1 0 1199 0 1 1632
box 0 0 30 49
use OR2X2  OR2X2_1779
timestamp 1516325494
transform -1 0 1248 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1318
timestamp 1516325494
transform -1 0 1267 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1033
timestamp 1516325494
transform -1 0 1286 0 1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_417
timestamp 1516325494
transform 1 0 1286 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_417
timestamp 1516325494
transform 1 0 1294 0 1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_21
timestamp 1516325494
transform -1 0 1317 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_21
timestamp 1516325494
transform -1 0 1332 0 1 1632
box 0 0 15 49
use NAND2X1  NAND2X1_161
timestamp 1516325494
transform 1 0 1332 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_385
timestamp 1516325494
transform 1 0 1347 0 1 1632
box 0 0 53 49
use MUX2X1  MUX2X1_161
timestamp 1516325494
transform -1 0 1430 0 1 1632
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_622
timestamp 1516325494
transform 1 0 1431 0 1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_892
timestamp 1516325494
transform 1 0 1484 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_837
timestamp 1516325494
transform -1 0 1529 0 1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_93
timestamp 1516325494
transform 1 0 1530 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_93
timestamp 1516325494
transform 1 0 1537 0 1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_482
timestamp 1516325494
transform 1 0 1552 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_482
timestamp 1516325494
transform 1 0 1560 0 1 1632
box 0 0 15 49
use OR2X2  OR2X2_1627
timestamp 1516325494
transform -1 0 1594 0 1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_334
timestamp 1516325494
transform 1 0 1594 0 1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_334
timestamp 1516325494
transform -1 0 1640 0 1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_481
timestamp 1516325494
transform -1 0 1648 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_481
timestamp 1516325494
transform -1 0 1662 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_719
timestamp 1516325494
transform -1 0 899 0 -1 1632
box 0 0 53 49
use FILL  FILL_OR2X2_150
timestamp 1516325494
transform 1 0 899 0 -1 1632
box 0 0 8 49
use OR2X2  OR2X2_150
timestamp 1516325494
transform 1 0 906 0 -1 1632
box 0 0 19 49
use FILL  FILL_OR2X2_151
timestamp 1516325494
transform -1 0 933 0 -1 1632
box 0 0 8 49
use OR2X2  OR2X2_151
timestamp 1516325494
transform -1 0 952 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_1867
timestamp 1516325494
transform 1 0 952 0 -1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_25
timestamp 1516325494
transform 1 0 971 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_25
timestamp 1516325494
transform -1 0 1016 0 -1 1632
box 0 0 15 49
use OR2X2  OR2X2_1743
timestamp 1516325494
transform -1 0 1036 0 -1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_569
timestamp 1516325494
transform 1 0 1036 0 -1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_473
timestamp 1516325494
transform 1 0 1089 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_473
timestamp 1516325494
transform -1 0 1134 0 -1 1632
box 0 0 30 49
use MUX2X1  MUX2X1_780
timestamp 1516325494
transform -1 0 1164 0 -1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_22
timestamp 1516325494
transform 1 0 1165 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_22
timestamp 1516325494
transform 1 0 1172 0 -1 1632
box 0 0 15 49
use FILL  FILL_AND2X2_156
timestamp 1516325494
transform -1 0 1196 0 -1 1632
box 0 0 8 49
use AND2X2  AND2X2_156
timestamp 1516325494
transform -1 0 1214 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1754
timestamp 1516325494
transform 1 0 1214 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_1875
timestamp 1516325494
transform -1 0 1252 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1755
timestamp 1516325494
transform -1 0 1271 0 -1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_314
timestamp 1516325494
transform 1 0 1271 0 -1 1632
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_89
timestamp 1516325494
transform 1 0 1324 0 -1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_153
timestamp 1516325494
transform 1 0 1378 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_153
timestamp 1516325494
transform 1 0 1393 0 -1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_608
timestamp 1516325494
transform -1 0 1431 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_608
timestamp 1516325494
transform -1 0 1446 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_458
timestamp 1516325494
transform -1 0 1454 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_458
timestamp 1516325494
transform -1 0 1469 0 -1 1632
box 0 0 15 49
use OR2X2  OR2X2_1416
timestamp 1516325494
transform -1 0 1488 0 -1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_820
timestamp 1516325494
transform 1 0 1488 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_820
timestamp 1516325494
transform 1 0 1495 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_551
timestamp 1516325494
transform -1 0 1519 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_551
timestamp 1516325494
transform -1 0 1533 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_173
timestamp 1516325494
transform 1 0 1533 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_173
timestamp 1516325494
transform 1 0 1541 0 -1 1632
box 0 0 15 49
use AND2X2  AND2X2_1620
timestamp 1516325494
transform -1 0 1575 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1423
timestamp 1516325494
transform -1 0 1594 0 -1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_398
timestamp 1516325494
transform 1 0 1594 0 -1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_174
timestamp 1516325494
transform 1 0 1647 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_250
timestamp 1516325494
transform -1 0 1671 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_250
timestamp 1516325494
transform -1 0 1685 0 1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_346
timestamp 1516325494
transform 1 0 1685 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_346
timestamp 1516325494
transform 1 0 1693 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_451
timestamp 1516325494
transform 1 0 1708 0 1 1632
box 0 0 53 49
use MUX2X1  MUX2X1_323
timestamp 1516325494
transform -1 0 1791 0 1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_323
timestamp 1516325494
transform -1 0 1807 0 1 1632
box 0 0 15 49
use OR2X2  OR2X2_1094
timestamp 1516325494
transform 1 0 1807 0 1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_387
timestamp 1516325494
transform 1 0 1826 0 1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_163
timestamp 1516325494
transform 1 0 1879 0 1 1632
box 0 0 15 49
use OR2X2  OR2X2_1093
timestamp 1516325494
transform 1 0 1894 0 1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_163
timestamp 1516325494
transform 1 0 1913 0 1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_543
timestamp 1516325494
transform 1 0 1944 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_543
timestamp 1516325494
transform 1 0 1959 0 1 1632
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_543
timestamp 1516325494
transform 1 0 1989 0 1 1632
box 0 0 53 49
use FILL  FILL_BUFX2_88
timestamp 1516325494
transform 1 0 2043 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_88
timestamp 1516325494
transform 1 0 2050 0 1 1632
box 0 0 15 49
use OR2X2  OR2X2_1087
timestamp 1516325494
transform 1 0 2065 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1363
timestamp 1516325494
transform 1 0 2084 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1086
timestamp 1516325494
transform -1 0 2122 0 1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_611
timestamp 1516325494
transform 1 0 2122 0 1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_881
timestamp 1516325494
transform 1 0 2176 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_826
timestamp 1516325494
transform -1 0 2221 0 1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_89
timestamp 1516325494
transform 1 0 2221 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_89
timestamp 1516325494
transform 1 0 2229 0 1 1632
box 0 0 15 49
use AND2X2  AND2X2_1362
timestamp 1516325494
transform -1 0 2263 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1117
timestamp 1516325494
transform -1 0 2282 0 1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_434
timestamp 1516325494
transform 1 0 2282 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_434
timestamp 1516325494
transform -1 0 2327 0 1 1632
box 0 0 30 49
use MUX2X1  MUX2X1_174
timestamp 1516325494
transform 1 0 1663 0 -1 1632
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_409
timestamp 1516325494
transform 1 0 1693 0 -1 1632
box 0 0 53 49
use FILL  FILL_BUFX2_127
timestamp 1516325494
transform 1 0 1746 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_127
timestamp 1516325494
transform 1 0 1754 0 -1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_53
timestamp 1516325494
transform 1 0 1769 0 -1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_437
timestamp 1516325494
transform 1 0 1822 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_437
timestamp 1516325494
transform -1 0 1867 0 -1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_39
timestamp 1516325494
transform 1 0 1868 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_39
timestamp 1516325494
transform 1 0 1875 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_515
timestamp 1516325494
transform -1 0 1899 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_515
timestamp 1516325494
transform -1 0 1913 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_717
timestamp 1516325494
transform 1 0 1913 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_717
timestamp 1516325494
transform 1 0 1921 0 -1 1632
box 0 0 15 49
use NAND2X1  NAND2X1_95
timestamp 1516325494
transform 1 0 1936 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_95
timestamp 1516325494
transform -1 0 1981 0 -1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_647
timestamp 1516325494
transform 1 0 1982 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_647
timestamp 1516325494
transform 1 0 1989 0 -1 1632
box 0 0 15 49
use NAND2X1  NAND2X1_515
timestamp 1516325494
transform 1 0 2005 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_515
timestamp 1516325494
transform -1 0 2050 0 -1 1632
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_35
timestamp 1516325494
transform 1 0 2050 0 -1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_419
timestamp 1516325494
transform 1 0 2103 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_419
timestamp 1516325494
transform -1 0 2149 0 -1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_716
timestamp 1516325494
transform 1 0 2149 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_716
timestamp 1516325494
transform 1 0 2157 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_498
timestamp 1516325494
transform -1 0 2180 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_498
timestamp 1516325494
transform -1 0 2194 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_724
timestamp 1516325494
transform 1 0 2195 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_724
timestamp 1516325494
transform 1 0 2202 0 -1 1632
box 0 0 15 49
use INVX1  INVX1_137
timestamp 1516325494
transform -1 0 2228 0 -1 1632
box 0 0 11 49
use FILL  FILL_BUFX2_427
timestamp 1516325494
transform 1 0 2229 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_427
timestamp 1516325494
transform 1 0 2236 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_4
timestamp 1516325494
transform 1 0 2252 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_4
timestamp 1516325494
transform -1 0 2297 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_402
timestamp 1516325494
transform 1 0 2297 0 -1 1632
box 0 0 30 49
use INVX1  INVX1_138
timestamp 1516325494
transform 1 0 2328 0 -1 1730
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_548
timestamp 1516325494
transform 1 0 2339 0 -1 1730
box 0 0 53 49
use MUX2X1  MUX2X1_452
timestamp 1516325494
transform -1 0 2422 0 -1 1730
box 0 0 30 49
use FILL  FILL_BUFX2_290
timestamp 1516325494
transform 1 0 2423 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_290
timestamp 1516325494
transform 1 0 2430 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_1704
timestamp 1516325494
transform -1 0 2464 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1531
timestamp 1516325494
transform -1 0 2483 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_594
timestamp 1516325494
transform 1 0 2483 0 -1 1730
box 0 0 53 49
use NAND2X1  NAND2X1_18
timestamp 1516325494
transform 1 0 2537 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_18
timestamp 1516325494
transform -1 0 2582 0 -1 1730
box 0 0 30 49
use FILL  FILL_BUFX2_822
timestamp 1516325494
transform 1 0 2582 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_822
timestamp 1516325494
transform 1 0 2590 0 -1 1730
box 0 0 15 49
use FILL  FILL_BUFX2_465
timestamp 1516325494
transform -1 0 2613 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_465
timestamp 1516325494
transform -1 0 2628 0 -1 1730
box 0 0 15 49
use FILL  FILL_BUFX2_502
timestamp 1516325494
transform 1 0 2628 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_502
timestamp 1516325494
transform 1 0 2635 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_36
timestamp 1516325494
transform -1 0 2681 0 -1 1730
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_644
timestamp 1516325494
transform -1 0 2734 0 -1 1730
box 0 0 53 49
use OR2X2  OR2X2_2008
timestamp 1516325494
transform -1 0 2753 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1767
timestamp 1516325494
transform -1 0 2772 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_213
timestamp 1516325494
transform 1 0 2772 0 -1 1730
box 0 0 53 49
use FILL  FILL_AND2X2_251
timestamp 1516325494
transform 1 0 2825 0 -1 1730
box 0 0 8 49
use AND2X2  AND2X2_251
timestamp 1516325494
transform 1 0 2833 0 -1 1730
box 0 0 19 49
use FILL  FILL_OR2X2_236
timestamp 1516325494
transform -1 0 2860 0 -1 1730
box 0 0 8 49
use OR2X2  OR2X2_236
timestamp 1516325494
transform -1 0 2879 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_381
timestamp 1516325494
transform -1 0 2898 0 -1 1730
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_181
timestamp 1516325494
transform 1 0 2898 0 -1 1730
box 0 0 53 49
use OR2X2  OR2X2_334
timestamp 1516325494
transform -1 0 2970 0 -1 1730
box 0 0 19 49
use NAND2X1  NAND2X1_612
timestamp 1516325494
transform 1 0 2970 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_612
timestamp 1516325494
transform -1 0 3015 0 -1 1730
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_196
timestamp 1516325494
transform -1 0 3068 0 -1 1730
box 0 0 53 49
use NAND2X1  NAND2X1_420
timestamp 1516325494
transform 1 0 2328 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_36
timestamp 1516325494
transform 1 0 2343 0 1 1632
box 0 0 53 49
use AND2X2  AND2X2_1382
timestamp 1516325494
transform -1 0 2415 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1111
timestamp 1516325494
transform -1 0 2434 0 1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_420
timestamp 1516325494
transform -1 0 2464 0 1 1632
box 0 0 30 49
use OR2X2  OR2X2_1532
timestamp 1516325494
transform -1 0 2483 0 1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_402
timestamp 1516325494
transform 1 0 2483 0 1 1632
box 0 0 15 49
use OR2X2  OR2X2_1114
timestamp 1516325494
transform 1 0 2499 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1922
timestamp 1516325494
transform 1 0 2518 0 1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_31
timestamp 1516325494
transform 1 0 2537 0 1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_31
timestamp 1516325494
transform -1 0 2582 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_607
timestamp 1516325494
transform -1 0 2635 0 1 1632
box 0 0 53 49
use OR2X2  OR2X2_1921
timestamp 1516325494
transform 1 0 2635 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_2003
timestamp 1516325494
transform -1 0 2673 0 1 1632
box 0 0 19 49
use OAI21X1  OAI21X1_20
timestamp 1516325494
transform 1 0 2673 0 1 1632
box 0 0 19 49
use INVX2  INVX2_9
timestamp 1516325494
transform -1 0 2703 0 1 1632
box 0 0 11 49
use FILL  FILL_BUFX2_370
timestamp 1516325494
transform 1 0 2704 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_370
timestamp 1516325494
transform 1 0 2711 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_50
timestamp 1516325494
transform -1 0 2757 0 1 1632
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_658
timestamp 1516325494
transform -1 0 2810 0 1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_629
timestamp 1516325494
transform 1 0 2810 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_629
timestamp 1516325494
transform -1 0 2855 0 1 1632
box 0 0 30 49
use AND2X2  AND2X2_1766
timestamp 1516325494
transform -1 0 2875 0 1 1632
box 0 0 19 49
use FILL  FILL_AND2X2_250
timestamp 1516325494
transform -1 0 2883 0 1 1632
box 0 0 8 49
use AND2X2  AND2X2_250
timestamp 1516325494
transform -1 0 2901 0 1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_245
timestamp 1516325494
transform 1 0 2901 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_245
timestamp 1516325494
transform -1 0 2947 0 1 1632
box 0 0 30 49
use AND2X2  AND2X2_325
timestamp 1516325494
transform -1 0 2966 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_355
timestamp 1516325494
transform 1 0 2966 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1881
timestamp 1516325494
transform -1 0 3004 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1927
timestamp 1516325494
transform -1 0 3023 0 1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_665
timestamp 1516325494
transform 1 0 3023 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_665
timestamp 1516325494
transform 1 0 3031 0 1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_111
timestamp 1516325494
transform 1 0 3046 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_111
timestamp 1516325494
transform 1 0 3053 0 1 1632
box 0 0 15 49
use FILL  FILL_OR2X2_3
timestamp 1516325494
transform -1 0 3077 0 -1 1730
box 0 0 8 49
use OR2X2  OR2X2_3
timestamp 1516325494
transform -1 0 3095 0 -1 1730
box 0 0 19 49
use NAND2X1  NAND2X1_580
timestamp 1516325494
transform 1 0 3095 0 -1 1730
box 0 0 15 49
use MUX2X1  MUX2X1_580
timestamp 1516325494
transform -1 0 3140 0 -1 1730
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_260
timestamp 1516325494
transform -1 0 3194 0 -1 1730
box 0 0 53 49
use OR2X2  OR2X2_1134
timestamp 1516325494
transform -1 0 3213 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1110
timestamp 1516325494
transform -1 0 3232 0 -1 1730
box 0 0 19 49
use FILL  FILL_BUFX2_837
timestamp 1516325494
transform -1 0 3240 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_837
timestamp 1516325494
transform -1 0 3255 0 -1 1730
box 0 0 15 49
use AND2X2  AND2X2_389
timestamp 1516325494
transform 1 0 3255 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_380
timestamp 1516325494
transform -1 0 3293 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_404
timestamp 1516325494
transform -1 0 3312 0 -1 1730
box 0 0 19 49
use FILL  FILL_BUFX2_770
timestamp 1516325494
transform -1 0 3320 0 -1 1730
box 0 0 8 49
use BUFX2  BUFX2_770
timestamp 1516325494
transform -1 0 3334 0 -1 1730
box 0 0 15 49
use OR2X2  OR2X2_310
timestamp 1516325494
transform -1 0 3354 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_329
timestamp 1516325494
transform -1 0 3373 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_2000
timestamp 1516325494
transform 1 0 3373 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_2007
timestamp 1516325494
transform -1 0 3411 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_2097
timestamp 1516325494
transform -1 0 3430 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1356
timestamp 1516325494
transform 1 0 3430 0 -1 1730
box 0 0 19 49
use FILL  FILL_OR2X2_2
timestamp 1516325494
transform -1 0 3457 0 -1 1730
box 0 0 8 49
use OR2X2  OR2X2_2
timestamp 1516325494
transform -1 0 3475 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_2112
timestamp 1516325494
transform 1 0 3475 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1379
timestamp 1516325494
transform 1 0 3494 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1109
timestamp 1516325494
transform -1 0 3532 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_379
timestamp 1516325494
transform -1 0 3551 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_405
timestamp 1516325494
transform -1 0 3570 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_406
timestamp 1516325494
transform -1 0 3589 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_2006
timestamp 1516325494
transform -1 0 3608 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_2098
timestamp 1516325494
transform -1 0 3627 0 -1 1730
box 0 0 19 49
use OR2X2  OR2X2_1108
timestamp 1516325494
transform -1 0 3646 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1381
timestamp 1516325494
transform 1 0 3646 0 -1 1730
box 0 0 19 49
use FILL  FILL_OR2X2_1
timestamp 1516325494
transform -1 0 3673 0 -1 1730
box 0 0 8 49
use OR2X2  OR2X2_1
timestamp 1516325494
transform -1 0 3692 0 -1 1730
box 0 0 19 49
use FILL  FILL_AND2X2_1
timestamp 1516325494
transform 1 0 3692 0 -1 1730
box 0 0 8 49
use AND2X2  AND2X2_1
timestamp 1516325494
transform 1 0 3699 0 -1 1730
box 0 0 19 49
use MUX2X1  MUX2X1_356
timestamp 1516325494
transform 1 0 3718 0 -1 1730
box 0 0 30 49
use NAND2X1  NAND2X1_356
timestamp 1516325494
transform -1 0 3764 0 -1 1730
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_324
timestamp 1516325494
transform -1 0 3817 0 -1 1730
box 0 0 53 49
use AND2X2  AND2X2_1183
timestamp 1516325494
transform -1 0 3836 0 -1 1730
box 0 0 19 49
use AND2X2  AND2X2_1182
timestamp 1516325494
transform 1 0 3836 0 -1 1730
box 0 0 19 49
use FILL  FILL_35_1
timestamp 1516325494
transform -1 0 3863 0 -1 1730
box 0 0 8 49
use FILL  FILL_35_2
timestamp 1516325494
transform -1 0 3871 0 -1 1730
box 0 0 8 49
use OR2X2  OR2X2_2019
timestamp 1516325494
transform 1 0 3069 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_2111
timestamp 1516325494
transform 1 0 3088 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_2018
timestamp 1516325494
transform -1 0 3126 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_2110
timestamp 1516325494
transform 1 0 3126 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1377
timestamp 1516325494
transform 1 0 3145 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1378
timestamp 1516325494
transform 1 0 3164 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1106
timestamp 1516325494
transform 1 0 3183 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1107
timestamp 1516325494
transform 1 0 3202 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1080
timestamp 1516325494
transform -1 0 3240 0 1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_196
timestamp 1516325494
transform 1 0 3240 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_196
timestamp 1516325494
transform -1 0 3285 0 1 1632
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_228
timestamp 1516325494
transform -1 0 3338 0 1 1632
box 0 0 53 49
use FILL  FILL_BUFX2_830
timestamp 1516325494
transform 1 0 3338 0 1 1632
box 0 0 8 49
use BUFX2  BUFX2_830
timestamp 1516325494
transform 1 0 3346 0 1 1632
box 0 0 15 49
use NAND2X1  NAND2X1_250
timestamp 1516325494
transform -1 0 3376 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_186
timestamp 1516325494
transform -1 0 3429 0 1 1632
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_434
timestamp 1516325494
transform -1 0 2381 0 -1 1632
box 0 0 53 49
use FILL  FILL_BUFX2_369
timestamp 1516325494
transform 1 0 2381 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_369
timestamp 1516325494
transform 1 0 2388 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_292
timestamp 1516325494
transform 1 0 2404 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_292
timestamp 1516325494
transform -1 0 2449 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_415
timestamp 1516325494
transform 1 0 2449 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_415
timestamp 1516325494
transform -1 0 2495 0 -1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_447
timestamp 1516325494
transform -1 0 2548 0 -1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_451
timestamp 1516325494
transform 1 0 2548 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_451
timestamp 1516325494
transform -1 0 2593 0 -1 1632
box 0 0 30 49
use FILL  FILL_BUFX2_91
timestamp 1516325494
transform -1 0 2602 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_91
timestamp 1516325494
transform -1 0 2616 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_255
timestamp 1516325494
transform 1 0 2616 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_255
timestamp 1516325494
transform -1 0 2662 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_826
timestamp 1516325494
transform -1 0 2670 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_826
timestamp 1516325494
transform -1 0 2685 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_90
timestamp 1516325494
transform -1 0 2693 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_90
timestamp 1516325494
transform -1 0 2707 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_368
timestamp 1516325494
transform -1 0 2716 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_368
timestamp 1516325494
transform -1 0 2730 0 -1 1632
box 0 0 15 49
use AND2X2  AND2X2_400
timestamp 1516325494
transform 1 0 2730 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_376
timestamp 1516325494
transform 1 0 2749 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_1996
timestamp 1516325494
transform 1 0 2768 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1915
timestamp 1516325494
transform 1 0 2787 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1917
timestamp 1516325494
transform 1 0 2806 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_378
timestamp 1516325494
transform 1 0 2825 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_377
timestamp 1516325494
transform -1 0 2863 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1916
timestamp 1516325494
transform -1 0 2882 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_402
timestamp 1516325494
transform -1 0 2901 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_1998
timestamp 1516325494
transform -1 0 2920 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_2108
timestamp 1516325494
transform 1 0 2920 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_2017
timestamp 1516325494
transform 1 0 2939 0 -1 1632
box 0 0 19 49
use AND2X2  AND2X2_2109
timestamp 1516325494
transform -1 0 2977 0 -1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_228
timestamp 1516325494
transform 1 0 2977 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_228
timestamp 1516325494
transform -1 0 3023 0 -1 1632
box 0 0 15 49
use AND2X2  AND2X2_1376
timestamp 1516325494
transform 1 0 3023 0 -1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_164
timestamp 1516325494
transform -1 0 3095 0 -1 1632
box 0 0 53 49
use AND2X2  AND2X2_1375
timestamp 1516325494
transform 1 0 3095 0 -1 1632
box 0 0 19 49
use OR2X2  OR2X2_1105
timestamp 1516325494
transform 1 0 3114 0 -1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_750
timestamp 1516325494
transform 1 0 3133 0 -1 1632
box 0 0 30 49
use OR2X2  OR2X2_1104
timestamp 1516325494
transform -1 0 3183 0 -1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_236
timestamp 1516325494
transform -1 0 3191 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_236
timestamp 1516325494
transform -1 0 3205 0 -1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_188
timestamp 1516325494
transform 1 0 3205 0 -1 1632
box 0 0 53 49
use OR2X2  OR2X2_366
timestamp 1516325494
transform -1 0 3278 0 -1 1632
box 0 0 19 49
use NAND2X1  NAND2X1_252
timestamp 1516325494
transform 1 0 3278 0 -1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_252
timestamp 1516325494
transform -1 0 3323 0 -1 1632
box 0 0 30 49
use INVX1  INVX1_279
timestamp 1516325494
transform 1 0 3323 0 -1 1632
box 0 0 11 49
use MUX2X1  MUX2X1_250
timestamp 1516325494
transform 1 0 3335 0 -1 1632
box 0 0 30 49
use OR2X2  OR2X2_365
timestamp 1516325494
transform -1 0 3384 0 -1 1632
box 0 0 19 49
use MUX2X1  MUX2X1_282
timestamp 1516325494
transform 1 0 3384 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_282
timestamp 1516325494
transform -1 0 3429 0 -1 1632
box 0 0 15 49
use OR2X2  OR2X2_1079
timestamp 1516325494
transform -1 0 3449 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_309
timestamp 1516325494
transform -1 0 3468 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_330
timestamp 1516325494
transform -1 0 3487 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1768
timestamp 1516325494
transform -1 0 3506 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1886
timestamp 1516325494
transform -1 0 3525 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1887
timestamp 1516325494
transform -1 0 3544 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_331
timestamp 1516325494
transform -1 0 3563 0 1 1632
box 0 0 19 49
use OR2X2  OR2X2_1078
timestamp 1516325494
transform -1 0 3582 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1357
timestamp 1516325494
transform 1 0 3582 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_1358
timestamp 1516325494
transform -1 0 3620 0 1 1632
box 0 0 19 49
use AND2X2  AND2X2_2099
timestamp 1516325494
transform -1 0 3639 0 1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_131
timestamp 1516325494
transform 1 0 3639 0 1 1632
box 0 0 53 49
use NAND2X1  NAND2X1_259
timestamp 1516325494
transform 1 0 3692 0 1 1632
box 0 0 15 49
use MUX2X1  MUX2X1_259
timestamp 1516325494
transform -1 0 3737 0 1 1632
box 0 0 30 49
use MUX2X1  MUX2X1_355
timestamp 1516325494
transform 1 0 3737 0 1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_355
timestamp 1516325494
transform -1 0 3783 0 1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_323
timestamp 1516325494
transform -1 0 3836 0 1 1632
box 0 0 53 49
use BUFX2  BUFX2_912
timestamp 1516325494
transform -1 0 3851 0 1 1632
box 0 0 15 49
use INVX1  INVX1_314
timestamp 1516325494
transform -1 0 3862 0 1 1632
box 0 0 11 49
use FILL  FILL_34_1
timestamp 1516325494
transform 1 0 3863 0 1 1632
box 0 0 8 49
use AND2X2  AND2X2_391
timestamp 1516325494
transform -1 0 3449 0 -1 1632
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_154
timestamp 1516325494
transform -1 0 3502 0 -1 1632
box 0 0 53 49
use MUX2X1  MUX2X1_378
timestamp 1516325494
transform 1 0 3502 0 -1 1632
box 0 0 30 49
use NAND2X1  NAND2X1_378
timestamp 1516325494
transform -1 0 3547 0 -1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_346
timestamp 1516325494
transform -1 0 3600 0 -1 1632
box 0 0 53 49
use FILL  FILL_AND2X2_211
timestamp 1516325494
transform -1 0 3609 0 -1 1632
box 0 0 8 49
use AND2X2  AND2X2_211
timestamp 1516325494
transform -1 0 3627 0 -1 1632
box 0 0 19 49
use FILL  FILL_BUFX2_831
timestamp 1516325494
transform 1 0 3627 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_831
timestamp 1516325494
transform 1 0 3635 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_189
timestamp 1516325494
transform -1 0 3658 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_189
timestamp 1516325494
transform -1 0 3673 0 -1 1632
box 0 0 15 49
use FILL  FILL_BUFX2_279
timestamp 1516325494
transform 1 0 3673 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_279
timestamp 1516325494
transform 1 0 3680 0 -1 1632
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_338
timestamp 1516325494
transform 1 0 3696 0 -1 1632
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_142
timestamp 1516325494
transform -1 0 3802 0 -1 1632
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_803
timestamp 1516325494
transform 1 0 3802 0 -1 1632
box 0 0 53 49
use FILL  FILL_33_1
timestamp 1516325494
transform -1 0 3863 0 -1 1632
box 0 0 8 49
use FILL  FILL_33_2
timestamp 1516325494
transform -1 0 3871 0 -1 1632
box 0 0 8 49
use BUFX2  BUFX2_881
timestamp 1516325494
transform 1 0 2 0 1 1533
box 0 0 15 49
use INVX1  INVX1_175
timestamp 1516325494
transform -1 0 28 0 1 1533
box 0 0 11 49
use OR2X2  OR2X2_837
timestamp 1516325494
transform -1 0 48 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_736
timestamp 1516325494
transform -1 0 67 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_869
timestamp 1516325494
transform -1 0 86 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1014
timestamp 1516325494
transform -1 0 105 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_847
timestamp 1516325494
transform -1 0 124 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_848
timestamp 1516325494
transform -1 0 143 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_898
timestamp 1516325494
transform 1 0 143 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_899
timestamp 1516325494
transform -1 0 181 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_900
timestamp 1516325494
transform 1 0 181 0 1 1533
box 0 0 19 49
use NAND3X1  NAND3X1_45
timestamp 1516325494
transform -1 0 219 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_868
timestamp 1516325494
transform -1 0 238 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_488
timestamp 1516325494
transform -1 0 257 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_432
timestamp 1516325494
transform -1 0 276 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_645
timestamp 1516325494
transform -1 0 291 0 1 1533
box 0 0 15 49
use AND2X2  AND2X2_476
timestamp 1516325494
transform -1 0 310 0 1 1533
box 0 0 19 49
use NAND3X1  NAND3X1_14
timestamp 1516325494
transform -1 0 329 0 1 1533
box 0 0 19 49
use NOR2X1  NOR2X1_18
timestamp 1516325494
transform -1 0 344 0 1 1533
box 0 0 15 49
use NAND3X1  NAND3X1_13
timestamp 1516325494
transform -1 0 363 0 1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_840
timestamp 1516325494
transform 1 0 363 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_840
timestamp 1516325494
transform 1 0 371 0 1 1533
box 0 0 15 49
use NAND3X1  NAND3X1_11
timestamp 1516325494
transform 1 0 386 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_642
timestamp 1516325494
transform -1 0 420 0 1 1533
box 0 0 15 49
use AND2X2  AND2X2_448
timestamp 1516325494
transform -1 0 439 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_937
timestamp 1516325494
transform -1 0 458 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_892
timestamp 1516325494
transform -1 0 477 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1088
timestamp 1516325494
transform -1 0 496 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_758
timestamp 1516325494
transform 1 0 496 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_706
timestamp 1516325494
transform 1 0 515 0 1 1533
box 0 0 15 49
use OR2X2  OR2X2_880
timestamp 1516325494
transform -1 0 549 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_705
timestamp 1516325494
transform -1 0 564 0 1 1533
box 0 0 15 49
use INVX1  INVX1_59
timestamp 1516325494
transform -1 0 575 0 1 1533
box 0 0 11 49
use AND2X2  AND2X2_757
timestamp 1516325494
transform -1 0 595 0 1 1533
box 0 0 19 49
use NAND3X1  NAND3X1_39
timestamp 1516325494
transform -1 0 614 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_632
timestamp 1516325494
transform -1 0 633 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_663
timestamp 1516325494
transform -1 0 648 0 1 1533
box 0 0 15 49
use NOR2X1  NOR2X1_19
timestamp 1516325494
transform 1 0 648 0 1 1533
box 0 0 15 49
use OR2X2  OR2X2_436
timestamp 1516325494
transform 1 0 663 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_884
timestamp 1516325494
transform -1 0 701 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_709
timestamp 1516325494
transform -1 0 716 0 1 1533
box 0 0 15 49
use NOR2X1  NOR2X1_35
timestamp 1516325494
transform 1 0 716 0 1 1533
box 0 0 15 49
use OR2X2  OR2X2_622
timestamp 1516325494
transform 1 0 732 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_602
timestamp 1516325494
transform 1 0 751 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_595
timestamp 1516325494
transform -1 0 789 0 1 1533
box 0 0 19 49
use NOR2X1  NOR2X1_32
timestamp 1516325494
transform -1 0 804 0 1 1533
box 0 0 15 49
use AOI21X1  AOI21X1_6
timestamp 1516325494
transform -1 0 823 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1064
timestamp 1516325494
transform 1 0 823 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1066
timestamp 1516325494
transform -1 0 861 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1065
timestamp 1516325494
transform -1 0 880 0 1 1533
box 0 0 19 49
use INVX1  INVX1_21
timestamp 1516325494
transform 1 0 880 0 1 1533
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_724
timestamp 1516325494
transform -1 0 944 0 1 1533
box 0 0 53 49
use INVX1  INVX1_154
timestamp 1516325494
transform 1 0 944 0 1 1533
box 0 0 11 49
use OR2X2  OR2X2_912
timestamp 1516325494
transform 1 0 956 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1116
timestamp 1516325494
transform 1 0 975 0 1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_601
timestamp 1516325494
transform -1 0 1047 0 1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_778
timestamp 1516325494
transform 1 0 1047 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_778
timestamp 1516325494
transform 1 0 1055 0 1 1533
box 0 0 15 49
use AND2X2  AND2X2_1868
timestamp 1516325494
transform 1 0 1070 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1745
timestamp 1516325494
transform -1 0 1108 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1866
timestamp 1516325494
transform 1 0 1108 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1889
timestamp 1516325494
transform -1 0 1146 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_332
timestamp 1516325494
transform -1 0 1165 0 1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_635
timestamp 1516325494
transform -1 0 1173 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_635
timestamp 1516325494
transform -1 0 1187 0 1 1533
box 0 0 15 49
use OR2X2  OR2X2_301
timestamp 1516325494
transform -1 0 1207 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_322
timestamp 1516325494
transform -1 0 1226 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_321
timestamp 1516325494
transform -1 0 1245 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1876
timestamp 1516325494
transform 1 0 1245 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1756
timestamp 1516325494
transform -1 0 1283 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1874
timestamp 1516325494
transform -1 0 1302 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_506
timestamp 1516325494
transform 1 0 1302 0 1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_506
timestamp 1516325494
transform -1 0 1347 0 1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_163
timestamp 1516325494
transform 1 0 1347 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_163
timestamp 1516325494
transform 1 0 1355 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_665
timestamp 1516325494
transform 1 0 1370 0 1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_57
timestamp 1516325494
transform 1 0 1423 0 1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_57
timestamp 1516325494
transform -1 0 1468 0 1 1533
box 0 0 30 49
use AND2X2  AND2X2_1873
timestamp 1516325494
transform -1 0 1488 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1752
timestamp 1516325494
transform -1 0 1507 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_935
timestamp 1516325494
transform 1 0 1507 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_377
timestamp 1516325494
transform 1 0 1522 0 1 1533
box 0 0 53 49
use MUX2X1  MUX2X1_880
timestamp 1516325494
transform 1 0 1575 0 1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_799
timestamp 1516325494
transform 1 0 1606 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_799
timestamp 1516325494
transform 1 0 1613 0 1 1533
box 0 0 15 49
use OR2X2  OR2X2_1753
timestamp 1516325494
transform -1 0 1647 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1422
timestamp 1516325494
transform -1 0 1666 0 1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_366
timestamp 1516325494
transform 1 0 1666 0 1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_185
timestamp 1516325494
transform 1 0 1720 0 1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_185
timestamp 1516325494
transform -1 0 1765 0 1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_924
timestamp 1516325494
transform 1 0 1765 0 1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_869
timestamp 1516325494
transform -1 0 1810 0 1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_762
timestamp 1516325494
transform 1 0 1811 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_762
timestamp 1516325494
transform 1 0 1818 0 1 1533
box 0 0 15 49
use OR2X2  OR2X2_839
timestamp 1516325494
transform -1 0 21 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_768
timestamp 1516325494
transform 1 0 21 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_746
timestamp 1516325494
transform 1 0 40 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_733
timestamp 1516325494
transform -1 0 78 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_732
timestamp 1516325494
transform -1 0 97 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_842
timestamp 1516325494
transform -1 0 116 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_682
timestamp 1516325494
transform 1 0 116 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_811
timestamp 1516325494
transform 1 0 135 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_730
timestamp 1516325494
transform -1 0 173 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_968
timestamp 1516325494
transform -1 0 192 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_967
timestamp 1516325494
transform -1 0 211 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_969
timestamp 1516325494
transform 1 0 211 0 -1 1533
box 0 0 19 49
use INVX1  INVX1_54
timestamp 1516325494
transform -1 0 241 0 -1 1533
box 0 0 11 49
use AND2X2  AND2X2_1025
timestamp 1516325494
transform 1 0 241 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_747
timestamp 1516325494
transform 1 0 260 0 -1 1533
box 0 0 19 49
use INVX1  INVX1_38
timestamp 1516325494
transform -1 0 290 0 -1 1533
box 0 0 11 49
use NAND3X1  NAND3X1_46
timestamp 1516325494
transform 1 0 291 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_889
timestamp 1516325494
transform 1 0 310 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_890
timestamp 1516325494
transform 1 0 329 0 -1 1533
box 0 0 19 49
use NAND3X1  NAND3X1_16
timestamp 1516325494
transform 1 0 348 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_652
timestamp 1516325494
transform -1 0 386 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_449
timestamp 1516325494
transform 1 0 386 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_934
timestamp 1516325494
transform -1 0 424 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_935
timestamp 1516325494
transform -1 0 443 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_936
timestamp 1516325494
transform 1 0 443 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_891
timestamp 1516325494
transform 1 0 462 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_482
timestamp 1516325494
transform 1 0 481 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_881
timestamp 1516325494
transform -1 0 519 0 -1 1533
box 0 0 19 49
use XOR2X1  XOR2X1_33
timestamp 1516325494
transform -1 0 553 0 -1 1533
box 0 0 34 49
use NOR2X1  NOR2X1_24
timestamp 1516325494
transform -1 0 568 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_542
timestamp 1516325494
transform 1 0 568 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_570
timestamp 1516325494
transform 1 0 587 0 -1 1533
box 0 0 19 49
use NOR2X1  NOR2X1_30
timestamp 1516325494
transform 1 0 606 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_585
timestamp 1516325494
transform 1 0 621 0 -1 1533
box 0 0 19 49
use XOR2X1  XOR2X1_28
timestamp 1516325494
transform -1 0 674 0 -1 1533
box 0 0 34 49
use AND2X2  AND2X2_705
timestamp 1516325494
transform -1 0 694 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_706
timestamp 1516325494
transform -1 0 713 0 -1 1533
box 0 0 19 49
use OAI21X1  OAI21X1_3
timestamp 1516325494
transform -1 0 732 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_593
timestamp 1516325494
transform -1 0 751 0 -1 1533
box 0 0 19 49
use NOR2X1  NOR2X1_36
timestamp 1516325494
transform 1 0 751 0 -1 1533
box 0 0 15 49
use AND2X2  AND2X2_704
timestamp 1516325494
transform -1 0 785 0 -1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_659
timestamp 1516325494
transform 1 0 785 0 -1 1533
box 0 0 15 49
use NOR2X1  NOR2X1_37
timestamp 1516325494
transform 1 0 800 0 -1 1533
box 0 0 15 49
use AND2X2  AND2X2_1067
timestamp 1516325494
transform 1 0 815 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1063
timestamp 1516325494
transform -1 0 853 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1062
timestamp 1516325494
transform -1 0 872 0 -1 1533
box 0 0 19 49
use INVX1  INVX1_17
timestamp 1516325494
transform 1 0 872 0 -1 1533
box 0 0 11 49
use FILL  FILL_BUFX2_316
timestamp 1516325494
transform -1 0 892 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_316
timestamp 1516325494
transform -1 0 906 0 -1 1533
box 0 0 15 49
use INVX1  INVX1_229
timestamp 1516325494
transform -1 0 917 0 -1 1533
box 0 0 11 49
use INVX1  INVX1_16
timestamp 1516325494
transform 1 0 918 0 -1 1533
box 0 0 11 49
use MUX2X1  MUX2X1_766
timestamp 1516325494
transform 1 0 929 0 -1 1533
box 0 0 30 49
use INVX1  INVX1_198
timestamp 1516325494
transform -1 0 971 0 -1 1533
box 0 0 11 49
use INVX1  INVX1_166
timestamp 1516325494
transform 1 0 971 0 -1 1533
box 0 0 11 49
use AND2X2  AND2X2_318
timestamp 1516325494
transform 1 0 982 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1741
timestamp 1516325494
transform -1 0 1020 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1865
timestamp 1516325494
transform -1 0 1039 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_317
timestamp 1516325494
transform 1 0 1039 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1751
timestamp 1516325494
transform -1 0 1077 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1763
timestamp 1516325494
transform 1 0 1077 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1764
timestamp 1516325494
transform -1 0 1115 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_303
timestamp 1516325494
transform -1 0 1134 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1748
timestamp 1516325494
transform -1 0 1153 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1322
timestamp 1516325494
transform 1 0 1153 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1036
timestamp 1516325494
transform 1 0 1172 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1319
timestamp 1516325494
transform -1 0 1210 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_2071
timestamp 1516325494
transform -1 0 1229 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1762
timestamp 1516325494
transform -1 0 1248 0 -1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_654
timestamp 1516325494
transform 1 0 1248 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_46
timestamp 1516325494
transform 1 0 1302 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_46
timestamp 1516325494
transform -1 0 1347 0 -1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_162
timestamp 1516325494
transform 1 0 1347 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_162
timestamp 1516325494
transform 1 0 1355 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_1761
timestamp 1516325494
transform -1 0 1389 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_302
timestamp 1516325494
transform -1 0 1408 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1880
timestamp 1516325494
transform -1 0 1427 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_324
timestamp 1516325494
transform -1 0 1446 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1879
timestamp 1516325494
transform 1 0 1446 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1616
timestamp 1516325494
transform -1 0 1484 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_548
timestamp 1516325494
transform -1 0 1492 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_548
timestamp 1516325494
transform -1 0 1507 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_1417
timestamp 1516325494
transform -1 0 1526 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_366
timestamp 1516325494
transform -1 0 1534 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_366
timestamp 1516325494
transform -1 0 1548 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_46
timestamp 1516325494
transform 1 0 1549 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_430
timestamp 1516325494
transform 1 0 1602 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_430
timestamp 1516325494
transform -1 0 1647 0 -1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_592
timestamp 1516325494
transform -1 0 1655 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_592
timestamp 1516325494
transform -1 0 1670 0 -1 1533
box 0 0 15 49
use AND2X2  AND2X2_2034
timestamp 1516325494
transform -1 0 1689 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1962
timestamp 1516325494
transform -1 0 1708 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1963
timestamp 1516325494
transform -1 0 1727 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_2036
timestamp 1516325494
transform -1 0 1746 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1965
timestamp 1516325494
transform -1 0 1765 0 -1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_384
timestamp 1516325494
transform 1 0 1765 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_942
timestamp 1516325494
transform 1 0 1818 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_1964
timestamp 1516325494
transform -1 0 1853 0 1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_456
timestamp 1516325494
transform 1 0 1853 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_456
timestamp 1516325494
transform 1 0 1860 0 1 1533
box 0 0 15 49
use NAND2X1  NAND2X1_352
timestamp 1516325494
transform 1 0 1875 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_480
timestamp 1516325494
transform 1 0 1891 0 1 1533
box 0 0 53 49
use MUX2X1  MUX2X1_352
timestamp 1516325494
transform -1 0 1974 0 1 1533
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_127
timestamp 1516325494
transform -1 0 2027 0 1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_321
timestamp 1516325494
transform 1 0 2027 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_321
timestamp 1516325494
transform 1 0 2035 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_470
timestamp 1516325494
transform -1 0 2058 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_470
timestamp 1516325494
transform -1 0 2073 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_797
timestamp 1516325494
transform 1 0 2073 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_797
timestamp 1516325494
transform 1 0 2081 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_515
timestamp 1516325494
transform -1 0 2149 0 1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_745
timestamp 1516325494
transform 1 0 2149 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_745
timestamp 1516325494
transform 1 0 2157 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_721
timestamp 1516325494
transform -1 0 2225 0 1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_800
timestamp 1516325494
transform -1 0 2233 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_800
timestamp 1516325494
transform -1 0 2248 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_634
timestamp 1516325494
transform -1 0 2256 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_634
timestamp 1516325494
transform -1 0 2270 0 1 1533
box 0 0 15 49
use INVX2  INVX2_36
timestamp 1516325494
transform -1 0 2282 0 1 1533
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_580
timestamp 1516325494
transform -1 0 2335 0 1 1533
box 0 0 53 49
use MUX2X1  MUX2X1_68
timestamp 1516325494
transform -1 0 2365 0 1 1533
box 0 0 30 49
use MUX2X1  MUX2X1_887
timestamp 1516325494
transform 1 0 1834 0 -1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_160
timestamp 1516325494
transform 1 0 1864 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_96
timestamp 1516325494
transform 1 0 1879 0 -1 1533
box 0 0 53 49
use MUX2X1  MUX2X1_160
timestamp 1516325494
transform -1 0 1962 0 -1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_846
timestamp 1516325494
transform 1 0 1963 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_846
timestamp 1516325494
transform 1 0 1970 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_416
timestamp 1516325494
transform 1 0 1986 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_192
timestamp 1516325494
transform 1 0 2039 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_192
timestamp 1516325494
transform -1 0 2084 0 -1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_537
timestamp 1516325494
transform 1 0 2084 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_537
timestamp 1516325494
transform 1 0 2100 0 -1 1533
box 0 0 53 49
use MUX2X1  MUX2X1_537
timestamp 1516325494
transform -1 0 2183 0 -1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_160
timestamp 1516325494
transform 1 0 2183 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_160
timestamp 1516325494
transform 1 0 2191 0 -1 1533
box 0 0 15 49
use AND2X2  AND2X2_1396
timestamp 1516325494
transform -1 0 2225 0 -1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_484
timestamp 1516325494
transform -1 0 2278 0 -1 1533
box 0 0 53 49
use OR2X2  OR2X2_1130
timestamp 1516325494
transform -1 0 2297 0 -1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_68
timestamp 1516325494
transform 1 0 2297 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_100
timestamp 1516325494
transform 1 0 2312 0 -1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_245
timestamp 1516325494
transform 1 0 2366 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_245
timestamp 1516325494
transform 1 0 2373 0 1 1533
box 0 0 15 49
use AND2X2  AND2X2_1361
timestamp 1516325494
transform -1 0 2407 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1112
timestamp 1516325494
transform -1 0 2426 0 1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_676
timestamp 1516325494
transform -1 0 2479 0 1 1533
box 0 0 53 49
use OR2X2  OR2X2_1084
timestamp 1516325494
transform -1 0 2499 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1083
timestamp 1516325494
transform -1 0 2518 0 1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_547
timestamp 1516325494
transform 1 0 2518 0 1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_761
timestamp 1516325494
transform 1 0 2571 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_761
timestamp 1516325494
transform 1 0 2578 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_181
timestamp 1516325494
transform -1 0 2602 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_181
timestamp 1516325494
transform -1 0 2616 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_191
timestamp 1516325494
transform -1 0 2669 0 1 1533
box 0 0 53 49
use OR2X2  OR2X2_2003
timestamp 1516325494
transform -1 0 2689 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_2094
timestamp 1516325494
transform -1 0 2708 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_401
timestamp 1516325494
transform 1 0 2708 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_2005
timestamp 1516325494
transform 1 0 2727 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1997
timestamp 1516325494
transform -1 0 2765 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_611
timestamp 1516325494
transform 1 0 2765 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_829
timestamp 1516325494
transform -1 0 2788 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_829
timestamp 1516325494
transform -1 0 2802 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_706
timestamp 1516325494
transform 1 0 2803 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_706
timestamp 1516325494
transform 1 0 2810 0 1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_381
timestamp 1516325494
transform 1 0 2825 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_381
timestamp 1516325494
transform 1 0 2833 0 1 1533
box 0 0 15 49
use AND2X2  AND2X2_403
timestamp 1516325494
transform 1 0 2848 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1999
timestamp 1516325494
transform -1 0 2886 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_2004
timestamp 1516325494
transform -1 0 2905 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_2096
timestamp 1516325494
transform -1 0 2924 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_2095
timestamp 1516325494
transform -1 0 2943 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1355
timestamp 1516325494
transform 1 0 2943 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1076
timestamp 1516325494
transform 1 0 2962 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1077
timestamp 1516325494
transform 1 0 2981 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1354
timestamp 1516325494
transform -1 0 3019 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_195
timestamp 1516325494
transform 1 0 3019 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_227
timestamp 1516325494
transform 1 0 3034 0 1 1533
box 0 0 53 49
use MUX2X1  MUX2X1_195
timestamp 1516325494
transform -1 0 3118 0 1 1533
box 0 0 30 49
use AND2X2  AND2X2_1607
timestamp 1516325494
transform 1 0 3118 0 1 1533
box 0 0 19 49
use AND2X2  AND2X2_1608
timestamp 1516325494
transform 1 0 3137 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1406
timestamp 1516325494
transform 1 0 3156 0 1 1533
box 0 0 19 49
use FILL  FILL_OR2X2_199
timestamp 1516325494
transform -1 0 3183 0 1 1533
box 0 0 8 49
use OR2X2  OR2X2_199
timestamp 1516325494
transform -1 0 3202 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_206
timestamp 1516325494
transform 1 0 3202 0 1 1533
box 0 0 15 49
use FILL  FILL_OR2X2_143
timestamp 1516325494
transform -1 0 3225 0 1 1533
box 0 0 8 49
use OR2X2  OR2X2_143
timestamp 1516325494
transform -1 0 3243 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1410
timestamp 1516325494
transform -1 0 3262 0 1 1533
box 0 0 19 49
use OR2X2  OR2X2_1407
timestamp 1516325494
transform -1 0 3281 0 1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_437
timestamp 1516325494
transform 1 0 3281 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_437
timestamp 1516325494
transform 1 0 3289 0 1 1533
box 0 0 15 49
use NAND2X1  NAND2X1_286
timestamp 1516325494
transform -1 0 3319 0 1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_286
timestamp 1516325494
transform -1 0 3349 0 1 1533
box 0 0 30 49
use MUX2X1  MUX2X1_382
timestamp 1516325494
transform 1 0 3350 0 1 1533
box 0 0 30 49
use AND2X2  AND2X2_390
timestamp 1516325494
transform -1 0 3399 0 1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_382
timestamp 1516325494
transform -1 0 3414 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_350
timestamp 1516325494
transform -1 0 3467 0 1 1533
box 0 0 53 49
use FILL  FILL_BUFX2_156
timestamp 1516325494
transform -1 0 3476 0 1 1533
box 0 0 8 49
use BUFX2  BUFX2_156
timestamp 1516325494
transform -1 0 3490 0 1 1533
box 0 0 15 49
use FILL  FILL_OR2X2_198
timestamp 1516325494
transform -1 0 3498 0 1 1533
box 0 0 8 49
use OR2X2  OR2X2_198
timestamp 1516325494
transform -1 0 3517 0 1 1533
box 0 0 19 49
use FILL  FILL_AND2X2_209
timestamp 1516325494
transform -1 0 3525 0 1 1533
box 0 0 8 49
use AND2X2  AND2X2_209
timestamp 1516325494
transform -1 0 3544 0 1 1533
box 0 0 19 49
use FILL  FILL_OR2X2_197
timestamp 1516325494
transform -1 0 3552 0 1 1533
box 0 0 8 49
use OR2X2  OR2X2_197
timestamp 1516325494
transform -1 0 3570 0 1 1533
box 0 0 19 49
use FILL  FILL_AND2X2_210
timestamp 1516325494
transform -1 0 3578 0 1 1533
box 0 0 8 49
use AND2X2  AND2X2_210
timestamp 1516325494
transform -1 0 3597 0 1 1533
box 0 0 19 49
use FILL  FILL_OR2X2_142
timestamp 1516325494
transform -1 0 3605 0 1 1533
box 0 0 8 49
use OR2X2  OR2X2_142
timestamp 1516325494
transform -1 0 3623 0 1 1533
box 0 0 19 49
use FILL  FILL_AND2X2_149
timestamp 1516325494
transform -1 0 3631 0 1 1533
box 0 0 8 49
use AND2X2  AND2X2_149
timestamp 1516325494
transform -1 0 3650 0 1 1533
box 0 0 19 49
use FILL  FILL_OR2X2_141
timestamp 1516325494
transform -1 0 3658 0 1 1533
box 0 0 8 49
use OR2X2  OR2X2_141
timestamp 1516325494
transform -1 0 3677 0 1 1533
box 0 0 19 49
use MUX2X1  MUX2X1_370
timestamp 1516325494
transform 1 0 3677 0 1 1533
box 0 0 30 49
use MUX2X1  MUX2X1_270
timestamp 1516325494
transform 1 0 3707 0 1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_270
timestamp 1516325494
transform -1 0 3752 0 1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_353
timestamp 1516325494
transform 1 0 3753 0 1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_353
timestamp 1516325494
transform -1 0 3798 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_321
timestamp 1516325494
transform -1 0 3851 0 1 1533
box 0 0 53 49
use BUFX2  BUFX2_875
timestamp 1516325494
transform -1 0 3866 0 1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_516
timestamp 1516325494
transform 1 0 2366 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_516
timestamp 1516325494
transform 1 0 2419 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_516
timestamp 1516325494
transform -1 0 2464 0 -1 1533
box 0 0 30 49
use OAI21X1  OAI21X1_49
timestamp 1516325494
transform 1 0 2464 0 -1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_388
timestamp 1516325494
transform 1 0 2483 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_388
timestamp 1516325494
transform -1 0 2529 0 -1 1533
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_420
timestamp 1516325494
transform -1 0 2582 0 -1 1533
box 0 0 53 49
use AND2X2  AND2X2_1365
timestamp 1516325494
transform -1 0 2601 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1088
timestamp 1516325494
transform -1 0 2620 0 -1 1533
box 0 0 19 49
use NAND2X1  NAND2X1_35
timestamp 1516325494
transform 1 0 2620 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_35
timestamp 1516325494
transform -1 0 2665 0 -1 1533
box 0 0 30 49
use OR2X2  OR2X2_911
timestamp 1516325494
transform -1 0 2685 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_348
timestamp 1516325494
transform -1 0 2693 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_348
timestamp 1516325494
transform -1 0 2707 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_639
timestamp 1516325494
transform 1 0 2708 0 -1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_639
timestamp 1516325494
transform -1 0 2753 0 -1 1533
box 0 0 15 49
use FILL  FILL_BUFX2_213
timestamp 1516325494
transform 1 0 2753 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_213
timestamp 1516325494
transform 1 0 2761 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_611
timestamp 1516325494
transform -1 0 2806 0 -1 1533
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_195
timestamp 1516325494
transform -1 0 2859 0 -1 1533
box 0 0 53 49
use AND2X2  AND2X2_1353
timestamp 1516325494
transform 1 0 2860 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1075
timestamp 1516325494
transform 1 0 2879 0 -1 1533
box 0 0 19 49
use MUX2X1  MUX2X1_607
timestamp 1516325494
transform 1 0 2898 0 -1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_607
timestamp 1516325494
transform -1 0 2943 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_287
timestamp 1516325494
transform -1 0 2996 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_579
timestamp 1516325494
transform 1 0 2996 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_579
timestamp 1516325494
transform -1 0 3042 0 -1 1533
box 0 0 30 49
use OAI21X1  OAI21X1_60
timestamp 1516325494
transform -1 0 3061 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_662
timestamp 1516325494
transform 1 0 3061 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_662
timestamp 1516325494
transform 1 0 3069 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_752
timestamp 1516325494
transform -1 0 3114 0 -1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_661
timestamp 1516325494
transform -1 0 3122 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_661
timestamp 1516325494
transform -1 0 3137 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_749
timestamp 1516325494
transform 1 0 3137 0 -1 1533
box 0 0 30 49
use FILL  FILL_BUFX2_549
timestamp 1516325494
transform -1 0 3175 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_549
timestamp 1516325494
transform -1 0 3190 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_206
timestamp 1516325494
transform 1 0 3190 0 -1 1533
box 0 0 30 49
use FILL  FILL_AND2X2_147
timestamp 1516325494
transform 1 0 3221 0 -1 1533
box 0 0 8 49
use AND2X2  AND2X2_147
timestamp 1516325494
transform 1 0 3228 0 -1 1533
box 0 0 19 49
use FILL  FILL_OR2X2_139
timestamp 1516325494
transform 1 0 3247 0 -1 1533
box 0 0 8 49
use OR2X2  OR2X2_139
timestamp 1516325494
transform 1 0 3255 0 -1 1533
box 0 0 19 49
use FILL  FILL_OR2X2_140
timestamp 1516325494
transform -1 0 3282 0 -1 1533
box 0 0 8 49
use OR2X2  OR2X2_140
timestamp 1516325494
transform -1 0 3300 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_556
timestamp 1516325494
transform -1 0 3308 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_556
timestamp 1516325494
transform -1 0 3323 0 -1 1533
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_158
timestamp 1516325494
transform -1 0 3376 0 -1 1533
box 0 0 53 49
use INVX1  INVX1_172
timestamp 1516325494
transform 1 0 3376 0 -1 1533
box 0 0 11 49
use OR2X2  OR2X2_1888
timestamp 1516325494
transform -1 0 3407 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1978
timestamp 1516325494
transform -1 0 3426 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_766
timestamp 1516325494
transform -1 0 3434 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_766
timestamp 1516325494
transform -1 0 3448 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_1530
timestamp 1516325494
transform -1 0 3468 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1979
timestamp 1516325494
transform -1 0 3487 0 -1 1533
box 0 0 19 49
use INVX1  INVX1_169
timestamp 1516325494
transform 1 0 3487 0 -1 1533
box 0 0 11 49
use OR2X2  OR2X2_1529
timestamp 1516325494
transform -1 0 3517 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1701
timestamp 1516325494
transform -1 0 3536 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1528
timestamp 1516325494
transform -1 0 3555 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1702
timestamp 1516325494
transform -1 0 3574 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1703
timestamp 1516325494
transform -1 0 3593 0 -1 1533
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_146
timestamp 1516325494
transform 1 0 3593 0 -1 1533
box 0 0 53 49
use NAND2X1  NAND2X1_274
timestamp 1516325494
transform 1 0 3646 0 -1 1533
box 0 0 15 49
use MUX2X1  MUX2X1_274
timestamp 1516325494
transform -1 0 3691 0 -1 1533
box 0 0 30 49
use NAND2X1  NAND2X1_370
timestamp 1516325494
transform 1 0 3692 0 -1 1533
box 0 0 15 49
use FILL  FILL_AND2X2_150
timestamp 1516325494
transform -1 0 3715 0 -1 1533
box 0 0 8 49
use AND2X2  AND2X2_150
timestamp 1516325494
transform -1 0 3734 0 -1 1533
box 0 0 19 49
use FILL  FILL_BUFX2_586
timestamp 1516325494
transform -1 0 3742 0 -1 1533
box 0 0 8 49
use BUFX2  BUFX2_586
timestamp 1516325494
transform -1 0 3756 0 -1 1533
box 0 0 15 49
use AND2X2  AND2X2_2055
timestamp 1516325494
transform -1 0 3775 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1302
timestamp 1516325494
transform 1 0 3775 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1018
timestamp 1516325494
transform 1 0 3794 0 -1 1533
box 0 0 19 49
use OR2X2  OR2X2_1019
timestamp 1516325494
transform -1 0 3832 0 -1 1533
box 0 0 19 49
use AND2X2  AND2X2_1298
timestamp 1516325494
transform -1 0 3851 0 -1 1533
box 0 0 19 49
use BUFX2  BUFX2_866
timestamp 1516325494
transform -1 0 3866 0 -1 1533
box 0 0 15 49
use OR2X2  OR2X2_732
timestamp 1516325494
transform -1 0 21 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_750
timestamp 1516325494
transform 1 0 21 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_707
timestamp 1516325494
transform -1 0 59 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_706
timestamp 1516325494
transform -1 0 78 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_837
timestamp 1516325494
transform -1 0 97 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_612
timestamp 1516325494
transform -1 0 116 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_712
timestamp 1516325494
transform -1 0 135 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_803
timestamp 1516325494
transform 1 0 135 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_866
timestamp 1516325494
transform 1 0 154 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_608
timestamp 1516325494
transform -1 0 192 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_804
timestamp 1516325494
transform 1 0 192 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_673
timestamp 1516325494
transform -1 0 226 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_852
timestamp 1516325494
transform 1 0 226 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_763
timestamp 1516325494
transform -1 0 264 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_798
timestamp 1516325494
transform -1 0 283 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_605
timestamp 1516325494
transform -1 0 302 0 1 1434
box 0 0 19 49
use NOR2X1  NOR2X1_53
timestamp 1516325494
transform -1 0 317 0 1 1434
box 0 0 15 49
use INVX1  INVX1_9
timestamp 1516325494
transform -1 0 328 0 1 1434
box 0 0 11 49
use OR2X2  OR2X2_744
timestamp 1516325494
transform 1 0 329 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1034
timestamp 1516325494
transform -1 0 367 0 1 1434
box 0 0 19 49
use NOR2X1  NOR2X1_49
timestamp 1516325494
transform -1 0 382 0 1 1434
box 0 0 15 49
use INVX1  INVX1_55
timestamp 1516325494
transform -1 0 393 0 1 1434
box 0 0 11 49
use AND2X2  AND2X2_1026
timestamp 1516325494
transform -1 0 412 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_550
timestamp 1516325494
transform -1 0 431 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_781
timestamp 1516325494
transform -1 0 450 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_772
timestamp 1516325494
transform -1 0 469 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_671
timestamp 1516325494
transform 1 0 469 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_546
timestamp 1516325494
transform -1 0 507 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_975
timestamp 1516325494
transform 1 0 507 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1022
timestamp 1516325494
transform 1 0 526 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_739
timestamp 1516325494
transform -1 0 564 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_418
timestamp 1516325494
transform -1 0 583 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_976
timestamp 1516325494
transform 1 0 583 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_977
timestamp 1516325494
transform -1 0 621 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_609
timestamp 1516325494
transform -1 0 640 0 1 1434
box 0 0 19 49
use NAND3X1  NAND3X1_26
timestamp 1516325494
transform -1 0 659 0 1 1434
box 0 0 19 49
use NAND3X1  NAND3X1_25
timestamp 1516325494
transform -1 0 678 0 1 1434
box 0 0 19 49
use AOI21X1  AOI21X1_2
timestamp 1516325494
transform -1 0 697 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_653
timestamp 1516325494
transform -1 0 712 0 1 1434
box 0 0 15 49
use INVX1  INVX1_61
timestamp 1516325494
transform -1 0 724 0 1 1434
box 0 0 11 49
use NAND2X1  NAND2X1_652
timestamp 1516325494
transform -1 0 739 0 1 1434
box 0 0 15 49
use NAND3X1  NAND3X1_28
timestamp 1516325494
transform -1 0 758 0 1 1434
box 0 0 19 49
use NOR2X1  NOR2X1_29
timestamp 1516325494
transform -1 0 773 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_638
timestamp 1516325494
transform 1 0 773 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_655
timestamp 1516325494
transform -1 0 807 0 1 1434
box 0 0 15 49
use XNOR2X1  XNOR2X1_7
timestamp 1516325494
transform 1 0 808 0 1 1434
box 0 0 34 49
use AND2X2  AND2X2_1058
timestamp 1516325494
transform 1 0 842 0 1 1434
box 0 0 19 49
use INVX1  INVX1_27
timestamp 1516325494
transform 1 0 861 0 1 1434
box 0 0 11 49
use MUX2X1  MUX2X1_770
timestamp 1516325494
transform 1 0 872 0 1 1434
box 0 0 30 49
use AND2X2  AND2X2_1061
timestamp 1516325494
transform -1 0 922 0 1 1434
box 0 0 19 49
use MUX2X1  MUX2X1_765
timestamp 1516325494
transform 1 0 922 0 1 1434
box 0 0 30 49
use INVX1  INVX1_13
timestamp 1516325494
transform 1 0 952 0 1 1434
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_720
timestamp 1516325494
transform -1 0 1016 0 1 1434
box 0 0 53 49
use MUX2X1  MUX2X1_778
timestamp 1516325494
transform 1 0 1017 0 1 1434
box 0 0 30 49
use OR2X2  OR2X2_298
timestamp 1516325494
transform 1 0 1047 0 1 1434
box 0 0 19 49
use INVX1  INVX1_224
timestamp 1516325494
transform -1 0 1077 0 1 1434
box 0 0 11 49
use OR2X2  OR2X2_300
timestamp 1516325494
transform 1 0 1077 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_304
timestamp 1516325494
transform 1 0 1096 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_305
timestamp 1516325494
transform -1 0 1134 0 1 1434
box 0 0 19 49
use MUX2X1  MUX2X1_809
timestamp 1516325494
transform -1 0 1164 0 1 1434
box 0 0 30 49
use OR2X2  OR2X2_1742
timestamp 1516325494
transform -1 0 1184 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_375
timestamp 1516325494
transform -1 0 1203 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1984
timestamp 1516325494
transform -1 0 1222 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_2073
timestamp 1516325494
transform -1 0 1241 0 1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_746
timestamp 1516325494
transform -1 0 1249 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_746
timestamp 1516325494
transform -1 0 1263 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_568
timestamp 1516325494
transform -1 0 1272 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_568
timestamp 1516325494
transform -1 0 1286 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_660
timestamp 1516325494
transform 1 0 1286 0 1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_52
timestamp 1516325494
transform 1 0 1340 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_52
timestamp 1516325494
transform -1 0 1385 0 1 1434
box 0 0 30 49
use AND2X2  AND2X2_2075
timestamp 1516325494
transform 1 0 1385 0 1 1434
box 0 0 19 49
use INVX1  INVX1_140
timestamp 1516325494
transform 1 0 1404 0 1 1434
box 0 0 11 49
use AND2X2  AND2X2_323
timestamp 1516325494
transform -1 0 1435 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1878
timestamp 1516325494
transform -1 0 1454 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1914
timestamp 1516325494
transform -1 0 1473 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1984
timestamp 1516325494
transform -1 0 1492 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1896
timestamp 1516325494
transform -1 0 1511 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1897
timestamp 1516325494
transform -1 0 1530 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_446
timestamp 1516325494
transform 1 0 1530 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_62
timestamp 1516325494
transform 1 0 1545 0 1 1434
box 0 0 53 49
use MUX2X1  MUX2X1_446
timestamp 1516325494
transform -1 0 1628 0 1 1434
box 0 0 30 49
use OAI21X1  OAI21X1_18
timestamp 1516325494
transform 1 0 1628 0 1 1434
box 0 0 19 49
use INVX2  INVX2_7
timestamp 1516325494
transform 1 0 1647 0 1 1434
box 0 0 11 49
use FILL  FILL_BUFX2_529
timestamp 1516325494
transform 1 0 1659 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_529
timestamp 1516325494
transform 1 0 1666 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_1272
timestamp 1516325494
transform -1 0 1701 0 1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_361
timestamp 1516325494
transform 1 0 1701 0 1 1434
box 0 0 53 49
use MUX2X1  MUX2X1_864
timestamp 1516325494
transform 1 0 1754 0 1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_919
timestamp 1516325494
transform 1 0 1784 0 1 1434
box 0 0 15 49
use OAI21X1  OAI21X1_37
timestamp 1516325494
transform 1 0 1799 0 1 1434
box 0 0 19 49
use INVX2  INVX2_26
timestamp 1516325494
transform 1 0 1818 0 1 1434
box 0 0 11 49
use NAND2X1  NAND2X1_734
timestamp 1516325494
transform -1 0 1845 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_137
timestamp 1516325494
transform 1 0 1845 0 1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_908
timestamp 1516325494
transform 1 0 1875 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_853
timestamp 1516325494
transform -1 0 1921 0 1 1434
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_638
timestamp 1516325494
transform 1 0 1921 0 1 1434
box 0 0 53 49
use AND2X2  AND2X2_1877
timestamp 1516325494
transform -1 0 1993 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1757
timestamp 1516325494
transform -1 0 2012 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1758
timestamp 1516325494
transform -1 0 2031 0 1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_25
timestamp 1516325494
transform 1 0 2031 0 1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_121
timestamp 1516325494
transform 1 0 2084 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_121
timestamp 1516325494
transform -1 0 2130 0 1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_548
timestamp 1516325494
transform -1 0 2145 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_548
timestamp 1516325494
transform -1 0 2175 0 1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_35
timestamp 1516325494
transform -1 0 2184 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_35
timestamp 1516325494
transform -1 0 2198 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_1129
timestamp 1516325494
transform 1 0 2198 0 1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_3
timestamp 1516325494
transform -1 0 2225 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_3
timestamp 1516325494
transform -1 0 2240 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_240
timestamp 1516325494
transform -1 0 2248 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_240
timestamp 1516325494
transform -1 0 2263 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_194
timestamp 1516325494
transform -1 0 2271 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_194
timestamp 1516325494
transform -1 0 2286 0 1 1434
box 0 0 15 49
use AND2X2  AND2X2_1394
timestamp 1516325494
transform -1 0 2305 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1127
timestamp 1516325494
transform -1 0 2324 0 1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_116
timestamp 1516325494
transform -1 0 2332 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_116
timestamp 1516325494
transform -1 0 2346 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_1128
timestamp 1516325494
transform -1 0 2366 0 1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_4
timestamp 1516325494
transform 1 0 2366 0 1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_100
timestamp 1516325494
transform 1 0 2419 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_100
timestamp 1516325494
transform -1 0 2464 0 1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_63
timestamp 1516325494
transform 1 0 2464 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_63
timestamp 1516325494
transform 1 0 2472 0 1 1434
box 0 0 15 49
use INVX2  INVX2_38
timestamp 1516325494
transform 1 0 2487 0 1 1434
box 0 0 11 49
use FILL  FILL_BUFX2_389
timestamp 1516325494
transform 1 0 2499 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_389
timestamp 1516325494
transform 1 0 2506 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_454
timestamp 1516325494
transform -1 0 2529 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_454
timestamp 1516325494
transform -1 0 2544 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_643
timestamp 1516325494
transform 1 0 2544 0 1 1434
box 0 0 53 49
use OR2X2  OR2X2_1089
timestamp 1516325494
transform -1 0 2616 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_483
timestamp 1516325494
transform -1 0 2631 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_223
timestamp 1516325494
transform 1 0 2632 0 1 1434
box 0 0 53 49
use AND2X2  AND2X2_2093
timestamp 1516325494
transform -1 0 2704 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_227
timestamp 1516325494
transform -1 0 2719 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_40
timestamp 1516325494
transform -1 0 2727 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_40
timestamp 1516325494
transform -1 0 2742 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_452
timestamp 1516325494
transform -1 0 2750 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_452
timestamp 1516325494
transform -1 0 2764 0 1 1434
box 0 0 15 49
use AND2X2  AND2X2_1352
timestamp 1516325494
transform 1 0 2765 0 1 1434
box 0 0 19 49
use MUX2X1  MUX2X1_254
timestamp 1516325494
transform 1 0 2784 0 1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_254
timestamp 1516325494
transform -1 0 2829 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_190
timestamp 1516325494
transform -1 0 2882 0 1 1434
box 0 0 53 49
use FILL  FILL_BUFX2_524
timestamp 1516325494
transform 1 0 2882 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_524
timestamp 1516325494
transform 1 0 2890 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_523
timestamp 1516325494
transform -1 0 2913 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_523
timestamp 1516325494
transform -1 0 2928 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_259
timestamp 1516325494
transform 1 0 2928 0 1 1434
box 0 0 53 49
use OR2X2  OR2X2_1890
timestamp 1516325494
transform -1 0 3000 0 1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_6
timestamp 1516325494
transform -1 0 3008 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_6
timestamp 1516325494
transform -1 0 3023 0 1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_337
timestamp 1516325494
transform 1 0 3023 0 1 1434
box 0 0 8 49
use BUFX2  BUFX2_337
timestamp 1516325494
transform 1 0 3031 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_367
timestamp 1516325494
transform -1 0 3065 0 1 1434
box 0 0 19 49
use OAI21X1  OAI21X1_59
timestamp 1516325494
transform -1 0 3084 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_594
timestamp 1516325494
transform -1 0 3099 0 1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_238
timestamp 1516325494
transform 1 0 3099 0 1 1434
box 0 0 53 49
use FILL  FILL_AND2X2_208
timestamp 1516325494
transform 1 0 3152 0 1 1434
box 0 0 8 49
use AND2X2  AND2X2_208
timestamp 1516325494
transform 1 0 3160 0 1 1434
box 0 0 19 49
use FILL  FILL_AND2X2_148
timestamp 1516325494
transform 1 0 3179 0 1 1434
box 0 0 8 49
use AND2X2  AND2X2_148
timestamp 1516325494
transform 1 0 3186 0 1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_590
timestamp 1516325494
transform 1 0 3205 0 1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_590
timestamp 1516325494
transform -1 0 3251 0 1 1434
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_270
timestamp 1516325494
transform 1 0 3251 0 1 1434
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_210
timestamp 1516325494
transform 1 0 3304 0 1 1434
box 0 0 53 49
use OR2X2  OR2X2_1889
timestamp 1516325494
transform -1 0 3376 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1977
timestamp 1516325494
transform -1 0 3395 0 1 1434
box 0 0 19 49
use FILL  FILL_OR2X2_138
timestamp 1516325494
transform -1 0 3403 0 1 1434
box 0 0 8 49
use OR2X2  OR2X2_138
timestamp 1516325494
transform -1 0 3422 0 1 1434
box 0 0 19 49
use FILL  FILL_AND2X2_145
timestamp 1516325494
transform -1 0 3430 0 1 1434
box 0 0 8 49
use AND2X2  AND2X2_145
timestamp 1516325494
transform -1 0 3449 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1405
timestamp 1516325494
transform -1 0 3468 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1605
timestamp 1516325494
transform -1 0 3487 0 1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_206
timestamp 1516325494
transform 1 0 3487 0 1 1434
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_174
timestamp 1516325494
transform 1 0 3540 0 1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_238
timestamp 1516325494
transform 1 0 3593 0 1 1434
box 0 0 15 49
use OR2X2  OR2X2_1409
timestamp 1516325494
transform -1 0 3627 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1609
timestamp 1516325494
transform -1 0 3646 0 1 1434
box 0 0 19 49
use FILL  FILL_AND2X2_151
timestamp 1516325494
transform 1 0 3646 0 1 1434
box 0 0 8 49
use AND2X2  AND2X2_151
timestamp 1516325494
transform 1 0 3654 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1611
timestamp 1516325494
transform 1 0 3673 0 1 1434
box 0 0 19 49
use OR2X2  OR2X2_1408
timestamp 1516325494
transform -1 0 3711 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_1610
timestamp 1516325494
transform -1 0 3730 0 1 1434
box 0 0 19 49
use AND2X2  AND2X2_2057
timestamp 1516325494
transform 1 0 3730 0 1 1434
box 0 0 19 49
use MUX2X1  MUX2X1_257
timestamp 1516325494
transform 1 0 3749 0 1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_257
timestamp 1516325494
transform -1 0 3794 0 1 1434
box 0 0 15 49
use AND2X2  AND2X2_1300
timestamp 1516325494
transform -1 0 3813 0 1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_129
timestamp 1516325494
transform -1 0 3866 0 1 1434
box 0 0 53 49
use FILL  FILL_BUFX2_303
timestamp 1516325494
transform -1 0 10 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_303
timestamp 1516325494
transform -1 0 25 0 -1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_302
timestamp 1516325494
transform -1 0 33 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_302
timestamp 1516325494
transform -1 0 47 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_770
timestamp 1516325494
transform -1 0 67 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_496
timestamp 1516325494
transform 1 0 67 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_965
timestamp 1516325494
transform 1 0 86 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_301
timestamp 1516325494
transform -1 0 113 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_301
timestamp 1516325494
transform -1 0 127 0 -1 1434
box 0 0 15 49
use OR2X2  OR2X2_802
timestamp 1516325494
transform 1 0 127 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_820
timestamp 1516325494
transform 1 0 146 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_83
timestamp 1516325494
transform 1 0 165 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_83
timestamp 1516325494
transform 1 0 173 0 -1 1434
box 0 0 15 49
use OR2X2  OR2X2_854
timestamp 1516325494
transform 1 0 188 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_943
timestamp 1516325494
transform -1 0 226 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_843
timestamp 1516325494
transform 1 0 226 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_843
timestamp 1516325494
transform 1 0 234 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_987
timestamp 1516325494
transform 1 0 249 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1033
timestamp 1516325494
transform -1 0 287 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_477
timestamp 1516325494
transform -1 0 306 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_478
timestamp 1516325494
transform 1 0 306 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_426
timestamp 1516325494
transform -1 0 344 0 -1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_644
timestamp 1516325494
transform -1 0 359 0 -1 1434
box 0 0 15 49
use AOI22X1  AOI22X1_1
timestamp 1516325494
transform -1 0 382 0 -1 1434
box 0 0 23 49
use OR2X2  OR2X2_558
timestamp 1516325494
transform 1 0 382 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_660
timestamp 1516325494
transform 1 0 401 0 -1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_649
timestamp 1516325494
transform -1 0 435 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_829
timestamp 1516325494
transform -1 0 454 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_300
timestamp 1516325494
transform -1 0 462 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_300
timestamp 1516325494
transform -1 0 477 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_481
timestamp 1516325494
transform 1 0 477 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1019
timestamp 1516325494
transform 1 0 496 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1020
timestamp 1516325494
transform -1 0 534 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_762
timestamp 1516325494
transform 1 0 534 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_610
timestamp 1516325494
transform -1 0 572 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_763
timestamp 1516325494
transform 1 0 572 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_522
timestamp 1516325494
transform -1 0 610 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_727
timestamp 1516325494
transform 1 0 610 0 -1 1434
box 0 0 19 49
use NOR2X1  NOR2X1_26
timestamp 1516325494
transform -1 0 644 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_764
timestamp 1516325494
transform 1 0 644 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_684
timestamp 1516325494
transform -1 0 682 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_683
timestamp 1516325494
transform -1 0 701 0 -1 1434
box 0 0 19 49
use NAND3X1  NAND3X1_29
timestamp 1516325494
transform -1 0 720 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_954
timestamp 1516325494
transform 1 0 720 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_577
timestamp 1516325494
transform -1 0 758 0 -1 1434
box 0 0 19 49
use AOI21X1  AOI21X1_5
timestamp 1516325494
transform -1 0 777 0 -1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_656
timestamp 1516325494
transform -1 0 792 0 -1 1434
box 0 0 15 49
use AOI21X1  AOI21X1_1
timestamp 1516325494
transform 1 0 792 0 -1 1434
box 0 0 19 49
use NOR2X1  NOR2X1_40
timestamp 1516325494
transform 1 0 811 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_1068
timestamp 1516325494
transform 1 0 827 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1059
timestamp 1516325494
transform 1 0 846 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1060
timestamp 1516325494
transform -1 0 884 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1085
timestamp 1516325494
transform 1 0 884 0 -1 1434
box 0 0 19 49
use INVX1  INVX1_158
timestamp 1516325494
transform 1 0 903 0 -1 1434
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_727
timestamp 1516325494
transform -1 0 967 0 -1 1434
box 0 0 53 49
use MUX2X1  MUX2X1_797
timestamp 1516325494
transform -1 0 997 0 -1 1434
box 0 0 30 49
use MUX2X1  MUX2X1_802
timestamp 1516325494
transform -1 0 1028 0 -1 1434
box 0 0 30 49
use INVX1  INVX1_200
timestamp 1516325494
transform -1 0 1039 0 -1 1434
box 0 0 11 49
use INVX1  INVX1_135
timestamp 1516325494
transform 1 0 1039 0 -1 1434
box 0 0 11 49
use OR2X2  OR2X2_443
timestamp 1516325494
transform -1 0 21 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_495
timestamp 1516325494
transform -1 0 40 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_645
timestamp 1516325494
transform 1 0 40 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_705
timestamp 1516325494
transform 1 0 59 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_735
timestamp 1516325494
transform -1 0 97 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_611
timestamp 1516325494
transform -1 0 116 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_869
timestamp 1516325494
transform 1 0 116 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_786
timestamp 1516325494
transform 1 0 135 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_702
timestamp 1516325494
transform -1 0 173 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_812
timestamp 1516325494
transform -1 0 192 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_747
timestamp 1516325494
transform -1 0 211 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_944
timestamp 1516325494
transform 1 0 211 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_813
timestamp 1516325494
transform 1 0 230 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_684
timestamp 1516325494
transform 1 0 249 0 1 1336
box 0 0 19 49
use INVX1  INVX1_20
timestamp 1516325494
transform -1 0 279 0 1 1336
box 0 0 11 49
use AND2X2  AND2X2_988
timestamp 1516325494
transform 1 0 279 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_520
timestamp 1516325494
transform 1 0 298 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_989
timestamp 1516325494
transform 1 0 317 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_641
timestamp 1516325494
transform 1 0 336 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_612
timestamp 1516325494
transform -1 0 374 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_611
timestamp 1516325494
transform 1 0 374 0 1 1336
box 0 0 19 49
use NAND2X1  NAND2X1_643
timestamp 1516325494
transform -1 0 408 0 1 1336
box 0 0 15 49
use INVX1  INVX1_15
timestamp 1516325494
transform -1 0 420 0 1 1336
box 0 0 11 49
use AND2X2  AND2X2_830
timestamp 1516325494
transform 1 0 420 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_945
timestamp 1516325494
transform 1 0 439 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_670
timestamp 1516325494
transform 1 0 458 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_831
timestamp 1516325494
transform -1 0 496 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_811
timestamp 1516325494
transform 1 0 496 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_993
timestamp 1516325494
transform 1 0 515 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_695
timestamp 1516325494
transform -1 0 553 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_849
timestamp 1516325494
transform 1 0 553 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1021
timestamp 1516325494
transform 1 0 572 0 1 1336
box 0 0 19 49
use FILL  FILL_BUFX2_81
timestamp 1516325494
transform 1 0 591 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_81
timestamp 1516325494
transform 1 0 599 0 1 1336
box 0 0 15 49
use OR2X2  OR2X2_777
timestamp 1516325494
transform -1 0 633 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_847
timestamp 1516325494
transform -1 0 652 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_631
timestamp 1516325494
transform -1 0 671 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_994
timestamp 1516325494
transform 1 0 671 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1002
timestamp 1516325494
transform 1 0 690 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_824
timestamp 1516325494
transform -1 0 728 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_796
timestamp 1516325494
transform -1 0 747 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_592
timestamp 1516325494
transform -1 0 766 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_957
timestamp 1516325494
transform -1 0 785 0 1 1336
box 0 0 19 49
use NAND2X1  NAND2X1_648
timestamp 1516325494
transform 1 0 785 0 1 1336
box 0 0 15 49
use NAND3X1  NAND3X1_18
timestamp 1516325494
transform 1 0 800 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_454
timestamp 1516325494
transform 1 0 819 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1056
timestamp 1516325494
transform 1 0 838 0 1 1336
box 0 0 19 49
use NOR2X1  NOR2X1_21
timestamp 1516325494
transform -1 0 872 0 1 1336
box 0 0 15 49
use AND2X2  AND2X2_1057
timestamp 1516325494
transform 1 0 872 0 1 1336
box 0 0 19 49
use INVX1  INVX1_30
timestamp 1516325494
transform 1 0 891 0 1 1336
box 0 0 11 49
use FILL  FILL_BUFX2_626
timestamp 1516325494
transform -1 0 911 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_626
timestamp 1516325494
transform -1 0 925 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_730
timestamp 1516325494
transform -1 0 978 0 1 1336
box 0 0 53 49
use MUX2X1  MUX2X1_758
timestamp 1516325494
transform 1 0 979 0 1 1336
box 0 0 30 49
use MUX2X1  MUX2X1_755
timestamp 1516325494
transform 1 0 1009 0 1 1336
box 0 0 30 49
use INVX1  INVX1_153
timestamp 1516325494
transform 1 0 1039 0 1 1336
box 0 0 11 49
use MUX2X1  MUX2X1_747
timestamp 1516325494
transform 1 0 1051 0 -1 1434
box 0 0 30 49
use OR2X2  OR2X2_299
timestamp 1516325494
transform -1 0 1100 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1044
timestamp 1516325494
transform -1 0 1119 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1871
timestamp 1516325494
transform -1 0 1138 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1043
timestamp 1516325494
transform -1 0 1157 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1749
timestamp 1516325494
transform -1 0 1176 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1042
timestamp 1516325494
transform -1 0 1195 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1986
timestamp 1516325494
transform -1 0 1214 0 -1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_313
timestamp 1516325494
transform 1 0 1214 0 -1 1434
box 0 0 53 49
use AND2X2  AND2X2_1985
timestamp 1516325494
transform -1 0 1286 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1598
timestamp 1516325494
transform -1 0 1305 0 -1 1434
box 0 0 19 49
use MUX2X1  MUX2X1_505
timestamp 1516325494
transform 1 0 1305 0 -1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_505
timestamp 1516325494
transform 1 0 1336 0 -1 1434
box 0 0 15 49
use OR2X2  OR2X2_1041
timestamp 1516325494
transform -1 0 1370 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1325
timestamp 1516325494
transform -1 0 1389 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1985
timestamp 1516325494
transform -1 0 1408 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1328
timestamp 1516325494
transform -1 0 1427 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_2077
timestamp 1516325494
transform -1 0 1446 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1746
timestamp 1516325494
transform -1 0 1465 0 -1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_633
timestamp 1516325494
transform 1 0 1465 0 -1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_903
timestamp 1516325494
transform 1 0 1518 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_848
timestamp 1516325494
transform -1 0 1563 0 -1 1434
box 0 0 30 49
use AND2X2  AND2X2_2035
timestamp 1516325494
transform 1 0 1564 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1966
timestamp 1516325494
transform 1 0 1583 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_2037
timestamp 1516325494
transform -1 0 1621 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1505
timestamp 1516325494
transform -1 0 1640 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1273
timestamp 1516325494
transform -1 0 1659 0 -1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_393
timestamp 1516325494
transform 1 0 1659 0 -1 1434
box 0 0 53 49
use AND2X2  AND2X2_427
timestamp 1516325494
transform 1 0 1712 0 -1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_169
timestamp 1516325494
transform 1 0 1731 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_169
timestamp 1516325494
transform 1 0 1746 0 -1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_448
timestamp 1516325494
transform -1 0 1785 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_448
timestamp 1516325494
transform -1 0 1799 0 -1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_631
timestamp 1516325494
transform 1 0 1799 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_631
timestamp 1516325494
transform 1 0 1807 0 -1 1434
box 0 0 15 49
use OR2X2  OR2X2_1905
timestamp 1516325494
transform 1 0 1822 0 -1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_137
timestamp 1516325494
transform 1 0 1841 0 -1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_73
timestamp 1516325494
transform 1 0 1856 0 -1 1434
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_94
timestamp 1516325494
transform 1 0 1910 0 -1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_158
timestamp 1516325494
transform 1 0 1963 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_158
timestamp 1516325494
transform 1 0 1978 0 -1 1434
box 0 0 30 49
use OR2X2  OR2X2_1759
timestamp 1516325494
transform -1 0 2027 0 -1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_641
timestamp 1516325494
transform 1 0 2027 0 -1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_569
timestamp 1516325494
transform 1 0 2081 0 -1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_505
timestamp 1516325494
transform 1 0 2096 0 -1 1434
box 0 0 53 49
use MUX2X1  MUX2X1_569
timestamp 1516325494
transform -1 0 2179 0 -1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_47
timestamp 1516325494
transform -1 0 2187 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_47
timestamp 1516325494
transform -1 0 2202 0 -1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_510
timestamp 1516325494
transform 1 0 2202 0 -1 1434
box 0 0 53 49
use OR2X2  OR2X2_1969
timestamp 1516325494
transform -1 0 2274 0 -1 1434
box 0 0 19 49
use MUX2X1  MUX2X1_576
timestamp 1516325494
transform 1 0 2274 0 -1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_576
timestamp 1516325494
transform -1 0 2320 0 -1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_512
timestamp 1516325494
transform -1 0 2373 0 -1 1434
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_128
timestamp 1516325494
transform 1 0 2373 0 -1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_96
timestamp 1516325494
transform 1 0 2426 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_96
timestamp 1516325494
transform -1 0 2472 0 -1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_429
timestamp 1516325494
transform -1 0 2480 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_429
timestamp 1516325494
transform -1 0 2495 0 -1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_30
timestamp 1516325494
transform -1 0 2503 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_30
timestamp 1516325494
transform -1 0 2517 0 -1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_675
timestamp 1516325494
transform 1 0 2518 0 -1 1434
box 0 0 53 49
use NAND2X1  NAND2X1_291
timestamp 1516325494
transform 1 0 2571 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_291
timestamp 1516325494
transform -1 0 2616 0 -1 1434
box 0 0 30 49
use MUX2X1  MUX2X1_483
timestamp 1516325494
transform -1 0 2646 0 -1 1434
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_291
timestamp 1516325494
transform -1 0 2700 0 -1 1434
box 0 0 53 49
use MUX2X1  MUX2X1_227
timestamp 1516325494
transform -1 0 2730 0 -1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_430
timestamp 1516325494
transform -1 0 2738 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_430
timestamp 1516325494
transform -1 0 2753 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_225
timestamp 1516325494
transform 1 0 2753 0 -1 1434
box 0 0 30 49
use NAND2X1  NAND2X1_225
timestamp 1516325494
transform -1 0 2799 0 -1 1434
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_161
timestamp 1516325494
transform -1 0 2852 0 -1 1434
box 0 0 53 49
use AND2X2  AND2X2_2044
timestamp 1516325494
transform 1 0 2852 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1287
timestamp 1516325494
transform 1 0 2871 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_560
timestamp 1516325494
transform 1 0 2890 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_560
timestamp 1516325494
transform 1 0 2898 0 -1 1434
box 0 0 15 49
use AND2X2  AND2X2_1973
timestamp 1516325494
transform 1 0 2913 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_385
timestamp 1516325494
transform 1 0 2932 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1974
timestamp 1516325494
transform 1 0 2951 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1885
timestamp 1516325494
transform 1 0 2970 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1887
timestamp 1516325494
transform -1 0 3008 0 -1 1434
box 0 0 19 49
use OAI21X1  OAI21X1_58
timestamp 1516325494
transform 1 0 3008 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1020
timestamp 1516325494
transform -1 0 3046 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_336
timestamp 1516325494
transform 1 0 3046 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_336
timestamp 1516325494
transform 1 0 3053 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_594
timestamp 1516325494
transform 1 0 3069 0 -1 1434
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_274
timestamp 1516325494
transform -1 0 3152 0 -1 1434
box 0 0 53 49
use FILL  FILL_BUFX2_338
timestamp 1516325494
transform -1 0 3160 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_338
timestamp 1516325494
transform -1 0 3175 0 -1 1434
box 0 0 15 49
use FILL  FILL_OR2X2_195
timestamp 1516325494
transform 1 0 3175 0 -1 1434
box 0 0 8 49
use OR2X2  OR2X2_195
timestamp 1516325494
transform 1 0 3183 0 -1 1434
box 0 0 19 49
use FILL  FILL_OR2X2_196
timestamp 1516325494
transform -1 0 3210 0 -1 1434
box 0 0 8 49
use OR2X2  OR2X2_196
timestamp 1516325494
transform -1 0 3228 0 -1 1434
box 0 0 19 49
use FILL  FILL_AND2X2_207
timestamp 1516325494
transform -1 0 3236 0 -1 1434
box 0 0 8 49
use AND2X2  AND2X2_207
timestamp 1516325494
transform -1 0 3255 0 -1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_242
timestamp 1516325494
transform 1 0 3255 0 -1 1434
box 0 0 53 49
use FILL  FILL_OR2X2_194
timestamp 1516325494
transform -1 0 3316 0 -1 1434
box 0 0 8 49
use OR2X2  OR2X2_194
timestamp 1516325494
transform -1 0 3335 0 -1 1434
box 0 0 19 49
use FILL  FILL_AND2X2_206
timestamp 1516325494
transform -1 0 3343 0 -1 1434
box 0 0 8 49
use AND2X2  AND2X2_206
timestamp 1516325494
transform -1 0 3361 0 -1 1434
box 0 0 19 49
use NAND2X1  NAND2X1_626
timestamp 1516325494
transform 1 0 3361 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_626
timestamp 1516325494
transform -1 0 3406 0 -1 1434
box 0 0 30 49
use FILL  FILL_AND2X2_205
timestamp 1516325494
transform -1 0 3415 0 -1 1434
box 0 0 8 49
use AND2X2  AND2X2_205
timestamp 1516325494
transform -1 0 3433 0 -1 1434
box 0 0 19 49
use FILL  FILL_AND2X2_146
timestamp 1516325494
transform -1 0 3441 0 -1 1434
box 0 0 8 49
use AND2X2  AND2X2_146
timestamp 1516325494
transform -1 0 3460 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_1606
timestamp 1516325494
transform -1 0 3479 0 -1 1434
box 0 0 19 49
use FILL  FILL_BUFX2_659
timestamp 1516325494
transform -1 0 3487 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_659
timestamp 1516325494
transform -1 0 3502 0 -1 1434
box 0 0 15 49
use NAND2X1  NAND2X1_622
timestamp 1516325494
transform 1 0 3502 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_622
timestamp 1516325494
transform -1 0 3547 0 -1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_455
timestamp 1516325494
transform -1 0 3555 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_455
timestamp 1516325494
transform -1 0 3570 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_238
timestamp 1516325494
transform 1 0 3570 0 -1 1434
box 0 0 30 49
use FILL  FILL_BUFX2_478
timestamp 1516325494
transform 1 0 3601 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_478
timestamp 1516325494
transform 1 0 3608 0 -1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_225
timestamp 1516325494
transform -1 0 3631 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_225
timestamp 1516325494
transform -1 0 3646 0 -1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_328
timestamp 1516325494
transform -1 0 3654 0 -1 1434
box 0 0 8 49
use BUFX2  BUFX2_328
timestamp 1516325494
transform -1 0 3669 0 -1 1434
box 0 0 15 49
use NAND2X1  NAND2X1_366
timestamp 1516325494
transform 1 0 3669 0 -1 1434
box 0 0 15 49
use MUX2X1  MUX2X1_366
timestamp 1516325494
transform -1 0 3714 0 -1 1434
box 0 0 30 49
use OR2X2  OR2X2_1979
timestamp 1516325494
transform -1 0 3734 0 -1 1434
box 0 0 19 49
use OR2X2  OR2X2_1978
timestamp 1516325494
transform -1 0 3753 0 -1 1434
box 0 0 19 49
use AND2X2  AND2X2_2059
timestamp 1516325494
transform -1 0 3772 0 -1 1434
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_799
timestamp 1516325494
transform 1 0 3772 0 -1 1434
box 0 0 53 49
use OR2X2  OR2X2_973
timestamp 1516325494
transform 1 0 3825 0 -1 1434
box 0 0 19 49
use INVX1  INVX1_315
timestamp 1516325494
transform -1 0 3855 0 -1 1434
box 0 0 11 49
use BUFX2  BUFX2_909
timestamp 1516325494
transform -1 0 3870 0 -1 1434
box 0 0 15 49
use FILL  FILL_BUFX2_850
timestamp 1516325494
transform -1 0 1059 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_850
timestamp 1516325494
transform -1 0 1073 0 1 1336
box 0 0 15 49
use OR2X2  OR2X2_1750
timestamp 1516325494
transform -1 0 1093 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_320
timestamp 1516325494
transform -1 0 1112 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_319
timestamp 1516325494
transform -1 0 1131 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1870
timestamp 1516325494
transform -1 0 1150 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1988
timestamp 1516325494
transform -1 0 1169 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1987
timestamp 1516325494
transform -1 0 1188 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_374
timestamp 1516325494
transform -1 0 1207 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_370
timestamp 1516325494
transform -1 0 1226 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_369
timestamp 1516325494
transform -1 0 1245 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_394
timestamp 1516325494
transform -1 0 1264 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1418
timestamp 1516325494
transform 1 0 1264 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1869
timestamp 1516325494
transform -1 0 1302 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1747
timestamp 1516325494
transform -1 0 1321 0 1 1336
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_57
timestamp 1516325494
transform 1 0 1321 0 1 1336
box 0 0 53 49
use NAND2X1  NAND2X1_441
timestamp 1516325494
transform 1 0 1374 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_441
timestamp 1516325494
transform -1 0 1419 0 1 1336
box 0 0 30 49
use FILL  FILL_BUFX2_94
timestamp 1516325494
transform -1 0 1427 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_94
timestamp 1516325494
transform -1 0 1442 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_441
timestamp 1516325494
transform 1 0 1442 0 1 1336
box 0 0 53 49
use NAND2X1  NAND2X1_409
timestamp 1516325494
transform 1 0 1495 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_409
timestamp 1516325494
transform -1 0 1541 0 1 1336
box 0 0 30 49
use FILL  FILL_BUFX2_445
timestamp 1516325494
transform -1 0 1549 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_445
timestamp 1516325494
transform -1 0 1564 0 1 1336
box 0 0 15 49
use NAND2X1  NAND2X1_930
timestamp 1516325494
transform -1 0 1579 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_875
timestamp 1516325494
transform 1 0 1579 0 1 1336
box 0 0 30 49
use OAI21X1  OAI21X1_36
timestamp 1516325494
transform -1 0 1628 0 1 1336
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_372
timestamp 1516325494
transform -1 0 1681 0 1 1336
box 0 0 53 49
use AND2X2  AND2X2_426
timestamp 1516325494
transform 1 0 1682 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1602
timestamp 1516325494
transform 1 0 1701 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_399
timestamp 1516325494
transform 1 0 1720 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1758
timestamp 1516325494
transform -1 0 1758 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1603
timestamp 1516325494
transform -1 0 1777 0 1 1336
box 0 0 19 49
use NAND2X1  NAND2X1_180
timestamp 1516325494
transform 1 0 1777 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_180
timestamp 1516325494
transform 1 0 1792 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_404
timestamp 1516325494
transform -1 0 1875 0 1 1336
box 0 0 53 49
use OR2X2  OR2X2_1362
timestamp 1516325494
transform -1 0 1894 0 1 1336
box 0 0 19 49
use FILL  FILL_BUFX2_12
timestamp 1516325494
transform 1 0 1894 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_12
timestamp 1516325494
transform 1 0 1902 0 1 1336
box 0 0 15 49
use NAND2X1  NAND2X1_922
timestamp 1516325494
transform 1 0 1917 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_867
timestamp 1516325494
transform 1 0 1932 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_364
timestamp 1516325494
transform -1 0 2016 0 1 1336
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_478
timestamp 1516325494
transform 1 0 2016 0 1 1336
box 0 0 53 49
use NAND2X1  NAND2X1_350
timestamp 1516325494
transform 1 0 2069 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_350
timestamp 1516325494
transform -1 0 2114 0 1 1336
box 0 0 30 49
use MUX2X1  MUX2X1_172
timestamp 1516325494
transform 1 0 2115 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_396
timestamp 1516325494
transform -1 0 2198 0 1 1336
box 0 0 53 49
use NAND2X1  NAND2X1_33
timestamp 1516325494
transform 1 0 2198 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_33
timestamp 1516325494
transform -1 0 2244 0 1 1336
box 0 0 30 49
use MUX2X1  MUX2X1_824
timestamp 1516325494
transform 1 0 2244 0 1 1336
box 0 0 30 49
use NAND2X1  NAND2X1_879
timestamp 1516325494
transform -1 0 2289 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_609
timestamp 1516325494
transform -1 0 2343 0 1 1336
box 0 0 53 49
use MUX2X1  MUX2X1_574
timestamp 1516325494
transform 1 0 2343 0 1 1336
box 0 0 30 49
use NAND2X1  NAND2X1_574
timestamp 1516325494
transform -1 0 2388 0 1 1336
box 0 0 15 49
use OR2X2  OR2X2_1909
timestamp 1516325494
transform 1 0 2388 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1970
timestamp 1516325494
transform -1 0 2426 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1994
timestamp 1516325494
transform -1 0 2445 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1910
timestamp 1516325494
transform -1 0 2464 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1327
timestamp 1516325494
transform -1 0 2483 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1040
timestamp 1516325494
transform -1 0 2502 0 1 1336
box 0 0 19 49
use FILL  FILL_BUFX2_53
timestamp 1516325494
transform 1 0 2502 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_53
timestamp 1516325494
transform 1 0 2510 0 1 1336
box 0 0 15 49
use FILL  FILL_BUFX2_145
timestamp 1516325494
transform 1 0 2525 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_145
timestamp 1516325494
transform 1 0 2533 0 1 1336
box 0 0 15 49
use FILL  FILL_BUFX2_136
timestamp 1516325494
transform 1 0 2548 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_136
timestamp 1516325494
transform 1 0 2556 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_97
timestamp 1516325494
transform -1 0 2624 0 1 1336
box 0 0 53 49
use OR2X2  OR2X2_1908
timestamp 1516325494
transform -1 0 2643 0 1 1336
box 0 0 19 49
use FILL  FILL_BUFX2_513
timestamp 1516325494
transform -1 0 2651 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_513
timestamp 1516325494
transform -1 0 2666 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_30
timestamp 1516325494
transform 1 0 2666 0 1 1336
box 0 0 53 49
use NAND2X1  NAND2X1_126
timestamp 1516325494
transform 1 0 2719 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_126
timestamp 1516325494
transform -1 0 2764 0 1 1336
box 0 0 30 49
use NAND2X1  NAND2X1_94
timestamp 1516325494
transform 1 0 2765 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_94
timestamp 1516325494
transform -1 0 2810 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_126
timestamp 1516325494
transform -1 0 2863 0 1 1336
box 0 0 53 49
use OR2X2  OR2X2_1980
timestamp 1516325494
transform -1 0 2882 0 1 1336
box 0 0 19 49
use FILL  FILL_BUFX2_530
timestamp 1516325494
transform -1 0 2890 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_530
timestamp 1516325494
transform -1 0 2905 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_163
timestamp 1516325494
transform -1 0 2958 0 1 1336
box 0 0 53 49
use FILL  FILL_BUFX2_161
timestamp 1516325494
transform -1 0 2966 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_161
timestamp 1516325494
transform -1 0 2981 0 1 1336
box 0 0 15 49
use AND2X2  AND2X2_1290
timestamp 1516325494
transform 1 0 2981 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1015
timestamp 1516325494
transform 1 0 3000 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1017
timestamp 1516325494
transform 1 0 3019 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_362
timestamp 1516325494
transform 1 0 3038 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_364
timestamp 1516325494
transform -1 0 3076 0 1 1336
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_193
timestamp 1516325494
transform -1 0 3129 0 1 1336
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_257
timestamp 1516325494
transform -1 0 3182 0 1 1336
box 0 0 53 49
use OR2X2  OR2X2_1886
timestamp 1516325494
transform -1 0 3202 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1976
timestamp 1516325494
transform -1 0 3221 0 1 1336
box 0 0 19 49
use FILL  FILL_BUFX2_383
timestamp 1516325494
transform -1 0 3229 0 1 1336
box 0 0 8 49
use BUFX2  BUFX2_383
timestamp 1516325494
transform -1 0 3243 0 1 1336
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_286
timestamp 1516325494
transform -1 0 3296 0 1 1336
box 0 0 53 49
use MUX2X1  MUX2X1_210
timestamp 1516325494
transform -1 0 3327 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_254
timestamp 1516325494
transform -1 0 3380 0 1 1336
box 0 0 53 49
use AND2X2  AND2X2_1700
timestamp 1516325494
transform 1 0 3380 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1526
timestamp 1516325494
transform 1 0 3399 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1698
timestamp 1516325494
transform 1 0 3418 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1527
timestamp 1516325494
transform 1 0 3437 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1525
timestamp 1516325494
transform -1 0 3475 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_1740
timestamp 1516325494
transform 1 0 3475 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1697
timestamp 1516325494
transform -1 0 3513 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_297
timestamp 1516325494
transform -1 0 3532 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_294
timestamp 1516325494
transform -1 0 3551 0 1 1336
box 0 0 19 49
use NAND2X1  NAND2X1_242
timestamp 1516325494
transform 1 0 3551 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_242
timestamp 1516325494
transform -1 0 3596 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_178
timestamp 1516325494
transform -1 0 3650 0 1 1336
box 0 0 53 49
use AND2X2  AND2X2_311
timestamp 1516325494
transform 1 0 3650 0 1 1336
box 0 0 19 49
use OR2X2  OR2X2_292
timestamp 1516325494
transform -1 0 3688 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_310
timestamp 1516325494
transform -1 0 3707 0 1 1336
box 0 0 19 49
use NAND2X1  NAND2X1_633
timestamp 1516325494
transform 1 0 3707 0 1 1336
box 0 0 15 49
use MUX2X1  MUX2X1_633
timestamp 1516325494
transform -1 0 3752 0 1 1336
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_217
timestamp 1516325494
transform -1 0 3806 0 1 1336
box 0 0 53 49
use OR2X2  OR2X2_1739
timestamp 1516325494
transform -1 0 3825 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1862
timestamp 1516325494
transform -1 0 3844 0 1 1336
box 0 0 19 49
use AND2X2  AND2X2_1863
timestamp 1516325494
transform -1 0 3863 0 1 1336
box 0 0 19 49
use FILL  FILL_28_1
timestamp 1516325494
transform 1 0 3863 0 1 1336
box 0 0 8 49
use OR2X2  OR2X2_646
timestamp 1516325494
transform -1 0 21 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_689
timestamp 1516325494
transform -1 0 40 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_580
timestamp 1516325494
transform 1 0 40 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_681
timestamp 1516325494
transform -1 0 78 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_802
timestamp 1516325494
transform -1 0 97 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_678
timestamp 1516325494
transform -1 0 116 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_610
timestamp 1516325494
transform -1 0 135 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_725
timestamp 1516325494
transform -1 0 154 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_693
timestamp 1516325494
transform 1 0 154 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_581
timestamp 1516325494
transform -1 0 192 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_767
timestamp 1516325494
transform -1 0 211 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_694
timestamp 1516325494
transform 1 0 211 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_676
timestamp 1516325494
transform -1 0 249 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_685
timestamp 1516325494
transform -1 0 268 0 -1 1335
box 0 0 19 49
use OAI21X1  OAI21X1_13
timestamp 1516325494
transform -1 0 287 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_841
timestamp 1516325494
transform -1 0 295 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_841
timestamp 1516325494
transform -1 0 310 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_80
timestamp 1516325494
transform -1 0 318 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_80
timestamp 1516325494
transform -1 0 332 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_651
timestamp 1516325494
transform 1 0 333 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_780
timestamp 1516325494
transform 1 0 352 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_651
timestamp 1516325494
transform -1 0 386 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_567
timestamp 1516325494
transform -1 0 405 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_494
timestamp 1516325494
transform -1 0 424 0 -1 1335
box 0 0 19 49
use NOR2X1  NOR2X1_22
timestamp 1516325494
transform 1 0 424 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_695
timestamp 1516325494
transform -1 0 458 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_761
timestamp 1516325494
transform -1 0 477 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_786
timestamp 1516325494
transform -1 0 496 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_697
timestamp 1516325494
transform -1 0 511 0 -1 1335
box 0 0 15 49
use NOR2X1  NOR2X1_34
timestamp 1516325494
transform -1 0 526 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_825
timestamp 1516325494
transform -1 0 545 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_842
timestamp 1516325494
transform 1 0 545 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_842
timestamp 1516325494
transform 1 0 553 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_761
timestamp 1516325494
transform 1 0 568 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_910
timestamp 1516325494
transform 1 0 587 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_82
timestamp 1516325494
transform -1 0 614 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_82
timestamp 1516325494
transform -1 0 629 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_493
timestamp 1516325494
transform -1 0 648 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_794
timestamp 1516325494
transform 1 0 648 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_787
timestamp 1516325494
transform 1 0 667 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_859
timestamp 1516325494
transform -1 0 705 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_668
timestamp 1516325494
transform 1 0 705 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_707
timestamp 1516325494
transform -1 0 743 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_955
timestamp 1516325494
transform 1 0 743 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_669
timestamp 1516325494
transform 1 0 762 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_795
timestamp 1516325494
transform 1 0 781 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_956
timestamp 1516325494
transform 1 0 800 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_512
timestamp 1516325494
transform -1 0 838 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_511
timestamp 1516325494
transform 1 0 838 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_647
timestamp 1516325494
transform -1 0 872 0 -1 1335
box 0 0 15 49
use NAND3X1  NAND3X1_17
timestamp 1516325494
transform -1 0 891 0 -1 1335
box 0 0 19 49
use XOR2X1  XOR2X1_32
timestamp 1516325494
transform -1 0 925 0 -1 1335
box 0 0 34 49
use OR2X2  OR2X2_513
timestamp 1516325494
transform -1 0 944 0 -1 1335
box 0 0 19 49
use NOR2X1  NOR2X1_23
timestamp 1516325494
transform -1 0 959 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_746
timestamp 1516325494
transform -1 0 990 0 -1 1335
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_735
timestamp 1516325494
transform -1 0 1043 0 -1 1335
box 0 0 53 49
use INVX1  INVX1_143
timestamp 1516325494
transform 1 0 1043 0 -1 1335
box 0 0 11 49
use FILL  FILL_BUFX2_212
timestamp 1516325494
transform 1 0 1055 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_212
timestamp 1516325494
transform 1 0 1062 0 -1 1335
box 0 0 15 49
use INVX1  INVX1_219
timestamp 1516325494
transform -1 0 1088 0 -1 1335
box 0 0 11 49
use AND2X2  AND2X2_1872
timestamp 1516325494
transform -1 0 1108 0 -1 1335
box 0 0 19 49
use FILL  FILL_AND2X2_154
timestamp 1516325494
transform -1 0 1116 0 -1 1335
box 0 0 8 49
use AND2X2  AND2X2_154
timestamp 1516325494
transform -1 0 1134 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1617
timestamp 1516325494
transform 1 0 1134 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1031
timestamp 1516325494
transform -1 0 1172 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1030
timestamp 1516325494
transform -1 0 1191 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1312
timestamp 1516325494
transform -1 0 1210 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_2066
timestamp 1516325494
transform 1 0 1210 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_395
timestamp 1516325494
transform -1 0 1248 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1987
timestamp 1516325494
transform 1 0 1248 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1900
timestamp 1516325494
transform 1 0 1267 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1756
timestamp 1516325494
transform -1 0 1305 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1599
timestamp 1516325494
transform -1 0 1324 0 -1 1335
box 0 0 19 49
use FILL  FILL_AND2X2_246
timestamp 1516325494
transform -1 0 1332 0 -1 1335
box 0 0 8 49
use AND2X2  AND2X2_246
timestamp 1516325494
transform -1 0 1351 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1759
timestamp 1516325494
transform 1 0 1351 0 -1 1335
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_308
timestamp 1516325494
transform 1 0 1370 0 -1 1335
box 0 0 53 49
use NAND2X1  NAND2X1_500
timestamp 1516325494
transform 1 0 1423 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_500
timestamp 1516325494
transform -1 0 1468 0 -1 1335
box 0 0 30 49
use OR2X2  OR2X2_1913
timestamp 1516325494
transform -1 0 1488 0 -1 1335
box 0 0 19 49
use MUX2X1  MUX2X1_436
timestamp 1516325494
transform -1 0 1518 0 -1 1335
box 0 0 30 49
use NAND2X1  NAND2X1_404
timestamp 1516325494
transform -1 0 1533 0 -1 1335
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_436
timestamp 1516325494
transform 1 0 1533 0 -1 1335
box 0 0 53 49
use MUX2X1  MUX2X1_404
timestamp 1516325494
transform -1 0 1617 0 -1 1335
box 0 0 30 49
use OR2X2  OR2X2_373
timestamp 1516325494
transform -1 0 1636 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_371
timestamp 1516325494
transform -1 0 1655 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_396
timestamp 1516325494
transform -1 0 1674 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_397
timestamp 1516325494
transform -1 0 1693 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1912
timestamp 1516325494
transform -1 0 1712 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1911
timestamp 1516325494
transform -1 0 1731 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1993
timestamp 1516325494
transform -1 0 1750 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_372
timestamp 1516325494
transform -1 0 1769 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_398
timestamp 1516325494
transform -1 0 1788 0 -1 1335
box 0 0 19 49
use OAI21X1  OAI21X1_42
timestamp 1516325494
transform 1 0 1788 0 -1 1335
box 0 0 19 49
use INVX2  INVX2_31
timestamp 1516325494
transform 1 0 1807 0 -1 1335
box 0 0 11 49
use AND2X2  AND2X2_399
timestamp 1516325494
transform 1 0 1818 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1995
timestamp 1516325494
transform 1 0 1837 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1990
timestamp 1516325494
transform 1 0 1856 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1574
timestamp 1516325494
transform -1 0 1894 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1904
timestamp 1516325494
transform -1 0 1913 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1363
timestamp 1516325494
transform -1 0 1932 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_218
timestamp 1516325494
transform 1 0 1932 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_218
timestamp 1516325494
transform 1 0 1940 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_736
timestamp 1516325494
transform 1 0 1955 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_736
timestamp 1516325494
transform 1 0 1963 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_1028
timestamp 1516325494
transform -1 0 1997 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_449
timestamp 1516325494
transform -1 0 2005 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_449
timestamp 1516325494
transform -1 0 2020 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_472
timestamp 1516325494
transform -1 0 2028 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_472
timestamp 1516325494
transform -1 0 2042 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_531
timestamp 1516325494
transform -1 0 2051 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_531
timestamp 1516325494
transform -1 0 2065 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_715
timestamp 1516325494
transform 1 0 2065 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_715
timestamp 1516325494
transform 1 0 2073 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_714
timestamp 1516325494
transform -1 0 2096 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_714
timestamp 1516325494
transform -1 0 2111 0 -1 1335
box 0 0 15 49
use NAND2X1  NAND2X1_172
timestamp 1516325494
transform 1 0 2111 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_1311
timestamp 1516325494
transform -1 0 2145 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1026
timestamp 1516325494
transform -1 0 2164 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1027
timestamp 1516325494
transform -1 0 2183 0 -1 1335
box 0 0 19 49
use MUX2X1  MUX2X1_556
timestamp 1516325494
transform 1 0 2183 0 -1 1335
box 0 0 30 49
use NAND2X1  NAND2X1_556
timestamp 1516325494
transform -1 0 2229 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_1369
timestamp 1516325494
transform -1 0 2248 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_2040
timestamp 1516325494
transform -1 0 2267 0 -1 1335
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_492
timestamp 1516325494
transform -1 0 2320 0 -1 1335
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_33
timestamp 1516325494
transform 1 0 2320 0 -1 1335
box 0 0 53 49
use NAND2X1  NAND2X1_417
timestamp 1516325494
transform 1 0 2373 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_417
timestamp 1516325494
transform -1 0 2418 0 -1 1335
box 0 0 30 49
use AND2X2  AND2X2_1992
timestamp 1516325494
transform -1 0 2438 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1907
timestamp 1516325494
transform -1 0 2457 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1039
timestamp 1516325494
transform 1 0 2457 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_65
timestamp 1516325494
transform -1 0 2491 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_65
timestamp 1516325494
transform -1 0 2521 0 -1 1335
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_542
timestamp 1516325494
transform 1 0 2521 0 -1 1335
box 0 0 53 49
use NAND2X1  NAND2X1_542
timestamp 1516325494
transform 1 0 2575 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_542
timestamp 1516325494
transform -1 0 2620 0 -1 1335
box 0 0 30 49
use OAI21X1  OAI21X1_23
timestamp 1516325494
transform 1 0 2620 0 -1 1335
box 0 0 19 49
use OAI21X1  OAI21X1_19
timestamp 1516325494
transform 1 0 2639 0 -1 1335
box 0 0 19 49
use INVX2  INVX2_8
timestamp 1516325494
transform 1 0 2658 0 -1 1335
box 0 0 11 49
use FILL  FILL_BUFX2_528
timestamp 1516325494
transform -1 0 2678 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_528
timestamp 1516325494
transform -1 0 2692 0 -1 1335
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_382
timestamp 1516325494
transform 1 0 2692 0 -1 1335
box 0 0 53 49
use FILL  FILL_BUFX2_712
timestamp 1516325494
transform 1 0 2746 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_712
timestamp 1516325494
transform 1 0 2753 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_713
timestamp 1516325494
transform -1 0 2776 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_713
timestamp 1516325494
transform -1 0 2791 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_170
timestamp 1516325494
transform -1 0 2799 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_170
timestamp 1516325494
transform -1 0 2814 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_1977
timestamp 1516325494
transform -1 0 2833 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1976
timestamp 1516325494
transform -1 0 2852 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1975
timestamp 1516325494
transform -1 0 2871 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_772
timestamp 1516325494
transform 1 0 2871 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_772
timestamp 1516325494
transform 1 0 2879 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_2047
timestamp 1516325494
transform -1 0 2913 0 -1 1335
box 0 0 19 49
use MUX2X1  MUX2X1_609
timestamp 1516325494
transform 1 0 2913 0 -1 1335
box 0 0 30 49
use NAND2X1  NAND2X1_609
timestamp 1516325494
transform 1 0 2943 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_1296
timestamp 1516325494
transform -1 0 2977 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_2053
timestamp 1516325494
transform -1 0 2996 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_386
timestamp 1516325494
transform 1 0 2996 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_577
timestamp 1516325494
transform 1 0 3015 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_577
timestamp 1516325494
transform -1 0 3061 0 -1 1335
box 0 0 30 49
use MUX2X1  MUX2X1_606
timestamp 1516325494
transform 1 0 3061 0 -1 1335
box 0 0 30 49
use NAND2X1  NAND2X1_606
timestamp 1516325494
transform -1 0 3106 0 -1 1335
box 0 0 15 49
use OR2X2  OR2X2_363
timestamp 1516325494
transform -1 0 3126 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_388
timestamp 1516325494
transform -1 0 3145 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_838
timestamp 1516325494
transform -1 0 3153 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_838
timestamp 1516325494
transform -1 0 3167 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_387
timestamp 1516325494
transform -1 0 3186 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1975
timestamp 1516325494
transform -1 0 3205 0 -1 1335
box 0 0 19 49
use MUX2X1  MUX2X1_601
timestamp 1516325494
transform 1 0 3205 0 -1 1335
box 0 0 30 49
use AND2X2  AND2X2_1699
timestamp 1516325494
transform 1 0 3236 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_210
timestamp 1516325494
transform 1 0 3255 0 -1 1335
box 0 0 15 49
use NAND2X1  NAND2X1_222
timestamp 1516325494
transform 1 0 3270 0 -1 1335
box 0 0 15 49
use FILL  FILL_BUFX2_446
timestamp 1516325494
transform 1 0 3285 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_446
timestamp 1516325494
transform 1 0 3293 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_222
timestamp 1516325494
transform -1 0 3338 0 -1 1335
box 0 0 30 49
use NAND2X1  NAND2X1_601
timestamp 1516325494
transform -1 0 3353 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_1861
timestamp 1516325494
transform 1 0 3354 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1736
timestamp 1516325494
transform 1 0 3373 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1860
timestamp 1516325494
transform -1 0 3411 0 -1 1335
box 0 0 19 49
use NAND2X1  NAND2X1_217
timestamp 1516325494
transform 1 0 3411 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_217
timestamp 1516325494
transform -1 0 3456 0 -1 1335
box 0 0 30 49
use OR2X2  OR2X2_1737
timestamp 1516325494
transform 1 0 3456 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1735
timestamp 1516325494
transform -1 0 3494 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1858
timestamp 1516325494
transform -1 0 3513 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1859
timestamp 1516325494
transform -1 0 3532 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_532
timestamp 1516325494
transform -1 0 3540 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_532
timestamp 1516325494
transform -1 0 3555 0 -1 1335
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_185
timestamp 1516325494
transform 1 0 3555 0 -1 1335
box 0 0 53 49
use NAND2X1  NAND2X1_249
timestamp 1516325494
transform 1 0 3608 0 -1 1335
box 0 0 15 49
use MUX2X1  MUX2X1_249
timestamp 1516325494
transform -1 0 3653 0 -1 1335
box 0 0 30 49
use AND2X2  AND2X2_2023
timestamp 1516325494
transform -1 0 3673 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_159
timestamp 1516325494
transform -1 0 3681 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_159
timestamp 1516325494
transform -1 0 3695 0 -1 1335
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_352
timestamp 1516325494
transform 1 0 3696 0 -1 1335
box 0 0 53 49
use AND2X2  AND2X2_1333
timestamp 1516325494
transform 1 0 3749 0 -1 1335
box 0 0 19 49
use FILL  FILL_BUFX2_484
timestamp 1516325494
transform 1 0 3768 0 -1 1335
box 0 0 8 49
use BUFX2  BUFX2_484
timestamp 1516325494
transform 1 0 3775 0 -1 1335
box 0 0 15 49
use AND2X2  AND2X2_2082
timestamp 1516325494
transform 1 0 3791 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_1864
timestamp 1516325494
transform 1 0 3810 0 -1 1335
box 0 0 19 49
use OR2X2  OR2X2_1738
timestamp 1516325494
transform -1 0 3848 0 -1 1335
box 0 0 19 49
use OAI21X1  OAI21X1_115
timestamp 1516325494
transform 1 0 3848 0 -1 1335
box 0 0 19 49
use AND2X2  AND2X2_836
timestamp 1516325494
transform -1 0 21 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_489
timestamp 1516325494
transform -1 0 40 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_688
timestamp 1516325494
transform -1 0 59 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_584
timestamp 1516325494
transform 1 0 59 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_920
timestamp 1516325494
transform 1 0 78 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_874
timestamp 1516325494
transform -1 0 116 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_838
timestamp 1516325494
transform 1 0 116 0 1 1237
box 0 0 19 49
use FILL  FILL_BUFX2_358
timestamp 1516325494
transform 1 0 135 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_358
timestamp 1516325494
transform 1 0 143 0 1 1237
box 0 0 15 49
use OAI21X1  OAI21X1_8
timestamp 1516325494
transform 1 0 158 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_677
timestamp 1516325494
transform 1 0 177 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_964
timestamp 1516325494
transform 1 0 196 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_785
timestamp 1516325494
transform -1 0 234 0 1 1237
box 0 0 19 49
use OAI21X1  OAI21X1_14
timestamp 1516325494
transform -1 0 253 0 1 1237
box 0 0 19 49
use NAND3X1  NAND3X1_27
timestamp 1516325494
transform 1 0 253 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_749
timestamp 1516325494
transform -1 0 291 0 1 1237
box 0 0 19 49
use NOR3X1  NOR3X1_4
timestamp 1516325494
transform 1 0 291 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_983
timestamp 1516325494
transform 1 0 310 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_814
timestamp 1516325494
transform -1 0 348 0 1 1237
box 0 0 19 49
use FILL  FILL_BUFX2_811
timestamp 1516325494
transform -1 0 356 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_811
timestamp 1516325494
transform -1 0 370 0 1 1237
box 0 0 15 49
use OAI21X1  OAI21X1_10
timestamp 1516325494
transform 1 0 371 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_691
timestamp 1516325494
transform 1 0 390 0 1 1237
box 0 0 19 49
use NAND3X1  NAND3X1_19
timestamp 1516325494
transform 1 0 409 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_513
timestamp 1516325494
transform -1 0 447 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_636
timestamp 1516325494
transform 1 0 447 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_568
timestamp 1516325494
transform -1 0 485 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_569
timestamp 1516325494
transform 1 0 485 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_549
timestamp 1516325494
transform -1 0 523 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_637
timestamp 1516325494
transform 1 0 523 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_778
timestamp 1516325494
transform -1 0 561 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_487
timestamp 1516325494
transform -1 0 580 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_754
timestamp 1516325494
transform 1 0 580 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_912
timestamp 1516325494
transform -1 0 618 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_913
timestamp 1516325494
transform 1 0 618 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_911
timestamp 1516325494
transform -1 0 656 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_595
timestamp 1516325494
transform -1 0 675 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_807
timestamp 1516325494
transform 1 0 675 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_972
timestamp 1516325494
transform -1 0 713 0 1 1237
box 0 0 19 49
use NAND3X1  NAND3X1_53
timestamp 1516325494
transform -1 0 732 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_789
timestamp 1516325494
transform 1 0 732 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_591
timestamp 1516325494
transform -1 0 770 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_722
timestamp 1516325494
transform -1 0 789 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_851
timestamp 1516325494
transform 1 0 789 0 1 1237
box 0 0 19 49
use FILL  FILL_BUFX2_355
timestamp 1516325494
transform 1 0 808 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_355
timestamp 1516325494
transform 1 0 815 0 1 1237
box 0 0 15 49
use OR2X2  OR2X2_793
timestamp 1516325494
transform -1 0 849 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1087
timestamp 1516325494
transform -1 0 868 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_879
timestamp 1516325494
transform -1 0 887 0 1 1237
box 0 0 19 49
use XOR2X1  XOR2X1_31
timestamp 1516325494
transform 1 0 887 0 1 1237
box 0 0 34 49
use AND2X2  AND2X2_1086
timestamp 1516325494
transform -1 0 941 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_877
timestamp 1516325494
transform -1 0 960 0 1 1237
box 0 0 19 49
use XOR2X1  XOR2X1_30
timestamp 1516325494
transform -1 0 994 0 1 1237
box 0 0 34 49
use XOR2X1  XOR2X1_29
timestamp 1516325494
transform 1 0 994 0 1 1237
box 0 0 34 49
use FILL  FILL_OR2X2_146
timestamp 1516325494
transform -1 0 1036 0 1 1237
box 0 0 8 49
use OR2X2  OR2X2_146
timestamp 1516325494
transform -1 0 1055 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_913
timestamp 1516325494
transform -1 0 1074 0 1 1237
box 0 0 19 49
use FILL  FILL_OR2X2_145
timestamp 1516325494
transform -1 0 1082 0 1 1237
box 0 0 8 49
use OR2X2  OR2X2_145
timestamp 1516325494
transform -1 0 1100 0 1 1237
box 0 0 19 49
use FILL  FILL_AND2X2_155
timestamp 1516325494
transform -1 0 1108 0 1 1237
box 0 0 8 49
use AND2X2  AND2X2_155
timestamp 1516325494
transform -1 0 1127 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1421
timestamp 1516325494
transform -1 0 1146 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1420
timestamp 1516325494
transform -1 0 1165 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1619
timestamp 1516325494
transform -1 0 1184 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1315
timestamp 1516325494
transform -1 0 1203 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2068
timestamp 1516325494
transform 1 0 1203 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1982
timestamp 1516325494
transform 1 0 1222 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1983
timestamp 1516325494
transform 1 0 1241 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_368
timestamp 1516325494
transform -1 0 1279 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_393
timestamp 1516325494
transform -1 0 1298 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1618
timestamp 1516325494
transform -1 0 1317 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1986
timestamp 1516325494
transform -1 0 1336 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1901
timestamp 1516325494
transform 1 0 1336 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1419
timestamp 1516325494
transform -1 0 1374 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1899
timestamp 1516325494
transform -1 0 1393 0 1 1237
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_302
timestamp 1516325494
transform 1 0 1393 0 1 1237
box 0 0 53 49
use NAND2X1  NAND2X1_494
timestamp 1516325494
transform 1 0 1446 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_494
timestamp 1516325494
transform -1 0 1491 0 1 1237
box 0 0 30 49
use NAND2X1  NAND2X1_436
timestamp 1516325494
transform 1 0 1492 0 1 1237
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_318
timestamp 1516325494
transform 1 0 1507 0 1 1237
box 0 0 53 49
use NAND2X1  NAND2X1_510
timestamp 1516325494
transform 1 0 1560 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_510
timestamp 1516325494
transform -1 0 1605 0 1 1237
box 0 0 30 49
use FILL  FILL_BUFX2_241
timestamp 1516325494
transform 1 0 1606 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_241
timestamp 1516325494
transform 1 0 1613 0 1 1237
box 0 0 15 49
use AND2X2  AND2X2_1991
timestamp 1516325494
transform 1 0 1628 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1989
timestamp 1516325494
transform 1 0 1647 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1906
timestamp 1516325494
transform 1 0 1666 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1973
timestamp 1516325494
transform 1 0 1685 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1972
timestamp 1516325494
transform -1 0 1723 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1971
timestamp 1516325494
transform -1 0 1742 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_429
timestamp 1516325494
transform 1 0 1742 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2041
timestamp 1516325494
transform -1 0 1780 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1982
timestamp 1516325494
transform -1 0 1799 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1893
timestamp 1516325494
transform -1 0 1818 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1314
timestamp 1516325494
transform -1 0 1837 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1029
timestamp 1516325494
transform -1 0 1856 0 1 1237
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_289
timestamp 1516325494
transform 1 0 1856 0 1 1237
box 0 0 53 49
use NAND2X1  NAND2X1_481
timestamp 1516325494
transform 1 0 1910 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_481
timestamp 1516325494
transform -1 0 1955 0 1 1237
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_574
timestamp 1516325494
transform 1 0 1955 0 1 1237
box 0 0 53 49
use NAND2X1  NAND2X1_478
timestamp 1516325494
transform 1 0 2008 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_478
timestamp 1516325494
transform -1 0 2054 0 1 1237
box 0 0 30 49
use OR2X2  OR2X2_1894
timestamp 1516325494
transform -1 0 2073 0 1 1237
box 0 0 19 49
use FILL  FILL_BUFX2_597
timestamp 1516325494
transform 1 0 2073 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_597
timestamp 1516325494
transform 1 0 2081 0 1 1237
box 0 0 15 49
use NAND2X1  NAND2X1_318
timestamp 1516325494
transform 1 0 2096 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_318
timestamp 1516325494
transform -1 0 2141 0 1 1237
box 0 0 30 49
use MUX2X1  MUX2X1_76
timestamp 1516325494
transform 1 0 2141 0 1 1237
box 0 0 30 49
use NAND2X1  NAND2X1_76
timestamp 1516325494
transform -1 0 2187 0 1 1237
box 0 0 15 49
use OR2X2  OR2X2_1370
timestamp 1516325494
transform 1 0 2187 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_1580
timestamp 1516325494
transform 1 0 2206 0 1 1237
box 0 0 19 49
use FILL  FILL_BUFX2_595
timestamp 1516325494
transform -1 0 2233 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_595
timestamp 1516325494
transform -1 0 2248 0 1 1237
box 0 0 15 49
use AND2X2  AND2X2_1308
timestamp 1516325494
transform -1 0 2267 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1023
timestamp 1516325494
transform -1 0 2286 0 1 1237
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_545
timestamp 1516325494
transform 1 0 2286 0 1 1237
box 0 0 53 49
use NAND2X1  NAND2X1_449
timestamp 1516325494
transform 1 0 2339 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_449
timestamp 1516325494
transform -1 0 2384 0 1 1237
box 0 0 30 49
use OR2X2  OR2X2_1024
timestamp 1516325494
transform -1 0 2404 0 1 1237
box 0 0 19 49
use NAND2X1  NAND2X1_289
timestamp 1516325494
transform 1 0 2404 0 1 1237
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_673
timestamp 1516325494
transform -1 0 2472 0 1 1237
box 0 0 53 49
use MUX2X1  MUX2X1_448
timestamp 1516325494
transform 1 0 2472 0 1 1237
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_64
timestamp 1516325494
transform 1 0 2502 0 1 1237
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_481
timestamp 1516325494
transform 1 0 2556 0 1 1237
box 0 0 53 49
use AND2X2  AND2X2_1988
timestamp 1516325494
transform -1 0 2628 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1903
timestamp 1516325494
transform -1 0 2647 0 1 1237
box 0 0 19 49
use INVX2  INVX2_12
timestamp 1516325494
transform 1 0 2647 0 1 1237
box 0 0 11 49
use OR2X2  OR2X2_1974
timestamp 1516325494
transform 1 0 2658 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1902
timestamp 1516325494
transform -1 0 2696 0 1 1237
box 0 0 19 49
use NAND2X1  NAND2X1_940
timestamp 1516325494
transform 1 0 2696 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_885
timestamp 1516325494
transform 1 0 2711 0 1 1237
box 0 0 30 49
use FILL  FILL_BUFX2_630
timestamp 1516325494
transform -1 0 2750 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_630
timestamp 1516325494
transform -1 0 2764 0 1 1237
box 0 0 15 49
use FILL  FILL_BUFX2_699
timestamp 1516325494
transform -1 0 2773 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_699
timestamp 1516325494
transform -1 0 2787 0 1 1237
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_288
timestamp 1516325494
transform 1 0 2787 0 1 1237
box 0 0 53 49
use MUX2X1  MUX2X1_608
timestamp 1516325494
transform 1 0 2841 0 1 1237
box 0 0 30 49
use NAND2X1  NAND2X1_608
timestamp 1516325494
transform -1 0 2886 0 1 1237
box 0 0 15 49
use OR2X2  OR2X2_1016
timestamp 1516325494
transform 1 0 2886 0 1 1237
box 0 0 19 49
use MUX2X1  MUX2X1_638
timestamp 1516325494
transform 1 0 2905 0 1 1237
box 0 0 30 49
use NAND2X1  NAND2X1_638
timestamp 1516325494
transform -1 0 2951 0 1 1237
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_222
timestamp 1516325494
transform -1 0 3004 0 1 1237
box 0 0 53 49
use MUX2X1  MUX2X1_578
timestamp 1516325494
transform -1 0 3034 0 1 1237
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_258
timestamp 1516325494
transform -1 0 3087 0 1 1237
box 0 0 53 49
use FILL  FILL_BUFX2_599
timestamp 1516325494
transform 1 0 3088 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_599
timestamp 1516325494
transform 1 0 3095 0 1 1237
box 0 0 15 49
use FILL  FILL_BUFX2_109
timestamp 1516325494
transform -1 0 3118 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_109
timestamp 1516325494
transform -1 0 3133 0 1 1237
box 0 0 15 49
use OAI21X1  OAI21X1_57
timestamp 1516325494
transform -1 0 3152 0 1 1237
box 0 0 19 49
use FILL  FILL_BUFX2_527
timestamp 1516325494
transform -1 0 3160 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_527
timestamp 1516325494
transform -1 0 3175 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_628
timestamp 1516325494
transform 1 0 3175 0 1 1237
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_212
timestamp 1516325494
transform -1 0 3258 0 1 1237
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_281
timestamp 1516325494
transform -1 0 3312 0 1 1237
box 0 0 53 49
use AND2X2  AND2X2_313
timestamp 1516325494
transform 1 0 3312 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2022
timestamp 1516325494
transform 1 0 3331 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_293
timestamp 1516325494
transform 1 0 3350 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_312
timestamp 1516325494
transform -1 0 3388 0 1 1237
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_249
timestamp 1516325494
transform 1 0 3388 0 1 1237
box 0 0 53 49
use OR2X2  OR2X2_1946
timestamp 1516325494
transform 1 0 3441 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1950
timestamp 1516325494
transform -1 0 3479 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1947
timestamp 1516325494
transform -1 0 3498 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1945
timestamp 1516325494
transform -1 0 3517 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2019
timestamp 1516325494
transform 1 0 3517 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_419
timestamp 1516325494
transform 1 0 3536 0 1 1237
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_192
timestamp 1516325494
transform 1 0 3555 0 1 1237
box 0 0 53 49
use OR2X2  OR2X2_1949
timestamp 1516325494
transform -1 0 3627 0 1 1237
box 0 0 19 49
use OR2X2  OR2X2_1948
timestamp 1516325494
transform -1 0 3646 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2025
timestamp 1516325494
transform -1 0 3665 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2024
timestamp 1516325494
transform -1 0 3684 0 1 1237
box 0 0 19 49
use MUX2X1  MUX2X1_384
timestamp 1516325494
transform 1 0 3684 0 1 1237
box 0 0 30 49
use NAND2X1  NAND2X1_288
timestamp 1516325494
transform 1 0 3715 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_288
timestamp 1516325494
transform -1 0 3760 0 1 1237
box 0 0 30 49
use FILL  FILL_BUFX2_281
timestamp 1516325494
transform -1 0 3768 0 1 1237
box 0 0 8 49
use BUFX2  BUFX2_281
timestamp 1516325494
transform -1 0 3783 0 1 1237
box 0 0 15 49
use AND2X2  AND2X2_1335
timestamp 1516325494
transform 1 0 3783 0 1 1237
box 0 0 19 49
use AND2X2  AND2X2_2084
timestamp 1516325494
transform 1 0 3802 0 1 1237
box 0 0 19 49
use NAND2X1  NAND2X1_354
timestamp 1516325494
transform 1 0 3821 0 1 1237
box 0 0 15 49
use MUX2X1  MUX2X1_354
timestamp 1516325494
transform -1 0 3866 0 1 1237
box 0 0 30 49
use OR2X2  OR2X2_647
timestamp 1516325494
transform 1 0 2 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_835
timestamp 1516325494
transform -1 0 40 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_704
timestamp 1516325494
transform -1 0 59 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_452
timestamp 1516325494
transform 1 0 59 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_453
timestamp 1516325494
transform 1 0 78 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_623
timestamp 1516325494
transform -1 0 116 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_958
timestamp 1516325494
transform 1 0 116 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_801
timestamp 1516325494
transform 1 0 135 0 -1 1236
box 0 0 19 49
use FILL  FILL_BUFX2_809
timestamp 1516325494
transform 1 0 154 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_809
timestamp 1516325494
transform 1 0 162 0 -1 1236
box 0 0 15 49
use INVX1  INVX1_5
timestamp 1516325494
transform 1 0 177 0 -1 1236
box 0 0 11 49
use FILL  FILL_BUFX2_810
timestamp 1516325494
transform -1 0 196 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_810
timestamp 1516325494
transform -1 0 211 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_940
timestamp 1516325494
transform -1 0 230 0 -1 1236
box 0 0 19 49
use NOR3X1  NOR3X1_5
timestamp 1516325494
transform 1 0 230 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_895
timestamp 1516325494
transform -1 0 268 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_678
timestamp 1516325494
transform 1 0 268 0 -1 1236
box 0 0 15 49
use OAI21X1  OAI21X1_12
timestamp 1516325494
transform -1 0 302 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_771
timestamp 1516325494
transform 1 0 302 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_650
timestamp 1516325494
transform 1 0 321 0 -1 1236
box 0 0 19 49
use INVX1  INVX1_12
timestamp 1516325494
transform -1 0 351 0 -1 1236
box 0 0 11 49
use FILL  FILL_BUFX2_808
timestamp 1516325494
transform -1 0 360 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_808
timestamp 1516325494
transform -1 0 374 0 -1 1236
box 0 0 15 49
use INVX1  INVX1_34
timestamp 1516325494
transform -1 0 385 0 -1 1236
box 0 0 11 49
use AND2X2  AND2X2_781
timestamp 1516325494
transform 1 0 386 0 -1 1236
box 0 0 19 49
use FILL  FILL_BUFX2_361
timestamp 1516325494
transform 1 0 405 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_361
timestamp 1516325494
transform 1 0 412 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_514
timestamp 1516325494
transform 1 0 428 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_536
timestamp 1516325494
transform 1 0 447 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_425
timestamp 1516325494
transform -1 0 485 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_463
timestamp 1516325494
transform -1 0 504 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_635
timestamp 1516325494
transform -1 0 523 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_662
timestamp 1516325494
transform 1 0 523 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_820
timestamp 1516325494
transform 1 0 542 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_694
timestamp 1516325494
transform -1 0 580 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_661
timestamp 1516325494
transform -1 0 599 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1040
timestamp 1516325494
transform -1 0 618 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_743
timestamp 1516325494
transform -1 0 637 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_753
timestamp 1516325494
transform -1 0 656 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_863
timestamp 1516325494
transform -1 0 675 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_860
timestamp 1516325494
transform -1 0 694 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_742
timestamp 1516325494
transform -1 0 713 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_886
timestamp 1516325494
transform -1 0 732 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_689
timestamp 1516325494
transform -1 0 747 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_1043
timestamp 1516325494
transform -1 0 766 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1041
timestamp 1516325494
transform -1 0 785 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_863
timestamp 1516325494
transform 1 0 785 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_721
timestamp 1516325494
transform -1 0 823 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_861
timestamp 1516325494
transform -1 0 842 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_792
timestamp 1516325494
transform -1 0 861 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_878
timestamp 1516325494
transform -1 0 880 0 -1 1236
box 0 0 19 49
use INVX1  INVX1_58
timestamp 1516325494
transform -1 0 891 0 -1 1236
box 0 0 11 49
use INVX1  INVX1_57
timestamp 1516325494
transform 1 0 891 0 -1 1236
box 0 0 11 49
use OR2X2  OR2X2_876
timestamp 1516325494
transform 1 0 903 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_471
timestamp 1516325494
transform -1 0 941 0 -1 1236
box 0 0 19 49
use NOR2X1  NOR2X1_20
timestamp 1516325494
transform -1 0 956 0 -1 1236
box 0 0 15 49
use INVX1  INVX1_35
timestamp 1516325494
transform 1 0 956 0 -1 1236
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_747
timestamp 1516325494
transform -1 0 1020 0 -1 1236
box 0 0 53 49
use NAND2X1  NAND2X1_750
timestamp 1516325494
transform -1 0 1035 0 -1 1236
box 0 0 15 49
use NAND3X1  NAND3X1_61
timestamp 1516325494
transform -1 0 1055 0 -1 1236
box 0 0 19 49
use FILL  FILL_OR2X2_144
timestamp 1516325494
transform -1 0 1063 0 -1 1236
box 0 0 8 49
use OR2X2  OR2X2_144
timestamp 1516325494
transform -1 0 1081 0 -1 1236
box 0 0 19 49
use FILL  FILL_AND2X2_153
timestamp 1516325494
transform -1 0 1089 0 -1 1236
box 0 0 8 49
use AND2X2  AND2X2_153
timestamp 1516325494
transform -1 0 1108 0 -1 1236
box 0 0 19 49
use FILL  FILL_AND2X2_152
timestamp 1516325494
transform -1 0 1116 0 -1 1236
box 0 0 8 49
use AND2X2  AND2X2_152
timestamp 1516325494
transform -1 0 1134 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1415
timestamp 1516325494
transform -1 0 1153 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1615
timestamp 1516325494
transform -1 0 1172 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1025
timestamp 1516325494
transform -1 0 1191 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1309
timestamp 1516325494
transform -1 0 1210 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1981
timestamp 1516325494
transform 1 0 1210 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_2064
timestamp 1516325494
transform -1 0 1248 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1983
timestamp 1516325494
transform -1 0 1267 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1895
timestamp 1516325494
transform 1 0 1267 0 -1 1236
box 0 0 19 49
use FILL  FILL_BUFX2_118
timestamp 1516325494
transform -1 0 1294 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_118
timestamp 1516325494
transform -1 0 1309 0 -1 1236
box 0 0 15 49
use OR2X2  OR2X2_1898
timestamp 1516325494
transform 1 0 1309 0 -1 1236
box 0 0 19 49
use FILL  FILL_OR2X2_231
timestamp 1516325494
transform 1 0 1328 0 -1 1236
box 0 0 8 49
use OR2X2  OR2X2_231
timestamp 1516325494
transform 1 0 1336 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1606
timestamp 1516325494
transform -1 0 1374 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1761
timestamp 1516325494
transform -1 0 1393 0 -1 1236
box 0 0 19 49
use FILL  FILL_AND2X2_247
timestamp 1516325494
transform -1 0 1401 0 -1 1236
box 0 0 8 49
use AND2X2  AND2X2_247
timestamp 1516325494
transform -1 0 1419 0 -1 1236
box 0 0 19 49
use INVX1  INVX1_231
timestamp 1516325494
transform -1 0 1430 0 -1 1236
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_52
timestamp 1516325494
transform 1 0 1431 0 -1 1236
box 0 0 53 49
use OR2X2  OR2X2_1597
timestamp 1516325494
transform 1 0 1484 0 -1 1236
box 0 0 19 49
use FILL  FILL_BUFX2_200
timestamp 1516325494
transform 1 0 1503 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_200
timestamp 1516325494
transform 1 0 1511 0 -1 1236
box 0 0 15 49
use OR2X2  OR2X2_1592
timestamp 1516325494
transform 1 0 1526 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1614
timestamp 1516325494
transform -1 0 1564 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1413
timestamp 1516325494
transform -1 0 1583 0 -1 1236
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_558
timestamp 1516325494
transform 1 0 1583 0 -1 1236
box 0 0 53 49
use NAND2X1  NAND2X1_462
timestamp 1516325494
transform 1 0 1636 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_462
timestamp 1516325494
transform -1 0 1681 0 -1 1236
box 0 0 30 49
use FILL  FILL_AND2X2_129
timestamp 1516325494
transform -1 0 1690 0 -1 1236
box 0 0 8 49
use AND2X2  AND2X2_129
timestamp 1516325494
transform -1 0 1708 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1581
timestamp 1516325494
transform -1 0 1727 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_401
timestamp 1516325494
transform -1 0 1746 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_400
timestamp 1516325494
transform -1 0 1765 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_2039
timestamp 1516325494
transform -1 0 1784 0 -1 1236
box 0 0 19 49
use MUX2X1  MUX2X1_329
timestamp 1516325494
transform 1 0 1784 0 -1 1236
box 0 0 30 49
use NAND2X1  NAND2X1_329
timestamp 1516325494
transform -1 0 1830 0 -1 1236
box 0 0 15 49
use OR2X2  OR2X2_1275
timestamp 1516325494
transform -1 0 1849 0 -1 1236
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_457
timestamp 1516325494
transform 1 0 1849 0 -1 1236
box 0 0 53 49
use OAI21X1  OAI21X1_26
timestamp 1516325494
transform 1 0 1902 0 -1 1236
box 0 0 19 49
use FILL  FILL_BUFX2_632
timestamp 1516325494
transform -1 0 1929 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_632
timestamp 1516325494
transform -1 0 1944 0 -1 1236
box 0 0 15 49
use OR2X2  OR2X2_1604
timestamp 1516325494
transform 1 0 1944 0 -1 1236
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_468
timestamp 1516325494
transform 1 0 1963 0 -1 1236
box 0 0 53 49
use NAND2X1  NAND2X1_340
timestamp 1516325494
transform 1 0 2016 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_340
timestamp 1516325494
transform -1 0 2061 0 -1 1236
box 0 0 30 49
use FILL  FILL_BUFX2_125
timestamp 1516325494
transform -1 0 2070 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_125
timestamp 1516325494
transform -1 0 2084 0 -1 1236
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_702
timestamp 1516325494
transform 1 0 2084 0 -1 1236
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_108
timestamp 1516325494
transform -1 0 2191 0 -1 1236
box 0 0 53 49
use NAND2X1  NAND2X1_553
timestamp 1516325494
transform 1 0 2191 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_553
timestamp 1516325494
transform -1 0 2236 0 -1 1236
box 0 0 30 49
use FILL  FILL_BUFX2_388
timestamp 1516325494
transform 1 0 2236 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_388
timestamp 1516325494
transform 1 0 2244 0 -1 1236
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_532
timestamp 1516325494
transform 1 0 2259 0 -1 1236
box 0 0 53 49
use OR2X2  OR2X2_1607
timestamp 1516325494
transform -1 0 2331 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_532
timestamp 1516325494
transform 1 0 2331 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_532
timestamp 1516325494
transform -1 0 2377 0 -1 1236
box 0 0 30 49
use FILL  FILL_BUFX2_633
timestamp 1516325494
transform 1 0 2377 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_633
timestamp 1516325494
transform 1 0 2385 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_289
timestamp 1516325494
transform 1 0 2400 0 -1 1236
box 0 0 30 49
use OR2X2  OR2X2_1967
timestamp 1516325494
transform 1 0 2430 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_544
timestamp 1516325494
transform 1 0 2449 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_544
timestamp 1516325494
transform -1 0 2494 0 -1 1236
box 0 0 30 49
use NAND2X1  NAND2X1_448
timestamp 1516325494
transform -1 0 2510 0 -1 1236
box 0 0 15 49
use NAND2X1  NAND2X1_62
timestamp 1516325494
transform 1 0 2510 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_62
timestamp 1516325494
transform -1 0 2555 0 -1 1236
box 0 0 30 49
use NAND2X1  NAND2X1_545
timestamp 1516325494
transform 1 0 2556 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_545
timestamp 1516325494
transform -1 0 2601 0 -1 1236
box 0 0 30 49
use MUX2X1  MUX2X1_190
timestamp 1516325494
transform 1 0 2601 0 -1 1236
box 0 0 30 49
use NAND2X1  NAND2X1_190
timestamp 1516325494
transform -1 0 2647 0 -1 1236
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_414
timestamp 1516325494
transform -1 0 2700 0 -1 1236
box 0 0 53 49
use FILL  FILL_BUFX2_392
timestamp 1516325494
transform -1 0 2708 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_392
timestamp 1516325494
transform -1 0 2723 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_193
timestamp 1516325494
transform 1 0 2723 0 -1 1236
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_225
timestamp 1516325494
transform -1 0 2806 0 -1 1236
box 0 0 53 49
use NAND2X1  NAND2X1_193
timestamp 1516325494
transform -1 0 2821 0 -1 1236
box 0 0 15 49
use FILL  FILL_BUFX2_836
timestamp 1516325494
transform 1 0 2822 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_836
timestamp 1516325494
transform 1 0 2829 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_2050
timestamp 1516325494
transform -1 0 2863 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1050
timestamp 1516325494
transform -1 0 2882 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1293
timestamp 1516325494
transform -1 0 2901 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1047
timestamp 1516325494
transform -1 0 2920 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1046
timestamp 1516325494
transform -1 0 2939 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1331
timestamp 1516325494
transform -1 0 2958 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1332
timestamp 1516325494
transform -1 0 2977 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1045
timestamp 1516325494
transform -1 0 2996 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_578
timestamp 1516325494
transform 1 0 2996 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_1329
timestamp 1516325494
transform -1 0 3031 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_2081
timestamp 1516325494
transform 1 0 3031 0 -1 1236
box 0 0 19 49
use MUX2X1  MUX2X1_610
timestamp 1516325494
transform 1 0 3050 0 -1 1236
box 0 0 30 49
use NAND2X1  NAND2X1_610
timestamp 1516325494
transform -1 0 3095 0 -1 1236
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_194
timestamp 1516325494
transform -1 0 3148 0 -1 1236
box 0 0 53 49
use AND2X2  AND2X2_1330
timestamp 1516325494
transform -1 0 3167 0 -1 1236
box 0 0 19 49
use MUX2X1  MUX2X1_212
timestamp 1516325494
transform 1 0 3167 0 -1 1236
box 0 0 30 49
use NAND2X1  NAND2X1_628
timestamp 1516325494
transform -1 0 3213 0 -1 1236
box 0 0 15 49
use NAND2X1  NAND2X1_212
timestamp 1516325494
transform -1 0 3228 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_1745
timestamp 1516325494
transform 1 0 3228 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1586
timestamp 1516325494
transform 1 0 3247 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1587
timestamp 1516325494
transform 1 0 3266 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1746
timestamp 1516325494
transform -1 0 3304 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1585
timestamp 1516325494
transform -1 0 3323 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1744
timestamp 1516325494
transform -1 0 3342 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_747
timestamp 1516325494
transform -1 0 3357 0 -1 1236
box 0 0 15 49
use FILL  FILL_AND2X2_236
timestamp 1516325494
transform 1 0 3357 0 -1 1236
box 0 0 8 49
use AND2X2  AND2X2_236
timestamp 1516325494
transform 1 0 3365 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_1743
timestamp 1516325494
transform -1 0 3403 0 -1 1236
box 0 0 19 49
use FILL  FILL_AND2X2_235
timestamp 1516325494
transform 1 0 3403 0 -1 1236
box 0 0 8 49
use AND2X2  AND2X2_235
timestamp 1516325494
transform 1 0 3411 0 -1 1236
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_180
timestamp 1516325494
transform 1 0 3430 0 -1 1236
box 0 0 53 49
use NAND2X1  NAND2X1_244
timestamp 1516325494
transform 1 0 3483 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_244
timestamp 1516325494
transform -1 0 3528 0 -1 1236
box 0 0 30 49
use AND2X2  AND2X2_2020
timestamp 1516325494
transform 1 0 3528 0 -1 1236
box 0 0 19 49
use FILL  FILL_BUFX2_391
timestamp 1516325494
transform -1 0 3555 0 -1 1236
box 0 0 8 49
use BUFX2  BUFX2_391
timestamp 1516325494
transform -1 0 3570 0 -1 1236
box 0 0 15 49
use OR2X2  OR2X2_394
timestamp 1516325494
transform -1 0 3589 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_415
timestamp 1516325494
transform 1 0 3589 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_256
timestamp 1516325494
transform 1 0 3608 0 -1 1236
box 0 0 15 49
use MUX2X1  MUX2X1_256
timestamp 1516325494
transform -1 0 3653 0 -1 1236
box 0 0 30 49
use OR2X2  OR2X2_393
timestamp 1516325494
transform -1 0 3673 0 -1 1236
box 0 0 19 49
use AND2X2  AND2X2_421
timestamp 1516325494
transform -1 0 3692 0 -1 1236
box 0 0 19 49
use NAND2X1  NAND2X1_384
timestamp 1516325494
transform 1 0 3692 0 -1 1236
box 0 0 15 49
use AND2X2  AND2X2_420
timestamp 1516325494
transform -1 0 3726 0 -1 1236
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_160
timestamp 1516325494
transform 1 0 3726 0 -1 1236
box 0 0 53 49
use OR2X2  OR2X2_1049
timestamp 1516325494
transform -1 0 3798 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1993
timestamp 1516325494
transform -1 0 3817 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1992
timestamp 1516325494
transform -1 0 3836 0 -1 1236
box 0 0 19 49
use OR2X2  OR2X2_1048
timestamp 1516325494
transform -1 0 3855 0 -1 1236
box 0 0 19 49
use INVX1  INVX1_302
timestamp 1516325494
transform -1 0 3866 0 -1 1236
box 0 0 11 49
use AND2X2  AND2X2_769
timestamp 1516325494
transform -1 0 21 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_768
timestamp 1516325494
transform -1 0 40 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_644
timestamp 1516325494
transform -1 0 59 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_510
timestamp 1516325494
transform 1 0 59 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_528
timestamp 1516325494
transform 1 0 78 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_807
timestamp 1516325494
transform -1 0 116 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_624
timestamp 1516325494
transform 1 0 116 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_963
timestamp 1516325494
transform -1 0 154 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_622
timestamp 1516325494
transform -1 0 173 0 1 1138
box 0 0 19 49
use AOI21X1  AOI21X1_9
timestamp 1516325494
transform -1 0 192 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_724
timestamp 1516325494
transform -1 0 211 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_711
timestamp 1516325494
transform -1 0 230 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_838
timestamp 1516325494
transform -1 0 249 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_708
timestamp 1516325494
transform -1 0 268 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_721
timestamp 1516325494
transform 1 0 268 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_679
timestamp 1516325494
transform -1 0 306 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_456
timestamp 1516325494
transform 1 0 306 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_858
timestamp 1516325494
transform -1 0 344 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_857
timestamp 1516325494
transform -1 0 363 0 1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_35
timestamp 1516325494
transform -1 0 382 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_416
timestamp 1516325494
transform -1 0 401 0 1 1138
box 0 0 19 49
use INVX1  INVX1_24
timestamp 1516325494
transform 1 0 401 0 1 1138
box 0 0 11 49
use OR2X2  OR2X2_461
timestamp 1516325494
transform 1 0 412 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_535
timestamp 1516325494
transform 1 0 431 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_417
timestamp 1516325494
transform -1 0 469 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_456
timestamp 1516325494
transform 1 0 469 0 1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_357
timestamp 1516325494
transform 1 0 488 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_357
timestamp 1516325494
transform 1 0 496 0 1 1138
box 0 0 15 49
use NAND3X1  NAND3X1_38
timestamp 1516325494
transform 1 0 511 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_717
timestamp 1516325494
transform 1 0 530 0 1 1138
box 0 0 19 49
use AOI21X1  AOI21X1_12
timestamp 1516325494
transform -1 0 568 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_718
timestamp 1516325494
transform 1 0 568 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_486
timestamp 1516325494
transform -1 0 606 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_562
timestamp 1516325494
transform -1 0 625 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_881
timestamp 1516325494
transform -1 0 644 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_630
timestamp 1516325494
transform 1 0 644 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_755
timestamp 1516325494
transform 1 0 663 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_594
timestamp 1516325494
transform -1 0 701 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_502
timestamp 1516325494
transform -1 0 720 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_588
timestamp 1516325494
transform 1 0 720 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_718
timestamp 1516325494
transform 1 0 739 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_792
timestamp 1516325494
transform -1 0 777 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_758
timestamp 1516325494
transform -1 0 796 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_901
timestamp 1516325494
transform -1 0 815 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_856
timestamp 1516325494
transform -1 0 834 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_946
timestamp 1516325494
transform 1 0 834 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1042
timestamp 1516325494
transform 1 0 853 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_809
timestamp 1516325494
transform -1 0 891 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_951
timestamp 1516325494
transform -1 0 910 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1036
timestamp 1516325494
transform 1 0 910 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_860
timestamp 1516325494
transform -1 0 948 0 1 1138
box 0 0 19 49
use XNOR2X1  XNOR2X1_4
timestamp 1516325494
transform 1 0 948 0 1 1138
box 0 0 34 49
use XNOR2X1  XNOR2X1_3
timestamp 1516325494
transform 1 0 982 0 1 1138
box 0 0 34 49
use MUX2X1  MUX2X1_799
timestamp 1516325494
transform -1 0 1047 0 1 1138
box 0 0 30 49
use MUX2X1  MUX2X1_786
timestamp 1516325494
transform -1 0 1077 0 1 1138
box 0 0 30 49
use INVX1  INVX1_208
timestamp 1516325494
transform -1 0 1088 0 1 1138
box 0 0 11 49
use FILL  FILL_OR2X2_235
timestamp 1516325494
transform -1 0 1097 0 1 1138
box 0 0 8 49
use OR2X2  OR2X2_235
timestamp 1516325494
transform -1 0 1115 0 1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_245
timestamp 1516325494
transform -1 0 1123 0 1 1138
box 0 0 8 49
use AND2X2  AND2X2_245
timestamp 1516325494
transform -1 0 1142 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1613
timestamp 1516325494
transform -1 0 1161 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1757
timestamp 1516325494
transform 1 0 1161 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1306
timestamp 1516325494
transform -1 0 1199 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_2062
timestamp 1516325494
transform 1 0 1199 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1600
timestamp 1516325494
transform 1 0 1218 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1601
timestamp 1516325494
transform 1 0 1237 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_392
timestamp 1516325494
transform -1 0 1275 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1981
timestamp 1516325494
transform -1 0 1294 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1613
timestamp 1516325494
transform 1 0 1294 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1614
timestamp 1516325494
transform -1 0 1332 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1612
timestamp 1516325494
transform -1 0 1351 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1611
timestamp 1516325494
transform -1 0 1370 0 1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_334
timestamp 1516325494
transform 1 0 1370 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_334
timestamp 1516325494
transform 1 0 1378 0 1 1138
box 0 0 15 49
use AND2X2  AND2X2_1763
timestamp 1516325494
transform -1 0 1412 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1612
timestamp 1516325494
transform -1 0 1431 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1412
timestamp 1516325494
transform -1 0 1450 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_430
timestamp 1516325494
transform 1 0 1450 0 1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_398
timestamp 1516325494
transform 1 0 1503 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_398
timestamp 1516325494
transform -1 0 1548 0 1 1138
box 0 0 30 49
use OR2X2  OR2X2_402
timestamp 1516325494
transform 1 0 1549 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_403
timestamp 1516325494
transform -1 0 1587 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1411
timestamp 1516325494
transform -1 0 1606 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_590
timestamp 1516325494
transform 1 0 1606 0 1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_14
timestamp 1516325494
transform 1 0 1659 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_14
timestamp 1516325494
transform -1 0 1704 0 1 1138
box 0 0 30 49
use OR2X2  OR2X2_1414
timestamp 1516325494
transform -1 0 1723 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_686
timestamp 1516325494
transform 1 0 1723 0 1 1138
box 0 0 53 49
use AND2X2  AND2X2_428
timestamp 1516325494
transform -1 0 1796 0 1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_302
timestamp 1516325494
transform 1 0 1796 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_302
timestamp 1516325494
transform -1 0 1841 0 1 1138
box 0 0 30 49
use AND2X2  AND2X2_1305
timestamp 1516325494
transform -1 0 1860 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1022
timestamp 1516325494
transform -1 0 1879 0 1 1138
box 0 0 19 49
use OAI21X1  OAI21X1_39
timestamp 1516325494
transform 1 0 1879 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_417
timestamp 1516325494
transform 1 0 1898 0 1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_385
timestamp 1516325494
transform 1 0 1951 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_385
timestamp 1516325494
transform -1 0 1997 0 1 1138
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_596
timestamp 1516325494
transform 1 0 1997 0 1 1138
box 0 0 53 49
use MUX2X1  MUX2X1_20
timestamp 1516325494
transform -1 0 2080 0 1 1138
box 0 0 30 49
use AND2X2  AND2X2_1760
timestamp 1516325494
transform -1 0 2100 0 1 1138
box 0 0 19 49
use MUX2X1  MUX2X1_843
timestamp 1516325494
transform -1 0 2130 0 1 1138
box 0 0 30 49
use MUX2X1  MUX2X1_1
timestamp 1516325494
transform 1 0 2130 0 1 1138
box 0 0 30 49
use NAND2X1  NAND2X1_1
timestamp 1516325494
transform -1 0 2175 0 1 1138
box 0 0 15 49
use OR2X2  OR2X2_703
timestamp 1516325494
transform -1 0 21 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_298
timestamp 1516325494
transform -1 0 29 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_298
timestamp 1516325494
transform -1 0 44 0 -1 1138
box 0 0 15 49
use AND2X2  AND2X2_638
timestamp 1516325494
transform 1 0 44 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_537
timestamp 1516325494
transform 1 0 63 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_354
timestamp 1516325494
transform 1 0 82 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_354
timestamp 1516325494
transform 1 0 89 0 -1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_360
timestamp 1516325494
transform -1 0 113 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_360
timestamp 1516325494
transform -1 0 127 0 -1 1138
box 0 0 15 49
use OR2X2  OR2X2_538
timestamp 1516325494
transform 1 0 127 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_868
timestamp 1516325494
transform -1 0 165 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_640
timestamp 1516325494
transform 1 0 165 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_607
timestamp 1516325494
transform 1 0 184 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1047
timestamp 1516325494
transform 1 0 203 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_874
timestamp 1516325494
transform -1 0 241 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_873
timestamp 1516325494
transform -1 0 260 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_817
timestamp 1516325494
transform 1 0 260 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_818
timestamp 1516325494
transform 1 0 279 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_295
timestamp 1516325494
transform -1 0 306 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_295
timestamp 1516325494
transform -1 0 321 0 -1 1138
box 0 0 15 49
use XOR2X1  XOR2X1_7
timestamp 1516325494
transform -1 0 355 0 -1 1138
box 0 0 34 49
use AND2X2  AND2X2_447
timestamp 1516325494
transform 1 0 355 0 -1 1138
box 0 0 19 49
use XOR2X1  XOR2X1_5
timestamp 1516325494
transform 1 0 374 0 -1 1138
box 0 0 34 49
use OR2X2  OR2X2_633
timestamp 1516325494
transform 1 0 409 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_356
timestamp 1516325494
transform -1 0 436 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_356
timestamp 1516325494
transform -1 0 450 0 -1 1138
box 0 0 15 49
use AND2X2  AND2X2_782
timestamp 1516325494
transform 1 0 450 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_634
timestamp 1516325494
transform 1 0 469 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_759
timestamp 1516325494
transform 1 0 488 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_760
timestamp 1516325494
transform 1 0 507 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_663
timestamp 1516325494
transform -1 0 545 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_785
timestamp 1516325494
transform -1 0 564 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_784
timestamp 1516325494
transform -1 0 583 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_660
timestamp 1516325494
transform -1 0 602 0 -1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_58
timestamp 1516325494
transform 1 0 602 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_557
timestamp 1516325494
transform 1 0 621 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_825
timestamp 1516325494
transform -1 0 659 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_297
timestamp 1516325494
transform -1 0 667 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_297
timestamp 1516325494
transform -1 0 682 0 -1 1138
box 0 0 15 49
use OR2X2  OR2X2_776
timestamp 1516325494
transform 1 0 682 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_930
timestamp 1516325494
transform -1 0 720 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_293
timestamp 1516325494
transform -1 0 728 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_293
timestamp 1516325494
transform -1 0 743 0 -1 1138
box 0 0 15 49
use OR2X2  OR2X2_775
timestamp 1516325494
transform -1 0 762 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_797
timestamp 1516325494
transform -1 0 781 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_796
timestamp 1516325494
transform -1 0 800 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_757
timestamp 1516325494
transform -1 0 819 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_846
timestamp 1516325494
transform 1 0 819 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1016
timestamp 1516325494
transform -1 0 857 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_672
timestamp 1516325494
transform 1 0 857 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_832
timestamp 1516325494
transform 1 0 876 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_831
timestamp 1516325494
transform -1 0 914 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_359
timestamp 1516325494
transform 1 0 914 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_359
timestamp 1516325494
transform 1 0 922 0 -1 1138
box 0 0 15 49
use AND2X2  AND2X2_999
timestamp 1516325494
transform -1 0 956 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1035
timestamp 1516325494
transform -1 0 975 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_655
timestamp 1516325494
transform 1 0 975 0 -1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_734
timestamp 1516325494
transform -1 0 1047 0 -1 1138
box 0 0 53 49
use INVX1  INVX1_33
timestamp 1516325494
transform 1 0 1047 0 -1 1138
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_733
timestamp 1516325494
transform -1 0 1111 0 -1 1138
box 0 0 53 49
use FILL  FILL_OR2X2_234
timestamp 1516325494
transform -1 0 1120 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_234
timestamp 1516325494
transform -1 0 1138 0 -1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_230
timestamp 1516325494
transform -1 0 1146 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_230
timestamp 1516325494
transform -1 0 1165 0 -1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_229
timestamp 1516325494
transform -1 0 1173 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_229
timestamp 1516325494
transform -1 0 1191 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_244
timestamp 1516325494
transform -1 0 1199 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_244
timestamp 1516325494
transform -1 0 1218 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1755
timestamp 1516325494
transform -1 0 1237 0 -1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_228
timestamp 1516325494
transform -1 0 1245 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_228
timestamp 1516325494
transform -1 0 1264 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_242
timestamp 1516325494
transform -1 0 1272 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_242
timestamp 1516325494
transform -1 0 1290 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_243
timestamp 1516325494
transform -1 0 1298 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_243
timestamp 1516325494
transform -1 0 1317 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1751
timestamp 1516325494
transform 1 0 1317 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_1595
timestamp 1516325494
transform -1 0 1355 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1753
timestamp 1516325494
transform -1 0 1374 0 -1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_233
timestamp 1516325494
transform -1 0 1382 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_233
timestamp 1516325494
transform -1 0 1400 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1506
timestamp 1516325494
transform -1 0 1419 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1888
timestamp 1516325494
transform -1 0 1438 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_1772
timestamp 1516325494
transform -1 0 1457 0 -1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_232
timestamp 1516325494
transform -1 0 1465 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_232
timestamp 1516325494
transform -1 0 1484 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_248
timestamp 1516325494
transform -1 0 1492 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_248
timestamp 1516325494
transform -1 0 1511 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1754
timestamp 1516325494
transform 1 0 1511 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1750
timestamp 1516325494
transform -1 0 1549 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1980
timestamp 1516325494
transform -1 0 1568 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_1892
timestamp 1516325494
transform -1 0 1587 0 -1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_446
timestamp 1516325494
transform 1 0 1587 0 -1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_414
timestamp 1516325494
transform 1 0 1640 0 -1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_414
timestamp 1516325494
transform -1 0 1685 0 -1 1138
box 0 0 30 49
use OR2X2  OR2X2_1891
timestamp 1516325494
transform -1 0 1704 0 -1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_30
timestamp 1516325494
transform 1 0 1704 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_606
timestamp 1516325494
transform 1 0 1720 0 -1 1138
box 0 0 53 49
use MUX2X1  MUX2X1_30
timestamp 1516325494
transform -1 0 1803 0 -1 1138
box 0 0 30 49
use AND2X2  AND2X2_1507
timestamp 1516325494
transform -1 0 1822 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_1274
timestamp 1516325494
transform -1 0 1841 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_27
timestamp 1516325494
transform -1 0 1849 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_27
timestamp 1516325494
transform -1 0 1864 0 -1 1138
box 0 0 15 49
use OR2X2  OR2X2_1591
timestamp 1516325494
transform -1 0 1883 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1752
timestamp 1516325494
transform -1 0 1902 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_1593
timestamp 1516325494
transform -1 0 1921 0 -1 1138
box 0 0 19 49
use OR2X2  OR2X2_1594
timestamp 1516325494
transform -1 0 1940 0 -1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_308
timestamp 1516325494
transform 1 0 1940 0 -1 1138
box 0 0 15 49
use NAND2X1  NAND2X1_20
timestamp 1516325494
transform 1 0 1955 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_692
timestamp 1516325494
transform 1 0 1970 0 -1 1138
box 0 0 53 49
use MUX2X1  MUX2X1_308
timestamp 1516325494
transform -1 0 2054 0 -1 1138
box 0 0 30 49
use INVX1  INVX1_136
timestamp 1516325494
transform -1 0 2065 0 -1 1138
box 0 0 11 49
use OR2X2  OR2X2_1596
timestamp 1516325494
transform -1 0 2084 0 -1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_898
timestamp 1516325494
transform 1 0 2084 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_628
timestamp 1516325494
transform 1 0 2100 0 -1 1138
box 0 0 53 49
use FILL  FILL_BUFX2_813
timestamp 1516325494
transform -1 0 2161 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_813
timestamp 1516325494
transform -1 0 2175 0 -1 1138
box 0 0 15 49
use OR2X2  OR2X2_1021
timestamp 1516325494
transform -1 0 2195 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_577
timestamp 1516325494
transform -1 0 2248 0 1 1138
box 0 0 53 49
use MUX2X1  MUX2X1_468
timestamp 1516325494
transform -1 0 2278 0 1 1138
box 0 0 30 49
use INVX2  INVX2_15
timestamp 1516325494
transform 1 0 2278 0 1 1138
box 0 0 11 49
use OR2X2  OR2X2_1605
timestamp 1516325494
transform -1 0 2309 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_1762
timestamp 1516325494
transform -1 0 2328 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_489
timestamp 1516325494
transform -1 0 2381 0 1 1138
box 0 0 53 49
use FILL  FILL_BUFX2_208
timestamp 1516325494
transform 1 0 2381 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_208
timestamp 1516325494
transform 1 0 2388 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_765
timestamp 1516325494
transform 1 0 2404 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_765
timestamp 1516325494
transform 1 0 2411 0 1 1138
box 0 0 15 49
use OR2X2  OR2X2_1608
timestamp 1516325494
transform -1 0 2445 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_2038
timestamp 1516325494
transform -1 0 2464 0 1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_116
timestamp 1516325494
transform 1 0 2464 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_116
timestamp 1516325494
transform -1 0 2510 0 1 1138
box 0 0 30 49
use OR2X2  OR2X2_1968
timestamp 1516325494
transform -1 0 2529 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_544
timestamp 1516325494
transform -1 0 2582 0 1 1138
box 0 0 53 49
use FILL  FILL_BUFX2_182
timestamp 1516325494
transform 1 0 2582 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_182
timestamp 1516325494
transform 1 0 2590 0 1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_670
timestamp 1516325494
transform -1 0 2658 0 1 1138
box 0 0 53 49
use NOR2X1  NOR2X1_14
timestamp 1516325494
transform -1 0 2673 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_10
timestamp 1516325494
transform -1 0 2688 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_1
timestamp 1516325494
transform -1 0 2704 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_8
timestamp 1516325494
transform -1 0 2719 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_12
timestamp 1516325494
transform -1 0 2734 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_11
timestamp 1516325494
transform -1 0 2749 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_174
timestamp 1516325494
transform -1 0 2764 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_596
timestamp 1516325494
transform 1 0 2765 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_596
timestamp 1516325494
transform 1 0 2772 0 1 1138
box 0 0 15 49
use INVX1  INVX1_1
timestamp 1516325494
transform 1 0 2787 0 1 1138
box 0 0 11 49
use NAND3X1  NAND3X1_9
timestamp 1516325494
transform 1 0 2799 0 1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_102
timestamp 1516325494
transform 1 0 2818 0 1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_1
timestamp 1516325494
transform 1 0 2837 0 1 1138
box 0 0 19 49
use NOR2X1  NOR2X1_17
timestamp 1516325494
transform 1 0 2856 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_248
timestamp 1516325494
transform -1 0 2879 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_248
timestamp 1516325494
transform -1 0 2894 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_5
timestamp 1516325494
transform 1 0 2894 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_6
timestamp 1516325494
transform 1 0 2909 0 1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_7
timestamp 1516325494
transform 1 0 2924 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_771
timestamp 1516325494
transform -1 0 2947 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_771
timestamp 1516325494
transform -1 0 2962 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_194
timestamp 1516325494
transform 1 0 2962 0 1 1138
box 0 0 30 49
use NAND2X1  NAND2X1_194
timestamp 1516325494
transform -1 0 3008 0 1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_226
timestamp 1516325494
transform -1 0 3061 0 1 1138
box 0 0 53 49
use AND2X2  AND2X2_2080
timestamp 1516325494
transform 1 0 3061 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1990
timestamp 1516325494
transform 1 0 3080 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1994
timestamp 1516325494
transform -1 0 3118 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1991
timestamp 1516325494
transform -1 0 3137 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_1989
timestamp 1516325494
transform -1 0 3156 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_2079
timestamp 1516325494
transform -1 0 3175 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_2078
timestamp 1516325494
transform -1 0 3194 0 1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_705
timestamp 1516325494
transform -1 0 3202 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_705
timestamp 1516325494
transform -1 0 3217 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_394
timestamp 1516325494
transform -1 0 3225 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_394
timestamp 1516325494
transform -1 0 3239 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_619
timestamp 1516325494
transform 1 0 3240 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_619
timestamp 1516325494
transform 1 0 3247 0 1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_244
timestamp 1516325494
transform -1 0 3315 0 1 1138
box 0 0 53 49
use FILL  FILL_AND2X2_237
timestamp 1516325494
transform 1 0 3316 0 1 1138
box 0 0 8 49
use AND2X2  AND2X2_237
timestamp 1516325494
transform 1 0 3323 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_418
timestamp 1516325494
transform 1 0 3342 0 1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_223
timestamp 1516325494
transform 1 0 3361 0 1 1138
box 0 0 8 49
use OR2X2  OR2X2_223
timestamp 1516325494
transform 1 0 3369 0 1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_224
timestamp 1516325494
transform 1 0 3388 0 1 1138
box 0 0 8 49
use OR2X2  OR2X2_224
timestamp 1516325494
transform 1 0 3395 0 1 1138
box 0 0 19 49
use FILL  FILL_OR2X2_222
timestamp 1516325494
transform 1 0 3414 0 1 1138
box 0 0 8 49
use OR2X2  OR2X2_222
timestamp 1516325494
transform 1 0 3422 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_2021
timestamp 1516325494
transform 1 0 3441 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_417
timestamp 1516325494
transform 1 0 3460 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_391
timestamp 1516325494
transform 1 0 3479 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_712
timestamp 1516325494
transform 1 0 3498 0 1 1138
box 0 0 53 49
use OR2X2  OR2X2_395
timestamp 1516325494
transform -1 0 3570 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_392
timestamp 1516325494
transform -1 0 3589 0 1 1138
box 0 0 19 49
use OR2X2  OR2X2_390
timestamp 1516325494
transform -1 0 3608 0 1 1138
box 0 0 19 49
use AND2X2  AND2X2_416
timestamp 1516325494
transform -1 0 3627 0 1 1138
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_224
timestamp 1516325494
transform 1 0 3627 0 1 1138
box 0 0 53 49
use MUX2X1  MUX2X1_640
timestamp 1516325494
transform 1 0 3680 0 1 1138
box 0 0 30 49
use NAND2X1  NAND2X1_640
timestamp 1516325494
transform 1 0 3711 0 1 1138
box 0 0 15 49
use INVX1  INVX1_266
timestamp 1516325494
transform 1 0 3726 0 1 1138
box 0 0 11 49
use FILL  FILL_BUFX2_834
timestamp 1516325494
transform -1 0 3745 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_834
timestamp 1516325494
transform -1 0 3760 0 1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_282
timestamp 1516325494
transform -1 0 3768 0 1 1138
box 0 0 8 49
use BUFX2  BUFX2_282
timestamp 1516325494
transform -1 0 3783 0 1 1138
box 0 0 15 49
use FILL  FILL_AND2X2_240
timestamp 1516325494
transform -1 0 3791 0 1 1138
box 0 0 8 49
use AND2X2  AND2X2_240
timestamp 1516325494
transform -1 0 3810 0 1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_276
timestamp 1516325494
transform 1 0 3810 0 1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_276
timestamp 1516325494
transform -1 0 3855 0 1 1138
box 0 0 30 49
use INVX1  INVX1_303
timestamp 1516325494
transform -1 0 3866 0 1 1138
box 0 0 11 49
use OR2X2  OR2X2_1279
timestamp 1516325494
transform 1 0 2176 0 -1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_468
timestamp 1516325494
transform 1 0 2195 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_564
timestamp 1516325494
transform 1 0 2210 0 -1 1138
box 0 0 53 49
use FILL  FILL_BUFX2_243
timestamp 1516325494
transform 1 0 2263 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_243
timestamp 1516325494
transform 1 0 2271 0 -1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_142
timestamp 1516325494
transform 1 0 2286 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_142
timestamp 1516325494
transform 1 0 2293 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_84
timestamp 1516325494
transform 1 0 2309 0 -1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_148
timestamp 1516325494
transform 1 0 2362 0 -1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_148
timestamp 1516325494
transform 1 0 2377 0 -1 1138
box 0 0 30 49
use FILL  FILL_BUFX2_796
timestamp 1516325494
transform 1 0 2407 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_796
timestamp 1516325494
transform 1 0 2415 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_20
timestamp 1516325494
transform 1 0 2430 0 -1 1138
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_32
timestamp 1516325494
transform 1 0 2483 0 -1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_128
timestamp 1516325494
transform 1 0 2537 0 -1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_128
timestamp 1516325494
transform -1 0 2582 0 -1 1138
box 0 0 30 49
use FILL  FILL_BUFX2_146
timestamp 1516325494
transform -1 0 2590 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_146
timestamp 1516325494
transform -1 0 2605 0 -1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_3
timestamp 1516325494
transform -1 0 2620 0 -1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_15
timestamp 1516325494
transform -1 0 2635 0 -1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_4
timestamp 1516325494
transform -1 0 2650 0 -1 1138
box 0 0 15 49
use NAND3X1  NAND3X1_7
timestamp 1516325494
transform -1 0 2670 0 -1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_6
timestamp 1516325494
transform -1 0 2689 0 -1 1138
box 0 0 19 49
use INVX1  INVX1_3
timestamp 1516325494
transform -1 0 2700 0 -1 1138
box 0 0 11 49
use NAND3X1  NAND3X1_10
timestamp 1516325494
transform -1 0 2719 0 -1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_103
timestamp 1516325494
transform -1 0 2738 0 -1 1138
box 0 0 19 49
use INVX1  INVX1_319
timestamp 1516325494
transform -1 0 2749 0 -1 1138
box 0 0 11 49
use INVX1  INVX1_322
timestamp 1516325494
transform -1 0 2760 0 -1 1138
box 0 0 11 49
use NAND3X1  NAND3X1_5
timestamp 1516325494
transform -1 0 2780 0 -1 1138
box 0 0 19 49
use NAND3X1  NAND3X1_4
timestamp 1516325494
transform -1 0 2799 0 -1 1138
box 0 0 19 49
use INVX1  INVX1_2
timestamp 1516325494
transform -1 0 2810 0 -1 1138
box 0 0 11 49
use MUX2X1  MUX2X1_512
timestamp 1516325494
transform -1 0 2840 0 -1 1138
box 0 0 30 49
use FILL  FILL_BUFX2_858
timestamp 1516325494
transform -1 0 2849 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_858
timestamp 1516325494
transform -1 0 2863 0 -1 1138
box 0 0 15 49
use NOR2X1  NOR2X1_9
timestamp 1516325494
transform 1 0 2863 0 -1 1138
box 0 0 15 49
use FILL  FILL_OR2X2_27
timestamp 1516325494
transform -1 0 2887 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_27
timestamp 1516325494
transform -1 0 2905 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_27
timestamp 1516325494
transform -1 0 2913 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_27
timestamp 1516325494
transform -1 0 2932 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_704
timestamp 1516325494
transform -1 0 2940 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_704
timestamp 1516325494
transform -1 0 2954 0 -1 1138
box 0 0 15 49
use FILL  FILL_AND2X2_28
timestamp 1516325494
transform -1 0 2963 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_28
timestamp 1516325494
transform -1 0 2981 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_380
timestamp 1516325494
transform -1 0 2989 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_380
timestamp 1516325494
transform -1 0 3004 0 -1 1138
box 0 0 15 49
use NAND2X1  NAND2X1_582
timestamp 1516325494
transform 1 0 3004 0 -1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_582
timestamp 1516325494
transform -1 0 3049 0 -1 1138
box 0 0 30 49
use FILL  FILL_BUFX2_396
timestamp 1516325494
transform 1 0 3050 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_396
timestamp 1516325494
transform 1 0 3057 0 -1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_108
timestamp 1516325494
transform -1 0 3080 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_108
timestamp 1516325494
transform -1 0 3095 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_253
timestamp 1516325494
transform 1 0 3095 0 -1 1138
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_162
timestamp 1516325494
transform 1 0 3148 0 -1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_226
timestamp 1516325494
transform 1 0 3202 0 -1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_226
timestamp 1516325494
transform -1 0 3247 0 -1 1138
box 0 0 30 49
use FILL  FILL_BUFX2_206
timestamp 1516325494
transform 1 0 3247 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_206
timestamp 1516325494
transform 1 0 3255 0 -1 1138
box 0 0 15 49
use OR2X2  OR2X2_1590
timestamp 1516325494
transform -1 0 3289 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_221
timestamp 1516325494
transform 1 0 3289 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_221
timestamp 1516325494
transform 1 0 3297 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1722
timestamp 1516325494
transform -1 0 3335 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_222
timestamp 1516325494
transform 1 0 3335 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_222
timestamp 1516325494
transform 1 0 3342 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_238
timestamp 1516325494
transform -1 0 3369 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_238
timestamp 1516325494
transform -1 0 3388 0 -1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_748
timestamp 1516325494
transform -1 0 3403 0 -1 1138
box 0 0 15 49
use FILL  FILL_OR2X2_227
timestamp 1516325494
transform -1 0 3411 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_227
timestamp 1516325494
transform -1 0 3430 0 -1 1138
box 0 0 19 49
use MUX2X1  MUX2X1_596
timestamp 1516325494
transform 1 0 3430 0 -1 1138
box 0 0 30 49
use NAND2X1  NAND2X1_596
timestamp 1516325494
transform -1 0 3475 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_276
timestamp 1516325494
transform -1 0 3528 0 -1 1138
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_256
timestamp 1516325494
transform 1 0 3528 0 -1 1138
box 0 0 53 49
use NAND2X1  NAND2X1_224
timestamp 1516325494
transform 1 0 3582 0 -1 1138
box 0 0 15 49
use MUX2X1  MUX2X1_224
timestamp 1516325494
transform -1 0 3627 0 -1 1138
box 0 0 30 49
use FILL  FILL_BUFX2_278
timestamp 1516325494
transform 1 0 3627 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_278
timestamp 1516325494
transform 1 0 3635 0 -1 1138
box 0 0 15 49
use FILL  FILL_OR2X2_226
timestamp 1516325494
transform -1 0 3658 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_226
timestamp 1516325494
transform -1 0 3677 0 -1 1138
box 0 0 19 49
use FILL  FILL_BUFX2_439
timestamp 1516325494
transform 1 0 3677 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_439
timestamp 1516325494
transform 1 0 3684 0 -1 1138
box 0 0 15 49
use FILL  FILL_BUFX2_413
timestamp 1516325494
transform -1 0 3707 0 -1 1138
box 0 0 8 49
use BUFX2  BUFX2_413
timestamp 1516325494
transform -1 0 3722 0 -1 1138
box 0 0 15 49
use FILL  FILL_OR2X2_225
timestamp 1516325494
transform -1 0 3730 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_225
timestamp 1516325494
transform -1 0 3749 0 -1 1138
box 0 0 19 49
use FILL  FILL_AND2X2_241
timestamp 1516325494
transform -1 0 3757 0 -1 1138
box 0 0 8 49
use AND2X2  AND2X2_241
timestamp 1516325494
transform -1 0 3775 0 -1 1138
box 0 0 19 49
use AND2X2  AND2X2_1748
timestamp 1516325494
transform -1 0 3794 0 -1 1138
box 0 0 19 49
use NAND2X1  NAND2X1_372
timestamp 1516325494
transform 1 0 3794 0 -1 1138
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_148
timestamp 1516325494
transform 1 0 3810 0 -1 1138
box 0 0 53 49
use FILL  FILL_23_1
timestamp 1516325494
transform -1 0 3871 0 -1 1138
box 0 0 8 49
use OR2X2  OR2X2_643
timestamp 1516325494
transform -1 0 21 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_509
timestamp 1516325494
transform 1 0 21 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_451
timestamp 1516325494
transform 1 0 40 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_619
timestamp 1516325494
transform -1 0 78 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_766
timestamp 1516325494
transform -1 0 97 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_914
timestamp 1516325494
transform -1 0 116 0 1 1039
box 0 0 19 49
use INVX2  INVX2_1
timestamp 1516325494
transform 1 0 116 0 1 1039
box 0 0 11 49
use OR2X2  OR2X2_731
timestamp 1516325494
transform -1 0 146 0 1 1039
box 0 0 19 49
use NOR3X1  NOR3X1_8
timestamp 1516325494
transform 1 0 146 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_527
timestamp 1516325494
transform 1 0 165 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_728
timestamp 1516325494
transform -1 0 203 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_843
timestamp 1516325494
transform 1 0 203 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1052
timestamp 1516325494
transform 1 0 222 0 1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_667
timestamp 1516325494
transform 1 0 241 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_667
timestamp 1516325494
transform 1 0 249 0 1 1039
box 0 0 15 49
use AOI21X1  AOI21X1_23
timestamp 1516325494
transform 1 0 264 0 1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_693
timestamp 1516325494
transform -1 0 298 0 1 1039
box 0 0 15 49
use AND2X2  AND2X2_982
timestamp 1516325494
transform -1 0 317 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1027
timestamp 1516325494
transform 1 0 317 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_776
timestamp 1516325494
transform -1 0 355 0 1 1039
box 0 0 19 49
use MUX2X1  MUX2X1_720
timestamp 1516325494
transform -1 0 385 0 1 1039
box 0 0 30 49
use AND2X2  AND2X2_1032
timestamp 1516325494
transform -1 0 405 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_470
timestamp 1516325494
transform 1 0 405 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_431
timestamp 1516325494
transform 1 0 424 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_818
timestamp 1516325494
transform -1 0 462 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_817
timestamp 1516325494
transform -1 0 481 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_690
timestamp 1516325494
transform -1 0 500 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_479
timestamp 1516325494
transform -1 0 519 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_543
timestamp 1516325494
transform -1 0 538 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_659
timestamp 1516325494
transform 1 0 538 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_819
timestamp 1516325494
transform -1 0 576 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_715
timestamp 1516325494
transform 1 0 576 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_850
timestamp 1516325494
transform -1 0 614 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_849
timestamp 1516325494
transform -1 0 633 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_600
timestamp 1516325494
transform 1 0 633 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_716
timestamp 1516325494
transform -1 0 671 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_714
timestamp 1516325494
transform 1 0 671 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_599
timestamp 1516325494
transform -1 0 709 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_708
timestamp 1516325494
transform 1 0 709 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_717
timestamp 1516325494
transform 1 0 728 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_711
timestamp 1516325494
transform -1 0 766 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_798
timestamp 1516325494
transform 1 0 766 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_788
timestamp 1516325494
transform 1 0 785 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_667
timestamp 1516325494
transform 1 0 804 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_741
timestamp 1516325494
transform -1 0 842 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_906
timestamp 1516325494
transform -1 0 861 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1000
timestamp 1516325494
transform 1 0 861 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1001
timestamp 1516325494
transform -1 0 899 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_774
timestamp 1516325494
transform -1 0 918 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_845
timestamp 1516325494
transform -1 0 937 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_926
timestamp 1516325494
transform -1 0 956 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_830
timestamp 1516325494
transform -1 0 975 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_998
timestamp 1516325494
transform -1 0 994 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1055
timestamp 1516325494
transform -1 0 1013 0 1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_666
timestamp 1516325494
transform 1 0 1013 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_666
timestamp 1516325494
transform 1 0 1020 0 1 1039
box 0 0 15 49
use INVX1  INVX1_29
timestamp 1516325494
transform 1 0 1036 0 1 1039
box 0 0 11 49
use INVX1  INVX1_28
timestamp 1516325494
transform 1 0 1047 0 1 1039
box 0 0 11 49
use MUX2X1  MUX2X1_796
timestamp 1516325494
transform -1 0 1088 0 1 1039
box 0 0 30 49
use INVX1  INVX1_146
timestamp 1516325494
transform 1 0 1089 0 1 1039
box 0 0 11 49
use FILL  FILL_BUFX2_62
timestamp 1516325494
transform -1 0 1108 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_62
timestamp 1516325494
transform -1 0 1123 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_779
timestamp 1516325494
transform 1 0 1123 0 1 1039
box 0 0 30 49
use MUX2X1  MUX2X1_783
timestamp 1516325494
transform 1 0 1153 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_139
timestamp 1516325494
transform 1 0 1184 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_139
timestamp 1516325494
transform 1 0 1191 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_749
timestamp 1516325494
transform -1 0 1215 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_749
timestamp 1516325494
transform -1 0 1229 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_273
timestamp 1516325494
transform 1 0 1229 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_273
timestamp 1516325494
transform 1 0 1237 0 1 1039
box 0 0 15 49
use OR2X2  OR2X2_1284
timestamp 1516325494
transform -1 0 1271 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1283
timestamp 1516325494
transform -1 0 1290 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1282
timestamp 1516325494
transform -1 0 1309 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1281
timestamp 1516325494
transform -1 0 1328 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1512
timestamp 1516325494
transform -1 0 1347 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1276
timestamp 1516325494
transform -1 0 1366 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1765
timestamp 1516325494
transform -1 0 1385 0 1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_249
timestamp 1516325494
transform 1 0 1385 0 1 1039
box 0 0 8 49
use AND2X2  AND2X2_249
timestamp 1516325494
transform 1 0 1393 0 1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_442
timestamp 1516325494
transform 1 0 1412 0 1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_410
timestamp 1516325494
transform 1 0 1465 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_410
timestamp 1516325494
transform -1 0 1510 0 1 1039
box 0 0 30 49
use AND2X2  AND2X2_1796
timestamp 1516325494
transform -1 0 1530 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1652
timestamp 1516325494
transform -1 0 1549 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1651
timestamp 1516325494
transform -1 0 1568 0 1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_598
timestamp 1516325494
transform 1 0 1568 0 1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_22
timestamp 1516325494
transform 1 0 1621 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_22
timestamp 1516325494
transform -1 0 1666 0 1 1039
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_438
timestamp 1516325494
transform 1 0 1666 0 1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_406
timestamp 1516325494
transform 1 0 1720 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_406
timestamp 1516325494
transform -1 0 1765 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_505
timestamp 1516325494
transform 1 0 1765 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_505
timestamp 1516325494
transform 1 0 1773 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_521
timestamp 1516325494
transform -1 0 1818 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_581
timestamp 1516325494
transform 1 0 1818 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_581
timestamp 1516325494
transform 1 0 1826 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_725
timestamp 1516325494
transform -1 0 1849 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_725
timestamp 1516325494
transform -1 0 1864 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_289
timestamp 1516325494
transform 1 0 1864 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_289
timestamp 1516325494
transform 1 0 1872 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_792
timestamp 1516325494
transform -1 0 1895 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_792
timestamp 1516325494
transform -1 0 1909 0 1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_509
timestamp 1516325494
transform 1 0 1910 0 1 1039
box 0 0 53 49
use MUX2X1  MUX2X1_524
timestamp 1516325494
transform 1 0 1963 0 1 1039
box 0 0 30 49
use OR2X2  OR2X2_1879
timestamp 1516325494
transform -1 0 2012 0 1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_573
timestamp 1516325494
transform 1 0 2012 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_573
timestamp 1516325494
transform -1 0 2057 0 1 1039
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_125
timestamp 1516325494
transform 1 0 2058 0 1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_93
timestamp 1516325494
transform 1 0 2111 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_93
timestamp 1516325494
transform -1 0 2156 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_814
timestamp 1516325494
transform -1 0 2165 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_814
timestamp 1516325494
transform -1 0 2179 0 1 1039
box 0 0 15 49
use AND2X2  AND2X2_1511
timestamp 1516325494
transform -1 0 2198 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1280
timestamp 1516325494
transform -1 0 2217 0 1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_546
timestamp 1516325494
transform -1 0 2232 0 1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_482
timestamp 1516325494
transform 1 0 2233 0 1 1039
box 0 0 53 49
use MUX2X1  MUX2X1_546
timestamp 1516325494
transform -1 0 2316 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_824
timestamp 1516325494
transform -1 0 2324 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_824
timestamp 1516325494
transform -1 0 2339 0 1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_105
timestamp 1516325494
transform 1 0 2339 0 1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_73
timestamp 1516325494
transform 1 0 2392 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_73
timestamp 1516325494
transform -1 0 2437 0 1 1039
box 0 0 30 49
use MUX2X1  MUX2X1_84
timestamp 1516325494
transform 1 0 2438 0 1 1039
box 0 0 30 49
use NAND2X1  NAND2X1_84
timestamp 1516325494
transform -1 0 2483 0 1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_116
timestamp 1516325494
transform -1 0 2536 0 1 1039
box 0 0 53 49
use OR2X2  OR2X2_1610
timestamp 1516325494
transform 1 0 2537 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1764
timestamp 1516325494
transform 1 0 2556 0 1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_434
timestamp 1516325494
transform 1 0 2575 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_434
timestamp 1516325494
transform 1 0 2582 0 1 1039
box 0 0 15 49
use NAND3X1  NAND3X1_3
timestamp 1516325494
transform -1 0 2616 0 1 1039
box 0 0 19 49
use MUX2X1  MUX2X1_564
timestamp 1516325494
transform 1 0 2616 0 1 1039
box 0 0 30 49
use NAND2X1  NAND2X1_564
timestamp 1516325494
transform -1 0 2662 0 1 1039
box 0 0 15 49
use OR2X2  OR2X2_1609
timestamp 1516325494
transform -1 0 2681 0 1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_500
timestamp 1516325494
transform -1 0 2734 0 1 1039
box 0 0 53 49
use NOR3X1  NOR3X1_33
timestamp 1516325494
transform -1 0 2753 0 1 1039
box 0 0 19 49
use INVX1  INVX1_321
timestamp 1516325494
transform -1 0 2764 0 1 1039
box 0 0 11 49
use NOR2X1  NOR2X1_2
timestamp 1516325494
transform 1 0 2765 0 1 1039
box 0 0 15 49
use NOR2X1  NOR2X1_13
timestamp 1516325494
transform -1 0 2795 0 1 1039
box 0 0 15 49
use NAND3X1  NAND3X1_8
timestamp 1516325494
transform 1 0 2795 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1014
timestamp 1516325494
transform -1 0 2833 0 1 1039
box 0 0 19 49
use NAND3X1  NAND3X1_2
timestamp 1516325494
transform -1 0 2852 0 1 1039
box 0 0 19 49
use NOR2X1  NOR2X1_16
timestamp 1516325494
transform 1 0 2852 0 1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_320
timestamp 1516325494
transform -1 0 2920 0 1 1039
box 0 0 53 49
use AND2X2  AND2X2_1423
timestamp 1516325494
transform 1 0 2920 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1166
timestamp 1516325494
transform -1 0 2958 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1424
timestamp 1516325494
transform -1 0 2977 0 1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_486
timestamp 1516325494
transform 1 0 2977 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_486
timestamp 1516325494
transform 1 0 2985 0 1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_262
timestamp 1516325494
transform 1 0 3000 0 1 1039
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_198
timestamp 1516325494
transform 1 0 3053 0 1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_614
timestamp 1516325494
transform 1 0 3107 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_614
timestamp 1516325494
transform -1 0 3152 0 1 1039
box 0 0 30 49
use MUX2X1  MUX2X1_221
timestamp 1516325494
transform -1 0 3182 0 1 1039
box 0 0 30 49
use OAI21X1  OAI21X1_55
timestamp 1516325494
transform 1 0 3183 0 1 1039
box 0 0 19 49
use OAI21X1  OAI21X1_56
timestamp 1516325494
transform 1 0 3202 0 1 1039
box 0 0 19 49
use OAI21X1  OAI21X1_54
timestamp 1516325494
transform -1 0 3240 0 1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_621
timestamp 1516325494
transform 1 0 3240 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_621
timestamp 1516325494
transform 1 0 3247 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_197
timestamp 1516325494
transform 1 0 3262 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_197
timestamp 1516325494
transform 1 0 3270 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_557
timestamp 1516325494
transform -1 0 3293 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_557
timestamp 1516325494
transform -1 0 3308 0 1 1039
box 0 0 15 49
use OR2X2  OR2X2_1556
timestamp 1516325494
transform -1 0 3327 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1723
timestamp 1516325494
transform -1 0 3346 0 1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_209
timestamp 1516325494
transform 1 0 3346 0 1 1039
box 0 0 8 49
use OR2X2  OR2X2_209
timestamp 1516325494
transform 1 0 3354 0 1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_223
timestamp 1516325494
transform 1 0 3373 0 1 1039
box 0 0 8 49
use AND2X2  AND2X2_223
timestamp 1516325494
transform 1 0 3380 0 1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_595
timestamp 1516325494
transform 1 0 3399 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_595
timestamp 1516325494
transform -1 0 3444 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_45
timestamp 1516325494
transform -1 0 3453 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_45
timestamp 1516325494
transform -1 0 3467 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_660
timestamp 1516325494
transform 1 0 3468 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_660
timestamp 1516325494
transform 1 0 3475 0 1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_171
timestamp 1516325494
transform -1 0 3498 0 1 1039
box 0 0 8 49
use BUFX2  BUFX2_171
timestamp 1516325494
transform -1 0 3513 0 1 1039
box 0 0 15 49
use NAND2X1  NAND2X1_211
timestamp 1516325494
transform 1 0 3513 0 1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_211
timestamp 1516325494
transform -1 0 3558 0 1 1039
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_243
timestamp 1516325494
transform -1 0 3612 0 1 1039
box 0 0 53 49
use AND2X2  AND2X2_1747
timestamp 1516325494
transform 1 0 3612 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1589
timestamp 1516325494
transform -1 0 3650 0 1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_239
timestamp 1516325494
transform 1 0 3650 0 1 1039
box 0 0 8 49
use AND2X2  AND2X2_239
timestamp 1516325494
transform 1 0 3658 0 1 1039
box 0 0 19 49
use MUX2X1  MUX2X1_627
timestamp 1516325494
transform -1 0 3707 0 1 1039
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_211
timestamp 1516325494
transform -1 0 3760 0 1 1039
box 0 0 53 49
use OR2X2  OR2X2_1588
timestamp 1516325494
transform -1 0 3779 0 1 1039
box 0 0 19 49
use AND2X2  AND2X2_1749
timestamp 1516325494
transform -1 0 3798 0 1 1039
box 0 0 19 49
use MUX2X1  MUX2X1_372
timestamp 1516325494
transform -1 0 3828 0 1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_294
timestamp 1516325494
transform 1 0 2 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_294
timestamp 1516325494
transform 1 0 10 0 -1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_299
timestamp 1516325494
transform 1 0 25 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_299
timestamp 1516325494
transform 1 0 32 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_621
timestamp 1516325494
transform 1 0 48 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_919
timestamp 1516325494
transform 1 0 67 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1003
timestamp 1516325494
transform 1 0 86 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_836
timestamp 1516325494
transform -1 0 124 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_745
timestamp 1516325494
transform -1 0 143 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_606
timestamp 1516325494
transform 1 0 143 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_723
timestamp 1516325494
transform -1 0 181 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_669
timestamp 1516325494
transform 1 0 181 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_669
timestamp 1516325494
transform 1 0 188 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_710
timestamp 1516325494
transform -1 0 222 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_842
timestamp 1516325494
transform -1 0 241 0 -1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_692
timestamp 1516325494
transform 1 0 241 0 -1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_719
timestamp 1516325494
transform -1 0 287 0 -1 1039
box 0 0 30 49
use AND2X2  AND2X2_682
timestamp 1516325494
transform -1 0 306 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_772
timestamp 1516325494
transform 1 0 306 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_649
timestamp 1516325494
transform 1 0 325 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_433
timestamp 1516325494
transform 1 0 344 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_478
timestamp 1516325494
transform 1 0 363 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_430
timestamp 1516325494
transform 1 0 382 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_856
timestamp 1516325494
transform -1 0 420 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_296
timestamp 1516325494
transform -1 0 428 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_296
timestamp 1516325494
transform -1 0 443 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_783
timestamp 1516325494
transform -1 0 462 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_569
timestamp 1516325494
transform 1 0 462 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_568
timestamp 1516325494
transform 1 0 481 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_667
timestamp 1516325494
transform 1 0 500 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_566
timestamp 1516325494
transform -1 0 538 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_548
timestamp 1516325494
transform 1 0 538 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_648
timestamp 1516325494
transform -1 0 576 0 -1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_660
timestamp 1516325494
transform 1 0 576 0 -1 1039
box 0 0 15 49
use NAND3X1  NAND3X1_33
timestamp 1516325494
transform 1 0 591 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_751
timestamp 1516325494
transform 1 0 610 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_629
timestamp 1516325494
transform 1 0 629 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_715
timestamp 1516325494
transform 1 0 648 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_716
timestamp 1516325494
transform 1 0 667 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_492
timestamp 1516325494
transform -1 0 705 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_700
timestamp 1516325494
transform 1 0 705 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_590
timestamp 1516325494
transform 1 0 724 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_703
timestamp 1516325494
transform -1 0 762 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_791
timestamp 1516325494
transform -1 0 781 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_852
timestamp 1516325494
transform 1 0 781 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_720
timestamp 1516325494
transform 1 0 800 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_884
timestamp 1516325494
transform 1 0 819 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_756
timestamp 1516325494
transform -1 0 857 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_904
timestamp 1516325494
transform -1 0 876 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_947
timestamp 1516325494
transform 1 0 876 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_929
timestamp 1516325494
transform 1 0 895 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_791
timestamp 1516325494
transform -1 0 933 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_950
timestamp 1516325494
transform -1 0 952 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_997
timestamp 1516325494
transform -1 0 971 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_829
timestamp 1516325494
transform -1 0 990 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_995
timestamp 1516325494
transform -1 0 1009 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_728
timestamp 1516325494
transform 1 0 1009 0 -1 1039
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_729
timestamp 1516325494
transform -1 0 1115 0 -1 1039
box 0 0 53 49
use INVX1  INVX1_218
timestamp 1516325494
transform -1 0 1126 0 -1 1039
box 0 0 11 49
use FILL  FILL_BUFX2_638
timestamp 1516325494
transform -1 0 1135 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_638
timestamp 1516325494
transform -1 0 1149 0 -1 1039
box 0 0 15 49
use INVX1  INVX1_201
timestamp 1516325494
transform -1 0 1161 0 -1 1039
box 0 0 11 49
use INVX1  INVX1_205
timestamp 1516325494
transform -1 0 1172 0 -1 1039
box 0 0 11 49
use AND2X2  AND2X2_272
timestamp 1516325494
transform -1 0 1191 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1797
timestamp 1516325494
transform 1 0 1191 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_801
timestamp 1516325494
transform -1 0 1218 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_801
timestamp 1516325494
transform -1 0 1233 0 -1 1039
box 0 0 15 49
use FILL  FILL_AND2X2_80
timestamp 1516325494
transform -1 0 1241 0 -1 1039
box 0 0 8 49
use AND2X2  AND2X2_80
timestamp 1516325494
transform -1 0 1260 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1504
timestamp 1516325494
transform 1 0 1260 0 -1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_39
timestamp 1516325494
transform -1 0 1287 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_39
timestamp 1516325494
transform -1 0 1305 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_2002
timestamp 1516325494
transform -1 0 1324 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1510
timestamp 1516325494
transform -1 0 1343 0 -1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_84
timestamp 1516325494
transform -1 0 1351 0 -1 1039
box 0 0 8 49
use AND2X2  AND2X2_84
timestamp 1516325494
transform -1 0 1370 0 -1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_78
timestamp 1516325494
transform 1 0 1370 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_78
timestamp 1516325494
transform 1 0 1378 0 -1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_83
timestamp 1516325494
transform -1 0 1405 0 -1 1039
box 0 0 8 49
use AND2X2  AND2X2_83
timestamp 1516325494
transform -1 0 1423 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_287
timestamp 1516325494
transform -1 0 1431 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_287
timestamp 1516325494
transform -1 0 1446 0 -1 1039
box 0 0 15 49
use FILL  FILL_AND2X2_81
timestamp 1516325494
transform -1 0 1454 0 -1 1039
box 0 0 8 49
use AND2X2  AND2X2_81
timestamp 1516325494
transform -1 0 1473 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_2092
timestamp 1516325494
transform 1 0 1473 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_1999
timestamp 1516325494
transform -1 0 1511 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_124
timestamp 1516325494
transform 1 0 1511 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_124
timestamp 1516325494
transform 1 0 1518 0 -1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_818
timestamp 1516325494
transform 1 0 1533 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_818
timestamp 1516325494
transform 1 0 1541 0 -1 1039
box 0 0 15 49
use AND2X2  AND2X2_1351
timestamp 1516325494
transform 1 0 1556 0 -1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_121
timestamp 1516325494
transform -1 0 1583 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_121
timestamp 1516325494
transform -1 0 1602 0 -1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_119
timestamp 1516325494
transform -1 0 1610 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_119
timestamp 1516325494
transform -1 0 1628 0 -1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_126
timestamp 1516325494
transform -1 0 1636 0 -1 1039
box 0 0 8 49
use AND2X2  AND2X2_126
timestamp 1516325494
transform -1 0 1655 0 -1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_120
timestamp 1516325494
transform -1 0 1663 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_120
timestamp 1516325494
transform -1 0 1682 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1579
timestamp 1516325494
transform -1 0 1701 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_1371
timestamp 1516325494
transform 1 0 1701 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1509
timestamp 1516325494
transform -1 0 1739 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_1277
timestamp 1516325494
transform -1 0 1758 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_55
timestamp 1516325494
transform -1 0 1766 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_55
timestamp 1516325494
transform -1 0 1780 0 -1 1039
box 0 0 15 49
use NAND2X1  NAND2X1_521
timestamp 1516325494
transform 1 0 1780 0 -1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_521
timestamp 1516325494
transform -1 0 1849 0 -1 1039
box 0 0 53 49
use FILL  FILL_BUFX2_497
timestamp 1516325494
transform -1 0 1857 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_497
timestamp 1516325494
transform -1 0 1871 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1654
timestamp 1516325494
transform -1 0 1891 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_694
timestamp 1516325494
transform 1 0 1891 0 -1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_310
timestamp 1516325494
transform 1 0 1944 0 -1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_310
timestamp 1516325494
transform -1 0 1989 0 -1 1039
box 0 0 30 49
use NAND2X1  NAND2X1_524
timestamp 1516325494
transform -1 0 2004 0 -1 1039
box 0 0 15 49
use AND2X2  AND2X2_1971
timestamp 1516325494
transform -1 0 2024 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_795
timestamp 1516325494
transform 1 0 2024 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_795
timestamp 1516325494
transform 1 0 2031 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1880
timestamp 1516325494
transform -1 0 2065 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_524
timestamp 1516325494
transform -1 0 2118 0 -1 1039
box 0 0 53 49
use FILL  FILL_BUFX2_720
timestamp 1516325494
transform 1 0 2119 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_720
timestamp 1516325494
transform 1 0 2126 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1068
timestamp 1516325494
transform -1 0 2160 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_2
timestamp 1516325494
transform 1 0 2160 0 -1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_98
timestamp 1516325494
transform 1 0 2214 0 -1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_98
timestamp 1516325494
transform -1 0 2259 0 -1 1039
box 0 0 30 49
use OR2X2  OR2X2_1069
timestamp 1516325494
transform 1 0 2259 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1350
timestamp 1516325494
transform -1 0 2297 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_504
timestamp 1516325494
transform 1 0 2297 0 -1 1039
box 0 0 53 49
use FILL  FILL_BUFX2_501
timestamp 1516325494
transform -1 0 2358 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_501
timestamp 1516325494
transform -1 0 2373 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1070
timestamp 1516325494
transform -1 0 2392 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_98
timestamp 1516325494
transform 1 0 2392 0 -1 1039
box 0 0 53 49
use OR2X2  OR2X2_1190
timestamp 1516325494
transform -1 0 2464 0 -1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_70
timestamp 1516325494
transform 1 0 2464 0 -1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_70
timestamp 1516325494
transform -1 0 2510 0 -1 1039
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_102
timestamp 1516325494
transform -1 0 2563 0 -1 1039
box 0 0 53 49
use FILL  FILL_BUFX2_36
timestamp 1516325494
transform 1 0 2563 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_36
timestamp 1516325494
transform 1 0 2571 0 -1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_10
timestamp 1516325494
transform -1 0 2594 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_10
timestamp 1516325494
transform -1 0 2609 0 -1 1039
box 0 0 15 49
use NAND3X1  NAND3X1_101
timestamp 1516325494
transform 1 0 2609 0 -1 1039
box 0 0 19 49
use FILL  FILL_BUFX2_700
timestamp 1516325494
transform -1 0 2636 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_700
timestamp 1516325494
transform -1 0 2650 0 -1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_848
timestamp 1516325494
transform -1 0 2659 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_848
timestamp 1516325494
transform -1 0 2673 0 -1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_861
timestamp 1516325494
transform 1 0 2673 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_861
timestamp 1516325494
transform 1 0 2681 0 -1 1039
box 0 0 15 49
use FILL  FILL_OR2X2_31
timestamp 1516325494
transform -1 0 2704 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_31
timestamp 1516325494
transform -1 0 2723 0 -1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_512
timestamp 1516325494
transform 1 0 2723 0 -1 1039
box 0 0 15 49
use INVX1  INVX1_320
timestamp 1516325494
transform 1 0 2738 0 -1 1039
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_278
timestamp 1516325494
transform -1 0 2802 0 -1 1039
box 0 0 53 49
use FILL  FILL_OR2X2_28
timestamp 1516325494
transform -1 0 2811 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_28
timestamp 1516325494
transform -1 0 2829 0 -1 1039
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_230
timestamp 1516325494
transform 1 0 2829 0 -1 1039
box 0 0 53 49
use MUX2X1  MUX2X1_198
timestamp 1516325494
transform 1 0 2882 0 -1 1039
box 0 0 30 49
use NAND2X1  NAND2X1_198
timestamp 1516325494
transform -1 0 2928 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1167
timestamp 1516325494
transform -1 0 2947 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_1170
timestamp 1516325494
transform 1 0 2947 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_1194
timestamp 1516325494
transform 1 0 2966 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1952
timestamp 1516325494
transform 1 0 2985 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_1856
timestamp 1516325494
transform 1 0 3004 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1953
timestamp 1516325494
transform -1 0 3042 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_373
timestamp 1516325494
transform 1 0 3042 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_372
timestamp 1516325494
transform 1 0 3061 0 -1 1039
box 0 0 19 49
use OR2X2  OR2X2_349
timestamp 1516325494
transform 1 0 3080 0 -1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_221
timestamp 1516325494
transform 1 0 3099 0 -1 1039
box 0 0 15 49
use NAND2X1  NAND2X1_605
timestamp 1516325494
transform 1 0 3114 0 -1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_605
timestamp 1516325494
transform -1 0 3159 0 -1 1039
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_285
timestamp 1516325494
transform 1 0 3160 0 -1 1039
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_707
timestamp 1516325494
transform 1 0 3213 0 -1 1039
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_275
timestamp 1516325494
transform 1 0 3266 0 -1 1039
box 0 0 53 49
use FILL  FILL_BUFX2_769
timestamp 1516325494
transform -1 0 3327 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_769
timestamp 1516325494
transform -1 0 3342 0 -1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_268
timestamp 1516325494
transform 1 0 3342 0 -1 1039
box 0 0 53 49
use MUX2X1  MUX2X1_265
timestamp 1516325494
transform 1 0 3395 0 -1 1039
box 0 0 30 49
use NAND2X1  NAND2X1_265
timestamp 1516325494
transform -1 0 3441 0 -1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_157
timestamp 1516325494
transform 1 0 3441 0 -1 1039
box 0 0 53 49
use NAND2X1  NAND2X1_285
timestamp 1516325494
transform 1 0 3494 0 -1 1039
box 0 0 15 49
use MUX2X1  MUX2X1_285
timestamp 1516325494
transform -1 0 3539 0 -1 1039
box 0 0 30 49
use FILL  FILL_BUFX2_585
timestamp 1516325494
transform -1 0 3548 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_585
timestamp 1516325494
transform -1 0 3562 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1169
timestamp 1516325494
transform -1 0 3582 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1425
timestamp 1516325494
transform -1 0 3601 0 -1 1039
box 0 0 19 49
use FILL  FILL_OR2X2_30
timestamp 1516325494
transform -1 0 3609 0 -1 1039
box 0 0 8 49
use OR2X2  OR2X2_30
timestamp 1516325494
transform -1 0 3627 0 -1 1039
box 0 0 19 49
use FILL  FILL_AND2X2_29
timestamp 1516325494
transform -1 0 3635 0 -1 1039
box 0 0 8 49
use AND2X2  AND2X2_29
timestamp 1516325494
transform -1 0 3654 0 -1 1039
box 0 0 19 49
use NAND2X1  NAND2X1_627
timestamp 1516325494
transform 1 0 3654 0 -1 1039
box 0 0 15 49
use FILL  FILL_BUFX2_588
timestamp 1516325494
transform -1 0 3677 0 -1 1039
box 0 0 8 49
use BUFX2  BUFX2_588
timestamp 1516325494
transform -1 0 3692 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_1168
timestamp 1516325494
transform -1 0 3711 0 -1 1039
box 0 0 19 49
use AND2X2  AND2X2_1427
timestamp 1516325494
transform -1 0 3730 0 -1 1039
box 0 0 19 49
use MUX2X1  MUX2X1_358
timestamp 1516325494
transform 1 0 3730 0 -1 1039
box 0 0 30 49
use NAND2X1  NAND2X1_358
timestamp 1516325494
transform -1 0 3775 0 -1 1039
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_326
timestamp 1516325494
transform -1 0 3828 0 -1 1039
box 0 0 53 49
use AND2X2  AND2X2_1190
timestamp 1516325494
transform -1 0 3848 0 1 1039
box 0 0 19 49
use OR2X2  OR2X2_1008
timestamp 1516325494
transform 1 0 3848 0 1 1039
box 0 0 19 49
use NOR2X1  NOR2X1_164
timestamp 1516325494
transform -1 0 3844 0 -1 1039
box 0 0 15 49
use INVX1  INVX1_310
timestamp 1516325494
transform 1 0 3844 0 -1 1039
box 0 0 11 49
use NOR2X1  NOR2X1_159
timestamp 1516325494
transform -1 0 3870 0 -1 1039
box 0 0 15 49
use OR2X2  OR2X2_583
timestamp 1516325494
transform -1 0 21 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_692
timestamp 1516325494
transform -1 0 40 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_867
timestamp 1516325494
transform 1 0 40 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_502
timestamp 1516325494
transform -1 0 78 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_525
timestamp 1516325494
transform -1 0 97 0 1 940
box 0 0 19 49
use NOR3X1  NOR3X1_7
timestamp 1516325494
transform 1 0 97 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1008
timestamp 1516325494
transform -1 0 135 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_442
timestamp 1516325494
transform -1 0 154 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_494
timestamp 1516325494
transform -1 0 173 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_579
timestamp 1516325494
transform -1 0 192 0 1 940
box 0 0 19 49
use FILL  FILL_BUFX2_759
timestamp 1516325494
transform -1 0 200 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_759
timestamp 1516325494
transform -1 0 215 0 1 940
box 0 0 15 49
use AND2X2  AND2X2_839
timestamp 1516325494
transform -1 0 234 0 1 940
box 0 0 19 49
use MUX2X1  MUX2X1_724
timestamp 1516325494
transform 1 0 234 0 1 940
box 0 0 30 49
use MUX2X1  MUX2X1_727
timestamp 1516325494
transform -1 0 294 0 1 940
box 0 0 30 49
use AND2X2  AND2X2_981
timestamp 1516325494
transform 1 0 295 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_816
timestamp 1516325494
transform -1 0 333 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_775
timestamp 1516325494
transform -1 0 352 0 1 940
box 0 0 19 49
use MUX2X1  MUX2X1_717
timestamp 1516325494
transform -1 0 382 0 1 940
box 0 0 30 49
use AND2X2  AND2X2_980
timestamp 1516325494
transform -1 0 401 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1031
timestamp 1516325494
transform 1 0 401 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1030
timestamp 1516325494
transform -1 0 439 0 1 940
box 0 0 19 49
use NAND3X1  NAND3X1_24
timestamp 1516325494
transform -1 0 458 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_689
timestamp 1516325494
transform -1 0 477 0 1 940
box 0 0 19 49
use NOR2X1  NOR2X1_25
timestamp 1516325494
transform 1 0 477 0 1 940
box 0 0 15 49
use OR2X2  OR2X2_567
timestamp 1516325494
transform -1 0 511 0 1 940
box 0 0 19 49
use AOI21X1  AOI21X1_3
timestamp 1516325494
transform 1 0 511 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_424
timestamp 1516325494
transform -1 0 549 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_459
timestamp 1516325494
transform -1 0 568 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_565
timestamp 1516325494
transform -1 0 587 0 1 940
box 0 0 19 49
use NOR3X1  NOR3X1_9
timestamp 1516325494
transform -1 0 606 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_422
timestamp 1516325494
transform -1 0 625 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_485
timestamp 1516325494
transform -1 0 644 0 1 940
box 0 0 19 49
use NOR3X1  NOR3X1_10
timestamp 1516325494
transform -1 0 663 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_458
timestamp 1516325494
transform -1 0 682 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_561
timestamp 1516325494
transform -1 0 701 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_754
timestamp 1516325494
transform -1 0 720 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_693
timestamp 1516325494
transform -1 0 739 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_821
timestamp 1516325494
transform -1 0 758 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_589
timestamp 1516325494
transform 1 0 758 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_824
timestamp 1516325494
transform -1 0 796 0 1 940
box 0 0 19 49
use FILL  FILL_BUFX2_754
timestamp 1516325494
transform 1 0 796 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_754
timestamp 1516325494
transform 1 0 804 0 1 940
box 0 0 15 49
use AND2X2  AND2X2_885
timestamp 1516325494
transform 1 0 819 0 1 940
box 0 0 19 49
use FILL  FILL_BUFX2_760
timestamp 1516325494
transform -1 0 846 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_760
timestamp 1516325494
transform -1 0 861 0 1 940
box 0 0 15 49
use AND2X2  AND2X2_855
timestamp 1516325494
transform -1 0 880 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_905
timestamp 1516325494
transform -1 0 899 0 1 940
box 0 0 19 49
use MUX2X1  MUX2X1_731
timestamp 1516325494
transform -1 0 929 0 1 940
box 0 0 30 49
use MUX2X1  MUX2X1_737
timestamp 1516325494
transform 1 0 929 0 1 940
box 0 0 30 49
use OR2X2  OR2X2_808
timestamp 1516325494
transform -1 0 979 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_970
timestamp 1516325494
transform -1 0 998 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_949
timestamp 1516325494
transform 1 0 998 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_790
timestamp 1516325494
transform -1 0 1036 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_948
timestamp 1516325494
transform 1 0 1036 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_971
timestamp 1516325494
transform -1 0 1074 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_996
timestamp 1516325494
transform -1 0 1093 0 1 940
box 0 0 19 49
use MUX2X1  MUX2X1_745
timestamp 1516325494
transform -1 0 1123 0 1 940
box 0 0 30 49
use MUX2X1  MUX2X1_757
timestamp 1516325494
transform -1 0 1153 0 1 940
box 0 0 30 49
use INVX1  INVX1_221
timestamp 1516325494
transform -1 0 1164 0 1 940
box 0 0 11 49
use MUX2X1  MUX2X1_789
timestamp 1516325494
transform -1 0 1195 0 1 940
box 0 0 30 49
use OR2X2  OR2X2_1655
timestamp 1516325494
transform -1 0 1214 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_221
timestamp 1516325494
transform -1 0 1222 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_221
timestamp 1516325494
transform -1 0 1241 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1799
timestamp 1516325494
transform -1 0 1260 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_273
timestamp 1516325494
transform -1 0 1279 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1270
timestamp 1516325494
transform 1 0 1279 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1271
timestamp 1516325494
transform -1 0 1317 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_2001
timestamp 1516325494
transform -1 0 1336 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_81
timestamp 1516325494
transform -1 0 1344 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_81
timestamp 1516325494
transform -1 0 1362 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_80
timestamp 1516325494
transform -1 0 1370 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_80
timestamp 1516325494
transform -1 0 1389 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_79
timestamp 1516325494
transform -1 0 1397 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_79
timestamp 1516325494
transform -1 0 1416 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_77
timestamp 1516325494
transform -1 0 1424 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_77
timestamp 1516325494
transform -1 0 1442 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_82
timestamp 1516325494
transform -1 0 1450 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_82
timestamp 1516325494
transform -1 0 1469 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_2000
timestamp 1516325494
transform -1 0 1488 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1508
timestamp 1516325494
transform -1 0 1507 0 1 940
box 0 0 19 49
use FILL  FILL_BUFX2_591
timestamp 1516325494
transform 1 0 1507 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_591
timestamp 1516325494
transform 1 0 1514 0 1 940
box 0 0 15 49
use OR2X2  OR2X2_1998
timestamp 1516325494
transform -1 0 1549 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_2090
timestamp 1516325494
transform -1 0 1568 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1071
timestamp 1516325494
transform -1 0 1587 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_2089
timestamp 1516325494
transform -1 0 1606 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_122
timestamp 1516325494
transform 1 0 1606 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_122
timestamp 1516325494
transform 1 0 1613 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1349
timestamp 1516325494
transform -1 0 1651 0 1 940
box 0 0 19 49
use INVX2  INVX2_25
timestamp 1516325494
transform 1 0 1651 0 1 940
box 0 0 11 49
use AND2X2  AND2X2_2091
timestamp 1516325494
transform -1 0 1682 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_128
timestamp 1516325494
transform -1 0 1690 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_128
timestamp 1516325494
transform -1 0 1708 0 1 940
box 0 0 19 49
use OAI21X1  OAI21X1_29
timestamp 1516325494
transform 1 0 1708 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_127
timestamp 1516325494
transform 1 0 1727 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_127
timestamp 1516325494
transform 1 0 1735 0 1 940
box 0 0 19 49
use FILL  FILL_BUFX2_487
timestamp 1516325494
transform 1 0 1754 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_487
timestamp 1516325494
transform 1 0 1761 0 1 940
box 0 0 15 49
use OR2X2  OR2X2_1368
timestamp 1516325494
transform 1 0 1777 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1578
timestamp 1516325494
transform 1 0 1796 0 1 940
box 0 0 19 49
use INVX2  INVX2_18
timestamp 1516325494
transform 1 0 1815 0 1 940
box 0 0 11 49
use OR2X2  OR2X2_1875
timestamp 1516325494
transform -1 0 1845 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1278
timestamp 1516325494
transform -1 0 1864 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1798
timestamp 1516325494
transform -1 0 1883 0 1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_93
timestamp 1516325494
transform 1 0 1883 0 1 940
box 0 0 53 49
use NAND2X1  NAND2X1_157
timestamp 1516325494
transform 1 0 1936 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_157
timestamp 1516325494
transform -1 0 1981 0 1 940
box 0 0 30 49
use INVX2  INVX2_28
timestamp 1516325494
transform 1 0 1982 0 1 940
box 0 0 11 49
use OR2X2  OR2X2_1367
timestamp 1516325494
transform -1 0 2012 0 1 940
box 0 0 19 49
use NAND2X1  NAND2X1_105
timestamp 1516325494
transform 1 0 2012 0 1 940
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_9
timestamp 1516325494
transform 1 0 2027 0 1 940
box 0 0 53 49
use MUX2X1  MUX2X1_105
timestamp 1516325494
transform -1 0 2111 0 1 940
box 0 0 30 49
use AND2X2  AND2X2_1348
timestamp 1516325494
transform -1 0 2130 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1067
timestamp 1516325494
transform -1 0 2149 0 1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_514
timestamp 1516325494
transform 1 0 2149 0 1 940
box 0 0 53 49
use NAND2X1  NAND2X1_514
timestamp 1516325494
transform 1 0 2202 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_514
timestamp 1516325494
transform -1 0 2247 0 1 940
box 0 0 30 49
use FILL  FILL_BUFX2_49
timestamp 1516325494
transform -1 0 2256 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_49
timestamp 1516325494
transform -1 0 2270 0 1 940
box 0 0 15 49
use OR2X2  OR2X2_1729
timestamp 1516325494
transform 1 0 2271 0 1 940
box 0 0 19 49
use NAND2X1  NAND2X1_568
timestamp 1516325494
transform 1 0 2290 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_568
timestamp 1516325494
transform -1 0 2335 0 1 940
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_120
timestamp 1516325494
transform 1 0 2335 0 1 940
box 0 0 53 49
use MUX2X1  MUX2X1_88
timestamp 1516325494
transform 1 0 2388 0 1 940
box 0 0 30 49
use NAND2X1  NAND2X1_88
timestamp 1516325494
transform 1 0 2419 0 1 940
box 0 0 15 49
use NAND2X1  NAND2X1_66
timestamp 1516325494
transform 1 0 2434 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_66
timestamp 1516325494
transform -1 0 2479 0 1 940
box 0 0 30 49
use AND2X2  AND2X2_744
timestamp 1516325494
transform -1 0 21 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_620
timestamp 1516325494
transform 1 0 21 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_619
timestamp 1516325494
transform -1 0 59 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_743
timestamp 1516325494
transform -1 0 78 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_615
timestamp 1516325494
transform 1 0 78 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_680
timestamp 1516325494
transform 1 0 97 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_618
timestamp 1516325494
transform -1 0 135 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_722
timestamp 1516325494
transform 1 0 135 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_803
timestamp 1516325494
transform -1 0 173 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_835
timestamp 1516325494
transform -1 0 192 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1006
timestamp 1516325494
transform -1 0 211 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1051
timestamp 1516325494
transform 1 0 211 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_872
timestamp 1516325494
transform -1 0 249 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_726
timestamp 1516325494
transform 1 0 249 0 -1 940
box 0 0 30 49
use OR2X2  OR2X2_521
timestamp 1516325494
transform -1 0 298 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_607
timestamp 1516325494
transform -1 0 317 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_455
timestamp 1516325494
transform -1 0 336 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1050
timestamp 1516325494
transform -1 0 355 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1049
timestamp 1516325494
transform -1 0 374 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_871
timestamp 1516325494
transform -1 0 393 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_681
timestamp 1516325494
transform -1 0 423 0 -1 940
box 0 0 30 49
use OR2X2  OR2X2_870
timestamp 1516325494
transform -1 0 443 0 -1 940
box 0 0 19 49
use AOI21X1  AOI21X1_27
timestamp 1516325494
transform -1 0 462 0 -1 940
box 0 0 19 49
use NAND3X1  NAND3X1_15
timestamp 1516325494
transform -1 0 481 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_757
timestamp 1516325494
transform -1 0 489 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_757
timestamp 1516325494
transform -1 0 503 0 -1 940
box 0 0 15 49
use INVX1  INVX1_11
timestamp 1516325494
transform 1 0 504 0 -1 940
box 0 0 11 49
use FILL  FILL_BUFX2_672
timestamp 1516325494
transform 1 0 515 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_672
timestamp 1516325494
transform 1 0 523 0 -1 940
box 0 0 15 49
use NAND3X1  NAND3X1_23
timestamp 1516325494
transform 1 0 538 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_566
timestamp 1516325494
transform 1 0 557 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_491
timestamp 1516325494
transform -1 0 595 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_646
timestamp 1516325494
transform 1 0 595 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_547
timestamp 1516325494
transform -1 0 633 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_558
timestamp 1516325494
transform -1 0 652 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_483
timestamp 1516325494
transform -1 0 671 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_598
timestamp 1516325494
transform -1 0 690 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_712
timestamp 1516325494
transform -1 0 709 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_647
timestamp 1516325494
transform -1 0 728 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_701
timestamp 1516325494
transform 1 0 728 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_628
timestamp 1516325494
transform -1 0 766 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_752
timestamp 1516325494
transform 1 0 766 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_702
timestamp 1516325494
transform -1 0 804 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_643
timestamp 1516325494
transform -1 0 834 0 -1 940
box 0 0 30 49
use OR2X2  OR2X2_692
timestamp 1516325494
transform -1 0 853 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_700
timestamp 1516325494
transform 1 0 853 0 -1 940
box 0 0 30 49
use OR2X2  OR2X2_719
timestamp 1516325494
transform -1 0 903 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_773
timestamp 1516325494
transform -1 0 922 0 -1 940
box 0 0 19 49
use INVX1  INVX1_50
timestamp 1516325494
transform 1 0 922 0 -1 940
box 0 0 11 49
use AND2X2  AND2X2_928
timestamp 1516325494
transform -1 0 952 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_723
timestamp 1516325494
transform -1 0 982 0 -1 940
box 0 0 30 49
use MUX2X1  MUX2X1_728
timestamp 1516325494
transform -1 0 1012 0 -1 940
box 0 0 30 49
use MUX2X1  MUX2X1_730
timestamp 1516325494
transform -1 0 1043 0 -1 940
box 0 0 30 49
use MUX2X1  MUX2X1_775
timestamp 1516325494
transform 1 0 1043 0 -1 940
box 0 0 30 49
use MUX2X1  MUX2X1_742
timestamp 1516325494
transform -1 0 1104 0 -1 940
box 0 0 30 49
use MUX2X1  MUX2X1_748
timestamp 1516325494
transform 1 0 1104 0 -1 940
box 0 0 30 49
use FILL  FILL_BUFX2_318
timestamp 1516325494
transform 1 0 1134 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_318
timestamp 1516325494
transform 1 0 1142 0 -1 940
box 0 0 15 49
use FILL  FILL_BUFX2_776
timestamp 1516325494
transform -1 0 1165 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_776
timestamp 1516325494
transform -1 0 1180 0 -1 940
box 0 0 15 49
use INVX1  INVX1_211
timestamp 1516325494
transform -1 0 1191 0 -1 940
box 0 0 11 49
use OR2X2  OR2X2_256
timestamp 1516325494
transform 1 0 1191 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_263
timestamp 1516325494
transform -1 0 1229 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1502
timestamp 1516325494
transform -1 0 1248 0 -1 940
box 0 0 19 49
use FILL  FILL_AND2X2_79
timestamp 1516325494
transform 1 0 1248 0 -1 940
box 0 0 8 49
use AND2X2  AND2X2_79
timestamp 1516325494
transform 1 0 1256 0 -1 940
box 0 0 19 49
use FILL  FILL_OR2X2_75
timestamp 1516325494
transform 1 0 1275 0 -1 940
box 0 0 8 49
use OR2X2  OR2X2_75
timestamp 1516325494
transform 1 0 1283 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1265
timestamp 1516325494
transform -1 0 1321 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1500
timestamp 1516325494
transform -1 0 1340 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_684
timestamp 1516325494
transform -1 0 1348 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_684
timestamp 1516325494
transform -1 0 1362 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1074
timestamp 1516325494
transform -1 0 1381 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1073
timestamp 1516325494
transform -1 0 1400 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_604
timestamp 1516325494
transform 1 0 1400 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_604
timestamp 1516325494
transform 1 0 1408 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1884
timestamp 1516325494
transform -1 0 1442 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1883
timestamp 1516325494
transform -1 0 1461 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1072
timestamp 1516325494
transform -1 0 1480 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1066
timestamp 1516325494
transform -1 0 1499 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1345
timestamp 1516325494
transform -1 0 1518 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1347
timestamp 1516325494
transform -1 0 1537 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_384
timestamp 1516325494
transform 1 0 1537 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1972
timestamp 1516325494
transform 1 0 1556 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1882
timestamp 1516325494
transform -1 0 1594 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1881
timestamp 1516325494
transform -1 0 1613 0 -1 940
box 0 0 19 49
use FILL  FILL_OR2X2_123
timestamp 1516325494
transform -1 0 1621 0 -1 940
box 0 0 8 49
use OR2X2  OR2X2_123
timestamp 1516325494
transform -1 0 1640 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1876
timestamp 1516325494
transform -1 0 1659 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1968
timestamp 1516325494
transform -1 0 1678 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_382
timestamp 1516325494
transform -1 0 1697 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_386
timestamp 1516325494
transform 1 0 1697 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_386
timestamp 1516325494
transform 1 0 1704 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1372
timestamp 1516325494
transform 1 0 1720 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1577
timestamp 1516325494
transform 1 0 1739 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1366
timestamp 1516325494
transform -1 0 1777 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1575
timestamp 1516325494
transform 1 0 1777 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1967
timestamp 1516325494
transform -1 0 1815 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1874
timestamp 1516325494
transform -1 0 1834 0 -1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_477
timestamp 1516325494
transform 1 0 1834 0 -1 940
box 0 0 53 49
use NAND2X1  NAND2X1_349
timestamp 1516325494
transform 1 0 1887 0 -1 940
box 0 0 15 49
use MUX2X1  MUX2X1_349
timestamp 1516325494
transform 1 0 1902 0 -1 940
box 0 0 30 49
use OR2X2  OR2X2_1664
timestamp 1516325494
transform -1 0 1951 0 -1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_470
timestamp 1516325494
transform 1 0 1951 0 -1 940
box 0 0 53 49
use NAND2X1  NAND2X1_342
timestamp 1516325494
transform 1 0 2005 0 -1 940
box 0 0 15 49
use MUX2X1  MUX2X1_342
timestamp 1516325494
transform -1 0 2050 0 -1 940
box 0 0 30 49
use FILL  FILL_BUFX2_738
timestamp 1516325494
transform 1 0 2050 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_738
timestamp 1516325494
transform 1 0 2058 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1653
timestamp 1516325494
transform -1 0 2092 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_847
timestamp 1516325494
transform 1 0 2092 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_847
timestamp 1516325494
transform 1 0 2100 0 -1 940
box 0 0 15 49
use INVX8  INVX8_1
timestamp 1516325494
transform 1 0 2115 0 -1 940
box 0 0 27 49
use DFFPOSX1  DFFPOSX1_566
timestamp 1516325494
transform 1 0 2141 0 -1 940
box 0 0 53 49
use NAND2X1  NAND2X1_470
timestamp 1516325494
transform 1 0 2195 0 -1 940
box 0 0 15 49
use MUX2X1  MUX2X1_470
timestamp 1516325494
transform -1 0 2240 0 -1 940
box 0 0 30 49
use FILL  FILL_BUFX2_51
timestamp 1516325494
transform -1 0 2248 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_51
timestamp 1516325494
transform -1 0 2263 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1727
timestamp 1516325494
transform -1 0 2282 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_645
timestamp 1516325494
transform 1 0 2282 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_645
timestamp 1516325494
transform 1 0 2290 0 -1 940
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_536
timestamp 1516325494
transform 1 0 2305 0 -1 940
box 0 0 53 49
use NAND2X1  NAND2X1_536
timestamp 1516325494
transform 1 0 2358 0 -1 940
box 0 0 15 49
use MUX2X1  MUX2X1_536
timestamp 1516325494
transform -1 0 2403 0 -1 940
box 0 0 30 49
use AND2X2  AND2X2_1856
timestamp 1516325494
transform -1 0 2423 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1730
timestamp 1516325494
transform 1 0 2423 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_387
timestamp 1516325494
transform 1 0 2442 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_387
timestamp 1516325494
transform 1 0 2449 0 -1 940
box 0 0 15 49
use NAND2X1  NAND2X1_86
timestamp 1516325494
transform 1 0 2464 0 -1 940
box 0 0 15 49
use FILL  FILL_BUFX2_66
timestamp 1516325494
transform 1 0 2480 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_66
timestamp 1516325494
transform 1 0 2487 0 1 940
box 0 0 15 49
use FILL  FILL_BUFX2_646
timestamp 1516325494
transform 1 0 2502 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_646
timestamp 1516325494
transform 1 0 2510 0 1 940
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_390
timestamp 1516325494
transform 1 0 2525 0 1 940
box 0 0 53 49
use MUX2X1  MUX2X1_166
timestamp 1516325494
transform -1 0 2608 0 1 940
box 0 0 30 49
use AND2X2  AND2X2_1503
timestamp 1516325494
transform -1 0 2628 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1268
timestamp 1516325494
transform -1 0 2647 0 1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_649
timestamp 1516325494
transform 1 0 2647 0 1 940
box 0 0 53 49
use NAND2X1  NAND2X1_41
timestamp 1516325494
transform 1 0 2700 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_41
timestamp 1516325494
transform -1 0 2745 0 1 940
box 0 0 30 49
use MUX2X1  MUX2X1_86
timestamp 1516325494
transform -1 0 2510 0 -1 940
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_70
timestamp 1516325494
transform -1 0 2563 0 -1 940
box 0 0 53 49
use FILL  FILL_BUFX2_270
timestamp 1516325494
transform 1 0 2563 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_270
timestamp 1516325494
transform 1 0 2571 0 -1 940
box 0 0 15 49
use AND2X2  AND2X2_1436
timestamp 1516325494
transform -1 0 2605 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1183
timestamp 1516325494
transform -1 0 2624 0 -1 940
box 0 0 19 49
use NAND2X1  NAND2X1_166
timestamp 1516325494
transform 1 0 2624 0 -1 940
box 0 0 15 49
use AND2X2  AND2X2_1344
timestamp 1516325494
transform -1 0 2658 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_48
timestamp 1516325494
transform -1 0 2666 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_48
timestamp 1516325494
transform -1 0 2681 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1062
timestamp 1516325494
transform -1 0 2700 0 -1 940
box 0 0 19 49
use NAND2X1  NAND2X1_912
timestamp 1516325494
transform 1 0 2700 0 -1 940
box 0 0 15 49
use MUX2X1  MUX2X1_857
timestamp 1516325494
transform -1 0 2745 0 -1 940
box 0 0 30 49
use FILL  FILL_BUFX2_464
timestamp 1516325494
transform 1 0 2746 0 1 940
box 0 0 8 49
use BUFX2  BUFX2_464
timestamp 1516325494
transform 1 0 2753 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_598
timestamp 1516325494
transform 1 0 2768 0 1 940
box 0 0 30 49
use NAND2X1  NAND2X1_598
timestamp 1516325494
transform -1 0 2814 0 1 940
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_246
timestamp 1516325494
transform 1 0 2814 0 1 940
box 0 0 53 49
use MUX2X1  MUX2X1_214
timestamp 1516325494
transform 1 0 2867 0 1 940
box 0 0 30 49
use FILL  FILL_OR2X2_26
timestamp 1516325494
transform -1 0 2906 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_26
timestamp 1516325494
transform -1 0 2924 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_25
timestamp 1516325494
transform -1 0 2932 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_25
timestamp 1516325494
transform -1 0 2951 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_26
timestamp 1516325494
transform -1 0 2959 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_26
timestamp 1516325494
transform -1 0 2977 0 1 940
box 0 0 19 49
use OR2X2  OR2X2_1165
timestamp 1516325494
transform -1 0 2996 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1422
timestamp 1516325494
transform -1 0 3015 0 1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_166
timestamp 1516325494
transform 1 0 3015 0 1 940
box 0 0 53 49
use MUX2X1  MUX2X1_230
timestamp 1516325494
transform 1 0 3069 0 1 940
box 0 0 30 49
use NAND2X1  NAND2X1_230
timestamp 1516325494
transform 1 0 3099 0 1 940
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_236
timestamp 1516325494
transform -1 0 3167 0 1 940
box 0 0 53 49
use NAND2X1  NAND2X1_204
timestamp 1516325494
transform -1 0 3182 0 1 940
box 0 0 15 49
use FILL  FILL_AND2X2_117
timestamp 1516325494
transform 1 0 3183 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_117
timestamp 1516325494
transform 1 0 3190 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1561
timestamp 1516325494
transform 1 0 3209 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_220
timestamp 1516325494
transform 1 0 3228 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_220
timestamp 1516325494
transform 1 0 3236 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_111
timestamp 1516325494
transform 1 0 3255 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_111
timestamp 1516325494
transform 1 0 3262 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1721
timestamp 1516325494
transform 1 0 3281 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_208
timestamp 1516325494
transform 1 0 3300 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_208
timestamp 1516325494
transform 1 0 3308 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_118
timestamp 1516325494
transform -1 0 3335 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_118
timestamp 1516325494
transform -1 0 3354 0 1 940
box 0 0 19 49
use FILL  FILL_OR2X2_210
timestamp 1516325494
transform 1 0 3354 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_210
timestamp 1516325494
transform 1 0 3361 0 1 940
box 0 0 19 49
use NAND2X1  NAND2X1_588
timestamp 1516325494
transform 1 0 3380 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_588
timestamp 1516325494
transform -1 0 3425 0 1 940
box 0 0 30 49
use FILL  FILL_OR2X2_213
timestamp 1516325494
transform -1 0 3434 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_213
timestamp 1516325494
transform -1 0 3452 0 1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_137
timestamp 1516325494
transform -1 0 3505 0 1 940
box 0 0 53 49
use MUX2X1  MUX2X1_361
timestamp 1516325494
transform 1 0 3506 0 1 940
box 0 0 30 49
use NAND2X1  NAND2X1_361
timestamp 1516325494
transform -1 0 3551 0 1 940
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_329
timestamp 1516325494
transform -1 0 3604 0 1 940
box 0 0 53 49
use AND2X2  AND2X2_375
timestamp 1516325494
transform -1 0 3623 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1955
timestamp 1516325494
transform -1 0 3642 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_224
timestamp 1516325494
transform 1 0 3642 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_224
timestamp 1516325494
transform 1 0 3650 0 1 940
box 0 0 19 49
use NAND2X1  NAND2X1_381
timestamp 1516325494
transform 1 0 3669 0 1 940
box 0 0 15 49
use MUX2X1  MUX2X1_381
timestamp 1516325494
transform -1 0 3714 0 1 940
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_349
timestamp 1516325494
transform -1 0 3768 0 1 940
box 0 0 53 49
use FILL  FILL_OR2X2_29
timestamp 1516325494
transform -1 0 3776 0 1 940
box 0 0 8 49
use OR2X2  OR2X2_29
timestamp 1516325494
transform -1 0 3794 0 1 940
box 0 0 19 49
use AND2X2  AND2X2_1426
timestamp 1516325494
transform -1 0 3813 0 1 940
box 0 0 19 49
use FILL  FILL_AND2X2_30
timestamp 1516325494
transform 1 0 3813 0 1 940
box 0 0 8 49
use AND2X2  AND2X2_30
timestamp 1516325494
transform 1 0 3821 0 1 940
box 0 0 19 49
use MUX2X1  MUX2X1_262
timestamp 1516325494
transform 1 0 3840 0 1 940
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_354
timestamp 1516325494
transform -1 0 2799 0 -1 940
box 0 0 53 49
use OR2X2  OR2X2_1182
timestamp 1516325494
transform -1 0 2818 0 -1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_358
timestamp 1516325494
transform -1 0 2871 0 -1 940
box 0 0 53 49
use AND2X2  AND2X2_1792
timestamp 1516325494
transform -1 0 2890 0 -1 940
box 0 0 19 49
use NAND2X1  NAND2X1_214
timestamp 1516325494
transform -1 0 2905 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_255
timestamp 1516325494
transform -1 0 2924 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_252
timestamp 1516325494
transform -1 0 2943 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_251
timestamp 1516325494
transform -1 0 2962 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_268
timestamp 1516325494
transform -1 0 2981 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_267
timestamp 1516325494
transform -1 0 3000 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1791
timestamp 1516325494
transform -1 0 3019 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1421
timestamp 1516325494
transform -1 0 3038 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1857
timestamp 1516325494
transform 1 0 3038 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1860
timestamp 1516325494
transform -1 0 3076 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_558
timestamp 1516325494
transform 1 0 3076 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_558
timestamp 1516325494
transform 1 0 3084 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_350
timestamp 1516325494
transform 1 0 3099 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_353
timestamp 1516325494
transform -1 0 3137 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_204
timestamp 1516325494
transform 1 0 3137 0 -1 940
box 0 0 30 49
use FILL  FILL_BUFX2_525
timestamp 1516325494
transform -1 0 3175 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_525
timestamp 1516325494
transform -1 0 3190 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1347
timestamp 1516325494
transform -1 0 3209 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_664
timestamp 1516325494
transform -1 0 3217 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_664
timestamp 1516325494
transform -1 0 3232 0 -1 940
box 0 0 15 49
use AND2X2  AND2X2_1720
timestamp 1516325494
transform 1 0 3232 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1346
timestamp 1516325494
transform -1 0 3270 0 -1 940
box 0 0 19 49
use FILL  FILL_BUFX2_415
timestamp 1516325494
transform -1 0 3278 0 -1 940
box 0 0 8 49
use BUFX2  BUFX2_415
timestamp 1516325494
transform -1 0 3293 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_1555
timestamp 1516325494
transform 1 0 3293 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1557
timestamp 1516325494
transform 1 0 3312 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1562
timestamp 1516325494
transform -1 0 3350 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_352
timestamp 1516325494
transform -1 0 3369 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_374
timestamp 1516325494
transform -1 0 3388 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_254
timestamp 1516325494
transform -1 0 3407 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_269
timestamp 1516325494
transform -1 0 3426 0 -1 940
box 0 0 19 49
use FILL  FILL_AND2X2_119
timestamp 1516325494
transform -1 0 3434 0 -1 940
box 0 0 8 49
use AND2X2  AND2X2_119
timestamp 1516325494
transform -1 0 3452 0 -1 940
box 0 0 19 49
use MUX2X1  MUX2X1_278
timestamp 1516325494
transform 1 0 3452 0 -1 940
box 0 0 30 49
use NAND2X1  NAND2X1_278
timestamp 1516325494
transform -1 0 3498 0 -1 940
box 0 0 15 49
use OR2X2  OR2X2_253
timestamp 1516325494
transform -1 0 3517 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_270
timestamp 1516325494
transform -1 0 3536 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1859
timestamp 1516325494
transform -1 0 3555 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1954
timestamp 1516325494
transform -1 0 3574 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_351
timestamp 1516325494
transform -1 0 3593 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_376
timestamp 1516325494
transform -1 0 3612 0 -1 940
box 0 0 19 49
use OR2X2  OR2X2_1858
timestamp 1516325494
transform -1 0 3631 0 -1 940
box 0 0 19 49
use AND2X2  AND2X2_1956
timestamp 1516325494
transform -1 0 3650 0 -1 940
box 0 0 19 49
use FILL  FILL_OR2X2_212
timestamp 1516325494
transform -1 0 3658 0 -1 940
box 0 0 8 49
use OR2X2  OR2X2_212
timestamp 1516325494
transform -1 0 3677 0 -1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_140
timestamp 1516325494
transform -1 0 3730 0 -1 940
box 0 0 53 49
use FILL  FILL_OR2X2_211
timestamp 1516325494
transform -1 0 3738 0 -1 940
box 0 0 8 49
use OR2X2  OR2X2_211
timestamp 1516325494
transform -1 0 3756 0 -1 940
box 0 0 19 49
use FILL  FILL_AND2X2_31
timestamp 1516325494
transform 1 0 3756 0 -1 940
box 0 0 8 49
use AND2X2  AND2X2_31
timestamp 1516325494
transform 1 0 3764 0 -1 940
box 0 0 19 49
use FILL  FILL_AND2X2_225
timestamp 1516325494
transform -1 0 3791 0 -1 940
box 0 0 8 49
use AND2X2  AND2X2_225
timestamp 1516325494
transform -1 0 3810 0 -1 940
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_147
timestamp 1516325494
transform 1 0 3810 0 -1 940
box 0 0 53 49
use FILL  FILL_19_1
timestamp 1516325494
transform -1 0 3871 0 -1 940
box 0 0 8 49
use AND2X2  AND2X2_637
timestamp 1516325494
transform -1 0 21 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_536
timestamp 1516325494
transform 1 0 21 0 1 842
box 0 0 19 49
use NOR3X1  NOR3X1_6
timestamp 1516325494
transform 1 0 40 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_742
timestamp 1516325494
transform -1 0 78 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_765
timestamp 1516325494
transform -1 0 97 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_918
timestamp 1516325494
transform -1 0 116 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_959
timestamp 1516325494
transform 1 0 116 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_800
timestamp 1516325494
transform 1 0 135 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_962
timestamp 1516325494
transform -1 0 173 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1007
timestamp 1516325494
transform 1 0 173 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_493
timestamp 1516325494
transform -1 0 211 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_609
timestamp 1516325494
transform -1 0 230 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_727
timestamp 1516325494
transform -1 0 249 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_773
timestamp 1516325494
transform 1 0 249 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_648
timestamp 1516325494
transform 1 0 268 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_608
timestamp 1516325494
transform -1 0 306 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_576
timestamp 1516325494
transform -1 0 325 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_680
timestamp 1516325494
transform -1 0 344 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_978
timestamp 1516325494
transform 1 0 344 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_815
timestamp 1516325494
transform 1 0 363 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_557
timestamp 1516325494
transform -1 0 401 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_405
timestamp 1516325494
transform -1 0 420 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_686
timestamp 1516325494
transform 1 0 420 0 1 842
box 0 0 30 49
use AND2X2  AND2X2_659
timestamp 1516325494
transform -1 0 469 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1048
timestamp 1516325494
transform -1 0 488 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_665
timestamp 1516325494
transform -1 0 507 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_666
timestamp 1516325494
transform -1 0 526 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_462
timestamp 1516325494
transform 1 0 526 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_706
timestamp 1516325494
transform -1 0 575 0 1 842
box 0 0 30 49
use MUX2X1  MUX2X1_685
timestamp 1516325494
transform -1 0 606 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_597
timestamp 1516325494
transform -1 0 625 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_710
timestamp 1516325494
transform -1 0 644 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_482
timestamp 1516325494
transform -1 0 663 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_553
timestamp 1516325494
transform -1 0 682 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_556
timestamp 1516325494
transform -1 0 701 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_713
timestamp 1516325494
transform -1 0 720 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_693
timestamp 1516325494
transform -1 0 750 0 1 842
box 0 0 30 49
use FILL  FILL_BUFX2_668
timestamp 1516325494
transform 1 0 751 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_668
timestamp 1516325494
transform 1 0 758 0 1 842
box 0 0 15 49
use NAND3X1  NAND3X1_34
timestamp 1516325494
transform -1 0 792 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_753
timestamp 1516325494
transform -1 0 811 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_789
timestamp 1516325494
transform 1 0 811 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_666
timestamp 1516325494
transform -1 0 849 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_822
timestamp 1516325494
transform -1 0 868 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_823
timestamp 1516325494
transform -1 0 887 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_853
timestamp 1516325494
transform 1 0 887 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_854
timestamp 1516325494
transform -1 0 925 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_882
timestamp 1516325494
transform 1 0 925 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_740
timestamp 1516325494
transform 1 0 944 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_883
timestamp 1516325494
transform -1 0 982 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_927
timestamp 1516325494
transform -1 0 1001 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_721
timestamp 1516325494
transform 1 0 1001 0 1 842
box 0 0 30 49
use MUX2X1  MUX2X1_733
timestamp 1516325494
transform -1 0 1062 0 1 842
box 0 0 30 49
use MUX2X1  MUX2X1_736
timestamp 1516325494
transform -1 0 1092 0 1 842
box 0 0 30 49
use MUX2X1  MUX2X1_744
timestamp 1516325494
transform -1 0 1123 0 1 842
box 0 0 30 49
use INVX1  INVX1_163
timestamp 1516325494
transform 1 0 1123 0 1 842
box 0 0 11 49
use MUX2X1  MUX2X1_763
timestamp 1516325494
transform 1 0 1134 0 1 842
box 0 0 30 49
use MUX2X1  MUX2X1_806
timestamp 1516325494
transform -1 0 1195 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_1674
timestamp 1516325494
transform -1 0 1214 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_258
timestamp 1516325494
transform 1 0 1214 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1584
timestamp 1516325494
transform -1 0 1252 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_262
timestamp 1516325494
transform -1 0 1271 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_260
timestamp 1516325494
transform 1 0 1271 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_261
timestamp 1516325494
transform -1 0 1309 0 1 842
box 0 0 19 49
use INVX1  INVX1_228
timestamp 1516325494
transform -1 0 1320 0 1 842
box 0 0 11 49
use AND2X2  AND2X2_1498
timestamp 1516325494
transform -1 0 1340 0 1 842
box 0 0 19 49
use FILL  FILL_OR2X2_76
timestamp 1516325494
transform 1 0 1340 0 1 842
box 0 0 8 49
use OR2X2  OR2X2_76
timestamp 1516325494
transform 1 0 1347 0 1 842
box 0 0 19 49
use FILL  FILL_OR2X2_38
timestamp 1516325494
transform -1 0 1374 0 1 842
box 0 0 8 49
use OR2X2  OR2X2_38
timestamp 1516325494
transform -1 0 1393 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1666
timestamp 1516325494
transform -1 0 1412 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1805
timestamp 1516325494
transform -1 0 1431 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_259
timestamp 1516325494
transform -1 0 1450 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_276
timestamp 1516325494
transform -1 0 1469 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_277
timestamp 1516325494
transform -1 0 1488 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1807
timestamp 1516325494
transform -1 0 1507 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_360
timestamp 1516325494
transform 1 0 1507 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_361
timestamp 1516325494
transform -1 0 1545 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_359
timestamp 1516325494
transform -1 0 1564 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_358
timestamp 1516325494
transform -1 0 1583 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_383
timestamp 1516325494
transform -1 0 1602 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1970
timestamp 1516325494
transform -1 0 1621 0 1 842
box 0 0 19 49
use FILL  FILL_BUFX2_324
timestamp 1516325494
transform 1 0 1621 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_324
timestamp 1516325494
transform 1 0 1628 0 1 842
box 0 0 15 49
use OR2X2  OR2X2_357
timestamp 1516325494
transform -1 0 1663 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_381
timestamp 1516325494
transform -1 0 1682 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1966
timestamp 1516325494
transform -1 0 1701 0 1 842
box 0 0 19 49
use FILL  FILL_BUFX2_364
timestamp 1516325494
transform 1 0 1701 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_364
timestamp 1516325494
transform 1 0 1708 0 1 842
box 0 0 15 49
use OR2X2  OR2X2_1373
timestamp 1516325494
transform 1 0 1723 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1374
timestamp 1516325494
transform -1 0 1761 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1576
timestamp 1516325494
transform -1 0 1780 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1365
timestamp 1516325494
transform -1 0 1799 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1364
timestamp 1516325494
transform -1 0 1818 0 1 842
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_76
timestamp 1516325494
transform 1 0 1818 0 1 842
box 0 0 53 49
use NAND2X1  NAND2X1_140
timestamp 1516325494
transform 1 0 1872 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_140
timestamp 1516325494
transform -1 0 1917 0 1 842
box 0 0 30 49
use AND2X2  AND2X2_1806
timestamp 1516325494
transform -1 0 1936 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1665
timestamp 1516325494
transform -1 0 1955 0 1 842
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_86
timestamp 1516325494
transform 1 0 1955 0 1 842
box 0 0 53 49
use NAND2X1  NAND2X1_150
timestamp 1516325494
transform 1 0 2008 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_150
timestamp 1516325494
transform -1 0 2054 0 1 842
box 0 0 30 49
use FILL  FILL_BUFX2_460
timestamp 1516325494
transform 1 0 2054 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_460
timestamp 1516325494
transform 1 0 2062 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_884
timestamp 1516325494
transform 1 0 2077 0 1 842
box 0 0 30 49
use NAND2X1  NAND2X1_939
timestamp 1516325494
transform -1 0 2122 0 1 842
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_381
timestamp 1516325494
transform -1 0 2175 0 1 842
box 0 0 53 49
use OR2X2  OR2X2_1872
timestamp 1516325494
transform 1 0 2176 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1965
timestamp 1516325494
transform -1 0 2214 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_566
timestamp 1516325494
transform 1 0 2214 0 1 842
box 0 0 30 49
use NAND2X1  NAND2X1_566
timestamp 1516325494
transform -1 0 2259 0 1 842
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_502
timestamp 1516325494
transform -1 0 2312 0 1 842
box 0 0 53 49
use OR2X2  OR2X2_1669
timestamp 1516325494
transform 1 0 2312 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1810
timestamp 1516325494
transform -1 0 2350 0 1 842
box 0 0 19 49
use FILL  FILL_BUFX2_37
timestamp 1516325494
transform -1 0 2358 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_37
timestamp 1516325494
transform -1 0 2373 0 1 842
box 0 0 15 49
use OR2X2  OR2X2_1670
timestamp 1516325494
transform -1 0 2392 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1873
timestamp 1516325494
transform -1 0 2411 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1442
timestamp 1516325494
transform -1 0 2430 0 1 842
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_118
timestamp 1516325494
transform 1 0 2430 0 1 842
box 0 0 53 49
use NAND2X1  NAND2X1_134
timestamp 1516325494
transform 1 0 2483 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_134
timestamp 1516325494
transform 1 0 2499 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_1189
timestamp 1516325494
transform -1 0 2548 0 1 842
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_486
timestamp 1516325494
transform 1 0 2548 0 1 842
box 0 0 53 49
use NAND2X1  NAND2X1_550
timestamp 1516325494
transform 1 0 2601 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_550
timestamp 1516325494
transform -1 0 2646 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_1063
timestamp 1516325494
transform -1 0 2666 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_162
timestamp 1516325494
transform -1 0 2696 0 1 842
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_386
timestamp 1516325494
transform -1 0 2749 0 1 842
box 0 0 53 49
use MUX2X1  MUX2X1_861
timestamp 1516325494
transform -1 0 2779 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_1650
timestamp 1516325494
transform -1 0 2799 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1647
timestamp 1516325494
transform -1 0 2818 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1645
timestamp 1516325494
transform -1 0 2837 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1789
timestamp 1516325494
transform -1 0 2856 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1646
timestamp 1516325494
transform -1 0 2875 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1790
timestamp 1516325494
transform -1 0 2894 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_266
timestamp 1516325494
transform -1 0 2913 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_250
timestamp 1516325494
transform 1 0 2913 0 1 842
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_214
timestamp 1516325494
transform 1 0 2932 0 1 842
box 0 0 53 49
use NAND2X1  NAND2X1_630
timestamp 1516325494
transform 1 0 2985 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_630
timestamp 1516325494
transform -1 0 3030 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_1855
timestamp 1516325494
transform -1 0 3050 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1950
timestamp 1516325494
transform -1 0 3069 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_371
timestamp 1516325494
transform 1 0 3069 0 1 842
box 0 0 19 49
use NAND2X1  NAND2X1_637
timestamp 1516325494
transform 1 0 3088 0 1 842
box 0 0 15 49
use OR2X2  OR2X2_348
timestamp 1516325494
transform -1 0 3122 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_370
timestamp 1516325494
transform -1 0 3141 0 1 842
box 0 0 19 49
use NAND2X1  NAND2X1_253
timestamp 1516325494
transform 1 0 3141 0 1 842
box 0 0 15 49
use OR2X2  OR2X2_1350
timestamp 1516325494
transform -1 0 3175 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1560
timestamp 1516325494
transform 1 0 3175 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1345
timestamp 1516325494
transform -1 0 3213 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1559
timestamp 1516325494
transform -1 0 3232 0 1 842
box 0 0 19 49
use FILL  FILL_OR2X2_115
timestamp 1516325494
transform -1 0 3240 0 1 842
box 0 0 8 49
use OR2X2  OR2X2_115
timestamp 1516325494
transform -1 0 3259 0 1 842
box 0 0 19 49
use FILL  FILL_OR2X2_112
timestamp 1516325494
transform -1 0 3267 0 1 842
box 0 0 8 49
use OR2X2  OR2X2_112
timestamp 1516325494
transform -1 0 3285 0 1 842
box 0 0 19 49
use FILL  FILL_BUFX2_310
timestamp 1516325494
transform -1 0 3293 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_310
timestamp 1516325494
transform -1 0 3308 0 1 842
box 0 0 15 49
use OR2X2  OR2X2_1560
timestamp 1516325494
transform -1 0 3327 0 1 842
box 0 0 19 49
use NAND2X1  NAND2X1_236
timestamp 1516325494
transform 1 0 3327 0 1 842
box 0 0 15 49
use MUX2X1  MUX2X1_236
timestamp 1516325494
transform -1 0 3372 0 1 842
box 0 0 30 49
use OR2X2  OR2X2_1349
timestamp 1516325494
transform -1 0 3392 0 1 842
box 0 0 19 49
use FILL  FILL_OR2X2_114
timestamp 1516325494
transform -1 0 3400 0 1 842
box 0 0 8 49
use OR2X2  OR2X2_114
timestamp 1516325494
transform -1 0 3418 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1495
timestamp 1516325494
transform -1 0 3437 0 1 842
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_150
timestamp 1516325494
transform -1 0 3490 0 1 842
box 0 0 53 49
use AND2X2  AND2X2_271
timestamp 1516325494
transform -1 0 3509 0 1 842
box 0 0 19 49
use FILL  FILL_AND2X2_75
timestamp 1516325494
transform -1 0 3517 0 1 842
box 0 0 8 49
use AND2X2  AND2X2_75
timestamp 1516325494
transform -1 0 3536 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1559
timestamp 1516325494
transform -1 0 3555 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1724
timestamp 1516325494
transform -1 0 3574 0 1 842
box 0 0 19 49
use FILL  FILL_AND2X2_120
timestamp 1516325494
transform -1 0 3582 0 1 842
box 0 0 8 49
use AND2X2  AND2X2_120
timestamp 1516325494
transform -1 0 3601 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1348
timestamp 1516325494
transform -1 0 3620 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1565
timestamp 1516325494
transform -1 0 3639 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1564
timestamp 1516325494
transform -1 0 3658 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_268
timestamp 1516325494
transform 1 0 3658 0 1 842
box 0 0 30 49
use NAND2X1  NAND2X1_268
timestamp 1516325494
transform -1 0 3703 0 1 842
box 0 0 15 49
use FILL  FILL_BUFX2_832
timestamp 1516325494
transform 1 0 3703 0 1 842
box 0 0 8 49
use BUFX2  BUFX2_832
timestamp 1516325494
transform 1 0 3711 0 1 842
box 0 0 15 49
use FILL  FILL_AND2X2_226
timestamp 1516325494
transform 1 0 3726 0 1 842
box 0 0 8 49
use AND2X2  AND2X2_226
timestamp 1516325494
transform 1 0 3734 0 1 842
box 0 0 19 49
use OR2X2  OR2X2_1558
timestamp 1516325494
transform -1 0 3772 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1726
timestamp 1516325494
transform -1 0 3791 0 1 842
box 0 0 19 49
use AND2X2  AND2X2_1725
timestamp 1516325494
transform -1 0 3810 0 1 842
box 0 0 19 49
use MUX2X1  MUX2X1_371
timestamp 1516325494
transform 1 0 3810 0 1 842
box 0 0 30 49
use NAND2X1  NAND2X1_371
timestamp 1516325494
transform -1 0 3855 0 1 842
box 0 0 15 49
use INVX1  INVX1_255
timestamp 1516325494
transform -1 0 3866 0 1 842
box 0 0 11 49
use FILL  FILL_BUFX2_671
timestamp 1516325494
transform -1 0 10 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_671
timestamp 1516325494
transform -1 0 25 0 -1 841
box 0 0 15 49
use OR2X2  OR2X2_535
timestamp 1516325494
transform -1 0 44 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_636
timestamp 1516325494
transform -1 0 63 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_758
timestamp 1516325494
transform 1 0 63 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_758
timestamp 1516325494
transform 1 0 70 0 -1 841
box 0 0 15 49
use AND2X2  AND2X2_806
timestamp 1516325494
transform -1 0 105 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_734
timestamp 1516325494
transform -1 0 124 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_870
timestamp 1516325494
transform -1 0 143 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_526
timestamp 1516325494
transform -1 0 162 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_621
timestamp 1516325494
transform -1 0 181 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_441
timestamp 1516325494
transform 1 0 181 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_726
timestamp 1516325494
transform -1 0 219 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_784
timestamp 1516325494
transform -1 0 238 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_939
timestamp 1516325494
transform -1 0 257 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_799
timestamp 1516325494
transform -1 0 276 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_960
timestamp 1516325494
transform -1 0 295 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_961
timestamp 1516325494
transform -1 0 314 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_681
timestamp 1516325494
transform -1 0 333 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_75
timestamp 1516325494
transform 1 0 333 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_75
timestamp 1516325494
transform 1 0 340 0 -1 841
box 0 0 15 49
use AND2X2  AND2X2_979
timestamp 1516325494
transform -1 0 374 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_834
timestamp 1516325494
transform -1 0 393 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1004
timestamp 1516325494
transform -1 0 412 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_672
timestamp 1516325494
transform -1 0 442 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_699
timestamp 1516325494
transform 1 0 443 0 -1 841
box 0 0 30 49
use OR2X2  OR2X2_421
timestamp 1516325494
transform -1 0 492 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_455
timestamp 1516325494
transform -1 0 511 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_671
timestamp 1516325494
transform 1 0 511 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_741
timestamp 1516325494
transform -1 0 572 0 -1 841
box 0 0 30 49
use OR2X2  OR2X2_855
timestamp 1516325494
transform -1 0 591 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1028
timestamp 1516325494
transform 1 0 591 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1005
timestamp 1516325494
transform -1 0 629 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1029
timestamp 1516325494
transform -1 0 648 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_732
timestamp 1516325494
transform -1 0 678 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_734
timestamp 1516325494
transform -1 0 708 0 -1 841
box 0 0 30 49
use FILL  FILL_BUFX2_79
timestamp 1516325494
transform -1 0 717 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_79
timestamp 1516325494
transform -1 0 731 0 -1 841
box 0 0 15 49
use OR2X2  OR2X2_484
timestamp 1516325494
transform -1 0 751 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_559
timestamp 1516325494
transform -1 0 770 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_729
timestamp 1516325494
transform -1 0 800 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_708
timestamp 1516325494
transform -1 0 830 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_642
timestamp 1516325494
transform 1 0 830 0 -1 841
box 0 0 30 49
use AND2X2  AND2X2_790
timestamp 1516325494
transform -1 0 880 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_710
timestamp 1516325494
transform -1 0 910 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_714
timestamp 1516325494
transform -1 0 940 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_644
timestamp 1516325494
transform -1 0 971 0 -1 841
box 0 0 30 49
use AND2X2  AND2X2_902
timestamp 1516325494
transform 1 0 971 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_755
timestamp 1516325494
transform -1 0 1009 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_903
timestamp 1516325494
transform -1 0 1028 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_743
timestamp 1516325494
transform -1 0 1058 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_735
timestamp 1516325494
transform 1 0 1058 0 -1 841
box 0 0 30 49
use OR2X2  OR2X2_1673
timestamp 1516325494
transform -1 0 1108 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1661
timestamp 1516325494
transform -1 0 1127 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1672
timestamp 1516325494
transform -1 0 1146 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1671
timestamp 1516325494
transform -1 0 1165 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1811
timestamp 1516325494
transform -1 0 1184 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_606
timestamp 1516325494
transform 1 0 1184 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_606
timestamp 1516325494
transform 1 0 1191 0 -1 841
box 0 0 15 49
use AND2X2  AND2X2_279
timestamp 1516325494
transform 1 0 1207 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_78
timestamp 1516325494
transform -1 0 1234 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_78
timestamp 1516325494
transform -1 0 1252 0 -1 841
box 0 0 19 49
use FILL  FILL_OR2X2_74
timestamp 1516325494
transform 1 0 1252 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_74
timestamp 1516325494
transform 1 0 1260 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_99
timestamp 1516325494
transform -1 0 1287 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_99
timestamp 1516325494
transform -1 0 1305 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_590
timestamp 1516325494
transform 1 0 1305 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_590
timestamp 1516325494
transform 1 0 1313 0 -1 841
box 0 0 15 49
use AND2X2  AND2X2_1535
timestamp 1516325494
transform -1 0 1347 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_331
timestamp 1516325494
transform 1 0 1347 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_331
timestamp 1516325494
transform 1 0 1355 0 -1 841
box 0 0 15 49
use FILL  FILL_BUFX2_96
timestamp 1516325494
transform -1 0 1378 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_96
timestamp 1516325494
transform -1 0 1393 0 -1 841
box 0 0 15 49
use FILL  FILL_OR2X2_37
timestamp 1516325494
transform -1 0 1401 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_37
timestamp 1516325494
transform -1 0 1419 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1857
timestamp 1516325494
transform -1 0 1438 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_309
timestamp 1516325494
transform -1 0 1457 0 -1 841
box 0 0 19 49
use FILL  FILL_OR2X2_36
timestamp 1516325494
transform -1 0 1465 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_36
timestamp 1516325494
transform -1 0 1484 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_39
timestamp 1516325494
transform -1 0 1492 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_39
timestamp 1516325494
transform -1 0 1511 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1443
timestamp 1516325494
transform 1 0 1511 0 -1 841
box 0 0 19 49
use FILL  FILL_OR2X2_35
timestamp 1516325494
transform -1 0 1538 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_35
timestamp 1516325494
transform -1 0 1556 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_37
timestamp 1516325494
transform -1 0 1564 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_37
timestamp 1516325494
transform -1 0 1583 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1186
timestamp 1516325494
transform -1 0 1602 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1439
timestamp 1516325494
transform -1 0 1621 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1437
timestamp 1516325494
transform -1 0 1640 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_36
timestamp 1516325494
transform -1 0 1648 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_36
timestamp 1516325494
transform -1 0 1666 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1804
timestamp 1516325494
transform -1 0 1685 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1663
timestamp 1516325494
transform -1 0 1704 0 -1 841
box 0 0 19 49
use MUX2X1  MUX2X1_108
timestamp 1516325494
transform 1 0 1704 0 -1 841
box 0 0 30 49
use NAND2X1  NAND2X1_108
timestamp 1516325494
transform -1 0 1750 0 -1 841
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_12
timestamp 1516325494
transform -1 0 1803 0 -1 841
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_406
timestamp 1516325494
transform 1 0 1803 0 -1 841
box 0 0 53 49
use NAND2X1  NAND2X1_332
timestamp 1516325494
transform 1 0 1856 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_332
timestamp 1516325494
transform 1 0 1872 0 -1 841
box 0 0 30 49
use NAND2X1  NAND2X1_182
timestamp 1516325494
transform 1 0 1902 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_182
timestamp 1516325494
transform 1 0 1917 0 -1 841
box 0 0 30 49
use AND2X2  AND2X2_630
timestamp 1516325494
transform 1 0 2 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_741
timestamp 1516325494
transform -1 0 40 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_439
timestamp 1516325494
transform -1 0 59 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_578
timestamp 1516325494
transform -1 0 78 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_687
timestamp 1516325494
transform -1 0 97 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_915
timestamp 1516325494
transform -1 0 116 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_873
timestamp 1516325494
transform 1 0 116 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_492
timestamp 1516325494
transform 1 0 135 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_764
timestamp 1516325494
transform -1 0 173 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_917
timestamp 1516325494
transform -1 0 192 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_620
timestamp 1516325494
transform -1 0 211 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_679
timestamp 1516325494
transform -1 0 230 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_938
timestamp 1516325494
transform -1 0 249 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_804
timestamp 1516325494
transform -1 0 268 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_774
timestamp 1516325494
transform -1 0 287 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_541
timestamp 1516325494
transform -1 0 295 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_541
timestamp 1516325494
transform -1 0 310 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_740
timestamp 1516325494
transform -1 0 340 0 1 743
box 0 0 30 49
use MUX2X1  MUX2X1_739
timestamp 1516325494
transform -1 0 370 0 1 743
box 0 0 30 49
use AND2X2  AND2X2_656
timestamp 1516325494
transform 1 0 371 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_471
timestamp 1516325494
transform 1 0 390 0 1 743
box 0 0 19 49
use NAND2X1  NAND2X1_641
timestamp 1516325494
transform 1 0 409 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_722
timestamp 1516325494
transform -1 0 454 0 1 743
box 0 0 30 49
use OR2X2  OR2X2_642
timestamp 1516325494
transform -1 0 473 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_377
timestamp 1516325494
transform 1 0 473 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_377
timestamp 1516325494
transform 1 0 481 0 1 743
box 0 0 15 49
use OR2X2  OR2X2_556
timestamp 1516325494
transform -1 0 515 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_452
timestamp 1516325494
transform -1 0 534 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_575
timestamp 1516325494
transform -1 0 553 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_678
timestamp 1516325494
transform 1 0 553 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_574
timestamp 1516325494
transform -1 0 591 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_596
timestamp 1516325494
transform 1 0 591 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_709
timestamp 1516325494
transform 1 0 610 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_627
timestamp 1516325494
transform 1 0 629 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_688
timestamp 1516325494
transform -1 0 667 0 1 743
box 0 0 19 49
use MUX2X1  MUX2X1_709
timestamp 1516325494
transform -1 0 697 0 1 743
box 0 0 30 49
use OR2X2  OR2X2_512
timestamp 1516325494
transform -1 0 716 0 1 743
box 0 0 19 49
use MUX2X1  MUX2X1_725
timestamp 1516325494
transform -1 0 746 0 1 743
box 0 0 30 49
use AND2X2  AND2X2_457
timestamp 1516325494
transform -1 0 766 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_420
timestamp 1516325494
transform -1 0 785 0 1 743
box 0 0 19 49
use INVX1  INVX1_22
timestamp 1516325494
transform 1 0 785 0 1 743
box 0 0 11 49
use AND2X2  AND2X2_560
timestamp 1516325494
transform -1 0 815 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_546
timestamp 1516325494
transform 1 0 815 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_546
timestamp 1516325494
transform 1 0 823 0 1 743
box 0 0 15 49
use OR2X2  OR2X2_423
timestamp 1516325494
transform -1 0 857 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_461
timestamp 1516325494
transform -1 0 876 0 1 743
box 0 0 19 49
use MUX2X1  MUX2X1_712
timestamp 1516325494
transform -1 0 906 0 1 743
box 0 0 30 49
use OR2X2  OR2X2_481
timestamp 1516325494
transform -1 0 925 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_554
timestamp 1516325494
transform -1 0 944 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_547
timestamp 1516325494
transform -1 0 952 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_547
timestamp 1516325494
transform -1 0 967 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_716
timestamp 1516325494
transform -1 0 997 0 1 743
box 0 0 30 49
use FILL  FILL_BUFX2_374
timestamp 1516325494
transform 1 0 998 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_374
timestamp 1516325494
transform 1 0 1005 0 1 743
box 0 0 15 49
use INVX1  INVX1_151
timestamp 1516325494
transform -1 0 1031 0 1 743
box 0 0 11 49
use FILL  FILL_BUFX2_372
timestamp 1516325494
transform 1 0 1032 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_372
timestamp 1516325494
transform 1 0 1039 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_72
timestamp 1516325494
transform 1 0 1055 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_72
timestamp 1516325494
transform 1 0 1062 0 1 743
box 0 0 15 49
use OAI21X1  OAI21X1_53
timestamp 1516325494
transform 1 0 1077 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1660
timestamp 1516325494
transform 1 0 1096 0 1 743
box 0 0 19 49
use INVX1  INVX1_145
timestamp 1516325494
transform -1 0 1126 0 1 743
box 0 0 11 49
use AND2X2  AND2X2_1801
timestamp 1516325494
transform -1 0 1146 0 1 743
box 0 0 19 49
use INVX1  INVX1_167
timestamp 1516325494
transform 1 0 1146 0 1 743
box 0 0 11 49
use OAI21X1  OAI21X1_51
timestamp 1516325494
transform 1 0 1157 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1809
timestamp 1516325494
transform -1 0 1195 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_333
timestamp 1516325494
transform 1 0 1195 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_333
timestamp 1516325494
transform 1 0 1203 0 1 743
box 0 0 15 49
use AND2X2  AND2X2_278
timestamp 1516325494
transform 1 0 1218 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_286
timestamp 1516325494
transform 1 0 1237 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_286
timestamp 1516325494
transform 1 0 1245 0 1 743
box 0 0 15 49
use FILL  FILL_OR2X2_92
timestamp 1516325494
transform -1 0 1268 0 1 743
box 0 0 8 49
use OR2X2  OR2X2_92
timestamp 1516325494
transform -1 0 1286 0 1 743
box 0 0 19 49
use FILL  FILL_AND2X2_77
timestamp 1516325494
transform -1 0 1294 0 1 743
box 0 0 8 49
use AND2X2  AND2X2_77
timestamp 1516325494
transform -1 0 1313 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1311
timestamp 1516325494
transform -1 0 1332 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1533
timestamp 1516325494
transform -1 0 1351 0 1 743
box 0 0 19 49
use FILL  FILL_AND2X2_98
timestamp 1516325494
transform -1 0 1359 0 1 743
box 0 0 8 49
use AND2X2  AND2X2_98
timestamp 1516325494
transform -1 0 1378 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1732
timestamp 1516325494
transform -1 0 1397 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1731
timestamp 1516325494
transform -1 0 1416 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1855
timestamp 1516325494
transform -1 0 1435 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_288
timestamp 1516325494
transform -1 0 1454 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_308
timestamp 1516325494
transform -1 0 1473 0 1 743
box 0 0 19 49
use FILL  FILL_AND2X2_38
timestamp 1516325494
transform -1 0 1481 0 1 743
box 0 0 8 49
use AND2X2  AND2X2_38
timestamp 1516325494
transform -1 0 1499 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1441
timestamp 1516325494
transform 1 0 1499 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1191
timestamp 1516325494
transform 1 0 1518 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1192
timestamp 1516325494
transform 1 0 1537 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1193
timestamp 1516325494
transform 1 0 1556 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_363
timestamp 1516325494
transform 1 0 1575 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_363
timestamp 1516325494
transform 1 0 1583 0 1 743
box 0 0 15 49
use AND2X2  AND2X2_1808
timestamp 1516325494
transform -1 0 1617 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_285
timestamp 1516325494
transform -1 0 1625 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_285
timestamp 1516325494
transform -1 0 1640 0 1 743
box 0 0 15 49
use OAI21X1  OAI21X1_50
timestamp 1516325494
transform 1 0 1640 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1668
timestamp 1516325494
transform -1 0 1678 0 1 743
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_22
timestamp 1516325494
transform 1 0 1678 0 1 743
box 0 0 53 49
use NAND2X1  NAND2X1_118
timestamp 1516325494
transform 1 0 1731 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_118
timestamp 1516325494
transform -1 0 1776 0 1 743
box 0 0 30 49
use OR2X2  OR2X2_1662
timestamp 1516325494
transform -1 0 1796 0 1 743
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_374
timestamp 1516325494
transform 1 0 1796 0 1 743
box 0 0 53 49
use NAND2X1  NAND2X1_932
timestamp 1516325494
transform 1 0 1849 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_877
timestamp 1516325494
transform -1 0 1894 0 1 743
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_460
timestamp 1516325494
transform -1 0 1947 0 1 743
box 0 0 53 49
use AND2X2  AND2X2_1969
timestamp 1516325494
transform -1 0 1967 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1877
timestamp 1516325494
transform -1 0 1986 0 -1 841
box 0 0 19 49
use NAND2X1  NAND2X1_541
timestamp 1516325494
transform 1 0 1986 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_541
timestamp 1516325494
transform -1 0 2031 0 -1 841
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_541
timestamp 1516325494
transform -1 0 2084 0 -1 841
box 0 0 53 49
use FILL  FILL_BUFX2_462
timestamp 1516325494
transform -1 0 2092 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_462
timestamp 1516325494
transform -1 0 2107 0 -1 841
box 0 0 15 49
use OR2X2  OR2X2_1878
timestamp 1516325494
transform -1 0 2126 0 -1 841
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_29
timestamp 1516325494
transform 1 0 2126 0 -1 841
box 0 0 53 49
use NAND2X1  NAND2X1_125
timestamp 1516325494
transform 1 0 2179 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_125
timestamp 1516325494
transform -1 0 2225 0 -1 841
box 0 0 30 49
use AND2X2  AND2X2_1438
timestamp 1516325494
transform -1 0 2244 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1854
timestamp 1516325494
transform -1 0 2263 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1728
timestamp 1516325494
transform -1 0 2282 0 -1 841
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_24
timestamp 1516325494
transform 1 0 2282 0 -1 841
box 0 0 53 49
use NAND2X1  NAND2X1_120
timestamp 1516325494
transform 1 0 2335 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_120
timestamp 1516325494
transform -1 0 2380 0 -1 841
box 0 0 30 49
use NAND2X1  NAND2X1_457
timestamp 1516325494
transform 1 0 2381 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_457
timestamp 1516325494
transform -1 0 2426 0 -1 841
box 0 0 30 49
use AND2X2  AND2X2_1534
timestamp 1516325494
transform -1 0 2445 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_739
timestamp 1516325494
transform -1 0 2453 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_739
timestamp 1516325494
transform -1 0 2468 0 -1 841
box 0 0 15 49
use OR2X2  OR2X2_1185
timestamp 1516325494
transform -1 0 2487 0 -1 841
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_413
timestamp 1516325494
transform 1 0 2487 0 -1 841
box 0 0 53 49
use NAND2X1  NAND2X1_189
timestamp 1516325494
transform 1 0 2540 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_189
timestamp 1516325494
transform -1 0 2586 0 -1 841
box 0 0 30 49
use FILL  FILL_BUFX2_390
timestamp 1516325494
transform 1 0 2586 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_390
timestamp 1516325494
transform 1 0 2594 0 -1 841
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_106
timestamp 1516325494
transform -1 0 2662 0 -1 841
box 0 0 53 49
use OR2X2  OR2X2_1309
timestamp 1516325494
transform -1 0 2681 0 -1 841
box 0 0 19 49
use NAND2X1  NAND2X1_162
timestamp 1516325494
transform -1 0 2696 0 -1 841
box 0 0 15 49
use NAND2X1  NAND2X1_554
timestamp 1516325494
transform 1 0 2696 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_554
timestamp 1516325494
transform -1 0 2741 0 -1 841
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_490
timestamp 1516325494
transform -1 0 2795 0 -1 841
box 0 0 53 49
use NAND2X1  NAND2X1_916
timestamp 1516325494
transform -1 0 2810 0 -1 841
box 0 0 15 49
use FILL  FILL_BUFX2_791
timestamp 1516325494
transform -1 0 2818 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_791
timestamp 1516325494
transform -1 0 2833 0 -1 841
box 0 0 15 49
use MUX2X1  MUX2X1_233
timestamp 1516325494
transform 1 0 2833 0 -1 841
box 0 0 30 49
use NAND2X1  NAND2X1_233
timestamp 1516325494
transform -1 0 2878 0 -1 841
box 0 0 15 49
use AND2X2  AND2X2_1490
timestamp 1516325494
transform -1 0 2898 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_70
timestamp 1516325494
transform -1 0 2906 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_70
timestamp 1516325494
transform -1 0 2924 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_265
timestamp 1516325494
transform -1 0 2943 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1260
timestamp 1516325494
transform -1 0 2962 0 -1 841
box 0 0 19 49
use FILL  FILL_BUFX2_774
timestamp 1516325494
transform -1 0 2970 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_774
timestamp 1516325494
transform -1 0 2985 0 -1 841
box 0 0 15 49
use FILL  FILL_BUFX2_703
timestamp 1516325494
transform 1 0 2985 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_703
timestamp 1516325494
transform 1 0 2993 0 -1 841
box 0 0 15 49
use FILL  FILL_BUFX2_459
timestamp 1516325494
transform 1 0 3008 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_459
timestamp 1516325494
transform 1 0 3015 0 -1 841
box 0 0 15 49
use AND2X2  AND2X2_1951
timestamp 1516325494
transform 1 0 3031 0 -1 841
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_221
timestamp 1516325494
transform 1 0 3050 0 -1 841
box 0 0 53 49
use MUX2X1  MUX2X1_637
timestamp 1516325494
transform -1 0 3133 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_253
timestamp 1516325494
transform 1 0 3133 0 -1 841
box 0 0 30 49
use MUX2X1  MUX2X1_620
timestamp 1516325494
transform 1 0 3164 0 -1 841
box 0 0 30 49
use NAND2X1  NAND2X1_620
timestamp 1516325494
transform -1 0 3209 0 -1 841
box 0 0 15 49
use FILL  FILL_AND2X2_116
timestamp 1516325494
transform 1 0 3209 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_116
timestamp 1516325494
transform 1 0 3217 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_115
timestamp 1516325494
transform 1 0 3236 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_115
timestamp 1516325494
transform 1 0 3243 0 -1 841
box 0 0 19 49
use FILL  FILL_OR2X2_110
timestamp 1516325494
transform 1 0 3262 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_110
timestamp 1516325494
transform 1 0 3270 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1259
timestamp 1516325494
transform -1 0 3308 0 -1 841
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_172
timestamp 1516325494
transform 1 0 3308 0 -1 841
box 0 0 53 49
use OR2X2  OR2X2_1649
timestamp 1516325494
transform -1 0 3380 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1563
timestamp 1516325494
transform -1 0 3399 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1258
timestamp 1516325494
transform -1 0 3418 0 -1 841
box 0 0 19 49
use OR2X2  OR2X2_1648
timestamp 1516325494
transform -1 0 3437 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1795
timestamp 1516325494
transform -1 0 3456 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1794
timestamp 1516325494
transform -1 0 3475 0 -1 841
box 0 0 19 49
use AND2X2  AND2X2_1496
timestamp 1516325494
transform -1 0 3494 0 -1 841
box 0 0 19 49
use FILL  FILL_OR2X2_71
timestamp 1516325494
transform -1 0 3502 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_71
timestamp 1516325494
transform -1 0 3521 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_76
timestamp 1516325494
transform -1 0 3529 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_76
timestamp 1516325494
transform -1 0 3547 0 -1 841
box 0 0 19 49
use FILL  FILL_OR2X2_113
timestamp 1516325494
transform -1 0 3555 0 -1 841
box 0 0 8 49
use OR2X2  OR2X2_113
timestamp 1516325494
transform -1 0 3574 0 -1 841
box 0 0 19 49
use FILL  FILL_AND2X2_121
timestamp 1516325494
transform -1 0 3582 0 -1 841
box 0 0 8 49
use AND2X2  AND2X2_121
timestamp 1516325494
transform -1 0 3601 0 -1 841
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_332
timestamp 1516325494
transform -1 0 3654 0 -1 841
box 0 0 53 49
use FILL  FILL_BUFX2_330
timestamp 1516325494
transform -1 0 3662 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_330
timestamp 1516325494
transform -1 0 3676 0 -1 841
box 0 0 15 49
use FILL  FILL_BUFX2_157
timestamp 1516325494
transform -1 0 3685 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_157
timestamp 1516325494
transform -1 0 3699 0 -1 841
box 0 0 15 49
use FILL  FILL_BUFX2_447
timestamp 1516325494
transform 1 0 3699 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_447
timestamp 1516325494
transform 1 0 3707 0 -1 841
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_331
timestamp 1516325494
transform -1 0 3775 0 -1 841
box 0 0 53 49
use FILL  FILL_BUFX2_423
timestamp 1516325494
transform -1 0 3783 0 -1 841
box 0 0 8 49
use BUFX2  BUFX2_423
timestamp 1516325494
transform -1 0 3798 0 -1 841
box 0 0 15 49
use NAND2X1  NAND2X1_275
timestamp 1516325494
transform 1 0 3798 0 -1 841
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_339
timestamp 1516325494
transform -1 0 3866 0 -1 841
box 0 0 53 49
use AND2X2  AND2X2_1499
timestamp 1516325494
transform 1 0 1948 0 1 743
box 0 0 19 49
use MUX2X1  MUX2X1_29
timestamp 1516325494
transform -1 0 1997 0 1 743
box 0 0 30 49
use FILL  FILL_BUFX2_480
timestamp 1516325494
transform 1 0 1997 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_480
timestamp 1516325494
transform 1 0 2005 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_269
timestamp 1516325494
transform 1 0 2020 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_269
timestamp 1516325494
transform 1 0 2027 0 1 743
box 0 0 15 49
use OR2X2  OR2X2_1263
timestamp 1516325494
transform -1 0 2062 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2074
timestamp 1516325494
transform -1 0 2081 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2076
timestamp 1516325494
transform -1 0 2100 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2072
timestamp 1516325494
transform -1 0 2119 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_495
timestamp 1516325494
transform -1 0 2127 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_495
timestamp 1516325494
transform -1 0 2141 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_198
timestamp 1516325494
transform 1 0 2141 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_198
timestamp 1516325494
transform 1 0 2149 0 1 743
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_454
timestamp 1516325494
transform -1 0 2217 0 1 743
box 0 0 53 49
use NAND2X1  NAND2X1_326
timestamp 1516325494
transform -1 0 2232 0 1 743
box 0 0 15 49
use OR2X2  OR2X2_1184
timestamp 1516325494
transform -1 0 2252 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1326
timestamp 1516325494
transform -1 0 2271 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1323
timestamp 1516325494
transform -1 0 2290 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1320
timestamp 1516325494
transform -1 0 2309 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1317
timestamp 1516325494
transform -1 0 2328 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_812
timestamp 1516325494
transform -1 0 2336 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_812
timestamp 1516325494
transform -1 0 2350 0 1 743
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_553
timestamp 1516325494
transform 1 0 2350 0 1 743
box 0 0 53 49
use FILL  FILL_BUFX2_186
timestamp 1516325494
transform -1 0 2412 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_186
timestamp 1516325494
transform -1 0 2426 0 1 743
box 0 0 15 49
use OR2X2  OR2X2_1310
timestamp 1516325494
transform 1 0 2426 0 1 743
box 0 0 19 49
use NAND2X1  NAND2X1_522
timestamp 1516325494
transform 1 0 2445 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_128
timestamp 1516325494
transform -1 0 2469 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_128
timestamp 1516325494
transform -1 0 2483 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_67
timestamp 1516325494
transform -1 0 2491 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_67
timestamp 1516325494
transform -1 0 2506 0 1 743
box 0 0 15 49
use NAND2X1  NAND2X1_74
timestamp 1516325494
transform 1 0 2506 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_74
timestamp 1516325494
transform -1 0 2551 0 1 743
box 0 0 30 49
use AND2X2  AND2X2_1316
timestamp 1516325494
transform -1 0 2571 0 1 743
box 0 0 19 49
use INVX1  INVX1_326
timestamp 1516325494
transform -1 0 2582 0 1 743
box 0 0 11 49
use FILL  FILL_BUFX2_272
timestamp 1516325494
transform -1 0 2590 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_272
timestamp 1516325494
transform -1 0 2605 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_493
timestamp 1516325494
transform -1 0 2613 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_493
timestamp 1516325494
transform -1 0 2628 0 1 743
box 0 0 15 49
use OR2X2  OR2X2_1269
timestamp 1516325494
transform -1 0 2647 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_475
timestamp 1516325494
transform 1 0 2647 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_475
timestamp 1516325494
transform 1 0 2654 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_201
timestamp 1516325494
transform 1 0 2670 0 1 743
box 0 0 30 49
use NAND2X1  NAND2X1_201
timestamp 1516325494
transform -1 0 2715 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_271
timestamp 1516325494
transform -1 0 2723 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_271
timestamp 1516325494
transform -1 0 2738 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_246
timestamp 1516325494
transform 1 0 2738 0 1 743
box 0 0 30 49
use NAND2X1  NAND2X1_246
timestamp 1516325494
transform -1 0 2783 0 1 743
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_169
timestamp 1516325494
transform 1 0 2784 0 1 743
box 0 0 53 49
use OR2X2  OR2X2_1255
timestamp 1516325494
transform 1 0 2837 0 1 743
box 0 0 19 49
use OR2X2  OR2X2_1257
timestamp 1516325494
transform 1 0 2856 0 1 743
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_182
timestamp 1516325494
transform -1 0 2928 0 1 743
box 0 0 53 49
use INVX1  INVX1_327
timestamp 1516325494
transform -1 0 2939 0 1 743
box 0 0 11 49
use AND2X2  AND2X2_2049
timestamp 1516325494
transform 1 0 2939 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2052
timestamp 1516325494
transform -1 0 2977 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2046
timestamp 1516325494
transform 1 0 2977 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1295
timestamp 1516325494
transform -1 0 3015 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1286
timestamp 1516325494
transform 1 0 3015 0 1 743
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_189
timestamp 1516325494
transform 1 0 3034 0 1 743
box 0 0 53 49
use AND2X2  AND2X2_1292
timestamp 1516325494
transform 1 0 3088 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_602
timestamp 1516325494
transform 1 0 3107 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_602
timestamp 1516325494
transform 1 0 3114 0 1 743
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_204
timestamp 1516325494
transform 1 0 3129 0 1 743
box 0 0 53 49
use AND2X2  AND2X2_1297
timestamp 1516325494
transform 1 0 3183 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1301
timestamp 1516325494
transform -1 0 3221 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1299
timestamp 1516325494
transform 1 0 3221 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_767
timestamp 1516325494
transform -1 0 3248 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_767
timestamp 1516325494
transform -1 0 3262 0 1 743
box 0 0 15 49
use AND2X2  AND2X2_1678
timestamp 1516325494
transform -1 0 3281 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1494
timestamp 1516325494
transform 1 0 3281 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2054
timestamp 1516325494
transform 1 0 3300 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2058
timestamp 1516325494
transform 1 0 3319 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_2056
timestamp 1516325494
transform 1 0 3338 0 1 743
box 0 0 19 49
use AND2X2  AND2X2_1793
timestamp 1516325494
transform 1 0 3357 0 1 743
box 0 0 19 49
use MUX2X1  MUX2X1_374
timestamp 1516325494
transform 1 0 3376 0 1 743
box 0 0 30 49
use NAND2X1  NAND2X1_374
timestamp 1516325494
transform -1 0 3422 0 1 743
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_342
timestamp 1516325494
transform -1 0 3475 0 1 743
box 0 0 53 49
use AND2X2  AND2X2_1540
timestamp 1516325494
transform -1 0 3494 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_533
timestamp 1516325494
transform 1 0 3494 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_533
timestamp 1516325494
transform 1 0 3502 0 1 743
box 0 0 15 49
use AND2X2  AND2X2_1680
timestamp 1516325494
transform -1 0 3536 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_535
timestamp 1516325494
transform -1 0 3544 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_535
timestamp 1516325494
transform -1 0 3559 0 1 743
box 0 0 15 49
use NAND2X1  NAND2X1_364
timestamp 1516325494
transform -1 0 3574 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_364
timestamp 1516325494
transform -1 0 3604 0 1 743
box 0 0 30 49
use FILL  FILL_BUFX2_329
timestamp 1516325494
transform 1 0 3604 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_329
timestamp 1516325494
transform 1 0 3612 0 1 743
box 0 0 15 49
use AND2X2  AND2X2_1542
timestamp 1516325494
transform 1 0 3627 0 1 743
box 0 0 19 49
use FILL  FILL_BUFX2_833
timestamp 1516325494
transform 1 0 3646 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_833
timestamp 1516325494
transform 1 0 3654 0 1 743
box 0 0 15 49
use FILL  FILL_BUFX2_158
timestamp 1516325494
transform -1 0 3677 0 1 743
box 0 0 8 49
use BUFX2  BUFX2_158
timestamp 1516325494
transform -1 0 3692 0 1 743
box 0 0 15 49
use NAND2X1  NAND2X1_363
timestamp 1516325494
transform 1 0 3692 0 1 743
box 0 0 15 49
use MUX2X1  MUX2X1_363
timestamp 1516325494
transform -1 0 3737 0 1 743
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_337
timestamp 1516325494
transform 1 0 3737 0 1 743
box 0 0 53 49
use INVX1  INVX1_265
timestamp 1516325494
transform 1 0 3791 0 1 743
box 0 0 11 49
use NAND2X1  NAND2X1_773
timestamp 1516325494
transform 1 0 3802 0 1 743
box 0 0 15 49
use INVX1  INVX1_267
timestamp 1516325494
transform 1 0 3817 0 1 743
box 0 0 11 49
use NAND2X1  NAND2X1_878
timestamp 1516325494
transform 1 0 3829 0 1 743
box 0 0 15 49
use NOR2X1  NOR2X1_173
timestamp 1516325494
transform 1 0 3844 0 1 743
box 0 0 15 49
use FILL  FILL_16_1
timestamp 1516325494
transform 1 0 3859 0 1 743
box 0 0 8 49
use OR2X2  OR2X2_582
timestamp 1516325494
transform -1 0 21 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_691
timestamp 1516325494
transform -1 0 40 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_485
timestamp 1516325494
transform 1 0 40 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_670
timestamp 1516325494
transform 1 0 59 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_670
timestamp 1516325494
transform 1 0 67 0 -1 742
box 0 0 15 49
use INVX2  INVX2_3
timestamp 1516325494
transform 1 0 82 0 -1 742
box 0 0 11 49
use FILL  FILL_BUFX2_756
timestamp 1516325494
transform -1 0 101 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_756
timestamp 1516325494
transform -1 0 116 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_733
timestamp 1516325494
transform -1 0 135 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_871
timestamp 1516325494
transform -1 0 154 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_872
timestamp 1516325494
transform -1 0 173 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_916
timestamp 1516325494
transform -1 0 192 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_893
timestamp 1516325494
transform 1 0 192 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_894
timestamp 1516325494
transform 1 0 211 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_748
timestamp 1516325494
transform 1 0 230 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_841
timestamp 1516325494
transform 1 0 249 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_78
timestamp 1516325494
transform 1 0 268 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_78
timestamp 1516325494
transform 1 0 276 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_738
timestamp 1516325494
transform 1 0 291 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_718
timestamp 1516325494
transform -1 0 351 0 -1 742
box 0 0 30 49
use OR2X2  OR2X2_404
timestamp 1516325494
transform 1 0 352 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_673
timestamp 1516325494
transform 1 0 371 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_667
timestamp 1516325494
transform -1 0 431 0 -1 742
box 0 0 30 49
use FILL  FILL_BUFX2_673
timestamp 1516325494
transform 1 0 431 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_673
timestamp 1516325494
transform 1 0 439 0 -1 742
box 0 0 15 49
use FILL  FILL_BUFX2_755
timestamp 1516325494
transform 1 0 454 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_755
timestamp 1516325494
transform 1 0 462 0 -1 742
box 0 0 15 49
use AND2X2  AND2X2_668
timestamp 1516325494
transform -1 0 496 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_658
timestamp 1516325494
transform -1 0 515 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_542
timestamp 1516325494
transform -1 0 534 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_474
timestamp 1516325494
transform -1 0 553 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_653
timestamp 1516325494
transform -1 0 583 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_654
timestamp 1516325494
transform -1 0 613 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_670
timestamp 1516325494
transform 1 0 614 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_668
timestamp 1516325494
transform -1 0 674 0 -1 742
box 0 0 30 49
use FILL  FILL_BUFX2_373
timestamp 1516325494
transform 1 0 675 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_373
timestamp 1516325494
transform 1 0 682 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_419
timestamp 1516325494
transform -1 0 716 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_669
timestamp 1516325494
transform -1 0 746 0 -1 742
box 0 0 30 49
use AND2X2  AND2X2_454
timestamp 1516325494
transform 1 0 747 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_453
timestamp 1516325494
transform 1 0 766 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_648
timestamp 1516325494
transform 1 0 785 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_645
timestamp 1516325494
transform 1 0 815 0 -1 742
box 0 0 30 49
use AND2X2  AND2X2_460
timestamp 1516325494
transform 1 0 846 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_646
timestamp 1516325494
transform 1 0 865 0 -1 742
box 0 0 30 49
use AND2X2  AND2X2_555
timestamp 1516325494
transform 1 0 895 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_641
timestamp 1516325494
transform 1 0 914 0 -1 742
box 0 0 30 49
use FILL  FILL_BUFX2_376
timestamp 1516325494
transform -1 0 952 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_376
timestamp 1516325494
transform -1 0 967 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_756
timestamp 1516325494
transform 1 0 967 0 -1 742
box 0 0 30 49
use OR2X2  OR2X2_1344
timestamp 1516325494
transform 1 0 998 0 -1 742
box 0 0 19 49
use FILL  FILL_OR2X2_176
timestamp 1516325494
transform -1 0 1025 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_176
timestamp 1516325494
transform -1 0 1043 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_189
timestamp 1516325494
transform -1 0 1051 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_189
timestamp 1516325494
transform -1 0 1070 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1673
timestamp 1516325494
transform -1 0 1089 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1314
timestamp 1516325494
transform -1 0 1108 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1313
timestamp 1516325494
transform -1 0 1127 0 -1 742
box 0 0 19 49
use FILL  FILL_OR2X2_93
timestamp 1516325494
transform -1 0 1135 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_93
timestamp 1516325494
transform -1 0 1153 0 -1 742
box 0 0 19 49
use BUFX2  BUFX2_873
timestamp 1516325494
transform -1 0 1168 0 -1 742
box 0 0 15 49
use FILL  FILL_OR2X2_91
timestamp 1516325494
transform -1 0 1177 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_91
timestamp 1516325494
transform -1 0 1195 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_97
timestamp 1516325494
transform -1 0 1203 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_97
timestamp 1516325494
transform -1 0 1222 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1312
timestamp 1516325494
transform -1 0 1241 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1306
timestamp 1516325494
transform -1 0 1260 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1531
timestamp 1516325494
transform -1 0 1279 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1529
timestamp 1516325494
transform -1 0 1298 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_96
timestamp 1516325494
transform -1 0 1306 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_96
timestamp 1516325494
transform -1 0 1324 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_95
timestamp 1516325494
transform 1 0 1324 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_95
timestamp 1516325494
transform 1 0 1332 0 -1 742
box 0 0 15 49
use AND2X2  AND2X2_1853
timestamp 1516325494
transform 1 0 1347 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1726
timestamp 1516325494
transform 1 0 1366 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1851
timestamp 1516325494
transform -1 0 1404 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_322
timestamp 1516325494
transform 1 0 1404 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_322
timestamp 1516325494
transform 1 0 1412 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_289
timestamp 1516325494
transform -1 0 1446 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_817
timestamp 1516325494
transform 1 0 1446 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_817
timestamp 1516325494
transform 1 0 1454 0 -1 742
box 0 0 15 49
use AND2X2  AND2X2_1440
timestamp 1516325494
transform 1 0 1469 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1187
timestamp 1516325494
transform -1 0 1507 0 -1 742
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_518
timestamp 1516325494
transform 1 0 1507 0 -1 742
box 0 0 53 49
use MUX2X1  MUX2X1_518
timestamp 1516325494
transform 1 0 1560 0 -1 742
box 0 0 30 49
use NAND2X1  NAND2X1_518
timestamp 1516325494
transform 1 0 1590 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_1667
timestamp 1516325494
transform -1 0 1625 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_52
timestamp 1516325494
transform -1 0 1633 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_52
timestamp 1516325494
transform -1 0 1647 0 -1 742
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_534
timestamp 1516325494
transform 1 0 1647 0 -1 742
box 0 0 53 49
use NAND2X1  NAND2X1_534
timestamp 1516325494
transform 1 0 1701 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_534
timestamp 1516325494
transform -1 0 1746 0 -1 742
box 0 0 30 49
use AND2X2  AND2X2_1346
timestamp 1516325494
transform -1 0 1765 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1065
timestamp 1516325494
transform -1 0 1784 0 -1 742
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_66
timestamp 1516325494
transform 1 0 1784 0 -1 742
box 0 0 53 49
use NAND2X1  NAND2X1_130
timestamp 1516325494
transform 1 0 1837 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_130
timestamp 1516325494
transform -1 0 1883 0 -1 742
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_605
timestamp 1516325494
transform 1 0 1883 0 -1 742
box 0 0 53 49
use NAND2X1  NAND2X1_29
timestamp 1516325494
transform 1 0 1936 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_1064
timestamp 1516325494
transform -1 0 1970 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_322
timestamp 1516325494
transform -1 0 2000 0 -1 742
box 0 0 30 49
use NAND2X1  NAND2X1_322
timestamp 1516325494
transform -1 0 2016 0 -1 742
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_450
timestamp 1516325494
transform -1 0 2069 0 -1 742
box 0 0 53 49
use FILL  FILL_BUFX2_815
timestamp 1516325494
transform 1 0 2069 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_815
timestamp 1516325494
transform 1 0 2077 0 -1 742
box 0 0 15 49
use AND2X2  AND2X2_2067
timestamp 1516325494
transform -1 0 2111 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_2061
timestamp 1516325494
transform -1 0 2130 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_2065
timestamp 1516325494
transform -1 0 2149 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_2070
timestamp 1516325494
transform -1 0 2168 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_2063
timestamp 1516325494
transform -1 0 2187 0 -1 742
box 0 0 19 49
use MUX2X1  MUX2X1_326
timestamp 1516325494
transform -1 0 2217 0 -1 742
box 0 0 30 49
use AND2X2  AND2X2_1313
timestamp 1516325494
transform -1 0 2236 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1310
timestamp 1516325494
transform -1 0 2255 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1489
timestamp 1516325494
transform 1 0 2255 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1672
timestamp 1516325494
transform -1 0 2293 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_54
timestamp 1516325494
transform -1 0 2301 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_54
timestamp 1516325494
transform -1 0 2316 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_1490
timestamp 1516325494
transform -1 0 2335 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1304
timestamp 1516325494
transform 1 0 2335 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1530
timestamp 1516325494
transform -1 0 2373 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_859
timestamp 1516325494
transform 1 0 2373 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_859
timestamp 1516325494
transform 1 0 2381 0 -1 742
box 0 0 15 49
use FILL  FILL_BUFX2_18
timestamp 1516325494
transform -1 0 2404 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_18
timestamp 1516325494
transform -1 0 2419 0 -1 742
box 0 0 15 49
use NAND2X1  NAND2X1_330
timestamp 1516325494
transform 1 0 2419 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_330
timestamp 1516325494
transform 1 0 2434 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_522
timestamp 1516325494
transform -1 0 2494 0 -1 742
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_458
timestamp 1516325494
transform 1 0 2495 0 -1 742
box 0 0 53 49
use AND2X2  AND2X2_1303
timestamp 1516325494
transform -1 0 2567 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_211
timestamp 1516325494
transform -1 0 2575 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_211
timestamp 1516325494
transform -1 0 2590 0 -1 742
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_88
timestamp 1516325494
transform 1 0 2590 0 -1 742
box 0 0 53 49
use AND2X2  AND2X2_2060
timestamp 1516325494
transform -1 0 2662 0 -1 742
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_233
timestamp 1516325494
transform -1 0 2715 0 -1 742
box 0 0 53 49
use FILL  FILL_AND2X2_72
timestamp 1516325494
transform -1 0 2723 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_72
timestamp 1516325494
transform -1 0 2742 0 -1 742
box 0 0 19 49
use FILL  FILL_OR2X2_73
timestamp 1516325494
transform -1 0 2750 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_73
timestamp 1516325494
transform -1 0 2768 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_71
timestamp 1516325494
transform 1 0 2768 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_71
timestamp 1516325494
transform 1 0 2776 0 -1 742
box 0 0 19 49
use FILL  FILL_OR2X2_68
timestamp 1516325494
transform 1 0 2795 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_68
timestamp 1516325494
transform 1 0 2803 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1492
timestamp 1516325494
transform -1 0 2841 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1491
timestamp 1516325494
transform -1 0 2860 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1256
timestamp 1516325494
transform -1 0 2879 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1493
timestamp 1516325494
transform -1 0 2898 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_379
timestamp 1516325494
transform -1 0 2906 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_379
timestamp 1516325494
transform -1 0 2920 0 -1 742
box 0 0 15 49
use AND2X2  AND2X2_2042
timestamp 1516325494
transform 1 0 2920 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_2043
timestamp 1516325494
transform -1 0 2958 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_393
timestamp 1516325494
transform -1 0 2966 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_393
timestamp 1516325494
transform -1 0 2981 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_1290
timestamp 1516325494
transform -1 0 3000 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_663
timestamp 1516325494
transform 1 0 3000 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_663
timestamp 1516325494
transform 1 0 3008 0 -1 742
box 0 0 15 49
use INVX1  INVX1_323
timestamp 1516325494
transform 1 0 3023 0 -1 742
box 0 0 11 49
use AND2X2  AND2X2_1285
timestamp 1516325494
transform 1 0 3034 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_603
timestamp 1516325494
transform 1 0 3053 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_603
timestamp 1516325494
transform 1 0 3061 0 -1 742
box 0 0 15 49
use AND2X2  AND2X2_1289
timestamp 1516325494
transform 1 0 3076 0 -1 742
box 0 0 19 49
use FILL  FILL_BUFX2_107
timestamp 1516325494
transform 1 0 3095 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_107
timestamp 1516325494
transform 1 0 3103 0 -1 742
box 0 0 15 49
use FILL  FILL_BUFX2_340
timestamp 1516325494
transform 1 0 3118 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_340
timestamp 1516325494
transform 1 0 3126 0 -1 742
box 0 0 15 49
use NOR2X1  NOR2X1_176
timestamp 1516325494
transform 1 0 3141 0 -1 742
box 0 0 15 49
use FILL  FILL_BUFX2_618
timestamp 1516325494
transform 1 0 3156 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_618
timestamp 1516325494
transform 1 0 3164 0 -1 742
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_708
timestamp 1516325494
transform -1 0 3232 0 -1 742
box 0 0 53 49
use NAND2X1  NAND2X1_749
timestamp 1516325494
transform -1 0 3247 0 -1 742
box 0 0 15 49
use OR2X2  OR2X2_1499
timestamp 1516325494
transform -1 0 3266 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1289
timestamp 1516325494
transform -1 0 3285 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1517
timestamp 1516325494
transform -1 0 3304 0 -1 742
box 0 0 19 49
use NOR2X1  NOR2X1_178
timestamp 1516325494
transform 1 0 3304 0 -1 742
box 0 0 15 49
use FILL  FILL_BUFX2_657
timestamp 1516325494
transform 1 0 3319 0 -1 742
box 0 0 8 49
use BUFX2  BUFX2_657
timestamp 1516325494
transform 1 0 3327 0 -1 742
box 0 0 15 49
use NAND2X1  NAND2X1_593
timestamp 1516325494
transform 1 0 3342 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_593
timestamp 1516325494
transform -1 0 3387 0 -1 742
box 0 0 30 49
use FILL  FILL_OR2X2_72
timestamp 1516325494
transform -1 0 3396 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_72
timestamp 1516325494
transform -1 0 3414 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1288
timestamp 1516325494
transform -1 0 3433 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1519
timestamp 1516325494
transform -1 0 3452 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1319
timestamp 1516325494
transform -1 0 3471 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1498
timestamp 1516325494
transform -1 0 3490 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1518
timestamp 1516325494
transform -1 0 3509 0 -1 742
box 0 0 19 49
use FILL  FILL_OR2X2_183
timestamp 1516325494
transform -1 0 3517 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_183
timestamp 1516325494
transform -1 0 3536 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_196
timestamp 1516325494
transform -1 0 3544 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_196
timestamp 1516325494
transform -1 0 3563 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1679
timestamp 1516325494
transform -1 0 3582 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_195
timestamp 1516325494
transform -1 0 3590 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_195
timestamp 1516325494
transform -1 0 3608 0 -1 742
box 0 0 19 49
use FILL  FILL_AND2X2_106
timestamp 1516325494
transform -1 0 3616 0 -1 742
box 0 0 8 49
use AND2X2  AND2X2_106
timestamp 1516325494
transform -1 0 3635 0 -1 742
box 0 0 19 49
use OR2X2  OR2X2_1318
timestamp 1516325494
transform -1 0 3654 0 -1 742
box 0 0 19 49
use AND2X2  AND2X2_1541
timestamp 1516325494
transform -1 0 3673 0 -1 742
box 0 0 19 49
use NAND2X1  NAND2X1_267
timestamp 1516325494
transform 1 0 3673 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_267
timestamp 1516325494
transform -1 0 3718 0 -1 742
box 0 0 30 49
use NAND2X1  NAND2X1_369
timestamp 1516325494
transform 1 0 3718 0 -1 742
box 0 0 15 49
use MUX2X1  MUX2X1_369
timestamp 1516325494
transform -1 0 3764 0 -1 742
box 0 0 30 49
use MUX2X1  MUX2X1_273
timestamp 1516325494
transform 1 0 3764 0 -1 742
box 0 0 30 49
use NAND2X1  NAND2X1_273
timestamp 1516325494
transform -1 0 3809 0 -1 742
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_145
timestamp 1516325494
transform -1 0 3863 0 -1 742
box 0 0 53 49
use FILL  FILL_15_1
timestamp 1516325494
transform -1 0 3871 0 -1 742
box 0 0 8 49
use OR2X2  OR2X2_450
timestamp 1516325494
transform 1 0 2 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_508
timestamp 1516325494
transform -1 0 40 0 1 644
box 0 0 19 49
use NAND3X1  NAND3X1_30
timestamp 1516325494
transform -1 0 59 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_690
timestamp 1516325494
transform -1 0 78 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_633
timestamp 1516325494
transform -1 0 97 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_488
timestamp 1516325494
transform -1 0 116 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_686
timestamp 1516325494
transform 1 0 116 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_524
timestamp 1516325494
transform -1 0 154 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_617
timestamp 1516325494
transform -1 0 173 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_616
timestamp 1516325494
transform -1 0 192 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_440
timestamp 1516325494
transform -1 0 211 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_491
timestamp 1516325494
transform -1 0 230 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_805
timestamp 1516325494
transform -1 0 249 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_709
timestamp 1516325494
transform -1 0 268 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_840
timestamp 1516325494
transform -1 0 287 0 1 644
box 0 0 19 49
use MUX2X1  MUX2X1_713
timestamp 1516325494
transform -1 0 317 0 1 644
box 0 0 30 49
use MUX2X1  MUX2X1_715
timestamp 1516325494
transform -1 0 347 0 1 644
box 0 0 30 49
use AND2X2  AND2X2_550
timestamp 1516325494
transform 1 0 348 0 1 644
box 0 0 19 49
use MUX2X1  MUX2X1_711
timestamp 1516325494
transform -1 0 397 0 1 644
box 0 0 30 49
use XOR2X1  XOR2X1_1
timestamp 1516325494
transform -1 0 431 0 1 644
box 0 0 34 49
use XOR2X1  XOR2X1_4
timestamp 1516325494
transform 1 0 431 0 1 644
box 0 0 34 49
use AND2X2  AND2X2_505
timestamp 1516325494
transform -1 0 21 0 -1 644
box 0 0 19 49
use NAND2X1  NAND2X1_658
timestamp 1516325494
transform -1 0 36 0 -1 644
box 0 0 15 49
use OR2X2  OR2X2_618
timestamp 1516325494
transform -1 0 55 0 -1 644
box 0 0 19 49
use NAND2X1  NAND2X1_657
timestamp 1516325494
transform -1 0 70 0 -1 644
box 0 0 15 49
use AND2X2  AND2X2_740
timestamp 1516325494
transform -1 0 89 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_523
timestamp 1516325494
transform -1 0 108 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_438
timestamp 1516325494
transform -1 0 127 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_487
timestamp 1516325494
transform -1 0 146 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_486
timestamp 1516325494
transform -1 0 165 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_679
timestamp 1516325494
transform 1 0 165 0 -1 644
box 0 0 30 49
use AND2X2  AND2X2_490
timestamp 1516325494
transform 1 0 196 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_678
timestamp 1516325494
transform -1 0 245 0 -1 644
box 0 0 30 49
use MUX2X1  MUX2X1_680
timestamp 1516325494
transform -1 0 275 0 -1 644
box 0 0 30 49
use FILL  FILL_BUFX2_542
timestamp 1516325494
transform 1 0 276 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_542
timestamp 1516325494
transform 1 0 283 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_666
timestamp 1516325494
transform -1 0 328 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_477
timestamp 1516325494
transform 1 0 329 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_549
timestamp 1516325494
transform -1 0 367 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_430
timestamp 1516325494
transform 1 0 367 0 -1 644
box 0 0 19 49
use INVX2  INVX2_4
timestamp 1516325494
transform -1 0 397 0 -1 644
box 0 0 11 49
use OR2X2  OR2X2_429
timestamp 1516325494
transform 1 0 397 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_469
timestamp 1516325494
transform -1 0 435 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_674
timestamp 1516325494
transform 1 0 435 0 -1 644
box 0 0 30 49
use AND2X2  AND2X2_669
timestamp 1516325494
transform -1 0 485 0 1 644
box 0 0 19 49
use FILL  FILL_BUFX2_375
timestamp 1516325494
transform 1 0 485 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_375
timestamp 1516325494
transform 1 0 492 0 1 644
box 0 0 15 49
use AND2X2  AND2X2_657
timestamp 1516325494
transform -1 0 526 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_676
timestamp 1516325494
transform 1 0 526 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_539
timestamp 1516325494
transform -1 0 564 0 1 644
box 0 0 19 49
use FILL  FILL_BUFX2_378
timestamp 1516325494
transform 1 0 564 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_378
timestamp 1516325494
transform 1 0 572 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_702
timestamp 1516325494
transform -1 0 617 0 1 644
box 0 0 30 49
use OR2X2  OR2X2_810
timestamp 1516325494
transform -1 0 637 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_850
timestamp 1516325494
transform -1 0 656 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_473
timestamp 1516325494
transform -1 0 675 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_541
timestamp 1516325494
transform -1 0 694 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_540
timestamp 1516325494
transform -1 0 713 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_451
timestamp 1516325494
transform -1 0 732 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_450
timestamp 1516325494
transform -1 0 751 0 1 644
box 0 0 19 49
use MUX2X1  MUX2X1_652
timestamp 1516325494
transform -1 0 781 0 1 644
box 0 0 30 49
use OR2X2  OR2X2_480
timestamp 1516325494
transform -1 0 800 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_551
timestamp 1516325494
transform 1 0 800 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_552
timestamp 1516325494
transform -1 0 838 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_665
timestamp 1516325494
transform -1 0 857 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_864
timestamp 1516325494
transform 1 0 857 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_828
timestamp 1516325494
transform 1 0 876 0 1 644
box 0 0 19 49
use FILL  FILL_BUFX2_371
timestamp 1516325494
transform 1 0 895 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_371
timestamp 1516325494
transform 1 0 903 0 1 644
box 0 0 15 49
use FILL  FILL_BUFX2_76
timestamp 1516325494
transform 1 0 918 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_76
timestamp 1516325494
transform 1 0 925 0 1 644
box 0 0 15 49
use FILL  FILL_BUFX2_544
timestamp 1516325494
transform -1 0 949 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_544
timestamp 1516325494
transform -1 0 963 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_801
timestamp 1516325494
transform 1 0 963 0 1 644
box 0 0 30 49
use MUX2X1  MUX2X1_794
timestamp 1516325494
transform 1 0 994 0 1 644
box 0 0 30 49
use INVX1  INVX1_144
timestamp 1516325494
transform 1 0 1024 0 1 644
box 0 0 11 49
use FILL  FILL_OR2X2_94
timestamp 1516325494
transform -1 0 1044 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_94
timestamp 1516325494
transform -1 0 1062 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1491
timestamp 1516325494
transform -1 0 1081 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1671
timestamp 1516325494
transform -1 0 1100 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_188
timestamp 1516325494
transform -1 0 1108 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_188
timestamp 1516325494
transform -1 0 1127 0 1 644
box 0 0 19 49
use FILL  FILL_OR2X2_220
timestamp 1516325494
transform 1 0 1127 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_220
timestamp 1516325494
transform 1 0 1134 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1581
timestamp 1516325494
transform 1 0 1153 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1524
timestamp 1516325494
transform -1 0 1191 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1582
timestamp 1516325494
transform 1 0 1191 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1583
timestamp 1516325494
transform 1 0 1210 0 1 644
box 0 0 19 49
use FILL  FILL_OR2X2_219
timestamp 1516325494
transform -1 0 1237 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_219
timestamp 1516325494
transform -1 0 1256 0 1 644
box 0 0 19 49
use FILL  FILL_OR2X2_218
timestamp 1516325494
transform -1 0 1264 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_218
timestamp 1516325494
transform -1 0 1283 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_234
timestamp 1516325494
transform -1 0 1291 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_234
timestamp 1516325494
transform -1 0 1309 0 1 644
box 0 0 19 49
use FILL  FILL_OR2X2_217
timestamp 1516325494
transform -1 0 1317 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_217
timestamp 1516325494
transform -1 0 1336 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_232
timestamp 1516325494
transform -1 0 1344 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_232
timestamp 1516325494
transform -1 0 1362 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1733
timestamp 1516325494
transform 1 0 1362 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1734
timestamp 1516325494
transform -1 0 1400 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_231
timestamp 1516325494
transform -1 0 1408 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_231
timestamp 1516325494
transform -1 0 1427 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_307
timestamp 1516325494
transform 1 0 1427 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_287
timestamp 1516325494
transform -1 0 1465 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_306
timestamp 1516325494
transform 1 0 1465 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1532
timestamp 1516325494
transform -1 0 1503 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1308
timestamp 1516325494
transform -1 0 1522 0 1 644
box 0 0 19 49
use NAND2X1  NAND2X1_106
timestamp 1516325494
transform 1 0 1522 0 1 644
box 0 0 15 49
use OR2X2  OR2X2_1307
timestamp 1516325494
transform -1 0 1556 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1188
timestamp 1516325494
transform -1 0 1575 0 1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_6
timestamp 1516325494
transform 1 0 1575 0 1 644
box 0 0 53 49
use NAND2X1  NAND2X1_102
timestamp 1516325494
transform 1 0 1628 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_102
timestamp 1516325494
transform -1 0 1674 0 1 644
box 0 0 30 49
use AND2X2  AND2X2_1528
timestamp 1516325494
transform -1 0 1693 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1850
timestamp 1516325494
transform -1 0 1712 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1501
timestamp 1516325494
transform -1 0 1731 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1266
timestamp 1516325494
transform -1 0 1750 0 1 644
box 0 0 19 49
use NAND2X1  NAND2X1_887
timestamp 1516325494
transform 1 0 1750 0 1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_617
timestamp 1516325494
transform 1 0 1765 0 1 644
box 0 0 53 49
use MUX2X1  MUX2X1_832
timestamp 1516325494
transform -1 0 1848 0 1 644
box 0 0 30 49
use OR2X2  OR2X2_1722
timestamp 1516325494
transform -1 0 1868 0 1 644
box 0 0 19 49
use FILL  FILL_BUFX2_13
timestamp 1516325494
transform 1 0 1868 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_13
timestamp 1516325494
transform 1 0 1875 0 1 644
box 0 0 15 49
use FILL  FILL_BUFX2_793
timestamp 1516325494
transform 1 0 1891 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_793
timestamp 1516325494
transform 1 0 1898 0 1 644
box 0 0 15 49
use OR2X2  OR2X2_1484
timestamp 1516325494
transform -1 0 1932 0 1 644
box 0 0 19 49
use NAND2X1  NAND2X1_336
timestamp 1516325494
transform 1 0 1932 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_336
timestamp 1516325494
transform -1 0 1978 0 1 644
box 0 0 30 49
use FILL  FILL_BUFX2_702
timestamp 1516325494
transform 1 0 1978 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_702
timestamp 1516325494
transform 1 0 1986 0 1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_464
timestamp 1516325494
transform -1 0 2054 0 1 644
box 0 0 53 49
use FILL  FILL_BUFX2_176
timestamp 1516325494
transform 1 0 2054 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_176
timestamp 1516325494
transform 1 0 2062 0 1 644
box 0 0 15 49
use FILL  FILL_BUFX2_438
timestamp 1516325494
transform -1 0 2085 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_438
timestamp 1516325494
transform -1 0 2099 0 1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_400
timestamp 1516325494
transform 1 0 2100 0 1 644
box 0 0 53 49
use NAND2X1  NAND2X1_176
timestamp 1516325494
transform 1 0 2153 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_176
timestamp 1516325494
transform -1 0 2198 0 1 644
box 0 0 30 49
use MUX2X1  MUX2X1_560
timestamp 1516325494
transform 1 0 2198 0 1 644
box 0 0 30 49
use NAND2X1  NAND2X1_560
timestamp 1516325494
transform -1 0 2244 0 1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_496
timestamp 1516325494
transform -1 0 2297 0 1 644
box 0 0 53 49
use AND2X2  AND2X2_1304
timestamp 1516325494
transform -1 0 2316 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1307
timestamp 1516325494
transform -1 0 2335 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1724
timestamp 1516325494
transform 1 0 2335 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1852
timestamp 1516325494
transform -1 0 2373 0 1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_472
timestamp 1516325494
transform -1 0 2426 0 1 644
box 0 0 53 49
use OR2X2  OR2X2_1305
timestamp 1516325494
transform -1 0 2445 0 1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_522
timestamp 1516325494
transform 1 0 2445 0 1 644
box 0 0 53 49
use MUX2X1  MUX2X1_650
timestamp 1516325494
transform -1 0 496 0 -1 644
box 0 0 30 49
use MUX2X1  MUX2X1_657
timestamp 1516325494
transform -1 0 526 0 -1 644
box 0 0 30 49
use MUX2X1  MUX2X1_651
timestamp 1516325494
transform -1 0 556 0 -1 644
box 0 0 30 49
use MUX2X1  MUX2X1_675
timestamp 1516325494
transform -1 0 587 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_623
timestamp 1516325494
transform 1 0 587 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_439
timestamp 1516325494
transform -1 0 625 0 -1 644
box 0 0 19 49
use FILL  FILL_BUFX2_698
timestamp 1516325494
transform -1 0 633 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_698
timestamp 1516325494
transform -1 0 648 0 -1 644
box 0 0 15 49
use AND2X2  AND2X2_642
timestamp 1516325494
transform -1 0 667 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_656
timestamp 1516325494
transform -1 0 697 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_587
timestamp 1516325494
transform 1 0 697 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_696
timestamp 1516325494
transform -1 0 735 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_574
timestamp 1516325494
transform -1 0 754 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_647
timestamp 1516325494
transform -1 0 784 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_408
timestamp 1516325494
transform -1 0 804 0 -1 644
box 0 0 19 49
use XOR2X1  XOR2X1_2
timestamp 1516325494
transform 1 0 804 0 -1 644
box 0 0 34 49
use XNOR2X1  XNOR2X1_2
timestamp 1516325494
transform 1 0 838 0 -1 644
box 0 0 34 49
use FILL  FILL_BUFX2_627
timestamp 1516325494
transform -1 0 880 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_627
timestamp 1516325494
transform -1 0 895 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_787
timestamp 1516325494
transform 1 0 895 0 -1 644
box 0 0 30 49
use INVX1  INVX1_209
timestamp 1516325494
transform -1 0 936 0 -1 644
box 0 0 11 49
use FILL  FILL_OR2X2_95
timestamp 1516325494
transform -1 0 945 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_95
timestamp 1516325494
transform -1 0 963 0 -1 644
box 0 0 19 49
use INVX1  INVX1_223
timestamp 1516325494
transform 1 0 963 0 -1 644
box 0 0 11 49
use INVX1  INVX1_216
timestamp 1516325494
transform 1 0 975 0 -1 644
box 0 0 11 49
use FILL  FILL_OR2X2_193
timestamp 1516325494
transform -1 0 994 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_193
timestamp 1516325494
transform -1 0 1013 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_177
timestamp 1516325494
transform -1 0 1021 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_177
timestamp 1516325494
transform -1 0 1039 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1492
timestamp 1516325494
transform -1 0 1058 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_203
timestamp 1516325494
transform -1 0 1066 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_203
timestamp 1516325494
transform -1 0 1085 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1740
timestamp 1516325494
transform -1 0 1104 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_233
timestamp 1516325494
transform 1 0 1104 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_233
timestamp 1516325494
transform 1 0 1112 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1694
timestamp 1516325494
transform 1 0 1131 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1742
timestamp 1516325494
transform 1 0 1150 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1486
timestamp 1516325494
transform -1 0 1188 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1669
timestamp 1516325494
transform -1 0 1207 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1667
timestamp 1516325494
transform -1 0 1226 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_175
timestamp 1516325494
transform -1 0 1234 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_175
timestamp 1516325494
transform -1 0 1252 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_186
timestamp 1516325494
transform -1 0 1260 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_186
timestamp 1516325494
transform -1 0 1279 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_187
timestamp 1516325494
transform -1 0 1287 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_187
timestamp 1516325494
transform -1 0 1305 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1576
timestamp 1516325494
transform -1 0 1324 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1736
timestamp 1516325494
transform -1 0 1343 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1738
timestamp 1516325494
transform -1 0 1362 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_290
timestamp 1516325494
transform 1 0 1362 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_291
timestamp 1516325494
transform -1 0 1400 0 -1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_602
timestamp 1516325494
transform 1 0 1400 0 -1 644
box 0 0 53 49
use NAND2X1  NAND2X1_26
timestamp 1516325494
transform 1 0 1454 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_26
timestamp 1516325494
transform -1 0 1499 0 -1 644
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_10
timestamp 1516325494
transform 1 0 1499 0 -1 644
box 0 0 53 49
use MUX2X1  MUX2X1_106
timestamp 1516325494
transform -1 0 1582 0 -1 644
box 0 0 30 49
use MUX2X1  MUX2X1_865
timestamp 1516325494
transform 1 0 1583 0 -1 644
box 0 0 30 49
use NAND2X1  NAND2X1_920
timestamp 1516325494
transform -1 0 1628 0 -1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_362
timestamp 1516325494
transform -1 0 1681 0 -1 644
box 0 0 53 49
use OR2X2  OR2X2_1302
timestamp 1516325494
transform -1 0 1701 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1668
timestamp 1516325494
transform -1 0 1720 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1485
timestamp 1516325494
transform -1 0 1739 0 -1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_80
timestamp 1516325494
transform 1 0 1739 0 -1 644
box 0 0 53 49
use NAND2X1  NAND2X1_144
timestamp 1516325494
transform 1 0 1792 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_144
timestamp 1516325494
transform 1 0 1807 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_1482
timestamp 1516325494
transform 1 0 1837 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1666
timestamp 1516325494
transform -1 0 1875 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1861
timestamp 1516325494
transform -1 0 1894 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1487
timestamp 1516325494
transform 1 0 1894 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1670
timestamp 1516325494
transform -1 0 1932 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1488
timestamp 1516325494
transform -1 0 1951 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1483
timestamp 1516325494
transform -1 0 1970 0 -1 644
box 0 0 19 49
use NAND2X1  NAND2X1_112
timestamp 1516325494
transform 1 0 1970 0 -1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_16
timestamp 1516325494
transform 1 0 1986 0 -1 644
box 0 0 53 49
use MUX2X1  MUX2X1_112
timestamp 1516325494
transform -1 0 2069 0 -1 644
box 0 0 30 49
use FILL  FILL_BUFX2_242
timestamp 1516325494
transform -1 0 2077 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_242
timestamp 1516325494
transform -1 0 2092 0 -1 644
box 0 0 15 49
use NAND2X1  NAND2X1_528
timestamp 1516325494
transform 1 0 2092 0 -1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_528
timestamp 1516325494
transform 1 0 2107 0 -1 644
box 0 0 53 49
use MUX2X1  MUX2X1_528
timestamp 1516325494
transform -1 0 2190 0 -1 644
box 0 0 30 49
use FILL  FILL_BUFX2_121
timestamp 1516325494
transform -1 0 2199 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_121
timestamp 1516325494
transform -1 0 2213 0 -1 644
box 0 0 15 49
use OR2X2  OR2X2_1957
timestamp 1516325494
transform -1 0 2233 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1739
timestamp 1516325494
transform -1 0 2252 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_1578
timestamp 1516325494
transform -1 0 2271 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_344
timestamp 1516325494
transform 1 0 2271 0 -1 644
box 0 0 30 49
use NAND2X1  NAND2X1_344
timestamp 1516325494
transform -1 0 2316 0 -1 644
box 0 0 15 49
use OR2X2  OR2X2_1959
timestamp 1516325494
transform -1 0 2335 0 -1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_399
timestamp 1516325494
transform 1 0 2335 0 -1 644
box 0 0 53 49
use NAND2X1  NAND2X1_175
timestamp 1516325494
transform 1 0 2388 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_175
timestamp 1516325494
transform 1 0 2404 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_1577
timestamp 1516325494
transform -1 0 2453 0 -1 644
box 0 0 19 49
use NAND2X1  NAND2X1_138
timestamp 1516325494
transform 1 0 2453 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_138
timestamp 1516325494
transform 1 0 2468 0 -1 644
box 0 0 30 49
use OR2X2  OR2X2_1725
timestamp 1516325494
transform -1 0 2518 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1735
timestamp 1516325494
transform -1 0 2537 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1573
timestamp 1516325494
transform -1 0 2556 0 1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_403
timestamp 1516325494
transform 1 0 2556 0 1 644
box 0 0 53 49
use NAND2X1  NAND2X1_179
timestamp 1516325494
transform 1 0 2609 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_179
timestamp 1516325494
transform -1 0 2654 0 1 644
box 0 0 30 49
use AND2X2  AND2X2_2069
timestamp 1516325494
transform -1 0 2673 0 1 644
box 0 0 19 49
use NAND2X1  NAND2X1_152
timestamp 1516325494
transform 1 0 2673 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_152
timestamp 1516325494
transform 1 0 2689 0 1 644
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_376
timestamp 1516325494
transform 1 0 2719 0 1 644
box 0 0 53 49
use NAND2X1  NAND2X1_934
timestamp 1516325494
transform 1 0 2772 0 1 644
box 0 0 15 49
use MUX2X1  MUX2X1_879
timestamp 1516325494
transform -1 0 2817 0 1 644
box 0 0 30 49
use FILL  FILL_OR2X2_70
timestamp 1516325494
transform 1 0 2818 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_70
timestamp 1516325494
transform 1 0 2825 0 1 644
box 0 0 19 49
use MUX2X1  MUX2X1_617
timestamp 1516325494
transform 1 0 2844 0 1 644
box 0 0 30 49
use NAND2X1  NAND2X1_617
timestamp 1516325494
transform -1 0 2890 0 1 644
box 0 0 15 49
use OR2X2  OR2X2_1710
timestamp 1516325494
transform -1 0 2909 0 1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_201
timestamp 1516325494
transform -1 0 2962 0 1 644
box 0 0 53 49
use MUX2X1  MUX2X1_243
timestamp 1516325494
transform 1 0 2962 0 1 644
box 0 0 30 49
use OR2X2  OR2X2_1287
timestamp 1516325494
transform -1 0 3012 0 1 644
box 0 0 19 49
use NAND2X1  NAND2X1_586
timestamp 1516325494
transform 1 0 3012 0 1 644
box 0 0 15 49
use OR2X2  OR2X2_1286
timestamp 1516325494
transform -1 0 3046 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1516
timestamp 1516325494
transform -1 0 3065 0 1 644
box 0 0 19 49
use OR2X2  OR2X2_1320
timestamp 1516325494
transform -1 0 3084 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1515
timestamp 1516325494
transform -1 0 3103 0 1 644
box 0 0 19 49
use FILL  FILL_BUFX2_339
timestamp 1516325494
transform 1 0 3103 0 1 644
box 0 0 8 49
use BUFX2  BUFX2_339
timestamp 1516325494
transform 1 0 3110 0 1 644
box 0 0 15 49
use NOR2X1  NOR2X1_175
timestamp 1516325494
transform -1 0 3141 0 1 644
box 0 0 15 49
use NAND2X1  NAND2X1_243
timestamp 1516325494
transform -1 0 3156 0 1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_179
timestamp 1516325494
transform -1 0 3209 0 1 644
box 0 0 53 49
use OR2X2  OR2X2_1500
timestamp 1516325494
transform -1 0 3228 0 1 644
box 0 0 19 49
use INVX1  INVX1_324
timestamp 1516325494
transform 1 0 3228 0 1 644
box 0 0 11 49
use AND2X2  AND2X2_1288
timestamp 1516325494
transform 1 0 3240 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1294
timestamp 1516325494
transform -1 0 3278 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1291
timestamp 1516325494
transform -1 0 3297 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_2045
timestamp 1516325494
transform -1 0 3316 0 1 644
box 0 0 19 49
use NOR2X1  NOR2X1_177
timestamp 1516325494
transform -1 0 3331 0 1 644
box 0 0 15 49
use OR2X2  OR2X2_1709
timestamp 1516325494
transform -1 0 3350 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_1839
timestamp 1516325494
transform -1 0 3369 0 1 644
box 0 0 19 49
use AND2X2  AND2X2_2048
timestamp 1516325494
transform -1 0 3388 0 1 644
box 0 0 19 49
use INVX1  INVX1_329
timestamp 1516325494
transform -1 0 3399 0 1 644
box 0 0 11 49
use NAND2X1  NAND2X1_362
timestamp 1516325494
transform -1 0 3414 0 1 644
box 0 0 15 49
use FILL  FILL_AND2X2_74
timestamp 1516325494
transform -1 0 3422 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_74
timestamp 1516325494
transform -1 0 3441 0 1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_273
timestamp 1516325494
transform -1 0 3494 0 1 644
box 0 0 53 49
use OR2X2  OR2X2_1708
timestamp 1516325494
transform 1 0 3494 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_89
timestamp 1516325494
transform 1 0 3513 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_89
timestamp 1516325494
transform 1 0 3521 0 1 644
box 0 0 19 49
use FILL  FILL_OR2X2_86
timestamp 1516325494
transform -1 0 3548 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_86
timestamp 1516325494
transform -1 0 3566 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_91
timestamp 1516325494
transform 1 0 3566 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_91
timestamp 1516325494
transform 1 0 3574 0 1 644
box 0 0 19 49
use FILL  FILL_OR2X2_85
timestamp 1516325494
transform -1 0 3601 0 1 644
box 0 0 8 49
use OR2X2  OR2X2_85
timestamp 1516325494
transform -1 0 3620 0 1 644
box 0 0 19 49
use FILL  FILL_AND2X2_90
timestamp 1516325494
transform -1 0 3628 0 1 644
box 0 0 8 49
use AND2X2  AND2X2_90
timestamp 1516325494
transform -1 0 3646 0 1 644
box 0 0 19 49
use MUX2X1  MUX2X1_266
timestamp 1516325494
transform 1 0 3646 0 1 644
box 0 0 30 49
use MUX2X1  MUX2X1_376
timestamp 1516325494
transform -1 0 3707 0 1 644
box 0 0 30 49
use NAND2X1  NAND2X1_266
timestamp 1516325494
transform -1 0 3722 0 1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_139
timestamp 1516325494
transform -1 0 3775 0 1 644
box 0 0 53 49
use INVX1  INVX1_264
timestamp 1516325494
transform 1 0 3775 0 1 644
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_138
timestamp 1516325494
transform -1 0 3840 0 1 644
box 0 0 53 49
use NAND3X1  NAND3X1_100
timestamp 1516325494
transform 1 0 3840 0 1 644
box 0 0 19 49
use FILL  FILL_14_1
timestamp 1516325494
transform 1 0 3859 0 1 644
box 0 0 8 49
use DFFPOSX1  DFFPOSX1_74
timestamp 1516325494
transform -1 0 2552 0 -1 644
box 0 0 53 49
use OR2X2  OR2X2_1572
timestamp 1516325494
transform -1 0 2571 0 -1 644
box 0 0 19 49
use FILL  FILL_BUFX2_1
timestamp 1516325494
transform -1 0 2579 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_1
timestamp 1516325494
transform -1 0 2593 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_531
timestamp 1516325494
transform 1 0 2594 0 -1 644
box 0 0 30 49
use NAND2X1  NAND2X1_531
timestamp 1516325494
transform -1 0 2639 0 -1 644
box 0 0 15 49
use FILL  FILL_BUFX2_463
timestamp 1516325494
transform 1 0 2639 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_463
timestamp 1516325494
transform 1 0 2647 0 -1 644
box 0 0 15 49
use INVX1  INVX1_330
timestamp 1516325494
transform 1 0 2662 0 -1 644
box 0 0 11 49
use FILL  FILL_BUFX2_44
timestamp 1516325494
transform 1 0 2673 0 -1 644
box 0 0 8 49
use BUFX2  BUFX2_44
timestamp 1516325494
transform 1 0 2681 0 -1 644
box 0 0 15 49
use FILL  FILL_OR2X2_69
timestamp 1516325494
transform -1 0 2704 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_69
timestamp 1516325494
transform -1 0 2723 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_73
timestamp 1516325494
transform -1 0 2731 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_73
timestamp 1516325494
transform -1 0 2749 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_87
timestamp 1516325494
transform -1 0 2757 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_87
timestamp 1516325494
transform -1 0 2776 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_84
timestamp 1516325494
transform -1 0 2784 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_84
timestamp 1516325494
transform -1 0 2803 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_83
timestamp 1516325494
transform -1 0 2811 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_83
timestamp 1516325494
transform -1 0 2829 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_88
timestamp 1516325494
transform -1 0 2837 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_88
timestamp 1516325494
transform -1 0 2856 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_87
timestamp 1516325494
transform -1 0 2864 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_87
timestamp 1516325494
transform -1 0 2882 0 -1 644
box 0 0 19 49
use NAND2X1  NAND2X1_585
timestamp 1516325494
transform 1 0 2882 0 -1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_234
timestamp 1516325494
transform 1 0 2898 0 -1 644
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_266
timestamp 1516325494
transform 1 0 2951 0 -1 644
box 0 0 53 49
use MUX2X1  MUX2X1_586
timestamp 1516325494
transform 1 0 3004 0 -1 644
box 0 0 30 49
use FILL  FILL_AND2X2_193
timestamp 1516325494
transform 1 0 3034 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_193
timestamp 1516325494
transform 1 0 3042 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1677
timestamp 1516325494
transform 1 0 3061 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_181
timestamp 1516325494
transform 1 0 3080 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_181
timestamp 1516325494
transform 1 0 3088 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_182
timestamp 1516325494
transform 1 0 3107 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_182
timestamp 1516325494
transform 1 0 3114 0 -1 644
box 0 0 19 49
use FILL  FILL_OR2X2_185
timestamp 1516325494
transform -1 0 3141 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_185
timestamp 1516325494
transform -1 0 3160 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_2051
timestamp 1516325494
transform 1 0 3160 0 -1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_705
timestamp 1516325494
transform 1 0 3179 0 -1 644
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_711
timestamp 1516325494
transform 1 0 3232 0 -1 644
box 0 0 53 49
use INVX1  INVX1_325
timestamp 1516325494
transform 1 0 3285 0 -1 644
box 0 0 11 49
use INVX1  INVX1_328
timestamp 1516325494
transform 1 0 3297 0 -1 644
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_330
timestamp 1516325494
transform 1 0 3308 0 -1 644
box 0 0 53 49
use MUX2X1  MUX2X1_362
timestamp 1516325494
transform 1 0 3361 0 -1 644
box 0 0 30 49
use FILL  FILL_OR2X2_184
timestamp 1516325494
transform -1 0 3400 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_184
timestamp 1516325494
transform -1 0 3418 0 -1 644
box 0 0 19 49
use OR2X2  OR2X2_281
timestamp 1516325494
transform -1 0 3437 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_301
timestamp 1516325494
transform -1 0 3456 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1841
timestamp 1516325494
transform 1 0 3456 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_300
timestamp 1516325494
transform -1 0 3494 0 -1 644
box 0 0 19 49
use AND2X2  AND2X2_1840
timestamp 1516325494
transform -1 0 3513 0 -1 644
box 0 0 19 49
use MUX2X1  MUX2X1_271
timestamp 1516325494
transform 1 0 3513 0 -1 644
box 0 0 30 49
use NAND2X1  NAND2X1_271
timestamp 1516325494
transform -1 0 3559 0 -1 644
box 0 0 15 49
use FILL  FILL_OR2X2_99
timestamp 1516325494
transform -1 0 3567 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_99
timestamp 1516325494
transform -1 0 3585 0 -1 644
box 0 0 19 49
use FILL  FILL_AND2X2_105
timestamp 1516325494
transform -1 0 3593 0 -1 644
box 0 0 8 49
use AND2X2  AND2X2_105
timestamp 1516325494
transform -1 0 3612 0 -1 644
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_344
timestamp 1516325494
transform 1 0 3612 0 -1 644
box 0 0 53 49
use NAND2X1  NAND2X1_376
timestamp 1516325494
transform 1 0 3665 0 -1 644
box 0 0 15 49
use NAND2X1  NAND2X1_280
timestamp 1516325494
transform 1 0 3680 0 -1 644
box 0 0 15 49
use MUX2X1  MUX2X1_280
timestamp 1516325494
transform -1 0 3726 0 -1 644
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_786
timestamp 1516325494
transform 1 0 3726 0 -1 644
box 0 0 53 49
use NOR2X1  NOR2X1_134
timestamp 1516325494
transform -1 0 3794 0 -1 644
box 0 0 15 49
use NOR2X1  NOR2X1_133
timestamp 1516325494
transform 1 0 3794 0 -1 644
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_787
timestamp 1516325494
transform -1 0 3863 0 -1 644
box 0 0 53 49
use FILL  FILL_13_1
timestamp 1516325494
transform -1 0 3871 0 -1 644
box 0 0 8 49
use OR2X2  OR2X2_532
timestamp 1516325494
transform -1 0 21 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_629
timestamp 1516325494
transform -1 0 40 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_739
timestamp 1516325494
transform 1 0 40 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_501
timestamp 1516325494
transform 1 0 59 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_447
timestamp 1516325494
transform -1 0 97 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_498
timestamp 1516325494
transform -1 0 116 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_497
timestamp 1516325494
transform -1 0 135 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_614
timestamp 1516325494
transform -1 0 154 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_613
timestamp 1516325494
transform -1 0 173 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_444
timestamp 1516325494
transform -1 0 192 0 1 545
box 0 0 19 49
use FILL  FILL_BUFX2_545
timestamp 1516325494
transform 1 0 192 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_545
timestamp 1516325494
transform 1 0 200 0 1 545
box 0 0 15 49
use FILL  FILL_BUFX2_74
timestamp 1516325494
transform 1 0 215 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_74
timestamp 1516325494
transform 1 0 222 0 1 545
box 0 0 15 49
use FILL  FILL_BUFX2_543
timestamp 1516325494
transform 1 0 238 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_543
timestamp 1516325494
transform 1 0 245 0 1 545
box 0 0 15 49
use AND2X2  AND2X2_545
timestamp 1516325494
transform -1 0 279 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_475
timestamp 1516325494
transform 1 0 279 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_544
timestamp 1516325494
transform -1 0 317 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_546
timestamp 1516325494
transform 1 0 317 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_655
timestamp 1516325494
transform 1 0 336 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_555
timestamp 1516325494
transform -1 0 374 0 1 545
box 0 0 19 49
use MUX2X1  MUX2X1_659
timestamp 1516325494
transform 1 0 374 0 1 545
box 0 0 30 49
use AND2X2  AND2X2_466
timestamp 1516325494
transform -1 0 424 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_427
timestamp 1516325494
transform -1 0 443 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_465
timestamp 1516325494
transform -1 0 462 0 1 545
box 0 0 19 49
use MUX2X1  MUX2X1_655
timestamp 1516325494
transform -1 0 492 0 1 545
box 0 0 30 49
use OR2X2  OR2X2_476
timestamp 1516325494
transform 1 0 492 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_548
timestamp 1516325494
transform -1 0 530 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_467
timestamp 1516325494
transform 1 0 530 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_428
timestamp 1516325494
transform -1 0 568 0 1 545
box 0 0 19 49
use MUX2X1  MUX2X1_676
timestamp 1516325494
transform -1 0 598 0 1 545
box 0 0 30 49
use AND2X2  AND2X2_468
timestamp 1516325494
transform -1 0 618 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_545
timestamp 1516325494
transform -1 0 637 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_816
timestamp 1516325494
transform 1 0 637 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_685
timestamp 1516325494
transform -1 0 675 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_664
timestamp 1516325494
transform 1 0 675 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_501
timestamp 1516325494
transform -1 0 713 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_725
timestamp 1516325494
transform -1 0 732 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_543
timestamp 1516325494
transform -1 0 751 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_410
timestamp 1516325494
transform -1 0 770 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_437
timestamp 1516325494
transform -1 0 789 0 1 545
box 0 0 19 49
use NAND3X1  NAND3X1_31
timestamp 1516325494
transform 1 0 789 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_436
timestamp 1516325494
transform -1 0 827 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_572
timestamp 1516325494
transform -1 0 846 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_495
timestamp 1516325494
transform 1 0 846 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_570
timestamp 1516325494
transform 1 0 865 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_497
timestamp 1516325494
transform -1 0 903 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_573
timestamp 1516325494
transform -1 0 922 0 1 545
box 0 0 19 49
use INVX1  INVX1_150
timestamp 1516325494
transform -1 0 933 0 1 545
box 0 0 11 49
use INVX1  INVX1_215
timestamp 1516325494
transform 1 0 933 0 1 545
box 0 0 11 49
use MUX2X1  MUX2X1_793
timestamp 1516325494
transform -1 0 974 0 1 545
box 0 0 30 49
use FILL  FILL_BUFX2_779
timestamp 1516325494
transform 1 0 975 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_779
timestamp 1516325494
transform 1 0 982 0 1 545
box 0 0 15 49
use FILL  FILL_OR2X2_192
timestamp 1516325494
transform -1 0 1006 0 1 545
box 0 0 8 49
use OR2X2  OR2X2_192
timestamp 1516325494
transform -1 0 1024 0 1 545
box 0 0 19 49
use FILL  FILL_OR2X2_191
timestamp 1516325494
transform -1 0 1032 0 1 545
box 0 0 8 49
use OR2X2  OR2X2_191
timestamp 1516325494
transform -1 0 1051 0 1 545
box 0 0 19 49
use FILL  FILL_OR2X2_190
timestamp 1516325494
transform -1 0 1059 0 1 545
box 0 0 8 49
use OR2X2  OR2X2_190
timestamp 1516325494
transform -1 0 1077 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_204
timestamp 1516325494
transform -1 0 1085 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_204
timestamp 1516325494
transform -1 0 1104 0 1 545
box 0 0 19 49
use OAI21X1  OAI21X1_52
timestamp 1516325494
transform 1 0 1104 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1696
timestamp 1516325494
transform 1 0 1123 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1521
timestamp 1516325494
transform 1 0 1142 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1523
timestamp 1516325494
transform 1 0 1161 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1522
timestamp 1516325494
transform -1 0 1199 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1552
timestamp 1516325494
transform -1 0 1218 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1516
timestamp 1516325494
transform -1 0 1237 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1690
timestamp 1516325494
transform -1 0 1256 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1692
timestamp 1516325494
transform -1 0 1275 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_202
timestamp 1516325494
transform 1 0 1275 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_202
timestamp 1516325494
transform 1 0 1283 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1693
timestamp 1516325494
transform -1 0 1321 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1644
timestamp 1516325494
transform -1 0 1340 0 1 545
box 0 0 19 49
use FILL  FILL_OR2X2_189
timestamp 1516325494
transform -1 0 1348 0 1 545
box 0 0 8 49
use OR2X2  OR2X2_189
timestamp 1516325494
transform -1 0 1366 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_201
timestamp 1516325494
transform -1 0 1374 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_201
timestamp 1516325494
transform -1 0 1393 0 1 545
box 0 0 19 49
use FILL  FILL_BUFX2_457
timestamp 1516325494
transform 1 0 1393 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_457
timestamp 1516325494
transform 1 0 1400 0 1 545
box 0 0 15 49
use OR2X2  OR2X2_1771
timestamp 1516325494
transform 1 0 1416 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1497
timestamp 1516325494
transform -1 0 1454 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1262
timestamp 1516325494
transform -1 0 1473 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1261
timestamp 1516325494
transform -1 0 1492 0 1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_585
timestamp 1516325494
transform 1 0 1492 0 1 545
box 0 0 53 49
use NAND2X1  NAND2X1_9
timestamp 1516325494
transform 1 0 1545 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_9
timestamp 1516325494
transform -1 0 1590 0 1 545
box 0 0 30 49
use MUX2X1  MUX2X1_872
timestamp 1516325494
transform -1 0 1620 0 1 545
box 0 0 30 49
use NAND2X1  NAND2X1_927
timestamp 1516325494
transform -1 0 1636 0 1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_369
timestamp 1516325494
transform -1 0 1689 0 1 545
box 0 0 53 49
use OR2X2  OR2X2_1512
timestamp 1516325494
transform 1 0 1689 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1723
timestamp 1516325494
transform -1 0 1727 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1689
timestamp 1516325494
transform -1 0 1746 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1303
timestamp 1516325494
transform -1 0 1765 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1334
timestamp 1516325494
transform -1 0 1784 0 1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_459
timestamp 1516325494
transform 1 0 1784 0 1 545
box 0 0 53 49
use NAND2X1  NAND2X1_331
timestamp 1516325494
transform 1 0 1837 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_331
timestamp 1516325494
transform -1 0 1883 0 1 545
box 0 0 30 49
use FILL  FILL_BUFX2_722
timestamp 1516325494
transform 1 0 1883 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_722
timestamp 1516325494
transform 1 0 1891 0 1 545
box 0 0 15 49
use OR2X2  OR2X2_1267
timestamp 1516325494
transform -1 0 1925 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1513
timestamp 1516325494
transform -1 0 1944 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1264
timestamp 1516325494
transform -1 0 1963 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1691
timestamp 1516325494
transform -1 0 1982 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1515
timestamp 1516325494
transform -1 0 2001 0 1 545
box 0 0 19 49
use NAND2X1  NAND2X1_145
timestamp 1516325494
transform -1 0 2016 0 1 545
box 0 0 15 49
use FILL  FILL_BUFX2_414
timestamp 1516325494
transform -1 0 2024 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_414
timestamp 1516325494
transform -1 0 2039 0 1 545
box 0 0 15 49
use NAND2X1  NAND2X1_177
timestamp 1516325494
transform 1 0 2039 0 1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_401
timestamp 1516325494
transform 1 0 2054 0 1 545
box 0 0 53 49
use MUX2X1  MUX2X1_177
timestamp 1516325494
transform -1 0 2137 0 1 545
box 0 0 30 49
use OR2X2  OR2X2_1514
timestamp 1516325494
transform -1 0 2157 0 1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_465
timestamp 1516325494
transform 1 0 2157 0 1 545
box 0 0 53 49
use NAND2X1  NAND2X1_337
timestamp 1516325494
transform 1 0 2210 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_337
timestamp 1516325494
transform -1 0 2255 0 1 545
box 0 0 30 49
use MUX2X1  MUX2X1_80
timestamp 1516325494
transform 1 0 2255 0 1 545
box 0 0 30 49
use NAND2X1  NAND2X1_80
timestamp 1516325494
transform -1 0 2301 0 1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_112
timestamp 1516325494
transform -1 0 2354 0 1 545
box 0 0 53 49
use FILL  FILL_BUFX2_752
timestamp 1516325494
transform 1 0 2354 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_752
timestamp 1516325494
transform 1 0 2362 0 1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_19
timestamp 1516325494
transform 1 0 2377 0 1 545
box 0 0 53 49
use NAND2X1  NAND2X1_115
timestamp 1516325494
transform 1 0 2430 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_115
timestamp 1516325494
transform -1 0 2475 0 1 545
box 0 0 30 49
use OR2X2  OR2X2_1453
timestamp 1516325494
transform 1 0 2476 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1643
timestamp 1516325494
transform 1 0 2495 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1737
timestamp 1516325494
transform 1 0 2514 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1574
timestamp 1516325494
transform -1 0 2552 0 1 545
box 0 0 19 49
use FILL  FILL_BUFX2_193
timestamp 1516325494
transform 1 0 2552 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_193
timestamp 1516325494
transform 1 0 2559 0 1 545
box 0 0 15 49
use OR2X2  OR2X2_1452
timestamp 1516325494
transform -1 0 2594 0 1 545
box 0 0 19 49
use FILL  FILL_BUFX2_506
timestamp 1516325494
transform 1 0 2594 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_506
timestamp 1516325494
transform 1 0 2601 0 1 545
box 0 0 15 49
use FILL  FILL_BUFX2_315
timestamp 1516325494
transform -1 0 2624 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_315
timestamp 1516325494
transform -1 0 2639 0 1 545
box 0 0 15 49
use FILL  FILL_BUFX2_411
timestamp 1516325494
transform 1 0 2639 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_411
timestamp 1516325494
transform 1 0 2647 0 1 545
box 0 0 15 49
use FILL  FILL_BUFX2_210
timestamp 1516325494
transform -1 0 2670 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_210
timestamp 1516325494
transform -1 0 2685 0 1 545
box 0 0 15 49
use NAND2X1  NAND2X1_925
timestamp 1516325494
transform 1 0 2685 0 1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_367
timestamp 1516325494
transform 1 0 2700 0 1 545
box 0 0 53 49
use MUX2X1  MUX2X1_870
timestamp 1516325494
transform -1 0 2783 0 1 545
box 0 0 30 49
use AND2X2  AND2X2_626
timestamp 1516325494
transform 1 0 2 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_529
timestamp 1516325494
transform -1 0 40 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_625
timestamp 1516325494
transform -1 0 59 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_530
timestamp 1516325494
transform -1 0 78 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_445
timestamp 1516325494
transform 1 0 78 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_533
timestamp 1516325494
transform -1 0 116 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_631
timestamp 1516325494
transform -1 0 135 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_632
timestamp 1516325494
transform -1 0 154 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_534
timestamp 1516325494
transform -1 0 173 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_635
timestamp 1516325494
transform -1 0 192 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_634
timestamp 1516325494
transform -1 0 211 0 -1 545
box 0 0 19 49
use FILL  FILL_BUFX2_73
timestamp 1516325494
transform 1 0 211 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_73
timestamp 1516325494
transform 1 0 219 0 -1 545
box 0 0 15 49
use AND2X2  AND2X2_653
timestamp 1516325494
transform -1 0 253 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_553
timestamp 1516325494
transform 1 0 253 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_654
timestamp 1516325494
transform -1 0 291 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_819
timestamp 1516325494
transform -1 0 310 0 -1 545
box 0 0 19 49
use MUX2X1  MUX2X1_658
timestamp 1516325494
transform 1 0 310 0 -1 545
box 0 0 30 49
use OR2X2  OR2X2_554
timestamp 1516325494
transform -1 0 359 0 -1 545
box 0 0 19 49
use XNOR2X1  XNOR2X1_1
timestamp 1516325494
transform -1 0 393 0 -1 545
box 0 0 34 49
use XOR2X1  XOR2X1_3
timestamp 1516325494
transform 1 0 393 0 -1 545
box 0 0 34 49
use AND2X2  AND2X2_464
timestamp 1516325494
transform 1 0 428 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_547
timestamp 1516325494
transform 1 0 447 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_537
timestamp 1516325494
transform 1 0 466 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_472
timestamp 1516325494
transform 1 0 485 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_538
timestamp 1516325494
transform -1 0 523 0 -1 545
box 0 0 19 49
use MUX2X1  MUX2X1_677
timestamp 1516325494
transform 1 0 523 0 -1 545
box 0 0 30 49
use MUX2X1  MUX2X1_649
timestamp 1516325494
transform -1 0 583 0 -1 545
box 0 0 30 49
use OR2X2  OR2X2_415
timestamp 1516325494
transform -1 0 602 0 -1 545
box 0 0 19 49
use FILL  FILL_BUFX2_77
timestamp 1516325494
transform 1 0 602 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_77
timestamp 1516325494
transform 1 0 610 0 -1 545
box 0 0 15 49
use AND2X2  AND2X2_750
timestamp 1516325494
transform 1 0 625 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_624
timestamp 1516325494
transform -1 0 663 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_862
timestamp 1516325494
transform -1 0 682 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_861
timestamp 1516325494
transform 1 0 682 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_411
timestamp 1516325494
transform -1 0 720 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_438
timestamp 1516325494
transform -1 0 739 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_431
timestamp 1516325494
transform -1 0 758 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_406
timestamp 1516325494
transform 1 0 758 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_434
timestamp 1516325494
transform -1 0 796 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_571
timestamp 1516325494
transform 1 0 796 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_496
timestamp 1516325494
transform 1 0 815 0 -1 545
box 0 0 19 49
use MUX2X1  MUX2X1_762
timestamp 1516325494
transform -1 0 864 0 -1 545
box 0 0 30 49
use INVX1  INVX1_149
timestamp 1516325494
transform -1 0 876 0 -1 545
box 0 0 11 49
use MUX2X1  MUX2X1_761
timestamp 1516325494
transform 1 0 876 0 -1 545
box 0 0 30 49
use OR2X2  OR2X2_1343
timestamp 1516325494
transform 1 0 906 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1342
timestamp 1516325494
transform -1 0 944 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1341
timestamp 1516325494
transform -1 0 963 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_1558
timestamp 1516325494
transform -1 0 982 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_1556
timestamp 1516325494
transform -1 0 1001 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_113
timestamp 1516325494
transform 1 0 1001 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_113
timestamp 1516325494
transform 1 0 1009 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1462
timestamp 1516325494
transform -1 0 1047 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_173
timestamp 1516325494
transform -1 0 1055 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_173
timestamp 1516325494
transform -1 0 1074 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_1648
timestamp 1516325494
transform 1 0 1074 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1461
timestamp 1516325494
transform 1 0 1093 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1336
timestamp 1516325494
transform -1 0 1131 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_1554
timestamp 1516325494
transform -1 0 1150 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_112
timestamp 1516325494
transform -1 0 1158 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_112
timestamp 1516325494
transform -1 0 1176 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_111
timestamp 1516325494
transform -1 0 1184 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_111
timestamp 1516325494
transform -1 0 1203 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1456
timestamp 1516325494
transform -1 0 1222 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_1646
timestamp 1516325494
transform -1 0 1241 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_172
timestamp 1516325494
transform -1 0 1249 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_172
timestamp 1516325494
transform -1 0 1267 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_171
timestamp 1516325494
transform -1 0 1275 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_171
timestamp 1516325494
transform -1 0 1294 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1517
timestamp 1516325494
transform 1 0 1294 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1518
timestamp 1516325494
transform -1 0 1332 0 -1 545
box 0 0 19 49
use NAND2X1  NAND2X1_113
timestamp 1516325494
transform 1 0 1332 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_113
timestamp 1516325494
transform -1 0 1377 0 -1 545
box 0 0 30 49
use AND2X2  AND2X2_1555
timestamp 1516325494
transform -1 0 1397 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1338
timestamp 1516325494
transform -1 0 1416 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1337
timestamp 1516325494
transform -1 0 1435 0 -1 545
box 0 0 19 49
use OAI21X1  OAI21X1_27
timestamp 1516325494
transform 1 0 1435 0 -1 545
box 0 0 19 49
use INVX2  INVX2_16
timestamp 1516325494
transform 1 0 1454 0 -1 545
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_363
timestamp 1516325494
transform 1 0 1465 0 -1 545
box 0 0 53 49
use AND2X2  AND2X2_1551
timestamp 1516325494
transform -1 0 1537 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1332
timestamp 1516325494
transform -1 0 1556 0 -1 545
box 0 0 19 49
use NAND2X1  NAND2X1_921
timestamp 1516325494
transform 1 0 1556 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_866
timestamp 1516325494
transform 1 0 1571 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_11
timestamp 1516325494
transform 1 0 1602 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_107
timestamp 1516325494
transform 1 0 1655 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_107
timestamp 1516325494
transform -1 0 1700 0 -1 545
box 0 0 30 49
use AND2X2  AND2X2_1553
timestamp 1516325494
transform -1 0 1720 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1335
timestamp 1516325494
transform -1 0 1739 0 -1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_75
timestamp 1516325494
transform 1 0 1739 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_139
timestamp 1516325494
transform 1 0 1792 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_139
timestamp 1516325494
transform 1 0 1807 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_368
timestamp 1516325494
transform 1 0 1837 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_926
timestamp 1516325494
transform 1 0 1891 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_871
timestamp 1516325494
transform -1 0 1936 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_681
timestamp 1516325494
transform 1 0 1936 0 -1 545
box 0 0 53 49
use MUX2X1  MUX2X1_145
timestamp 1516325494
transform 1 0 1989 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_81
timestamp 1516325494
transform -1 0 2073 0 -1 545
box 0 0 53 49
use FILL  FILL_BUFX2_790
timestamp 1516325494
transform 1 0 2073 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_790
timestamp 1516325494
transform 1 0 2081 0 -1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_113
timestamp 1516325494
transform 1 0 2096 0 -1 545
box 0 0 53 49
use AND2X2  AND2X2_1647
timestamp 1516325494
transform -1 0 2168 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1458
timestamp 1516325494
transform -1 0 2187 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1457
timestamp 1516325494
transform -1 0 2206 0 -1 545
box 0 0 19 49
use NAND2X1  NAND2X1_111
timestamp 1516325494
transform 1 0 2206 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_111
timestamp 1516325494
transform -1 0 2251 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_527
timestamp 1516325494
transform 1 0 2252 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_527
timestamp 1516325494
transform 1 0 2305 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_527
timestamp 1516325494
transform -1 0 2350 0 -1 545
box 0 0 30 49
use AND2X2  AND2X2_1645
timestamp 1516325494
transform -1 0 2369 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1454
timestamp 1516325494
transform -1 0 2388 0 -1 545
box 0 0 19 49
use FILL  FILL_BUFX2_514
timestamp 1516325494
transform 1 0 2388 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_514
timestamp 1516325494
transform 1 0 2396 0 -1 545
box 0 0 15 49
use NAND2X1  NAND2X1_335
timestamp 1516325494
transform 1 0 2411 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_335
timestamp 1516325494
transform -1 0 2456 0 -1 545
box 0 0 30 49
use MUX2X1  MUX2X1_339
timestamp 1516325494
transform -1 0 2487 0 -1 545
box 0 0 30 49
use NAND2X1  NAND2X1_339
timestamp 1516325494
transform -1 0 2502 0 -1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_467
timestamp 1516325494
transform -1 0 2555 0 -1 545
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_371
timestamp 1516325494
transform 1 0 2556 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_929
timestamp 1516325494
transform 1 0 2609 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_874
timestamp 1516325494
transform 1 0 2624 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_297
timestamp 1516325494
transform 1 0 2654 0 -1 545
box 0 0 53 49
use FILL  FILL_BUFX2_167
timestamp 1516325494
transform -1 0 2716 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_167
timestamp 1516325494
transform -1 0 2730 0 -1 545
box 0 0 15 49
use FILL  FILL_BUFX2_311
timestamp 1516325494
transform -1 0 2738 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_311
timestamp 1516325494
transform -1 0 2753 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_240
timestamp 1516325494
transform 1 0 2753 0 -1 545
box 0 0 30 49
use OR2X2  OR2X2_283
timestamp 1516325494
transform -1 0 2803 0 1 545
box 0 0 19 49
use FILL  FILL_BUFX2_753
timestamp 1516325494
transform -1 0 2811 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_753
timestamp 1516325494
transform -1 0 2825 0 1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_531
timestamp 1516325494
transform -1 0 2878 0 1 545
box 0 0 53 49
use FILL  FILL_BUFX2_313
timestamp 1516325494
transform -1 0 2887 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_313
timestamp 1516325494
transform -1 0 2901 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_585
timestamp 1516325494
transform -1 0 2931 0 1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_265
timestamp 1516325494
transform -1 0 2985 0 1 545
box 0 0 53 49
use FILL  FILL_AND2X2_86
timestamp 1516325494
transform 1 0 2985 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_86
timestamp 1516325494
transform 1 0 2993 0 1 545
box 0 0 19 49
use FILL  FILL_OR2X2_82
timestamp 1516325494
transform -1 0 3020 0 1 545
box 0 0 8 49
use OR2X2  OR2X2_82
timestamp 1516325494
transform -1 0 3038 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_85
timestamp 1516325494
transform -1 0 3046 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_85
timestamp 1516325494
transform -1 0 3065 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1513
timestamp 1516325494
transform 1 0 3065 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1285
timestamp 1516325494
transform -1 0 3103 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1514
timestamp 1516325494
transform -1 0 3122 0 1 545
box 0 0 19 49
use NAND2X1  NAND2X1_202
timestamp 1516325494
transform 1 0 3122 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_202
timestamp 1516325494
transform -1 0 3167 0 1 545
box 0 0 30 49
use FILL  FILL_BUFX2_526
timestamp 1516325494
transform -1 0 3175 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_526
timestamp 1516325494
transform -1 0 3190 0 1 545
box 0 0 15 49
use OR2X2  OR2X2_1497
timestamp 1516325494
transform 1 0 3190 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1496
timestamp 1516325494
transform -1 0 3228 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1676
timestamp 1516325494
transform 1 0 3228 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_192
timestamp 1516325494
transform 1 0 3247 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_192
timestamp 1516325494
transform 1 0 3255 0 1 545
box 0 0 19 49
use FILL  FILL_BUFX2_426
timestamp 1516325494
transform -1 0 3282 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_426
timestamp 1516325494
transform -1 0 3296 0 1 545
box 0 0 15 49
use NAND2X1  NAND2X1_209
timestamp 1516325494
transform 1 0 3297 0 1 545
box 0 0 15 49
use MUX2X1  MUX2X1_209
timestamp 1516325494
transform -1 0 3342 0 1 545
box 0 0 30 49
use FILL  FILL_BUFX2_839
timestamp 1516325494
transform 1 0 3342 0 1 545
box 0 0 8 49
use BUFX2  BUFX2_839
timestamp 1516325494
transform 1 0 3350 0 1 545
box 0 0 15 49
use OR2X2  OR2X2_1469
timestamp 1516325494
transform -1 0 3384 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1655
timestamp 1516325494
transform -1 0 3403 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_194
timestamp 1516325494
transform -1 0 3411 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_194
timestamp 1516325494
transform -1 0 3430 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_282
timestamp 1516325494
transform -1 0 3449 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_299
timestamp 1516325494
transform -1 0 3468 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_179
timestamp 1516325494
transform -1 0 3476 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_179
timestamp 1516325494
transform -1 0 3494 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1632
timestamp 1516325494
transform 1 0 3494 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1439
timestamp 1516325494
transform -1 0 3532 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1468
timestamp 1516325494
transform -1 0 3551 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1656
timestamp 1516325494
transform -1 0 3570 0 1 545
box 0 0 19 49
use NAND2X1  NAND2X1_368
timestamp 1516325494
transform -1 0 3585 0 1 545
box 0 0 15 49
use AND2X2  AND2X2_1657
timestamp 1516325494
transform -1 0 3604 0 1 545
box 0 0 19 49
use FILL  FILL_OR2X2_169
timestamp 1516325494
transform -1 0 3612 0 1 545
box 0 0 8 49
use OR2X2  OR2X2_169
timestamp 1516325494
transform -1 0 3631 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_180
timestamp 1516325494
transform -1 0 3639 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_180
timestamp 1516325494
transform -1 0 3658 0 1 545
box 0 0 19 49
use FILL  FILL_AND2X2_165
timestamp 1516325494
transform 1 0 3658 0 1 545
box 0 0 8 49
use AND2X2  AND2X2_165
timestamp 1516325494
transform 1 0 3665 0 1 545
box 0 0 19 49
use NAND2X1  NAND2X1_367
timestamp 1516325494
transform -1 0 3699 0 1 545
box 0 0 15 49
use AND2X2  AND2X2_1634
timestamp 1516325494
transform 1 0 3699 0 1 545
box 0 0 19 49
use OR2X2  OR2X2_1438
timestamp 1516325494
transform -1 0 3737 0 1 545
box 0 0 19 49
use AND2X2  AND2X2_1633
timestamp 1516325494
transform 1 0 3737 0 1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_143
timestamp 1516325494
transform -1 0 3809 0 1 545
box 0 0 53 49
use NAND2X1  NAND2X1_240
timestamp 1516325494
transform -1 0 2799 0 -1 545
box 0 0 15 49
use NAND2X1  NAND2X1_248
timestamp 1516325494
transform 1 0 2799 0 -1 545
box 0 0 15 49
use FILL  FILL_BUFX2_424
timestamp 1516325494
transform 1 0 2814 0 -1 545
box 0 0 8 49
use BUFX2  BUFX2_424
timestamp 1516325494
transform 1 0 2822 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_248
timestamp 1516325494
transform -1 0 2867 0 -1 545
box 0 0 30 49
use MUX2X1  MUX2X1_234
timestamp 1516325494
transform 1 0 2867 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_170
timestamp 1516325494
transform -1 0 2951 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_234
timestamp 1516325494
transform -1 0 2966 0 -1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_202
timestamp 1516325494
transform 1 0 2966 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_618
timestamp 1516325494
transform 1 0 3019 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_618
timestamp 1516325494
transform -1 0 3064 0 -1 545
box 0 0 30 49
use AND2X2  AND2X2_1674
timestamp 1516325494
transform 1 0 3065 0 -1 545
box 0 0 19 49
use AND2X2  AND2X2_1675
timestamp 1516325494
transform 1 0 3084 0 -1 545
box 0 0 19 49
use OR2X2  OR2X2_1495
timestamp 1516325494
transform 1 0 3103 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_191
timestamp 1516325494
transform 1 0 3122 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_191
timestamp 1516325494
transform 1 0 3129 0 -1 545
box 0 0 19 49
use FILL  FILL_OR2X2_180
timestamp 1516325494
transform -1 0 3156 0 -1 545
box 0 0 8 49
use OR2X2  OR2X2_180
timestamp 1516325494
transform -1 0 3175 0 -1 545
box 0 0 19 49
use FILL  FILL_AND2X2_190
timestamp 1516325494
transform -1 0 3183 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_190
timestamp 1516325494
transform -1 0 3202 0 -1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_241
timestamp 1516325494
transform 1 0 3202 0 -1 545
box 0 0 53 49
use NAND2X1  NAND2X1_241
timestamp 1516325494
transform 1 0 3255 0 -1 545
box 0 0 15 49
use MUX2X1  MUX2X1_241
timestamp 1516325494
transform -1 0 3300 0 -1 545
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_177
timestamp 1516325494
transform -1 0 3353 0 -1 545
box 0 0 53 49
use DFFNEGX1  DFFNEGX1_1
timestamp 1516325494
transform 1 0 3354 0 -1 545
box 0 0 57 49
use FILL  FILL_OR2X2_170
timestamp 1516325494
transform -1 0 3419 0 -1 545
box 0 0 8 49
use OR2X2  OR2X2_170
timestamp 1516325494
transform -1 0 3437 0 -1 545
box 0 0 19 49
use MUX2X1  MUX2X1_272
timestamp 1516325494
transform 1 0 3437 0 -1 545
box 0 0 30 49
use NAND2X1  NAND2X1_272
timestamp 1516325494
transform -1 0 3483 0 -1 545
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_144
timestamp 1516325494
transform -1 0 3536 0 -1 545
box 0 0 53 49
use MUX2X1  MUX2X1_368
timestamp 1516325494
transform 1 0 3536 0 -1 545
box 0 0 30 49
use MUX2X1  MUX2X1_367
timestamp 1516325494
transform 1 0 3566 0 -1 545
box 0 0 30 49
use FILL  FILL_AND2X2_166
timestamp 1516325494
transform 1 0 3597 0 -1 545
box 0 0 8 49
use AND2X2  AND2X2_166
timestamp 1516325494
transform 1 0 3604 0 -1 545
box 0 0 19 49
use FILL  FILL_OR2X2_155
timestamp 1516325494
transform -1 0 3631 0 -1 545
box 0 0 8 49
use OR2X2  OR2X2_155
timestamp 1516325494
transform -1 0 3650 0 -1 545
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_768
timestamp 1516325494
transform 1 0 3650 0 -1 545
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_769
timestamp 1516325494
transform -1 0 3756 0 -1 545
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_717
timestamp 1516325494
transform 1 0 3756 0 -1 545
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_152
timestamp 1516325494
transform -1 0 3863 0 1 545
box 0 0 53 49
use FILL  FILL_12_1
timestamp 1516325494
transform 1 0 3863 0 1 545
box 0 0 8 49
use DFFPOSX1  DFFPOSX1_753
timestamp 1516325494
transform -1 0 3863 0 -1 545
box 0 0 53 49
use FILL  FILL_11_1
timestamp 1516325494
transform -1 0 3871 0 -1 545
box 0 0 8 49
use OR2X2  OR2X2_448
timestamp 1516325494
transform -1 0 21 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_503
timestamp 1516325494
transform -1 0 40 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_531
timestamp 1516325494
transform -1 0 59 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_627
timestamp 1516325494
transform -1 0 78 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_628
timestamp 1516325494
transform -1 0 97 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_504
timestamp 1516325494
transform -1 0 116 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_449
timestamp 1516325494
transform -1 0 135 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_506
timestamp 1516325494
transform -1 0 154 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_834
timestamp 1516325494
transform 1 0 154 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_541
timestamp 1516325494
transform -1 0 192 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_738
timestamp 1516325494
transform 1 0 192 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_617
timestamp 1516325494
transform -1 0 230 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_843
timestamp 1516325494
transform -1 0 249 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_598
timestamp 1516325494
transform 1 0 249 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_801
timestamp 1516325494
transform 1 0 268 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_673
timestamp 1516325494
transform -1 0 306 0 1 446
box 0 0 19 49
use FILL  FILL_BUFX2_697
timestamp 1516325494
transform 1 0 306 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_697
timestamp 1516325494
transform 1 0 314 0 1 446
box 0 0 15 49
use OR2X2  OR2X2_639
timestamp 1516325494
transform 1 0 329 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_767
timestamp 1516325494
transform 1 0 348 0 1 446
box 0 0 19 49
use NAND3X1  NAND3X1_42
timestamp 1516325494
transform -1 0 386 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_470
timestamp 1516325494
transform 1 0 386 0 1 446
box 0 0 19 49
use NAND3X1  NAND3X1_57
timestamp 1516325494
transform -1 0 424 0 1 446
box 0 0 19 49
use NOR2X1  NOR2X1_28
timestamp 1516325494
transform 1 0 424 0 1 446
box 0 0 15 49
use OR2X2  OR2X2_573
timestamp 1516325494
transform 1 0 439 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_564
timestamp 1516325494
transform 1 0 458 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_562
timestamp 1516325494
transform -1 0 496 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_561
timestamp 1516325494
transform -1 0 515 0 1 446
box 0 0 19 49
use NAND3X1  NAND3X1_32
timestamp 1516325494
transform 1 0 515 0 1 446
box 0 0 19 49
use NOR2X1  NOR2X1_33
timestamp 1516325494
transform -1 0 549 0 1 446
box 0 0 15 49
use AND2X2  AND2X2_815
timestamp 1516325494
transform 1 0 549 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_686
timestamp 1516325494
transform 1 0 568 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_687
timestamp 1516325494
transform 1 0 587 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_645
timestamp 1516325494
transform 1 0 606 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_601
timestamp 1516325494
transform 1 0 625 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_726
timestamp 1516325494
transform 1 0 644 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_724
timestamp 1516325494
transform 1 0 663 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_699
timestamp 1516325494
transform 1 0 682 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_435
timestamp 1516325494
transform 1 0 701 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_409
timestamp 1516325494
transform -1 0 739 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_432
timestamp 1516325494
transform -1 0 758 0 1 446
box 0 0 19 49
use INVX1  INVX1_4
timestamp 1516325494
transform -1 0 769 0 1 446
box 0 0 11 49
use AND2X2  AND2X2_433
timestamp 1516325494
transform -1 0 789 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_576
timestamp 1516325494
transform -1 0 808 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_586
timestamp 1516325494
transform -1 0 827 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_697
timestamp 1516325494
transform -1 0 846 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1494
timestamp 1516325494
transform -1 0 865 0 1 446
box 0 0 19 49
use MUX2X1  MUX2X1_792
timestamp 1516325494
transform -1 0 895 0 1 446
box 0 0 30 49
use MUX2X1  MUX2X1_788
timestamp 1516325494
transform 1 0 895 0 1 446
box 0 0 30 49
use FILL  FILL_OR2X2_179
timestamp 1516325494
transform -1 0 933 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_179
timestamp 1516325494
transform -1 0 952 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_107
timestamp 1516325494
transform -1 0 960 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_107
timestamp 1516325494
transform -1 0 979 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1464
timestamp 1516325494
transform -1 0 998 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1463
timestamp 1516325494
transform -1 0 1017 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_106
timestamp 1516325494
transform -1 0 1025 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_106
timestamp 1516325494
transform -1 0 1043 0 1 446
box 0 0 19 49
use FILL  FILL_AND2X2_114
timestamp 1516325494
transform -1 0 1051 0 1 446
box 0 0 8 49
use AND2X2  AND2X2_114
timestamp 1516325494
transform -1 0 1070 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_162
timestamp 1516325494
transform -1 0 1078 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_162
timestamp 1516325494
transform -1 0 1096 0 1 446
box 0 0 19 49
use AND2X2  AND2X2_1650
timestamp 1516325494
transform -1 0 1115 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1997
timestamp 1516325494
transform 1 0 1115 0 1 446
box 0 0 19 49
use FILL  FILL_AND2X2_174
timestamp 1516325494
transform -1 0 1142 0 1 446
box 0 0 8 49
use AND2X2  AND2X2_174
timestamp 1516325494
transform -1 0 1161 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_105
timestamp 1516325494
transform -1 0 1169 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_105
timestamp 1516325494
transform -1 0 1188 0 1 446
box 0 0 19 49
use FILL  FILL_BUFX2_566
timestamp 1516325494
transform -1 0 1196 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_566
timestamp 1516325494
transform -1 0 1210 0 1 446
box 0 0 15 49
use FILL  FILL_BUFX2_274
timestamp 1516325494
transform 1 0 1210 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_274
timestamp 1516325494
transform 1 0 1218 0 1 446
box 0 0 15 49
use FILL  FILL_OR2X2_161
timestamp 1516325494
transform -1 0 1241 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_161
timestamp 1516325494
transform -1 0 1260 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1871
timestamp 1516325494
transform 1 0 1260 0 1 446
box 0 0 19 49
use FILL  FILL_BUFX2_277
timestamp 1516325494
transform -1 0 1287 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_277
timestamp 1516325494
transform -1 0 1301 0 1 446
box 0 0 15 49
use AND2X2  AND2X2_378
timestamp 1516325494
transform 1 0 1302 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_354
timestamp 1516325494
transform 1 0 1321 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_398
timestamp 1516325494
transform 1 0 1340 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_356
timestamp 1516325494
transform 1 0 1359 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_17
timestamp 1516325494
transform 1 0 1378 0 1 446
box 0 0 53 49
use OAI21X1  OAI21X1_41
timestamp 1516325494
transform 1 0 1431 0 1 446
box 0 0 19 49
use INVX2  INVX2_30
timestamp 1516325494
transform 1 0 1450 0 1 446
box 0 0 11 49
use NAND2X1  NAND2X1_523
timestamp 1516325494
transform 1 0 1461 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_529
timestamp 1516325494
transform 1 0 1476 0 1 446
box 0 0 53 49
use NAND2X1  NAND2X1_529
timestamp 1516325494
transform 1 0 1530 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_529
timestamp 1516325494
transform -1 0 1575 0 1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_425
timestamp 1516325494
transform 1 0 1575 0 1 446
box 0 0 53 49
use NAND2X1  NAND2X1_393
timestamp 1516325494
transform 1 0 1628 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_393
timestamp 1516325494
transform -1 0 1674 0 1 446
box 0 0 30 49
use NAND2X1  NAND2X1_184
timestamp 1516325494
transform -1 0 1689 0 1 446
box 0 0 15 49
use OR2X2  OR2X2_1333
timestamp 1516325494
transform -1 0 1708 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_408
timestamp 1516325494
transform -1 0 1761 0 1 446
box 0 0 53 49
use FILL  FILL_BUFX2_312
timestamp 1516325494
transform 1 0 1761 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_312
timestamp 1516325494
transform 1 0 1769 0 1 446
box 0 0 15 49
use FILL  FILL_BUFX2_190
timestamp 1516325494
transform -1 0 1792 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_190
timestamp 1516325494
transform -1 0 1807 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_394
timestamp 1516325494
transform 1 0 1807 0 1 446
box 0 0 53 49
use NAND2X1  NAND2X1_170
timestamp 1516325494
transform 1 0 1860 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_170
timestamp 1516325494
transform -1 0 1905 0 1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_41
timestamp 1516325494
transform 1 0 1906 0 1 446
box 0 0 53 49
use NAND2X1  NAND2X1_425
timestamp 1516325494
transform 1 0 1959 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_425
timestamp 1516325494
transform -1 0 2004 0 1 446
box 0 0 30 49
use NAND2X1  NAND2X1_297
timestamp 1516325494
transform 1 0 2005 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_297
timestamp 1516325494
transform -1 0 2050 0 1 446
box 0 0 30 49
use AND2X2  AND2X2_1695
timestamp 1516325494
transform -1 0 2069 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1520
timestamp 1516325494
transform -1 0 2088 0 1 446
box 0 0 19 49
use FILL  FILL_BUFX2_23
timestamp 1516325494
transform 1 0 2088 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_23
timestamp 1516325494
transform 1 0 2096 0 1 446
box 0 0 15 49
use NAND2X1  NAND2X1_81
timestamp 1516325494
transform 1 0 2111 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_81
timestamp 1516325494
transform -1 0 2156 0 1 446
box 0 0 30 49
use AND2X2  AND2X2_1741
timestamp 1516325494
transform -1 0 2176 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1580
timestamp 1516325494
transform -1 0 2195 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_15
timestamp 1516325494
transform 1 0 2195 0 1 446
box 0 0 53 49
use FILL  FILL_BUFX2_352
timestamp 1516325494
transform -1 0 2256 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_352
timestamp 1516325494
transform -1 0 2270 0 1 446
box 0 0 15 49
use OR2X2  OR2X2_1579
timestamp 1516325494
transform -1 0 2290 0 1 446
box 0 0 19 49
use FILL  FILL_BUFX2_33
timestamp 1516325494
transform 1 0 2290 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_33
timestamp 1516325494
transform 1 0 2297 0 1 446
box 0 0 15 49
use NAND2X1  NAND2X1_563
timestamp 1516325494
transform 1 0 2312 0 1 446
box 0 0 15 49
use OR2X2  OR2X2_446
timestamp 1516325494
transform -1 0 21 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_499
timestamp 1516325494
transform -1 0 40 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_500
timestamp 1516325494
transform -1 0 59 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_437
timestamp 1516325494
transform -1 0 78 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_484
timestamp 1516325494
transform -1 0 97 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_483
timestamp 1516325494
transform -1 0 116 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_507
timestamp 1516325494
transform 1 0 116 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_674
timestamp 1516325494
transform 1 0 135 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_675
timestamp 1516325494
transform 1 0 154 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_614
timestamp 1516325494
transform 1 0 173 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_519
timestamp 1516325494
transform 1 0 192 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_599
timestamp 1516325494
transform -1 0 230 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_515
timestamp 1516325494
transform 1 0 230 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_514
timestamp 1516325494
transform -1 0 268 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_597
timestamp 1516325494
transform -1 0 287 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_596
timestamp 1516325494
transform -1 0 306 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_696
timestamp 1516325494
transform 1 0 306 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_696
timestamp 1516325494
transform 1 0 314 0 -1 446
box 0 0 15 49
use AND2X2  AND2X2_516
timestamp 1516325494
transform -1 0 348 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_515
timestamp 1516325494
transform -1 0 367 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_457
timestamp 1516325494
transform 1 0 367 0 -1 446
box 0 0 19 49
use AOI21X1  AOI21X1_4
timestamp 1516325494
transform 1 0 386 0 -1 446
box 0 0 19 49
use MUX2X1  MUX2X1_664
timestamp 1516325494
transform -1 0 435 0 -1 446
box 0 0 30 49
use MUX2X1  MUX2X1_665
timestamp 1516325494
transform 1 0 435 0 -1 446
box 0 0 30 49
use MUX2X1  MUX2X1_663
timestamp 1516325494
transform -1 0 496 0 -1 446
box 0 0 30 49
use AND2X2  AND2X2_480
timestamp 1516325494
transform 1 0 496 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_434
timestamp 1516325494
transform 1 0 515 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_435
timestamp 1516325494
transform -1 0 553 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_479
timestamp 1516325494
transform 1 0 553 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_563
timestamp 1516325494
transform -1 0 591 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_814
timestamp 1516325494
transform -1 0 610 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_695
timestamp 1516325494
transform 1 0 610 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_695
timestamp 1516325494
transform 1 0 618 0 -1 446
box 0 0 15 49
use OR2X2  OR2X2_544
timestamp 1516325494
transform -1 0 652 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_584
timestamp 1516325494
transform -1 0 671 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_398
timestamp 1516325494
transform -1 0 679 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_398
timestamp 1516325494
transform -1 0 693 0 -1 446
box 0 0 15 49
use AND2X2  AND2X2_643
timestamp 1516325494
transform -1 0 713 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_658
timestamp 1516325494
transform 1 0 713 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_407
timestamp 1516325494
transform -1 0 751 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_577
timestamp 1516325494
transform -1 0 770 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_575
timestamp 1516325494
transform 1 0 770 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_498
timestamp 1516325494
transform 1 0 789 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_698
timestamp 1516325494
transform 1 0 808 0 -1 446
box 0 0 19 49
use INVX1  INVX1_210
timestamp 1516325494
transform 1 0 827 0 -1 446
box 0 0 11 49
use OR2X2  OR2X2_1493
timestamp 1516325494
transform 1 0 838 0 -1 446
box 0 0 19 49
use OAI21X1  OAI21X1_32
timestamp 1516325494
transform 1 0 857 0 -1 446
box 0 0 19 49
use INVX2  INVX2_21
timestamp 1516325494
transform 1 0 876 0 -1 446
box 0 0 11 49
use INVX1  INVX1_214
timestamp 1516325494
transform -1 0 898 0 -1 446
box 0 0 11 49
use FILL  FILL_OR2X2_165
timestamp 1516325494
transform -1 0 907 0 -1 446
box 0 0 8 49
use OR2X2  OR2X2_165
timestamp 1516325494
transform -1 0 925 0 -1 446
box 0 0 19 49
use FILL  FILL_OR2X2_164
timestamp 1516325494
transform -1 0 933 0 -1 446
box 0 0 8 49
use OR2X2  OR2X2_164
timestamp 1516325494
transform -1 0 952 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_570
timestamp 1516325494
transform 1 0 952 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_570
timestamp 1516325494
transform 1 0 960 0 -1 446
box 0 0 15 49
use FILL  FILL_OR2X2_163
timestamp 1516325494
transform -1 0 983 0 -1 446
box 0 0 8 49
use OR2X2  OR2X2_163
timestamp 1516325494
transform -1 0 1001 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_582
timestamp 1516325494
transform 1 0 1001 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_582
timestamp 1516325494
transform 1 0 1009 0 -1 446
box 0 0 15 49
use OAI21X1  OAI21X1_46
timestamp 1516325494
transform 1 0 1024 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_257
timestamp 1516325494
transform 1 0 1043 0 -1 446
box 0 0 19 49
use INVX2  INVX2_35
timestamp 1516325494
transform 1 0 1062 0 -1 446
box 0 0 11 49
use AND2X2  AND2X2_2086
timestamp 1516325494
transform -1 0 1093 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1995
timestamp 1516325494
transform 1 0 1093 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_2085
timestamp 1516325494
transform -1 0 1131 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1337
timestamp 1516325494
transform 1 0 1131 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1055
timestamp 1516325494
transform -1 0 1169 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1339
timestamp 1516325494
transform -1 0 1188 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1721
timestamp 1516325494
transform 1 0 1188 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1958
timestamp 1516325494
transform -1 0 1226 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1865
timestamp 1516325494
transform -1 0 1245 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1960
timestamp 1516325494
transform -1 0 1264 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_580
timestamp 1516325494
transform -1 0 1272 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_580
timestamp 1516325494
transform -1 0 1286 0 -1 446
box 0 0 15 49
use AND2X2  AND2X2_377
timestamp 1516325494
transform 1 0 1286 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_422
timestamp 1516325494
transform -1 0 1324 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_396
timestamp 1516325494
transform 1 0 1324 0 -1 446
box 0 0 19 49
use OAI21X1  OAI21X1_28
timestamp 1516325494
transform 1 0 1343 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_2027
timestamp 1516325494
transform 1 0 1362 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1955
timestamp 1516325494
transform 1 0 1381 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1961
timestamp 1516325494
transform 1 0 1400 0 -1 446
box 0 0 19 49
use INVX2  INVX2_17
timestamp 1516325494
transform 1 0 1419 0 -1 446
box 0 0 11 49
use NAND2X1  NAND2X1_738
timestamp 1516325494
transform 1 0 1431 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_750
timestamp 1516325494
transform -1 0 1454 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_750
timestamp 1516325494
transform -1 0 1469 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_523
timestamp 1516325494
transform -1 0 1499 0 -1 446
box 0 0 30 49
use FILL  FILL_BUFX2_292
timestamp 1516325494
transform 1 0 1499 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_292
timestamp 1516325494
transform 1 0 1507 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_615
timestamp 1516325494
transform -1 0 1530 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_615
timestamp 1516325494
transform -1 0 1545 0 -1 446
box 0 0 15 49
use NAND2X1  NAND2X1_726
timestamp 1516325494
transform 1 0 1545 0 -1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_395
timestamp 1516325494
transform 1 0 1560 0 -1 446
box 0 0 53 49
use NAND2X1  NAND2X1_171
timestamp 1516325494
transform 1 0 1613 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_171
timestamp 1516325494
transform 1 0 1628 0 -1 446
box 0 0 30 49
use MUX2X1  MUX2X1_184
timestamp 1516325494
transform -1 0 1689 0 -1 446
box 0 0 30 49
use FILL  FILL_BUFX2_353
timestamp 1516325494
transform 1 0 1689 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_353
timestamp 1516325494
transform 1 0 1697 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_614
timestamp 1516325494
transform 1 0 1712 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_614
timestamp 1516325494
transform 1 0 1720 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_825
timestamp 1516325494
transform -1 0 1765 0 -1 446
box 0 0 30 49
use FILL  FILL_BUFX2_237
timestamp 1516325494
transform -1 0 1773 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_237
timestamp 1516325494
transform -1 0 1788 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_43
timestamp 1516325494
transform 1 0 1788 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_43
timestamp 1516325494
transform 1 0 1796 0 -1 446
box 0 0 15 49
use AND2X2  AND2X2_1957
timestamp 1516325494
transform -1 0 1830 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_723
timestamp 1516325494
transform 1 0 1830 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_723
timestamp 1516325494
transform 1 0 1837 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_555
timestamp 1516325494
transform 1 0 1853 0 -1 446
box 0 0 30 49
use NAND2X1  NAND2X1_555
timestamp 1516325494
transform -1 0 1898 0 -1 446
box 0 0 15 49
use AND2X2  AND2X2_1557
timestamp 1516325494
transform -1 0 1917 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1339
timestamp 1516325494
transform -1 0 1936 0 -1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_497
timestamp 1516325494
transform 1 0 1936 0 -1 446
box 0 0 53 49
use OR2X2  OR2X2_1519
timestamp 1516325494
transform 1 0 1989 0 -1 446
box 0 0 19 49
use NAND2X1  NAND2X1_561
timestamp 1516325494
transform 1 0 2008 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_561
timestamp 1516325494
transform -1 0 2054 0 -1 446
box 0 0 30 49
use OR2X2  OR2X2_1340
timestamp 1516325494
transform -1 0 2073 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1649
timestamp 1516325494
transform -1 0 2092 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1460
timestamp 1516325494
transform -1 0 2111 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1459
timestamp 1516325494
transform -1 0 2130 0 -1 446
box 0 0 19 49
use NAND2X1  NAND2X1_559
timestamp 1516325494
transform 1 0 2130 0 -1 446
box 0 0 15 49
use NAND2X1  NAND2X1_79
timestamp 1516325494
transform 1 0 2145 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_559
timestamp 1516325494
transform -1 0 2190 0 -1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_111
timestamp 1516325494
transform 1 0 2191 0 -1 446
box 0 0 53 49
use MUX2X1  MUX2X1_79
timestamp 1516325494
transform -1 0 2274 0 -1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_701
timestamp 1516325494
transform -1 0 2327 0 -1 446
box 0 0 53 49
use MUX2X1  MUX2X1_563
timestamp 1516325494
transform -1 0 2358 0 1 446
box 0 0 30 49
use OR2X2  OR2X2_1455
timestamp 1516325494
transform -1 0 2377 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_463
timestamp 1516325494
transform 1 0 2377 0 1 446
box 0 0 53 49
use MUX2X1  MUX2X1_83
timestamp 1516325494
transform 1 0 2430 0 1 446
box 0 0 30 49
use NAND2X1  NAND2X1_83
timestamp 1516325494
transform -1 0 2476 0 1 446
box 0 0 15 49
use FILL  FILL_BUFX2_71
timestamp 1516325494
transform 1 0 2476 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_71
timestamp 1516325494
transform 1 0 2483 0 1 446
box 0 0 15 49
use OR2X2  OR2X2_1575
timestamp 1516325494
transform 1 0 2499 0 1 446
box 0 0 19 49
use NAND2X1  NAND2X1_147
timestamp 1516325494
transform 1 0 2518 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_83
timestamp 1516325494
transform 1 0 2533 0 1 446
box 0 0 53 49
use MUX2X1  MUX2X1_147
timestamp 1516325494
transform 1 0 2586 0 1 446
box 0 0 30 49
use MUX2X1  MUX2X1_489
timestamp 1516325494
transform 1 0 2616 0 1 446
box 0 0 30 49
use NAND2X1  NAND2X1_489
timestamp 1516325494
transform -1 0 2662 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_767
timestamp 1516325494
transform 1 0 2662 0 1 446
box 0 0 53 49
use FILL  FILL_BUFX2_351
timestamp 1516325494
transform -1 0 2723 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_351
timestamp 1516325494
transform -1 0 2738 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_176
timestamp 1516325494
transform -1 0 2791 0 1 446
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_184
timestamp 1516325494
transform 1 0 2791 0 1 446
box 0 0 53 49
use FILL  FILL_OR2X2_166
timestamp 1516325494
transform 1 0 2844 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_166
timestamp 1516325494
transform 1 0 2852 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1440
timestamp 1516325494
transform -1 0 2890 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_168
timestamp 1516325494
transform 1 0 2890 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_168
timestamp 1516325494
transform 1 0 2898 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_171
timestamp 1516325494
transform -1 0 2925 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_171
timestamp 1516325494
transform -1 0 2943 0 1 446
box 0 0 19 49
use OR2X2  OR2X2_1470
timestamp 1516325494
transform -1 0 2962 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_167
timestamp 1516325494
transform -1 0 2970 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_167
timestamp 1516325494
transform -1 0 2989 0 1 446
box 0 0 19 49
use FILL  FILL_BUFX2_183
timestamp 1516325494
transform -1 0 2997 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_183
timestamp 1516325494
transform -1 0 3011 0 1 446
box 0 0 15 49
use FILL  FILL_AND2X2_178
timestamp 1516325494
transform -1 0 3020 0 1 446
box 0 0 8 49
use AND2X2  AND2X2_178
timestamp 1516325494
transform -1 0 3038 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_272
timestamp 1516325494
transform 1 0 3038 0 1 446
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_209
timestamp 1516325494
transform 1 0 3091 0 1 446
box 0 0 53 49
use NAND2X1  NAND2X1_625
timestamp 1516325494
transform 1 0 3145 0 1 446
box 0 0 15 49
use MUX2X1  MUX2X1_625
timestamp 1516325494
transform -1 0 3190 0 1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_762
timestamp 1516325494
transform 1 0 3190 0 1 446
box 0 0 53 49
use INVX8  INVX8_2
timestamp 1516325494
transform -1 0 3270 0 1 446
box 0 0 27 49
use FILL  FILL_OR2X2_100
timestamp 1516325494
transform -1 0 3278 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_100
timestamp 1516325494
transform -1 0 3297 0 1 446
box 0 0 19 49
use FILL  FILL_AND2X2_104
timestamp 1516325494
transform -1 0 3305 0 1 446
box 0 0 8 49
use AND2X2  AND2X2_104
timestamp 1516325494
transform -1 0 3323 0 1 446
box 0 0 19 49
use FILL  FILL_OR2X2_156
timestamp 1516325494
transform -1 0 3331 0 1 446
box 0 0 8 49
use OR2X2  OR2X2_156
timestamp 1516325494
transform -1 0 3350 0 1 446
box 0 0 19 49
use FILL  FILL_AND2X2_164
timestamp 1516325494
transform -1 0 3358 0 1 446
box 0 0 8 49
use AND2X2  AND2X2_164
timestamp 1516325494
transform -1 0 3376 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_713
timestamp 1516325494
transform -1 0 3429 0 1 446
box 0 0 53 49
use FILL  FILL_BUFX2_165
timestamp 1516325494
transform 1 0 3430 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_165
timestamp 1516325494
transform 1 0 3437 0 1 446
box 0 0 15 49
use FILL  FILL_BUFX2_175
timestamp 1516325494
transform -1 0 3460 0 1 446
box 0 0 8 49
use BUFX2  BUFX2_175
timestamp 1516325494
transform -1 0 3475 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_336
timestamp 1516325494
transform 1 0 3475 0 1 446
box 0 0 53 49
use FILL  FILL_AND2X2_181
timestamp 1516325494
transform 1 0 3528 0 1 446
box 0 0 8 49
use AND2X2  AND2X2_181
timestamp 1516325494
transform 1 0 3536 0 1 446
box 0 0 19 49
use INVX1  INVX1_248
timestamp 1516325494
transform 1 0 3555 0 1 446
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_335
timestamp 1516325494
transform -1 0 3619 0 1 446
box 0 0 53 49
use NOR2X1  NOR2X1_113
timestamp 1516325494
transform 1 0 3620 0 1 446
box 0 0 15 49
use AOI22X1  AOI22X1_2
timestamp 1516325494
transform 1 0 3635 0 1 446
box 0 0 23 49
use AOI21X1  AOI21X1_33
timestamp 1516325494
transform 1 0 3658 0 1 446
box 0 0 19 49
use NOR2X1  NOR2X1_118
timestamp 1516325494
transform 1 0 3677 0 1 446
box 0 0 15 49
use NOR2X1  NOR2X1_117
timestamp 1516325494
transform 1 0 3692 0 1 446
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_771
timestamp 1516325494
transform -1 0 3760 0 1 446
box 0 0 53 49
use NAND2X1  NAND2X1_762
timestamp 1516325494
transform -1 0 3775 0 1 446
box 0 0 15 49
use OAI21X1  OAI21X1_93
timestamp 1516325494
transform 1 0 3775 0 1 446
box 0 0 19 49
use AOI21X1  AOI21X1_38
timestamp 1516325494
transform 1 0 3794 0 1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_777
timestamp 1516325494
transform -1 0 3866 0 1 446
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_499
timestamp 1516325494
transform 1 0 2328 0 -1 446
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_107
timestamp 1516325494
transform 1 0 2381 0 -1 446
box 0 0 53 49
use NAND2X1  NAND2X1_75
timestamp 1516325494
transform 1 0 2434 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_75
timestamp 1516325494
transform -1 0 2479 0 -1 446
box 0 0 30 49
use FILL  FILL_BUFX2_227
timestamp 1516325494
transform 1 0 2480 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_227
timestamp 1516325494
transform 1 0 2487 0 -1 446
box 0 0 15 49
use NAND2X1  NAND2X1_143
timestamp 1516325494
transform 1 0 2502 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_143
timestamp 1516325494
transform -1 0 2548 0 -1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_115
timestamp 1516325494
transform -1 0 2601 0 -1 446
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_310
timestamp 1516325494
transform -1 0 2654 0 -1 446
box 0 0 53 49
use FILL  FILL_BUFX2_598
timestamp 1516325494
transform 1 0 2654 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_598
timestamp 1516325494
transform 1 0 2662 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_217
timestamp 1516325494
transform 1 0 2677 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_217
timestamp 1516325494
transform 1 0 2685 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_38
timestamp 1516325494
transform 1 0 2700 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_38
timestamp 1516325494
transform 1 0 2708 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_624
timestamp 1516325494
transform 1 0 2723 0 -1 446
box 0 0 30 49
use NAND2X1  NAND2X1_624
timestamp 1516325494
transform -1 0 2768 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_613
timestamp 1516325494
transform 1 0 2768 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_613
timestamp 1516325494
transform 1 0 2776 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_616
timestamp 1516325494
transform -1 0 2799 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_616
timestamp 1516325494
transform -1 0 2814 0 -1 446
box 0 0 15 49
use FILL  FILL_AND2X2_175
timestamp 1516325494
transform 1 0 2814 0 -1 446
box 0 0 8 49
use AND2X2  AND2X2_175
timestamp 1516325494
transform 1 0 2822 0 -1 446
box 0 0 19 49
use FILL  FILL_AND2X2_176
timestamp 1516325494
transform 1 0 2841 0 -1 446
box 0 0 8 49
use AND2X2  AND2X2_176
timestamp 1516325494
transform 1 0 2848 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1652
timestamp 1516325494
transform 1 0 2867 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1651
timestamp 1516325494
transform 1 0 2886 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1465
timestamp 1516325494
transform 1 0 2905 0 -1 446
box 0 0 19 49
use FILL  FILL_OR2X2_157
timestamp 1516325494
transform -1 0 2932 0 -1 446
box 0 0 8 49
use OR2X2  OR2X2_157
timestamp 1516325494
transform -1 0 2951 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1467
timestamp 1516325494
transform -1 0 2970 0 -1 446
box 0 0 19 49
use FILL  FILL_AND2X2_177
timestamp 1516325494
transform -1 0 2978 0 -1 446
box 0 0 8 49
use AND2X2  AND2X2_177
timestamp 1516325494
transform -1 0 2996 0 -1 446
box 0 0 19 49
use OR2X2  OR2X2_1466
timestamp 1516325494
transform -1 0 3015 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1654
timestamp 1516325494
transform -1 0 3034 0 -1 446
box 0 0 19 49
use AND2X2  AND2X2_1653
timestamp 1516325494
transform -1 0 3053 0 -1 446
box 0 0 19 49
use NAND2X1  NAND2X1_592
timestamp 1516325494
transform 1 0 3053 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_592
timestamp 1516325494
transform -1 0 3099 0 -1 446
box 0 0 30 49
use FILL  FILL_OR2X2_101
timestamp 1516325494
transform -1 0 3107 0 -1 446
box 0 0 8 49
use OR2X2  OR2X2_101
timestamp 1516325494
transform -1 0 3126 0 -1 446
box 0 0 19 49
use NAND2X1  NAND2X1_208
timestamp 1516325494
transform 1 0 3126 0 -1 446
box 0 0 15 49
use MUX2X1  MUX2X1_208
timestamp 1516325494
transform -1 0 3171 0 -1 446
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_240
timestamp 1516325494
transform -1 0 3224 0 -1 446
box 0 0 53 49
use NAND3X1  NAND3X1_75
timestamp 1516325494
transform -1 0 3243 0 -1 446
box 0 0 19 49
use AOI21X1  AOI21X1_41
timestamp 1516325494
transform -1 0 3262 0 -1 446
box 0 0 19 49
use NAND3X1  NAND3X1_79
timestamp 1516325494
transform 1 0 3262 0 -1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_765
timestamp 1516325494
transform 1 0 3281 0 -1 446
box 0 0 53 49
use AOI21X1  AOI21X1_44
timestamp 1516325494
transform -1 0 3354 0 -1 446
box 0 0 19 49
use NAND2X1  NAND2X1_771
timestamp 1516325494
transform -1 0 3369 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_518
timestamp 1516325494
transform 1 0 3369 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_518
timestamp 1516325494
transform 1 0 3376 0 -1 446
box 0 0 15 49
use NAND3X1  NAND3X1_76
timestamp 1516325494
transform 1 0 3392 0 -1 446
box 0 0 19 49
use FILL  FILL_BUFX2_519
timestamp 1516325494
transform -1 0 3419 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_519
timestamp 1516325494
transform -1 0 3433 0 -1 446
box 0 0 15 49
use AOI21X1  AOI21X1_42
timestamp 1516325494
transform -1 0 3452 0 -1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_718
timestamp 1516325494
transform 1 0 3452 0 -1 446
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_752
timestamp 1516325494
transform 1 0 3506 0 -1 446
box 0 0 53 49
use OAI21X1  OAI21X1_89
timestamp 1516325494
transform 1 0 3559 0 -1 446
box 0 0 19 49
use AOI21X1  AOI21X1_48
timestamp 1516325494
transform 1 0 3578 0 -1 446
box 0 0 19 49
use OAI21X1  OAI21X1_96
timestamp 1516325494
transform -1 0 3616 0 -1 446
box 0 0 19 49
use AOI21X1  AOI21X1_30
timestamp 1516325494
transform -1 0 3635 0 -1 446
box 0 0 19 49
use NOR3X1  NOR3X1_12
timestamp 1516325494
transform 1 0 3635 0 -1 446
box 0 0 19 49
use OAI21X1  OAI21X1_90
timestamp 1516325494
transform 1 0 3654 0 -1 446
box 0 0 19 49
use AOI21X1  AOI21X1_32
timestamp 1516325494
transform 1 0 3673 0 -1 446
box 0 0 19 49
use NOR2X1  NOR2X1_115
timestamp 1516325494
transform 1 0 3692 0 -1 446
box 0 0 15 49
use OAI21X1  OAI21X1_88
timestamp 1516325494
transform -1 0 3726 0 -1 446
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_772
timestamp 1516325494
transform -1 0 3779 0 -1 446
box 0 0 53 49
use NOR2X1  NOR2X1_110
timestamp 1516325494
transform -1 0 3794 0 -1 446
box 0 0 15 49
use FILL  FILL_BUFX2_520
timestamp 1516325494
transform -1 0 3802 0 -1 446
box 0 0 8 49
use BUFX2  BUFX2_520
timestamp 1516325494
transform -1 0 3817 0 -1 446
box 0 0 15 49
use NOR2X1  NOR2X1_171
timestamp 1516325494
transform -1 0 3832 0 -1 446
box 0 0 15 49
use NOR2X1  NOR2X1_169
timestamp 1516325494
transform -1 0 3847 0 -1 446
box 0 0 15 49
use NOR2X1  NOR2X1_168
timestamp 1516325494
transform -1 0 3863 0 -1 446
box 0 0 15 49
use FILL  FILL_9_1
timestamp 1516325494
transform -1 0 3871 0 -1 446
box 0 0 8 49
use OR2X2  OR2X2_540
timestamp 1516325494
transform -1 0 21 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_639
timestamp 1516325494
transform -1 0 40 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_539
timestamp 1516325494
transform -1 0 59 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_800
timestamp 1516325494
transform 1 0 59 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_799
timestamp 1516325494
transform -1 0 97 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_606
timestamp 1516325494
transform 1 0 97 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_864
timestamp 1516325494
transform -1 0 135 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_604
timestamp 1516325494
transform 1 0 135 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_701
timestamp 1516325494
transform -1 0 173 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_832
timestamp 1516325494
transform -1 0 192 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_460
timestamp 1516325494
transform -1 0 211 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_520
timestamp 1516325494
transform -1 0 230 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_459
timestamp 1516325494
transform -1 0 249 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_519
timestamp 1516325494
transform -1 0 268 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_458
timestamp 1516325494
transform -1 0 287 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_518
timestamp 1516325494
transform -1 0 306 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_517
timestamp 1516325494
transform -1 0 325 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_677
timestamp 1516325494
transform 1 0 325 0 1 348
box 0 0 19 49
use MUX2X1  MUX2X1_694
timestamp 1516325494
transform 1 0 344 0 1 348
box 0 0 30 49
use MUX2X1  MUX2X1_662
timestamp 1516325494
transform 1 0 374 0 1 348
box 0 0 30 49
use FILL  FILL_BUFX2_687
timestamp 1516325494
transform -1 0 413 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_687
timestamp 1516325494
transform -1 0 427 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_690
timestamp 1516325494
transform -1 0 436 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_690
timestamp 1516325494
transform -1 0 450 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_749
timestamp 1516325494
transform 1 0 450 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_625
timestamp 1516325494
transform 1 0 469 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_626
timestamp 1516325494
transform 1 0 488 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_748
timestamp 1516325494
transform -1 0 526 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_572
timestamp 1516325494
transform -1 0 534 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_572
timestamp 1516325494
transform -1 0 549 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_446
timestamp 1516325494
transform 1 0 549 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_783
timestamp 1516325494
transform 1 0 568 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_657
timestamp 1516325494
transform -1 0 606 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_678
timestamp 1516325494
transform -1 0 614 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_678
timestamp 1516325494
transform -1 0 629 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_441
timestamp 1516325494
transform -1 0 648 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_733
timestamp 1516325494
transform -1 0 656 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_733
timestamp 1516325494
transform -1 0 671 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_581
timestamp 1516325494
transform 1 0 671 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_500
timestamp 1516325494
transform -1 0 709 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_580
timestamp 1516325494
transform -1 0 728 0 1 348
box 0 0 19 49
use FILL  FILL_OR2X2_178
timestamp 1516325494
transform 1 0 728 0 1 348
box 0 0 8 49
use OR2X2  OR2X2_178
timestamp 1516325494
transform 1 0 735 0 1 348
box 0 0 19 49
use FILL  FILL_OR2X2_108
timestamp 1516325494
transform 1 0 754 0 1 348
box 0 0 8 49
use OR2X2  OR2X2_108
timestamp 1516325494
transform 1 0 762 0 1 348
box 0 0 19 49
use FILL  FILL_OR2X2_109
timestamp 1516325494
transform -1 0 789 0 1 348
box 0 0 8 49
use OR2X2  OR2X2_109
timestamp 1516325494
transform -1 0 808 0 1 348
box 0 0 19 49
use FILL  FILL_OR2X2_216
timestamp 1516325494
transform 1 0 808 0 1 348
box 0 0 8 49
use OR2X2  OR2X2_216
timestamp 1516325494
transform 1 0 815 0 1 348
box 0 0 19 49
use OAI21X1  OAI21X1_33
timestamp 1516325494
transform -1 0 853 0 1 348
box 0 0 19 49
use INVX2  INVX2_22
timestamp 1516325494
transform 1 0 853 0 1 348
box 0 0 11 49
use FILL  FILL_BUFX2_58
timestamp 1516325494
transform 1 0 865 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_58
timestamp 1516325494
transform 1 0 872 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_61
timestamp 1516325494
transform -1 0 895 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_61
timestamp 1516325494
transform -1 0 910 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_275
timestamp 1516325494
transform -1 0 929 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1803
timestamp 1516325494
transform 1 0 929 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_137
timestamp 1516325494
transform 1 0 948 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_137
timestamp 1516325494
transform 1 0 956 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_140
timestamp 1516325494
transform -1 0 979 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_140
timestamp 1516325494
transform -1 0 994 0 1 348
box 0 0 15 49
use NAND2X1  NAND2X1_743
timestamp 1516325494
transform 1 0 994 0 1 348
box 0 0 15 49
use OAI21X1  OAI21X1_34
timestamp 1516325494
transform -1 0 1028 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_802
timestamp 1516325494
transform 1 0 1028 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_802
timestamp 1516325494
transform 1 0 1036 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_274
timestamp 1516325494
transform -1 0 1070 0 1 348
box 0 0 19 49
use INVX2  INVX2_23
timestamp 1516325494
transform 1 0 1070 0 1 348
box 0 0 11 49
use FILL  FILL_BUFX2_636
timestamp 1516325494
transform -1 0 1089 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_636
timestamp 1516325494
transform -1 0 1104 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_303
timestamp 1516325494
transform 1 0 1104 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1061
timestamp 1516325494
transform 1 0 1123 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1715
timestamp 1516325494
transform 1 0 1142 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1843
timestamp 1516325494
transform -1 0 1180 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1720
timestamp 1516325494
transform 1 0 1180 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_302
timestamp 1516325494
transform 1 0 1199 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_284
timestamp 1516325494
transform 1 0 1218 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_286
timestamp 1516325494
transform 1 0 1237 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_425
timestamp 1516325494
transform -1 0 1275 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_397
timestamp 1516325494
transform 1 0 1275 0 1 348
box 0 0 19 49
use FILL  FILL_AND2X2_122
timestamp 1516325494
transform -1 0 1302 0 1 348
box 0 0 8 49
use AND2X2  AND2X2_122
timestamp 1516325494
transform -1 0 1321 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_423
timestamp 1516325494
transform -1 0 1340 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_2033
timestamp 1516325494
transform 1 0 1340 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1960
timestamp 1516325494
transform 1 0 1359 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_2029
timestamp 1516325494
transform -1 0 1397 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_420
timestamp 1516325494
transform -1 0 1405 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_420
timestamp 1516325494
transform -1 0 1419 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_1566
timestamp 1516325494
transform -1 0 1438 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1351
timestamp 1516325494
transform -1 0 1457 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1352
timestamp 1516325494
transform -1 0 1476 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_523
timestamp 1516325494
transform 1 0 1476 0 1 348
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_428
timestamp 1516325494
transform 1 0 1530 0 1 348
box 0 0 53 49
use NAND2X1  NAND2X1_396
timestamp 1516325494
transform 1 0 1583 0 1 348
box 0 0 15 49
use MUX2X1  MUX2X1_396
timestamp 1516325494
transform -1 0 1628 0 1 348
box 0 0 30 49
use NAND2X1  NAND2X1_12
timestamp 1516325494
transform 1 0 1628 0 1 348
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_588
timestamp 1516325494
transform 1 0 1644 0 1 348
box 0 0 53 49
use MUX2X1  MUX2X1_12
timestamp 1516325494
transform -1 0 1727 0 1 348
box 0 0 30 49
use NAND2X1  NAND2X1_880
timestamp 1516325494
transform 1 0 1727 0 1 348
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_610
timestamp 1516325494
transform 1 0 1742 0 1 348
box 0 0 53 49
use FILL  FILL_BUFX2_119
timestamp 1516325494
transform -1 0 1804 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_119
timestamp 1516325494
transform -1 0 1818 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_226
timestamp 1516325494
transform -1 0 1826 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_226
timestamp 1516325494
transform -1 0 1841 0 1 348
box 0 0 15 49
use OR2X2  OR2X2_1862
timestamp 1516325494
transform -1 0 1860 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_491
timestamp 1516325494
transform -1 0 1913 0 1 348
box 0 0 53 49
use NAND2X1  NAND2X1_413
timestamp 1516325494
transform 1 0 1913 0 1 348
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_445
timestamp 1516325494
transform 1 0 1929 0 1 348
box 0 0 53 49
use MUX2X1  MUX2X1_413
timestamp 1516325494
transform -1 0 2012 0 1 348
box 0 0 30 49
use OR2X2  OR2X2_1954
timestamp 1516325494
transform -1 0 2031 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_704
timestamp 1516325494
transform 1 0 2031 0 1 348
box 0 0 53 49
use NAND2X1  NAND2X1_320
timestamp 1516325494
transform 1 0 2084 0 1 348
box 0 0 15 49
use MUX2X1  MUX2X1_320
timestamp 1516325494
transform -1 0 2130 0 1 348
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_495
timestamp 1516325494
transform 1 0 2130 0 1 348
box 0 0 53 49
use FILL  FILL_BUFX2_494
timestamp 1516325494
transform -1 0 2191 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_494
timestamp 1516325494
transform -1 0 2206 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_70
timestamp 1516325494
transform 1 0 2206 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_70
timestamp 1516325494
transform 1 0 2214 0 1 348
box 0 0 15 49
use AND2X2  AND2X2_1959
timestamp 1516325494
transform -1 0 2248 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1864
timestamp 1516325494
transform -1 0 2267 0 1 348
box 0 0 19 49
use MUX2X1  MUX2X1_317
timestamp 1516325494
transform 1 0 2267 0 1 348
box 0 0 30 49
use AND2X2  AND2X2_2032
timestamp 1516325494
transform -1 0 2316 0 1 348
box 0 0 19 49
use NAND2X1  NAND2X1_317
timestamp 1516325494
transform 1 0 2316 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_132
timestamp 1516325494
transform 1 0 2331 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_132
timestamp 1516325494
transform 1 0 2339 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_468
timestamp 1516325494
transform 1 0 2354 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_468
timestamp 1516325494
transform 1 0 2362 0 1 348
box 0 0 15 49
use FILL  FILL_BUFX2_308
timestamp 1516325494
transform -1 0 2385 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_308
timestamp 1516325494
transform -1 0 2400 0 1 348
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_79
timestamp 1516325494
transform 1 0 2400 0 1 348
box 0 0 53 49
use AND2X2  AND2X2_1802
timestamp 1516325494
transform -1 0 2472 0 1 348
box 0 0 19 49
use FILL  FILL_BUFX2_653
timestamp 1516325494
transform -1 0 2480 0 1 348
box 0 0 8 49
use BUFX2  BUFX2_653
timestamp 1516325494
transform -1 0 2495 0 1 348
box 0 0 15 49
use OR2X2  OR2X2_1659
timestamp 1516325494
transform -1 0 2514 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1800
timestamp 1516325494
transform -1 0 2533 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1657
timestamp 1516325494
transform -1 0 2552 0 1 348
box 0 0 19 49
use NAND2X1  NAND2X1_502
timestamp 1516325494
transform 1 0 2552 0 1 348
box 0 0 15 49
use MUX2X1  MUX2X1_502
timestamp 1516325494
transform -1 0 2597 0 1 348
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_54
timestamp 1516325494
transform 1 0 2597 0 1 348
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_208
timestamp 1516325494
transform 1 0 2651 0 1 348
box 0 0 53 49
use OR2X2  OR2X2_280
timestamp 1516325494
transform -1 0 2723 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_278
timestamp 1516325494
transform -1 0 2742 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_295
timestamp 1516325494
transform -1 0 2761 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1835
timestamp 1516325494
transform -1 0 2780 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1707
timestamp 1516325494
transform -1 0 2799 0 1 348
box 0 0 19 49
use FILL  FILL_AND2X2_161
timestamp 1516325494
transform 1 0 2799 0 1 348
box 0 0 8 49
use AND2X2  AND2X2_161
timestamp 1516325494
transform 1 0 2806 0 1 348
box 0 0 19 49
use FILL  FILL_OR2X2_154
timestamp 1516325494
transform 1 0 2825 0 1 348
box 0 0 8 49
use OR2X2  OR2X2_154
timestamp 1516325494
transform 1 0 2833 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1629
timestamp 1516325494
transform 1 0 2852 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1437
timestamp 1516325494
transform -1 0 2890 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1435
timestamp 1516325494
transform -1 0 2909 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1628
timestamp 1516325494
transform -1 0 2928 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1536
timestamp 1516325494
transform 1 0 2928 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1315
timestamp 1516325494
transform 1 0 2947 0 1 348
box 0 0 19 49
use OR2X2  OR2X2_1317
timestamp 1516325494
transform 1 0 2966 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1537
timestamp 1516325494
transform -1 0 3004 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_171
timestamp 1516325494
transform 1 0 3004 0 1 348
box 0 0 53 49
use MUX2X1  MUX2X1_235
timestamp 1516325494
transform -1 0 3087 0 1 348
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_759
timestamp 1516325494
transform -1 0 3141 0 1 348
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_706
timestamp 1516325494
transform 1 0 3141 0 1 348
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_764
timestamp 1516325494
transform 1 0 3194 0 1 348
box 0 0 53 49
use NAND3X1  NAND3X1_77
timestamp 1516325494
transform 1 0 3247 0 1 348
box 0 0 19 49
use AOI21X1  AOI21X1_43
timestamp 1516325494
transform -1 0 3285 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_714
timestamp 1516325494
transform 1 0 3285 0 1 348
box 0 0 53 49
use INVX1  INVX1_241
timestamp 1516325494
transform 1 0 3338 0 1 348
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_709
timestamp 1516325494
transform 1 0 3350 0 1 348
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_763
timestamp 1516325494
transform 1 0 3403 0 1 348
box 0 0 53 49
use INVX1  INVX1_262
timestamp 1516325494
transform 1 0 3456 0 1 348
box 0 0 11 49
use NAND3X1  NAND3X1_74
timestamp 1516325494
transform 1 0 3468 0 1 348
box 0 0 19 49
use INVX1  INVX1_242
timestamp 1516325494
transform -1 0 3498 0 1 348
box 0 0 11 49
use NAND3X1  NAND3X1_78
timestamp 1516325494
transform -1 0 3517 0 1 348
box 0 0 19 49
use NAND2X1  NAND2X1_767
timestamp 1516325494
transform -1 0 3532 0 1 348
box 0 0 15 49
use NOR3X1  NOR3X1_25
timestamp 1516325494
transform 1 0 3532 0 1 348
box 0 0 19 49
use NAND2X1  NAND2X1_772
timestamp 1516325494
transform 1 0 3551 0 1 348
box 0 0 15 49
use NOR2X1  NOR2X1_132
timestamp 1516325494
transform 1 0 3566 0 1 348
box 0 0 15 49
use AOI21X1  AOI21X1_31
timestamp 1516325494
transform 1 0 3582 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_770
timestamp 1516325494
transform -1 0 3654 0 1 348
box 0 0 53 49
use NOR2X1  NOR2X1_114
timestamp 1516325494
transform 1 0 3654 0 1 348
box 0 0 15 49
use INVX1  INVX1_245
timestamp 1516325494
transform 1 0 3669 0 1 348
box 0 0 11 49
use NOR3X1  NOR3X1_24
timestamp 1516325494
transform 1 0 3680 0 1 348
box 0 0 19 49
use NOR2X1  NOR2X1_170
timestamp 1516325494
transform -1 0 3714 0 1 348
box 0 0 15 49
use AOI21X1  AOI21X1_37
timestamp 1516325494
transform 1 0 3715 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1129
timestamp 1516325494
transform -1 0 3753 0 1 348
box 0 0 19 49
use AND2X2  AND2X2_1133
timestamp 1516325494
transform -1 0 3772 0 1 348
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_778
timestamp 1516325494
transform -1 0 3825 0 1 348
box 0 0 53 49
use NOR2X1  NOR2X1_158
timestamp 1516325494
transform 1 0 3825 0 1 348
box 0 0 15 49
use INVX1  INVX1_316
timestamp 1516325494
transform -1 0 3851 0 1 348
box 0 0 11 49
use INVX1  INVX1_304
timestamp 1516325494
transform -1 0 3862 0 1 348
box 0 0 11 49
use FILL  FILL_8_1
timestamp 1516325494
transform 1 0 3863 0 1 348
box 0 0 8 49
use MUX2X1  MUX2X1_691
timestamp 1516325494
transform 1 0 2 0 -1 347
box 0 0 30 49
use MUX2X1  MUX2X1_690
timestamp 1516325494
transform -1 0 62 0 -1 347
box 0 0 30 49
use MUX2X1  MUX2X1_692
timestamp 1516325494
transform 1 0 2 0 1 249
box 0 0 30 49
use MUX2X1  MUX2X1_707
timestamp 1516325494
transform 1 0 32 0 1 249
box 0 0 30 49
use MUX2X1  MUX2X1_688
timestamp 1516325494
transform 1 0 63 0 -1 347
box 0 0 30 49
use AND2X2  AND2X2_865
timestamp 1516325494
transform 1 0 93 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_728
timestamp 1516325494
transform 1 0 112 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_729
timestamp 1516325494
transform 1 0 131 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_720
timestamp 1516325494
transform -1 0 169 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_700
timestamp 1516325494
transform -1 0 188 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_525
timestamp 1516325494
transform -1 0 207 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_524
timestamp 1516325494
transform -1 0 226 0 -1 347
box 0 0 19 49
use FILL  FILL_BUFX2_688
timestamp 1516325494
transform 1 0 226 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_688
timestamp 1516325494
transform 1 0 234 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_641
timestamp 1516325494
transform 1 0 249 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_640
timestamp 1516325494
transform -1 0 287 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_522
timestamp 1516325494
transform -1 0 306 0 -1 347
box 0 0 19 49
use MUX2X1  MUX2X1_697
timestamp 1516325494
transform -1 0 336 0 -1 347
box 0 0 30 49
use FILL  FILL_BUFX2_689
timestamp 1516325494
transform 1 0 336 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_689
timestamp 1516325494
transform 1 0 344 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_734
timestamp 1516325494
transform 1 0 359 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_734
timestamp 1516325494
transform 1 0 367 0 -1 347
box 0 0 15 49
use AND2X2  AND2X2_583
timestamp 1516325494
transform -1 0 401 0 -1 347
box 0 0 19 49
use MUX2X1  MUX2X1_661
timestamp 1516325494
transform 1 0 401 0 -1 347
box 0 0 30 49
use AND2X2  AND2X2_590
timestamp 1516325494
transform 1 0 431 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_585
timestamp 1516325494
transform 1 0 450 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_505
timestamp 1516325494
transform 1 0 469 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_507
timestamp 1516325494
transform 1 0 488 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_593
timestamp 1516325494
transform 1 0 507 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_511
timestamp 1516325494
transform -1 0 545 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_656
timestamp 1516325494
transform 1 0 545 0 -1 347
box 0 0 19 49
use MUX2X1  MUX2X1_704
timestamp 1516325494
transform 1 0 564 0 -1 347
box 0 0 30 49
use MUX2X1  MUX2X1_705
timestamp 1516325494
transform 1 0 595 0 -1 347
box 0 0 30 49
use MUX2X1  MUX2X1_703
timestamp 1516325494
transform 1 0 625 0 -1 347
box 0 0 30 49
use AND2X2  AND2X2_440
timestamp 1516325494
transform -1 0 675 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_578
timestamp 1516325494
transform 1 0 675 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_579
timestamp 1516325494
transform 1 0 694 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_499
timestamp 1516325494
transform 1 0 713 0 -1 347
box 0 0 19 49
use INVX1  INVX1_181
timestamp 1516325494
transform -1 0 743 0 -1 347
box 0 0 11 49
use OR2X2  OR2X2_1481
timestamp 1516325494
transform -1 0 762 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1475
timestamp 1516325494
transform -1 0 781 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1659
timestamp 1516325494
transform -1 0 800 0 -1 347
box 0 0 19 49
use FILL  FILL_OR2X2_214
timestamp 1516325494
transform -1 0 808 0 -1 347
box 0 0 8 49
use OR2X2  OR2X2_214
timestamp 1516325494
transform -1 0 827 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_730
timestamp 1516325494
transform -1 0 842 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_637
timestamp 1516325494
transform 1 0 842 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_637
timestamp 1516325494
transform 1 0 849 0 -1 347
box 0 0 15 49
use NAND2X1  NAND2X1_729
timestamp 1516325494
transform 1 0 865 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_803
timestamp 1516325494
transform 1 0 880 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_803
timestamp 1516325494
transform 1 0 887 0 -1 347
box 0 0 15 49
use FILL  FILL_AND2X2_228
timestamp 1516325494
transform -1 0 911 0 -1 347
box 0 0 8 49
use AND2X2  AND2X2_228
timestamp 1516325494
transform -1 0 929 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_731
timestamp 1516325494
transform 1 0 929 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1571
timestamp 1516325494
transform -1 0 963 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1565
timestamp 1516325494
transform -1 0 982 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1730
timestamp 1516325494
transform -1 0 1001 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1728
timestamp 1516325494
transform -1 0 1020 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_2087
timestamp 1516325494
transform 1 0 1020 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1996
timestamp 1516325494
transform 1 0 1039 0 -1 347
box 0 0 19 49
use FILL  FILL_BUFX2_126
timestamp 1516325494
transform 1 0 1058 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_126
timestamp 1516325494
transform 1 0 1066 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1060
timestamp 1516325494
transform 1 0 1081 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1341
timestamp 1516325494
transform -1 0 1119 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1845
timestamp 1516325494
transform 1 0 1119 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1870
timestamp 1516325494
transform 1 0 1138 0 -1 347
box 0 0 19 49
use FILL  FILL_BUFX2_654
timestamp 1516325494
transform 1 0 1157 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_654
timestamp 1516325494
transform 1 0 1165 0 -1 347
box 0 0 15 49
use AND2X2  AND2X2_1847
timestamp 1516325494
transform -1 0 1199 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_285
timestamp 1516325494
transform 1 0 1199 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_304
timestamp 1516325494
transform -1 0 1237 0 -1 347
box 0 0 19 49
use FILL  FILL_OR2X2_118
timestamp 1516325494
transform -1 0 1245 0 -1 347
box 0 0 8 49
use OR2X2  OR2X2_118
timestamp 1516325494
transform -1 0 1264 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_424
timestamp 1516325494
transform -1 0 1283 0 -1 347
box 0 0 19 49
use FILL  FILL_OR2X2_116
timestamp 1516325494
transform -1 0 1291 0 -1 347
box 0 0 8 49
use OR2X2  OR2X2_116
timestamp 1516325494
transform -1 0 1309 0 -1 347
box 0 0 19 49
use FILL  FILL_AND2X2_123
timestamp 1516325494
transform -1 0 1317 0 -1 347
box 0 0 8 49
use AND2X2  AND2X2_123
timestamp 1516325494
transform -1 0 1336 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_2031
timestamp 1516325494
transform 1 0 1336 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1338
timestamp 1516325494
transform -1 0 1374 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_725
timestamp 1516325494
transform -1 0 1389 0 -1 347
box 0 0 15 49
use AND2X2  AND2X2_1567
timestamp 1516325494
transform 1 0 1389 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1569
timestamp 1516325494
transform 1 0 1408 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1355
timestamp 1516325494
transform 1 0 1427 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1361
timestamp 1516325494
transform 1 0 1446 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1054
timestamp 1516325494
transform -1 0 1484 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_724
timestamp 1516325494
transform -1 0 1499 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_309
timestamp 1516325494
transform 1 0 1499 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_309
timestamp 1516325494
transform 1 0 1507 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_825
timestamp 1516325494
transform 1 0 1522 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_825
timestamp 1516325494
transform 1 0 1530 0 -1 347
box 0 0 15 49
use AND2X2  AND2X2_1340
timestamp 1516325494
transform -1 0 1564 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1057
timestamp 1516325494
transform -1 0 1583 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_739
timestamp 1516325494
transform 1 0 1583 0 -1 347
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_34
timestamp 1516325494
transform 1 0 1598 0 -1 347
box 0 0 53 49
use NAND2X1  NAND2X1_418
timestamp 1516325494
transform 1 0 1651 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_418
timestamp 1516325494
transform -1 0 1696 0 -1 347
box 0 0 30 49
use FILL  FILL_BUFX2_345
timestamp 1516325494
transform 1 0 1697 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_345
timestamp 1516325494
transform 1 0 1704 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1056
timestamp 1516325494
transform -1 0 1739 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_290
timestamp 1516325494
transform 1 0 1739 0 -1 347
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_674
timestamp 1516325494
transform 1 0 1754 0 -1 347
box 0 0 53 49
use MUX2X1  MUX2X1_290
timestamp 1516325494
transform -1 0 1837 0 -1 347
box 0 0 30 49
use FILL  FILL_BUFX2_350
timestamp 1516325494
transform 1 0 1837 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_350
timestamp 1516325494
transform 1 0 1845 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_435
timestamp 1516325494
transform -1 0 1868 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_435
timestamp 1516325494
transform -1 0 1883 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_701
timestamp 1516325494
transform 1 0 1883 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_701
timestamp 1516325494
transform 1 0 1891 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1353
timestamp 1516325494
transform -1 0 1925 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1568
timestamp 1516325494
transform -1 0 1944 0 -1 347
box 0 0 19 49
use FILL  FILL_BUFX2_220
timestamp 1516325494
transform -1 0 1952 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_220
timestamp 1516325494
transform -1 0 1966 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1354
timestamp 1516325494
transform -1 0 1986 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_2028
timestamp 1516325494
transform -1 0 2005 0 -1 347
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_684
timestamp 1516325494
transform 1 0 2005 0 -1 347
box 0 0 53 49
use NAND2X1  NAND2X1_300
timestamp 1516325494
transform 1 0 2058 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_300
timestamp 1516325494
transform -1 0 2103 0 -1 347
box 0 0 30 49
use FILL  FILL_BUFX2_288
timestamp 1516325494
transform -1 0 2111 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_288
timestamp 1516325494
transform -1 0 2126 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_821
timestamp 1516325494
transform 1 0 2126 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_821
timestamp 1516325494
transform 1 0 2134 0 -1 347
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_51
timestamp 1516325494
transform 1 0 2149 0 -1 347
box 0 0 53 49
use AND2X2  AND2X2_2030
timestamp 1516325494
transform -1 0 2221 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1956
timestamp 1516325494
transform -1 0 2240 0 -1 347
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_640
timestamp 1516325494
transform 1 0 2240 0 -1 347
box 0 0 53 49
use FILL  FILL_BUFX2_123
timestamp 1516325494
transform -1 0 2301 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_123
timestamp 1516325494
transform -1 0 2316 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1958
timestamp 1516325494
transform -1 0 2335 0 -1 347
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_672
timestamp 1516325494
transform 1 0 2335 0 -1 347
box 0 0 53 49
use NAND2X1  NAND2X1_64
timestamp 1516325494
transform 1 0 2388 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_64
timestamp 1516325494
transform -1 0 2434 0 -1 347
box 0 0 30 49
use FILL  FILL_BUFX2_496
timestamp 1516325494
transform -1 0 2442 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_496
timestamp 1516325494
transform -1 0 2457 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1658
timestamp 1516325494
transform 1 0 2457 0 -1 347
box 0 0 19 49
use FILL  FILL_BUFX2_135
timestamp 1516325494
transform -1 0 2484 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_135
timestamp 1516325494
transform -1 0 2498 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_349
timestamp 1516325494
transform -1 0 2507 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_349
timestamp 1516325494
transform -1 0 2521 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_1656
timestamp 1516325494
transform -1 0 2540 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1716
timestamp 1516325494
transform 1 0 2540 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1846
timestamp 1516325494
transform -1 0 2578 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1717
timestamp 1516325494
transform -1 0 2597 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_438
timestamp 1516325494
transform 1 0 2597 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_438
timestamp 1516325494
transform -1 0 2643 0 -1 347
box 0 0 30 49
use FILL  FILL_BUFX2_751
timestamp 1516325494
transform -1 0 2651 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_751
timestamp 1516325494
transform -1 0 2666 0 -1 347
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_56
timestamp 1516325494
transform 1 0 2666 0 -1 347
box 0 0 53 49
use NAND2X1  NAND2X1_440
timestamp 1516325494
transform 1 0 2719 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_440
timestamp 1516325494
transform -1 0 2764 0 -1 347
box 0 0 30 49
use AND2X2  AND2X2_296
timestamp 1516325494
transform -1 0 2784 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1705
timestamp 1516325494
transform 1 0 2784 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1836
timestamp 1516325494
transform -1 0 2822 0 -1 347
box 0 0 19 49
use FILL  FILL_OR2X2_152
timestamp 1516325494
transform -1 0 2830 0 -1 347
box 0 0 8 49
use OR2X2  OR2X2_152
timestamp 1516325494
transform -1 0 2848 0 -1 347
box 0 0 19 49
use FILL  FILL_AND2X2_160
timestamp 1516325494
transform -1 0 2856 0 -1 347
box 0 0 8 49
use AND2X2  AND2X2_160
timestamp 1516325494
transform -1 0 2875 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_1436
timestamp 1516325494
transform -1 0 2894 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1631
timestamp 1516325494
transform -1 0 2913 0 -1 347
box 0 0 19 49
use FILL  FILL_OR2X2_153
timestamp 1516325494
transform -1 0 2921 0 -1 347
box 0 0 8 49
use OR2X2  OR2X2_153
timestamp 1516325494
transform -1 0 2939 0 -1 347
box 0 0 19 49
use FILL  FILL_AND2X2_163
timestamp 1516325494
transform -1 0 2947 0 -1 347
box 0 0 8 49
use AND2X2  AND2X2_163
timestamp 1516325494
transform -1 0 2966 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_591
timestamp 1516325494
transform 1 0 2966 0 -1 347
box 0 0 15 49
use FILL  FILL_AND2X2_100
timestamp 1516325494
transform 1 0 2981 0 -1 347
box 0 0 8 49
use AND2X2  AND2X2_100
timestamp 1516325494
transform 1 0 2989 0 -1 347
box 0 0 19 49
use FILL  FILL_OR2X2_96
timestamp 1516325494
transform -1 0 3016 0 -1 347
box 0 0 8 49
use OR2X2  OR2X2_96
timestamp 1516325494
transform -1 0 3034 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_235
timestamp 1516325494
transform 1 0 3034 0 -1 347
box 0 0 15 49
use FILL  FILL_AND2X2_101
timestamp 1516325494
transform -1 0 3058 0 -1 347
box 0 0 8 49
use AND2X2  AND2X2_101
timestamp 1516325494
transform -1 0 3076 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_619
timestamp 1516325494
transform 1 0 3076 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_619
timestamp 1516325494
transform -1 0 3121 0 -1 347
box 0 0 30 49
use AND2X2  AND2X2_1137
timestamp 1516325494
transform -1 0 3141 0 -1 347
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_235
timestamp 1516325494
transform 1 0 3141 0 -1 347
box 0 0 53 49
use NAND2X1  NAND2X1_203
timestamp 1516325494
transform 1 0 3194 0 -1 347
box 0 0 15 49
use MUX2X1  MUX2X1_203
timestamp 1516325494
transform -1 0 3239 0 -1 347
box 0 0 30 49
use AND2X2  AND2X2_1140
timestamp 1516325494
transform 1 0 3240 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1165
timestamp 1516325494
transform 1 0 3259 0 -1 347
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_760
timestamp 1516325494
transform 1 0 3278 0 -1 347
box 0 0 53 49
use AND2X2  AND2X2_1161
timestamp 1516325494
transform 1 0 3331 0 -1 347
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_756
timestamp 1516325494
transform 1 0 3350 0 -1 347
box 0 0 53 49
use OAI21X1  OAI21X1_95
timestamp 1516325494
transform -1 0 3422 0 -1 347
box 0 0 19 49
use NOR2X1  NOR2X1_130
timestamp 1516325494
transform -1 0 3437 0 -1 347
box 0 0 15 49
use FILL  FILL_BUFX2_233
timestamp 1516325494
transform 1 0 3437 0 -1 347
box 0 0 8 49
use BUFX2  BUFX2_233
timestamp 1516325494
transform 1 0 3445 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_935
timestamp 1516325494
transform -1 0 3479 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_769
timestamp 1516325494
transform -1 0 3494 0 -1 347
box 0 0 15 49
use AND2X2  AND2X2_1122
timestamp 1516325494
transform 1 0 3494 0 -1 347
box 0 0 19 49
use NAND3X1  NAND3X1_65
timestamp 1516325494
transform 1 0 3513 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_755
timestamp 1516325494
transform 1 0 3532 0 -1 347
box 0 0 15 49
use NAND3X1  NAND3X1_66
timestamp 1516325494
transform -1 0 3566 0 -1 347
box 0 0 19 49
use NAND3X1  NAND3X1_67
timestamp 1516325494
transform 1 0 3566 0 -1 347
box 0 0 19 49
use OAI21X1  OAI21X1_87
timestamp 1516325494
transform -1 0 3604 0 -1 347
box 0 0 19 49
use NOR2X1  NOR2X1_116
timestamp 1516325494
transform -1 0 3619 0 -1 347
box 0 0 15 49
use OR2X2  OR2X2_915
timestamp 1516325494
transform -1 0 3639 0 -1 347
box 0 0 19 49
use NAND2X1  NAND2X1_770
timestamp 1516325494
transform -1 0 3654 0 -1 347
box 0 0 15 49
use INVX1  INVX1_244
timestamp 1516325494
transform -1 0 3665 0 -1 347
box 0 0 11 49
use NAND3X1  NAND3X1_64
timestamp 1516325494
transform -1 0 3684 0 -1 347
box 0 0 19 49
use NOR2X1  NOR2X1_122
timestamp 1516325494
transform 1 0 3684 0 -1 347
box 0 0 15 49
use INVX1  INVX1_243
timestamp 1516325494
transform -1 0 3710 0 -1 347
box 0 0 11 49
use AND2X2  AND2X2_1123
timestamp 1516325494
transform 1 0 3711 0 -1 347
box 0 0 19 49
use OAI21X1  OAI21X1_91
timestamp 1516325494
transform 1 0 3730 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_917
timestamp 1516325494
transform -1 0 3768 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1127
timestamp 1516325494
transform -1 0 3787 0 -1 347
box 0 0 19 49
use OR2X2  OR2X2_924
timestamp 1516325494
transform -1 0 3806 0 -1 347
box 0 0 19 49
use AND2X2  AND2X2_1132
timestamp 1516325494
transform 1 0 3806 0 -1 347
box 0 0 19 49
use NOR3X1  NOR3X1_20
timestamp 1516325494
transform -1 0 3844 0 -1 347
box 0 0 19 49
use NOR2X1  NOR2X1_166
timestamp 1516325494
transform -1 0 3859 0 -1 347
box 0 0 15 49
use FILL  FILL_7_1
timestamp 1516325494
transform -1 0 3867 0 -1 347
box 0 0 8 49
use MUX2X1  MUX2X1_689
timestamp 1516325494
transform 1 0 63 0 1 249
box 0 0 30 49
use AND2X2  AND2X2_528
timestamp 1516325494
transform -1 0 112 0 1 249
box 0 0 19 49
use MUX2X1  MUX2X1_687
timestamp 1516325494
transform -1 0 142 0 1 249
box 0 0 30 49
use OR2X2  OR2X2_603
timestamp 1516325494
transform -1 0 162 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_833
timestamp 1516325494
transform 1 0 162 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_464
timestamp 1516325494
transform 1 0 181 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_465
timestamp 1516325494
transform 1 0 200 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_521
timestamp 1516325494
transform -1 0 238 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_765
timestamp 1516325494
transform 1 0 238 0 1 249
box 0 0 19 49
use MUX2X1  MUX2X1_696
timestamp 1516325494
transform 1 0 257 0 1 249
box 0 0 30 49
use FILL  FILL_BUFX2_399
timestamp 1516325494
transform 1 0 287 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_399
timestamp 1516325494
transform 1 0 295 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_698
timestamp 1516325494
transform -1 0 340 0 1 249
box 0 0 30 49
use AND2X2  AND2X2_582
timestamp 1516325494
transform 1 0 340 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_504
timestamp 1516325494
transform 1 0 359 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_503
timestamp 1516325494
transform -1 0 397 0 1 249
box 0 0 19 49
use MUX2X1  MUX2X1_660
timestamp 1516325494
transform 1 0 397 0 1 249
box 0 0 30 49
use AND2X2  AND2X2_591
timestamp 1516325494
transform 1 0 428 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_509
timestamp 1516325494
transform 1 0 447 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_586
timestamp 1516325494
transform -1 0 485 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_506
timestamp 1516325494
transform -1 0 504 0 1 249
box 0 0 19 49
use MUX2X1  MUX2X1_701
timestamp 1516325494
transform -1 0 534 0 1 249
box 0 0 30 49
use OR2X2  OR2X2_414
timestamp 1516325494
transform -1 0 553 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_442
timestamp 1516325494
transform -1 0 572 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_444
timestamp 1516325494
transform -1 0 591 0 1 249
box 0 0 19 49
use INVX1  INVX1_182
timestamp 1516325494
transform -1 0 602 0 1 249
box 0 0 11 49
use AND2X2  AND2X2_644
timestamp 1516325494
transform 1 0 602 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_412
timestamp 1516325494
transform -1 0 640 0 1 249
box 0 0 19 49
use FILL  FILL_OR2X2_174
timestamp 1516325494
transform 1 0 640 0 1 249
box 0 0 8 49
use OR2X2  OR2X2_174
timestamp 1516325494
transform 1 0 648 0 1 249
box 0 0 19 49
use FILL  FILL_OR2X2_172
timestamp 1516325494
transform -1 0 675 0 1 249
box 0 0 8 49
use OR2X2  OR2X2_172
timestamp 1516325494
transform -1 0 694 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_183
timestamp 1516325494
transform -1 0 702 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_183
timestamp 1516325494
transform -1 0 720 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_182
timestamp 1516325494
transform -1 0 728 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_182
timestamp 1516325494
transform -1 0 747 0 1 249
box 0 0 19 49
use FILL  FILL_OR2X2_188
timestamp 1516325494
transform 1 0 747 0 1 249
box 0 0 8 49
use OR2X2  OR2X2_188
timestamp 1516325494
transform 1 0 754 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1661
timestamp 1516325494
transform -1 0 792 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_227
timestamp 1516325494
transform -1 0 800 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_227
timestamp 1516325494
transform -1 0 819 0 1 249
box 0 0 19 49
use FILL  FILL_OR2X2_215
timestamp 1516325494
transform -1 0 827 0 1 249
box 0 0 8 49
use OR2X2  OR2X2_215
timestamp 1516325494
transform -1 0 846 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_229
timestamp 1516325494
transform -1 0 854 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_229
timestamp 1516325494
transform -1 0 872 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1511
timestamp 1516325494
transform 1 0 872 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_230
timestamp 1516325494
transform -1 0 899 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_230
timestamp 1516325494
transform -1 0 918 0 1 249
box 0 0 19 49
use FILL  FILL_BUFX2_682
timestamp 1516325494
transform -1 0 926 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_682
timestamp 1516325494
transform -1 0 940 0 1 249
box 0 0 15 49
use AND2X2  AND2X2_1732
timestamp 1516325494
transform 1 0 941 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1570
timestamp 1516325494
transform -1 0 979 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1734
timestamp 1516325494
transform 1 0 979 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1729
timestamp 1516325494
transform -1 0 1017 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1563
timestamp 1516325494
transform -1 0 1036 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_2088
timestamp 1516325494
transform -1 0 1055 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1343
timestamp 1516325494
transform 1 0 1055 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1964
timestamp 1516325494
transform -1 0 1093 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_380
timestamp 1516325494
transform 1 0 1093 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_355
timestamp 1516325494
transform 1 0 1112 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_379
timestamp 1516325494
transform -1 0 1150 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1962
timestamp 1516325494
transform -1 0 1169 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1849
timestamp 1516325494
transform -1 0 1188 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_305
timestamp 1516325494
transform 1 0 1188 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_125
timestamp 1516325494
transform -1 0 1215 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_125
timestamp 1516325494
transform -1 0 1233 0 1 249
box 0 0 19 49
use FILL  FILL_OR2X2_117
timestamp 1516325494
transform 1 0 1233 0 1 249
box 0 0 8 49
use OR2X2  OR2X2_117
timestamp 1516325494
transform 1 0 1241 0 1 249
box 0 0 19 49
use FILL  FILL_AND2X2_124
timestamp 1516325494
transform -1 0 1268 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_124
timestamp 1516325494
transform -1 0 1286 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1573
timestamp 1516325494
transform 1 0 1286 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1571
timestamp 1516325494
transform 1 0 1305 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1360
timestamp 1516325494
transform 1 0 1324 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1336
timestamp 1516325494
transform -1 0 1362 0 1 249
box 0 0 19 49
use FILL  FILL_BUFX2_29
timestamp 1516325494
transform -1 0 1370 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_29
timestamp 1516325494
transform -1 0 1385 0 1 249
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_595
timestamp 1516325494
transform 1 0 1385 0 1 249
box 0 0 53 49
use NAND2X1  NAND2X1_19
timestamp 1516325494
transform 1 0 1438 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_19
timestamp 1516325494
transform -1 0 1484 0 1 249
box 0 0 30 49
use FILL  FILL_BUFX2_205
timestamp 1516325494
transform -1 0 1492 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_205
timestamp 1516325494
transform -1 0 1507 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_2
timestamp 1516325494
transform 1 0 1507 0 1 249
box 0 0 30 49
use NAND2X1  NAND2X1_2
timestamp 1516325494
transform -1 0 1552 0 1 249
box 0 0 15 49
use OR2X2  OR2X2_1051
timestamp 1516325494
transform -1 0 1571 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_578
timestamp 1516325494
transform -1 0 1624 0 1 249
box 0 0 53 49
use AND2X2  AND2X2_1658
timestamp 1516325494
transform -1 0 1644 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1471
timestamp 1516325494
transform -1 0 1663 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1472
timestamp 1516325494
transform -1 0 1682 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_432
timestamp 1516325494
transform 1 0 1682 0 1 249
box 0 0 53 49
use NAND2X1  NAND2X1_400
timestamp 1516325494
transform 1 0 1735 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_400
timestamp 1516325494
transform -1 0 1780 0 1 249
box 0 0 30 49
use AND2X2  AND2X2_1660
timestamp 1516325494
transform -1 0 1799 0 1 249
box 0 0 19 49
use MUX2X1  MUX2X1_460
timestamp 1516325494
transform 1 0 1799 0 1 249
box 0 0 30 49
use NAND2X1  NAND2X1_460
timestamp 1516325494
transform -1 0 1845 0 1 249
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_556
timestamp 1516325494
transform -1 0 1898 0 1 249
box 0 0 53 49
use NAND2X1  NAND2X1_464
timestamp 1516325494
transform -1 0 1913 0 1 249
box 0 0 15 49
use OR2X2  OR2X2_1473
timestamp 1516325494
transform -1 0 1932 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_560
timestamp 1516325494
transform -1 0 1985 0 1 249
box 0 0 53 49
use FILL  FILL_BUFX2_425
timestamp 1516325494
transform -1 0 1994 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_425
timestamp 1516325494
transform -1 0 2008 0 1 249
box 0 0 15 49
use FILL  FILL_BUFX2_652
timestamp 1516325494
transform -1 0 2016 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_652
timestamp 1516325494
transform -1 0 2031 0 1 249
box 0 0 15 49
use OR2X2  OR2X2_1953
timestamp 1516325494
transform -1 0 2050 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_576
timestamp 1516325494
transform 1 0 2050 0 1 249
box 0 0 53 49
use NAND2X1  NAND2X1_480
timestamp 1516325494
transform 1 0 2103 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_480
timestamp 1516325494
transform -1 0 2149 0 1 249
box 0 0 30 49
use AND2X2  AND2X2_1731
timestamp 1516325494
transform -1 0 2168 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1567
timestamp 1516325494
transform -1 0 2187 0 1 249
box 0 0 19 49
use NAND2X1  NAND2X1_435
timestamp 1516325494
transform 1 0 2187 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_435
timestamp 1516325494
transform -1 0 2232 0 1 249
box 0 0 30 49
use NAND2X1  NAND2X1_477
timestamp 1516325494
transform 1 0 2233 0 1 249
box 0 0 15 49
use OR2X2  OR2X2_1863
timestamp 1516325494
transform -1 0 2267 0 1 249
box 0 0 19 49
use NAND2X1  NAND2X1_910
timestamp 1516325494
transform 1 0 2267 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_855
timestamp 1516325494
transform -1 0 2312 0 1 249
box 0 0 30 49
use FILL  FILL_BUFX2_655
timestamp 1516325494
transform -1 0 2320 0 1 249
box 0 0 8 49
use BUFX2  BUFX2_655
timestamp 1516325494
transform -1 0 2335 0 1 249
box 0 0 15 49
use OR2X2  OR2X2_1508
timestamp 1516325494
transform -1 0 2354 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_657
timestamp 1516325494
transform 1 0 2354 0 1 249
box 0 0 53 49
use NAND2X1  NAND2X1_49
timestamp 1516325494
transform 1 0 2407 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_49
timestamp 1516325494
transform -1 0 2453 0 1 249
box 0 0 30 49
use NAND2X1  NAND2X1_54
timestamp 1516325494
transform -1 0 2468 0 1 249
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_662
timestamp 1516325494
transform 1 0 2468 0 1 249
box 0 0 53 49
use MUX2X1  MUX2X1_54
timestamp 1516325494
transform -1 0 2551 0 1 249
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_630
timestamp 1516325494
transform 1 0 2552 0 1 249
box 0 0 53 49
use NAND2X1  NAND2X1_900
timestamp 1516325494
transform 1 0 2605 0 1 249
box 0 0 15 49
use MUX2X1  MUX2X1_845
timestamp 1516325494
transform -1 0 2650 0 1 249
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_216
timestamp 1516325494
transform 1 0 2651 0 1 249
box 0 0 53 49
use MUX2X1  MUX2X1_632
timestamp 1516325494
transform 1 0 2704 0 1 249
box 0 0 30 49
use NAND2X1  NAND2X1_632
timestamp 1516325494
transform -1 0 2749 0 1 249
box 0 0 15 49
use OR2X2  OR2X2_279
timestamp 1516325494
transform -1 0 2768 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_297
timestamp 1516325494
transform -1 0 2787 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1706
timestamp 1516325494
transform -1 0 2806 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1838
timestamp 1516325494
transform -1 0 2825 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1837
timestamp 1516325494
transform -1 0 2844 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1630
timestamp 1516325494
transform 1 0 2844 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_271
timestamp 1516325494
transform -1 0 2916 0 1 249
box 0 0 53 49
use AND2X2  AND2X2_1539
timestamp 1516325494
transform 1 0 2917 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_1316
timestamp 1516325494
transform 1 0 2936 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1538
timestamp 1516325494
transform -1 0 2974 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_203
timestamp 1516325494
transform 1 0 2974 0 1 249
box 0 0 53 49
use OR2X2  OR2X2_929
timestamp 1516325494
transform -1 0 3046 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_758
timestamp 1516325494
transform 1 0 3046 0 1 249
box 0 0 53 49
use AND2X2  AND2X2_1138
timestamp 1516325494
transform -1 0 3118 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1135
timestamp 1516325494
transform 1 0 3118 0 1 249
box 0 0 19 49
use AOI22X1  AOI22X1_3
timestamp 1516325494
transform -1 0 3160 0 1 249
box 0 0 23 49
use AND2X2  AND2X2_1136
timestamp 1516325494
transform -1 0 3179 0 1 249
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_757
timestamp 1516325494
transform 1 0 3179 0 1 249
box 0 0 53 49
use NOR2X1  NOR2X1_124
timestamp 1516325494
transform 1 0 3232 0 1 249
box 0 0 15 49
use AOI22X1  AOI22X1_4
timestamp 1516325494
transform -1 0 3270 0 1 249
box 0 0 23 49
use AND2X2  AND2X2_1166
timestamp 1516325494
transform -1 0 3289 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_928
timestamp 1516325494
transform -1 0 3308 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1175
timestamp 1516325494
transform -1 0 3327 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_944
timestamp 1516325494
transform -1 0 3346 0 1 249
box 0 0 19 49
use OAI21X1  OAI21X1_94
timestamp 1516325494
transform -1 0 3365 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1160
timestamp 1516325494
transform -1 0 3384 0 1 249
box 0 0 19 49
use NOR2X1  NOR2X1_125
timestamp 1516325494
transform 1 0 3384 0 1 249
box 0 0 15 49
use OAI21X1  OAI21X1_86
timestamp 1516325494
transform -1 0 3418 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1134
timestamp 1516325494
transform -1 0 3437 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_927
timestamp 1516325494
transform -1 0 3456 0 1 249
box 0 0 19 49
use OR2X2  OR2X2_916
timestamp 1516325494
transform -1 0 3475 0 1 249
box 0 0 19 49
use INVX1  INVX1_239
timestamp 1516325494
transform 1 0 3475 0 1 249
box 0 0 11 49
use NAND3X1  NAND3X1_73
timestamp 1516325494
transform -1 0 3506 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1155
timestamp 1516325494
transform -1 0 3525 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1154
timestamp 1516325494
transform -1 0 3544 0 1 249
box 0 0 19 49
use NOR3X1  NOR3X1_11
timestamp 1516325494
transform -1 0 3563 0 1 249
box 0 0 19 49
use AOI21X1  AOI21X1_28
timestamp 1516325494
transform 1 0 3563 0 1 249
box 0 0 19 49
use NAND2X1  NAND2X1_752
timestamp 1516325494
transform 1 0 3582 0 1 249
box 0 0 15 49
use NAND2X1  NAND2X1_757
timestamp 1516325494
transform 1 0 3597 0 1 249
box 0 0 15 49
use INVX1  INVX1_247
timestamp 1516325494
transform -1 0 3623 0 1 249
box 0 0 11 49
use OR2X2  OR2X2_914
timestamp 1516325494
transform 1 0 3623 0 1 249
box 0 0 19 49
use OAI21X1  OAI21X1_85
timestamp 1516325494
transform -1 0 3661 0 1 249
box 0 0 19 49
use NAND2X1  NAND2X1_751
timestamp 1516325494
transform -1 0 3676 0 1 249
box 0 0 15 49
use NOR2X1  NOR2X1_106
timestamp 1516325494
transform 1 0 3677 0 1 249
box 0 0 15 49
use NAND3X1  NAND3X1_63
timestamp 1516325494
transform -1 0 3711 0 1 249
box 0 0 19 49
use NAND3X1  NAND3X1_62
timestamp 1516325494
transform -1 0 3730 0 1 249
box 0 0 19 49
use INVX1  INVX1_237
timestamp 1516325494
transform 1 0 3730 0 1 249
box 0 0 11 49
use AOI21X1  AOI21X1_34
timestamp 1516325494
transform 1 0 3741 0 1 249
box 0 0 19 49
use AND2X2  AND2X2_1128
timestamp 1516325494
transform -1 0 3779 0 1 249
box 0 0 19 49
use NAND2X1  NAND2X1_758
timestamp 1516325494
transform -1 0 3794 0 1 249
box 0 0 15 49
use NAND3X1  NAND3X1_68
timestamp 1516325494
transform -1 0 3813 0 1 249
box 0 0 19 49
use INVX1  INVX1_236
timestamp 1516325494
transform -1 0 3824 0 1 249
box 0 0 11 49
use INVX1  INVX1_235
timestamp 1516325494
transform -1 0 3836 0 1 249
box 0 0 11 49
use INVX1  INVX1_253
timestamp 1516325494
transform -1 0 3847 0 1 249
box 0 0 11 49
use BUFX2  BUFX2_871
timestamp 1516325494
transform -1 0 3863 0 1 249
box 0 0 15 49
use FILL  FILL_6_1
timestamp 1516325494
transform 1 0 3863 0 1 249
box 0 0 8 49
use AND2X2  AND2X2_735
timestamp 1516325494
transform -1 0 21 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_600
timestamp 1516325494
transform 1 0 21 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_516
timestamp 1516325494
transform 1 0 40 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_601
timestamp 1516325494
transform -1 0 78 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_529
timestamp 1516325494
transform 1 0 78 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_466
timestamp 1516325494
transform 1 0 97 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_532
timestamp 1516325494
transform 1 0 116 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_531
timestamp 1516325494
transform 1 0 135 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_467
timestamp 1516325494
transform 1 0 154 0 -1 248
box 0 0 19 49
use FILL  FILL_BUFX2_735
timestamp 1516325494
transform 1 0 173 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_735
timestamp 1516325494
transform 1 0 181 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_731
timestamp 1516325494
transform -1 0 204 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_731
timestamp 1516325494
transform -1 0 218 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_526
timestamp 1516325494
transform 1 0 219 0 -1 248
box 0 0 19 49
use INVX1  INVX1_19
timestamp 1516325494
transform 1 0 238 0 -1 248
box 0 0 11 49
use AND2X2  AND2X2_534
timestamp 1516325494
transform -1 0 268 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_766
timestamp 1516325494
transform 1 0 268 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_462
timestamp 1516325494
transform -1 0 306 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_523
timestamp 1516325494
transform -1 0 325 0 -1 248
box 0 0 19 49
use MUX2X1  MUX2X1_682
timestamp 1516325494
transform 1 0 325 0 -1 248
box 0 0 30 49
use FILL  FILL_BUFX2_680
timestamp 1516325494
transform 1 0 355 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_680
timestamp 1516325494
transform 1 0 363 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_730
timestamp 1516325494
transform -1 0 386 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_730
timestamp 1516325494
transform -1 0 401 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_662
timestamp 1516325494
transform 1 0 401 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_663
timestamp 1516325494
transform -1 0 439 0 -1 248
box 0 0 19 49
use FILL  FILL_BUFX2_574
timestamp 1516325494
transform -1 0 447 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_574
timestamp 1516325494
transform -1 0 462 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_592
timestamp 1516325494
transform 1 0 462 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_510
timestamp 1516325494
transform 1 0 481 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_445
timestamp 1516325494
transform 1 0 500 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_588
timestamp 1516325494
transform -1 0 538 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_587
timestamp 1516325494
transform -1 0 557 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_413
timestamp 1516325494
transform -1 0 576 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_443
timestamp 1516325494
transform -1 0 595 0 -1 248
box 0 0 19 49
use FILL  FILL_BUFX2_681
timestamp 1516325494
transform -1 0 603 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_681
timestamp 1516325494
transform -1 0 617 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_732
timestamp 1516325494
transform 1 0 618 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_732
timestamp 1516325494
transform 1 0 625 0 -1 248
box 0 0 15 49
use FILL  FILL_OR2X2_173
timestamp 1516325494
transform -1 0 648 0 -1 248
box 0 0 8 49
use OR2X2  OR2X2_173
timestamp 1516325494
transform -1 0 667 0 -1 248
box 0 0 19 49
use FILL  FILL_AND2X2_185
timestamp 1516325494
transform -1 0 675 0 -1 248
box 0 0 8 49
use AND2X2  AND2X2_185
timestamp 1516325494
transform -1 0 694 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1665
timestamp 1516325494
transform 1 0 694 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1480
timestamp 1516325494
transform 1 0 713 0 -1 248
box 0 0 19 49
use FILL  FILL_OR2X2_186
timestamp 1516325494
transform 1 0 732 0 -1 248
box 0 0 8 49
use OR2X2  OR2X2_186
timestamp 1516325494
transform 1 0 739 0 -1 248
box 0 0 19 49
use FILL  FILL_OR2X2_187
timestamp 1516325494
transform -1 0 766 0 -1 248
box 0 0 8 49
use OR2X2  OR2X2_187
timestamp 1516325494
transform -1 0 785 0 -1 248
box 0 0 19 49
use FILL  FILL_AND2X2_200
timestamp 1516325494
transform -1 0 793 0 -1 248
box 0 0 8 49
use AND2X2  AND2X2_200
timestamp 1516325494
transform -1 0 811 0 -1 248
box 0 0 19 49
use FILL  FILL_AND2X2_197
timestamp 1516325494
transform -1 0 819 0 -1 248
box 0 0 8 49
use AND2X2  AND2X2_197
timestamp 1516325494
transform -1 0 838 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1682
timestamp 1516325494
transform 1 0 838 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1505
timestamp 1516325494
transform 1 0 857 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1510
timestamp 1516325494
transform -1 0 895 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1688
timestamp 1516325494
transform -1 0 914 0 -1 248
box 0 0 19 49
use FILL  FILL_BUFX2_747
timestamp 1516325494
transform 1 0 914 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_747
timestamp 1516325494
transform 1 0 922 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_748
timestamp 1516325494
transform -1 0 945 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_748
timestamp 1516325494
transform -1 0 959 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_691
timestamp 1516325494
transform 1 0 960 0 -1 248
box 0 0 53 49
use OR2X2  OR2X2_1564
timestamp 1516325494
transform -1 0 1032 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_307
timestamp 1516325494
transform 1 0 1032 0 -1 248
box 0 0 15 49
use MUX2X1  MUX2X1_307
timestamp 1516325494
transform -1 0 1077 0 -1 248
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_563
timestamp 1516325494
transform 1 0 1077 0 -1 248
box 0 0 53 49
use NAND2X1  NAND2X1_467
timestamp 1516325494
transform 1 0 1131 0 -1 248
box 0 0 15 49
use MUX2X1  MUX2X1_467
timestamp 1516325494
transform -1 0 1176 0 -1 248
box 0 0 30 49
use AND2X2  AND2X2_1727
timestamp 1516325494
transform -1 0 1195 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1562
timestamp 1516325494
transform -1 0 1214 0 -1 248
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_435
timestamp 1516325494
transform 1 0 1214 0 -1 248
box 0 0 53 49
use NAND2X1  NAND2X1_403
timestamp 1516325494
transform 1 0 1267 0 -1 248
box 0 0 15 49
use MUX2X1  MUX2X1_403
timestamp 1516325494
transform -1 0 1313 0 -1 248
box 0 0 30 49
use FILL  FILL_BUFX2_436
timestamp 1516325494
transform 1 0 1313 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_436
timestamp 1516325494
transform 1 0 1321 0 -1 248
box 0 0 15 49
use OR2X2  OR2X2_1561
timestamp 1516325494
transform -1 0 1355 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1052
timestamp 1516325494
transform -1 0 1374 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_386
timestamp 1516325494
transform 1 0 1374 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_418
timestamp 1516325494
transform 1 0 1389 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_386
timestamp 1516325494
transform -1 0 1472 0 -1 248
box 0 0 30 49
use OR2X2  OR2X2_615
timestamp 1516325494
transform 1 0 2 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_737
timestamp 1516325494
transform 1 0 21 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_616
timestamp 1516325494
transform 1 0 40 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_736
timestamp 1516325494
transform -1 0 78 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_605
timestamp 1516325494
transform 1 0 78 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_518
timestamp 1516325494
transform -1 0 116 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_602
timestamp 1516325494
transform -1 0 135 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_719
timestamp 1516325494
transform 1 0 135 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_572
timestamp 1516325494
transform 1 0 154 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_672
timestamp 1516325494
transform -1 0 192 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_573
timestamp 1516325494
transform 1 0 192 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_573
timestamp 1516325494
transform 1 0 200 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_683
timestamp 1516325494
transform -1 0 245 0 1 150
box 0 0 30 49
use OR2X2  OR2X2_469
timestamp 1516325494
transform 1 0 245 0 1 150
box 0 0 19 49
use MUX2X1  MUX2X1_695
timestamp 1516325494
transform 1 0 264 0 1 150
box 0 0 30 49
use MUX2X1  MUX2X1_684
timestamp 1516325494
transform 1 0 295 0 1 150
box 0 0 30 49
use FILL  FILL_BUFX2_400
timestamp 1516325494
transform 1 0 325 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_400
timestamp 1516325494
transform 1 0 333 0 1 150
box 0 0 15 49
use FILL  FILL_BUFX2_679
timestamp 1516325494
transform 1 0 348 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_679
timestamp 1516325494
transform 1 0 355 0 1 150
box 0 0 15 49
use FILL  FILL_BUFX2_575
timestamp 1516325494
transform -1 0 379 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_575
timestamp 1516325494
transform -1 0 393 0 1 150
box 0 0 15 49
use AND2X2  AND2X2_664
timestamp 1516325494
transform -1 0 412 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_559
timestamp 1516325494
transform -1 0 431 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_401
timestamp 1516325494
transform -1 0 439 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_401
timestamp 1516325494
transform -1 0 454 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_560
timestamp 1516325494
transform -1 0 473 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_661
timestamp 1516325494
transform -1 0 492 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_589
timestamp 1516325494
transform -1 0 511 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_508
timestamp 1516325494
transform -1 0 530 0 1 150
box 0 0 19 49
use FILL  FILL_OR2X2_90
timestamp 1516325494
transform 1 0 530 0 1 150
box 0 0 8 49
use OR2X2  OR2X2_90
timestamp 1516325494
transform 1 0 538 0 1 150
box 0 0 19 49
use FILL  FILL_OR2X2_104
timestamp 1516325494
transform 1 0 557 0 1 150
box 0 0 8 49
use OR2X2  OR2X2_104
timestamp 1516325494
transform 1 0 564 0 1 150
box 0 0 19 49
use FILL  FILL_OR2X2_160
timestamp 1516325494
transform 1 0 583 0 1 150
box 0 0 8 49
use OR2X2  OR2X2_160
timestamp 1516325494
transform 1 0 591 0 1 150
box 0 0 19 49
use INVX1  INVX1_176
timestamp 1516325494
transform -1 0 621 0 1 150
box 0 0 11 49
use OR2X2  OR2X2_1445
timestamp 1516325494
transform 1 0 621 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1451
timestamp 1516325494
transform 1 0 640 0 1 150
box 0 0 19 49
use INVX1  INVX1_168
timestamp 1516325494
transform -1 0 670 0 1 150
box 0 0 11 49
use FILL  FILL_AND2X2_184
timestamp 1516325494
transform -1 0 679 0 1 150
box 0 0 8 49
use AND2X2  AND2X2_184
timestamp 1516325494
transform -1 0 697 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1663
timestamp 1516325494
transform 1 0 697 0 1 150
box 0 0 19 49
use FILL  FILL_AND2X2_198
timestamp 1516325494
transform -1 0 724 0 1 150
box 0 0 8 49
use AND2X2  AND2X2_198
timestamp 1516325494
transform -1 0 743 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1684
timestamp 1516325494
transform 1 0 743 0 1 150
box 0 0 19 49
use FILL  FILL_AND2X2_199
timestamp 1516325494
transform -1 0 770 0 1 150
box 0 0 8 49
use AND2X2  AND2X2_199
timestamp 1516325494
transform -1 0 789 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1683
timestamp 1516325494
transform -1 0 808 0 1 150
box 0 0 19 49
use FILL  FILL_OR2X2_34
timestamp 1516325494
transform 1 0 808 0 1 150
box 0 0 8 49
use OR2X2  OR2X2_34
timestamp 1516325494
transform 1 0 815 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_685
timestamp 1516325494
transform 1 0 834 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_685
timestamp 1516325494
transform 1 0 842 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_1504
timestamp 1516325494
transform -1 0 876 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1686
timestamp 1516325494
transform 1 0 876 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_689
timestamp 1516325494
transform 1 0 895 0 1 150
box 0 0 53 49
use NAND2X1  NAND2X1_305
timestamp 1516325494
transform 1 0 948 0 1 150
box 0 0 15 49
use NAND2X1  NAND2X1_472
timestamp 1516325494
transform -1 0 978 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_305
timestamp 1516325494
transform -1 0 1009 0 1 150
box 0 0 30 49
use NAND2X1  NAND2X1_465
timestamp 1516325494
transform 1 0 1009 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_465
timestamp 1516325494
transform -1 0 1054 0 1 150
box 0 0 30 49
use OR2X2  OR2X2_1713
timestamp 1516325494
transform 1 0 1055 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_24
timestamp 1516325494
transform 1 0 1074 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_24
timestamp 1516325494
transform 1 0 1081 0 1 150
box 0 0 15 49
use AND2X2  AND2X2_1844
timestamp 1516325494
transform -1 0 1115 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1714
timestamp 1516325494
transform -1 0 1134 0 1 150
box 0 0 19 49
use NAND2X1  NAND2X1_312
timestamp 1516325494
transform 1 0 1134 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_312
timestamp 1516325494
transform -1 0 1180 0 1 150
box 0 0 30 49
use OR2X2  OR2X2_1712
timestamp 1516325494
transform 1 0 1180 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1842
timestamp 1516325494
transform 1 0 1199 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1711
timestamp 1516325494
transform -1 0 1237 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_600
timestamp 1516325494
transform 1 0 1237 0 1 150
box 0 0 53 49
use NAND2X1  NAND2X1_24
timestamp 1516325494
transform 1 0 1290 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_24
timestamp 1516325494
transform -1 0 1335 0 1 150
box 0 0 30 49
use OR2X2  OR2X2_1053
timestamp 1516325494
transform 1 0 1336 0 1 150
box 0 0 19 49
use NAND2X1  NAND2X1_450
timestamp 1516325494
transform 1 0 1355 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_1059
timestamp 1516325494
transform 1 0 1370 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_546
timestamp 1516325494
transform 1 0 1389 0 1 150
box 0 0 53 49
use MUX2X1  MUX2X1_450
timestamp 1516325494
transform -1 0 1472 0 1 150
box 0 0 30 49
use FILL  FILL_BUFX2_512
timestamp 1516325494
transform -1 0 1481 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_512
timestamp 1516325494
transform -1 0 1495 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_764
timestamp 1516325494
transform 1 0 1495 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_764
timestamp 1516325494
transform 1 0 1503 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_28
timestamp 1516325494
transform -1 0 1526 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_28
timestamp 1516325494
transform -1 0 1541 0 -1 248
box 0 0 15 49
use INVX2  INVX2_5
timestamp 1516325494
transform 1 0 1541 0 -1 248
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_656
timestamp 1516325494
transform 1 0 1552 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_48
timestamp 1516325494
transform 1 0 1606 0 -1 248
box 0 0 30 49
use NAND2X1  NAND2X1_48
timestamp 1516325494
transform 1 0 1636 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_592
timestamp 1516325494
transform 1 0 1651 0 -1 248
box 0 0 53 49
use NAND2X1  NAND2X1_16
timestamp 1516325494
transform 1 0 1704 0 -1 248
box 0 0 15 49
use MUX2X1  MUX2X1_16
timestamp 1516325494
transform -1 0 1750 0 -1 248
box 0 0 30 49
use FILL  FILL_BUFX2_474
timestamp 1516325494
transform 1 0 1750 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_474
timestamp 1516325494
transform 1 0 1758 0 -1 248
box 0 0 15 49
use OR2X2  OR2X2_1951
timestamp 1516325494
transform 1 0 1773 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_2026
timestamp 1516325494
transform -1 0 1811 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1952
timestamp 1516325494
transform -1 0 1830 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_32
timestamp 1516325494
transform 1 0 1830 0 -1 248
box 0 0 15 49
use MUX2X1  MUX2X1_32
timestamp 1516325494
transform -1 0 1875 0 -1 248
box 0 0 30 49
use MUX2X1  MUX2X1_464
timestamp 1516325494
transform 1 0 1875 0 -1 248
box 0 0 30 49
use MUX2X1  MUX2X1_17
timestamp 1516325494
transform 1 0 1906 0 -1 248
box 0 0 30 49
use NAND2X1  NAND2X1_17
timestamp 1516325494
transform -1 0 1951 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_508
timestamp 1516325494
transform -1 0 1959 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_508
timestamp 1516325494
transform -1 0 1974 0 -1 248
box 0 0 15 49
use NAND2X1  NAND2X1_416
timestamp 1516325494
transform 1 0 1974 0 -1 248
box 0 0 15 49
use MUX2X1  MUX2X1_416
timestamp 1516325494
transform -1 0 2019 0 -1 248
box 0 0 30 49
use OR2X2  OR2X2_1566
timestamp 1516325494
transform 1 0 2020 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_897
timestamp 1516325494
transform 1 0 2039 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_627
timestamp 1516325494
transform 1 0 2054 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_842
timestamp 1516325494
transform -1 0 2137 0 -1 248
box 0 0 30 49
use FILL  FILL_BUFX2_718
timestamp 1516325494
transform 1 0 2138 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_718
timestamp 1516325494
transform 1 0 2145 0 -1 248
box 0 0 15 49
use FILL  FILL_BUFX2_763
timestamp 1516325494
transform -1 0 2168 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_763
timestamp 1516325494
transform -1 0 2183 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_573
timestamp 1516325494
transform 1 0 2183 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_477
timestamp 1516325494
transform -1 0 2266 0 -1 248
box 0 0 30 49
use FILL  FILL_BUFX2_17
timestamp 1516325494
transform 1 0 2267 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_17
timestamp 1516325494
transform 1 0 2274 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_1342
timestamp 1516325494
transform 1 0 1473 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1058
timestamp 1516325494
transform -1 0 1511 0 1 150
box 0 0 19 49
use MUX2X1  MUX2X1_56
timestamp 1516325494
transform 1 0 1511 0 1 150
box 0 0 30 49
use NAND2X1  NAND2X1_56
timestamp 1516325494
transform -1 0 1556 0 1 150
box 0 0 15 49
use AND2X2  AND2X2_1664
timestamp 1516325494
transform 1 0 1556 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1478
timestamp 1516325494
transform -1 0 1594 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_664
timestamp 1516325494
transform -1 0 1647 0 1 150
box 0 0 53 49
use OR2X2  OR2X2_1718
timestamp 1516325494
transform 1 0 1647 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1848
timestamp 1516325494
transform -1 0 1685 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_15
timestamp 1516325494
transform -1 0 1693 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_15
timestamp 1516325494
transform -1 0 1708 0 1 150
box 0 0 15 49
use AND2X2  AND2X2_1572
timestamp 1516325494
transform -1 0 1727 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1358
timestamp 1516325494
transform -1 0 1746 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_652
timestamp 1516325494
transform 1 0 1746 0 1 150
box 0 0 53 49
use NAND2X1  NAND2X1_44
timestamp 1516325494
transform 1 0 1799 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_44
timestamp 1516325494
transform -1 0 1845 0 1 150
box 0 0 30 49
use OR2X2  OR2X2_1474
timestamp 1516325494
transform -1 0 1864 0 1 150
box 0 0 19 49
use NAND2X1  NAND2X1_304
timestamp 1516325494
transform -1 0 1879 0 1 150
box 0 0 15 49
use AND2X2  AND2X2_1570
timestamp 1516325494
transform 1 0 1879 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_608
timestamp 1516325494
transform -1 0 1951 0 1 150
box 0 0 53 49
use MUX2X1  MUX2X1_304
timestamp 1516325494
transform -1 0 1981 0 1 150
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_688
timestamp 1516325494
transform -1 0 2035 0 1 150
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_593
timestamp 1516325494
transform -1 0 2088 0 1 150
box 0 0 53 49
use OR2X2  OR2X2_1501
timestamp 1516325494
transform 1 0 2088 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1681
timestamp 1516325494
transform -1 0 2126 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_594
timestamp 1516325494
transform 1 0 2126 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_594
timestamp 1516325494
transform 1 0 2134 0 1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_448
timestamp 1516325494
transform -1 0 2202 0 1 150
box 0 0 53 49
use OR2X2  OR2X2_1324
timestamp 1516325494
transform -1 0 2221 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_683
timestamp 1516325494
transform 1 0 2221 0 1 150
box 0 0 53 49
use NAND2X1  NAND2X1_299
timestamp 1516325494
transform 1 0 2274 0 1 150
box 0 0 15 49
use FILL  FILL_BUFX2_719
timestamp 1516325494
transform -1 0 2298 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_719
timestamp 1516325494
transform -1 0 2312 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_1687
timestamp 1516325494
transform -1 0 2331 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1509
timestamp 1516325494
transform -1 0 2350 0 -1 248
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_305
timestamp 1516325494
transform 1 0 2350 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_497
timestamp 1516325494
transform -1 0 2434 0 -1 248
box 0 0 30 49
use FILL  FILL_BUFX2_314
timestamp 1516325494
transform 1 0 2434 0 -1 248
box 0 0 8 49
use BUFX2  BUFX2_314
timestamp 1516325494
transform 1 0 2442 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_1963
timestamp 1516325494
transform -1 0 2476 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_1869
timestamp 1516325494
transform -1 0 2495 0 -1 248
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_669
timestamp 1516325494
transform -1 0 2548 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_509
timestamp 1516325494
transform 1 0 2548 0 -1 248
box 0 0 30 49
use NAND2X1  NAND2X1_509
timestamp 1516325494
transform -1 0 2593 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_317
timestamp 1516325494
transform -1 0 2647 0 -1 248
box 0 0 53 49
use NAND2X1  NAND2X1_902
timestamp 1516325494
transform 1 0 2647 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_632
timestamp 1516325494
transform 1 0 2662 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_847
timestamp 1516325494
transform -1 0 2745 0 -1 248
box 0 0 30 49
use AND2X2  AND2X2_298
timestamp 1516325494
transform 1 0 2746 0 -1 248
box 0 0 19 49
use MUX2X1  MUX2X1_623
timestamp 1516325494
transform 1 0 2765 0 -1 248
box 0 0 30 49
use NAND2X1  NAND2X1_623
timestamp 1516325494
transform -1 0 2810 0 -1 248
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_207
timestamp 1516325494
transform -1 0 2863 0 -1 248
box 0 0 53 49
use MUX2X1  MUX2X1_591
timestamp 1516325494
transform 1 0 2863 0 -1 248
box 0 0 30 49
use FILL  FILL_AND2X2_162
timestamp 1516325494
transform 1 0 2894 0 -1 248
box 0 0 8 49
use AND2X2  AND2X2_162
timestamp 1516325494
transform 1 0 2901 0 -1 248
box 0 0 19 49
use FILL  FILL_AND2X2_103
timestamp 1516325494
transform 1 0 2920 0 -1 248
box 0 0 8 49
use AND2X2  AND2X2_103
timestamp 1516325494
transform 1 0 2928 0 -1 248
box 0 0 19 49
use FILL  FILL_OR2X2_97
timestamp 1516325494
transform 1 0 2947 0 -1 248
box 0 0 8 49
use OR2X2  OR2X2_97
timestamp 1516325494
transform 1 0 2955 0 -1 248
box 0 0 19 49
use FILL  FILL_AND2X2_102
timestamp 1516325494
transform -1 0 2982 0 -1 248
box 0 0 8 49
use AND2X2  AND2X2_102
timestamp 1516325494
transform -1 0 3000 0 -1 248
box 0 0 19 49
use FILL  FILL_OR2X2_98
timestamp 1516325494
transform 1 0 3000 0 -1 248
box 0 0 8 49
use OR2X2  OR2X2_98
timestamp 1516325494
transform 1 0 3008 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1139
timestamp 1516325494
transform 1 0 3027 0 -1 248
box 0 0 19 49
use XOR2X1  XOR2X1_63
timestamp 1516325494
transform -1 0 3080 0 -1 248
box 0 0 34 49
use AND2X2  AND2X2_1173
timestamp 1516325494
transform -1 0 3099 0 -1 248
box 0 0 19 49
use NOR2X1  NOR2X1_123
timestamp 1516325494
transform -1 0 3114 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_1142
timestamp 1516325494
transform 1 0 3114 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1143
timestamp 1516325494
transform 1 0 3133 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_930
timestamp 1516325494
transform -1 0 3171 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1141
timestamp 1516325494
transform -1 0 3190 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1172
timestamp 1516325494
transform -1 0 3209 0 -1 248
box 0 0 19 49
use XOR2X1  XOR2X1_66
timestamp 1516325494
transform -1 0 3243 0 -1 248
box 0 0 34 49
use AND2X2  AND2X2_1169
timestamp 1516325494
transform -1 0 3262 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_948
timestamp 1516325494
transform -1 0 3281 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_950
timestamp 1516325494
transform -1 0 3300 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1176
timestamp 1516325494
transform -1 0 3319 0 -1 248
box 0 0 19 49
use MUX2X1  MUX2X1_811
timestamp 1516325494
transform -1 0 3349 0 -1 248
box 0 0 30 49
use AND2X2  AND2X2_1164
timestamp 1516325494
transform -1 0 3369 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1168
timestamp 1516325494
transform -1 0 3388 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_943
timestamp 1516325494
transform -1 0 3407 0 -1 248
box 0 0 19 49
use INVX1  INVX1_257
timestamp 1516325494
transform -1 0 3418 0 -1 248
box 0 0 11 49
use OR2X2  OR2X2_926
timestamp 1516325494
transform -1 0 3437 0 -1 248
box 0 0 19 49
use OR2X2  OR2X2_925
timestamp 1516325494
transform -1 0 3456 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1163
timestamp 1516325494
transform -1 0 3475 0 -1 248
box 0 0 19 49
use AND2X2  AND2X2_1162
timestamp 1516325494
transform -1 0 3494 0 -1 248
box 0 0 19 49
use AOI22X1  AOI22X1_5
timestamp 1516325494
transform -1 0 3517 0 -1 248
box 0 0 23 49
use NAND2X1  NAND2X1_768
timestamp 1516325494
transform -1 0 3532 0 -1 248
box 0 0 15 49
use NAND2X1  NAND2X1_766
timestamp 1516325494
transform -1 0 3547 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_1126
timestamp 1516325494
transform -1 0 3566 0 -1 248
box 0 0 19 49
use AOI21X1  AOI21X1_45
timestamp 1516325494
transform 1 0 3566 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_756
timestamp 1516325494
transform 1 0 3585 0 -1 248
box 0 0 15 49
use AND2X2  AND2X2_1125
timestamp 1516325494
transform -1 0 3620 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_759
timestamp 1516325494
transform -1 0 3635 0 -1 248
box 0 0 15 49
use NOR3X1  NOR3X1_13
timestamp 1516325494
transform 1 0 3635 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_761
timestamp 1516325494
transform 1 0 3654 0 -1 248
box 0 0 15 49
use NOR3X1  NOR3X1_22
timestamp 1516325494
transform -1 0 3688 0 -1 248
box 0 0 19 49
use NOR2X1  NOR2X1_121
timestamp 1516325494
transform -1 0 3703 0 -1 248
box 0 0 15 49
use NAND3X1  NAND3X1_69
timestamp 1516325494
transform 1 0 3703 0 -1 248
box 0 0 19 49
use NAND3X1  NAND3X1_72
timestamp 1516325494
transform 1 0 3722 0 -1 248
box 0 0 19 49
use NAND2X1  NAND2X1_760
timestamp 1516325494
transform -1 0 3756 0 -1 248
box 0 0 15 49
use INVX1  INVX1_249
timestamp 1516325494
transform -1 0 3767 0 -1 248
box 0 0 11 49
use NOR3X1  NOR3X1_21
timestamp 1516325494
transform 1 0 3768 0 -1 248
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_780
timestamp 1516325494
transform 1 0 3787 0 -1 248
box 0 0 53 49
use AND2X2  AND2X2_1229
timestamp 1516325494
transform -1 0 3859 0 -1 248
box 0 0 19 49
use FILL  FILL_5_1
timestamp 1516325494
transform -1 0 3867 0 -1 248
box 0 0 8 49
use MUX2X1  MUX2X1_299
timestamp 1516325494
transform -1 0 2320 0 1 150
box 0 0 30 49
use FILL  FILL_BUFX2_418
timestamp 1516325494
transform 1 0 2320 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_418
timestamp 1516325494
transform 1 0 2328 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_1719
timestamp 1516325494
transform -1 0 2362 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1507
timestamp 1516325494
transform 1 0 2362 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1685
timestamp 1516325494
transform 1 0 2381 0 1 150
box 0 0 19 49
use NAND2X1  NAND2X1_497
timestamp 1516325494
transform 1 0 2400 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_1506
timestamp 1516325494
transform -1 0 2434 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_503
timestamp 1516325494
transform 1 0 2434 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_503
timestamp 1516325494
transform 1 0 2442 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_1867
timestamp 1516325494
transform 1 0 2457 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1961
timestamp 1516325494
transform 1 0 2476 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_443
timestamp 1516325494
transform -1 0 2503 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_443
timestamp 1516325494
transform -1 0 2517 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_61
timestamp 1516325494
transform 1 0 2518 0 1 150
box 0 0 30 49
use NAND2X1  NAND2X1_61
timestamp 1516325494
transform -1 0 2563 0 1 150
box 0 0 15 49
use OR2X2  OR2X2_1868
timestamp 1516325494
transform -1 0 2582 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_1866
timestamp 1516325494
transform -1 0 2601 0 1 150
box 0 0 19 49
use FILL  FILL_BUFX2_509
timestamp 1516325494
transform 1 0 2601 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_509
timestamp 1516325494
transform 1 0 2609 0 1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_312
timestamp 1516325494
transform 1 0 2624 0 1 150
box 0 0 53 49
use FILL  FILL_BUFX2_467
timestamp 1516325494
transform 1 0 2677 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_467
timestamp 1516325494
transform 1 0 2685 0 1 150
box 0 0 15 49
use FILL  FILL_BUFX2_479
timestamp 1516325494
transform -1 0 2708 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_479
timestamp 1516325494
transform -1 0 2723 0 1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_766
timestamp 1516325494
transform 1 0 2723 0 1 150
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_248
timestamp 1516325494
transform 1 0 2776 0 1 150
box 0 0 53 49
use NAND2X1  NAND2X1_216
timestamp 1516325494
transform 1 0 2829 0 1 150
box 0 0 15 49
use FILL  FILL_BUFX2_8
timestamp 1516325494
transform -1 0 2852 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_8
timestamp 1516325494
transform -1 0 2867 0 1 150
box 0 0 15 49
use NAND2X1  NAND2X1_207
timestamp 1516325494
transform -1 0 2882 0 1 150
box 0 0 15 49
use MUX2X1  MUX2X1_587
timestamp 1516325494
transform 1 0 2882 0 1 150
box 0 0 30 49
use NAND2X1  NAND2X1_587
timestamp 1516325494
transform -1 0 2928 0 1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_716
timestamp 1516325494
transform 1 0 2928 0 1 150
box 0 0 53 49
use AND2X2  AND2X2_1180
timestamp 1516325494
transform -1 0 3000 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1170
timestamp 1516325494
transform 1 0 3000 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1178
timestamp 1516325494
transform -1 0 3038 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1174
timestamp 1516325494
transform -1 0 3057 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_949
timestamp 1516325494
transform -1 0 3076 0 1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_761
timestamp 1516325494
transform 1 0 3076 0 1 150
box 0 0 53 49
use AND2X2  AND2X2_1144
timestamp 1516325494
transform -1 0 3148 0 1 150
box 0 0 19 49
use XOR2X1  XOR2X1_65
timestamp 1516325494
transform 1 0 3148 0 1 150
box 0 0 34 49
use AND2X2  AND2X2_1171
timestamp 1516325494
transform 1 0 3183 0 1 150
box 0 0 19 49
use XOR2X1  XOR2X1_67
timestamp 1516325494
transform -1 0 3236 0 1 150
box 0 0 34 49
use NOR2X1  NOR2X1_128
timestamp 1516325494
transform 1 0 3236 0 1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_774
timestamp 1516325494
transform -1 0 3304 0 1 150
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_776
timestamp 1516325494
transform 1 0 3304 0 1 150
box 0 0 53 49
use AND2X2  AND2X2_1124
timestamp 1516325494
transform -1 0 3376 0 1 150
box 0 0 19 49
use NAND2X1  NAND2X1_753
timestamp 1516325494
transform -1 0 3391 0 1 150
box 0 0 15 49
use AOI21X1  AOI21X1_29
timestamp 1516325494
transform -1 0 3411 0 1 150
box 0 0 19 49
use MUX2X1  MUX2X1_813
timestamp 1516325494
transform -1 0 3441 0 1 150
box 0 0 30 49
use FILL  FILL_BUFX2_187
timestamp 1516325494
transform 1 0 3441 0 1 150
box 0 0 8 49
use BUFX2  BUFX2_187
timestamp 1516325494
transform 1 0 3449 0 1 150
box 0 0 15 49
use AOI21X1  AOI21X1_39
timestamp 1516325494
transform -1 0 3483 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_947
timestamp 1516325494
transform -1 0 3502 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_945
timestamp 1516325494
transform -1 0 3521 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_946
timestamp 1516325494
transform -1 0 3540 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_1167
timestamp 1516325494
transform -1 0 3559 0 1 150
box 0 0 19 49
use NOR2X1  NOR2X1_111
timestamp 1516325494
transform 1 0 3559 0 1 150
box 0 0 15 49
use INVX1  INVX1_238
timestamp 1516325494
transform 1 0 3574 0 1 150
box 0 0 11 49
use AOI21X1  AOI21X1_47
timestamp 1516325494
transform 1 0 3585 0 1 150
box 0 0 19 49
use AOI21X1  AOI21X1_46
timestamp 1516325494
transform 1 0 3604 0 1 150
box 0 0 19 49
use NOR3X1  NOR3X1_29
timestamp 1516325494
transform 1 0 3623 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_952
timestamp 1516325494
transform 1 0 3642 0 1 150
box 0 0 19 49
use NOR2X1  NOR2X1_112
timestamp 1516325494
transform 1 0 3661 0 1 150
box 0 0 15 49
use OAI21X1  OAI21X1_92
timestamp 1516325494
transform 1 0 3677 0 1 150
box 0 0 19 49
use INVX1  INVX1_240
timestamp 1516325494
transform -1 0 3707 0 1 150
box 0 0 11 49
use NOR2X1  NOR2X1_120
timestamp 1516325494
transform 1 0 3707 0 1 150
box 0 0 15 49
use NAND3X1  NAND3X1_71
timestamp 1516325494
transform 1 0 3722 0 1 150
box 0 0 19 49
use AOI21X1  AOI21X1_36
timestamp 1516325494
transform 1 0 3741 0 1 150
box 0 0 19 49
use AOI21X1  AOI21X1_35
timestamp 1516325494
transform -1 0 3779 0 1 150
box 0 0 19 49
use INVX1  INVX1_256
timestamp 1516325494
transform 1 0 3779 0 1 150
box 0 0 11 49
use NAND3X1  NAND3X1_70
timestamp 1516325494
transform -1 0 3810 0 1 150
box 0 0 19 49
use NOR3X1  NOR3X1_16
timestamp 1516325494
transform -1 0 3829 0 1 150
box 0 0 19 49
use NOR3X1  NOR3X1_17
timestamp 1516325494
transform 1 0 3829 0 1 150
box 0 0 19 49
use OR2X2  OR2X2_920
timestamp 1516325494
transform 1 0 3848 0 1 150
box 0 0 19 49
use AND2X2  AND2X2_734
timestamp 1516325494
transform 1 0 2 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_517
timestamp 1516325494
transform -1 0 40 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_604
timestamp 1516325494
transform -1 0 59 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_603
timestamp 1516325494
transform -1 0 78 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_673
timestamp 1516325494
transform 1 0 78 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_571
timestamp 1516325494
transform 1 0 97 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_674
timestamp 1516325494
transform 1 0 116 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_675
timestamp 1516325494
transform 1 0 135 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_530
timestamp 1516325494
transform 1 0 154 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_533
timestamp 1516325494
transform 1 0 173 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_468
timestamp 1516325494
transform 1 0 192 0 -1 150
box 0 0 19 49
use FILL  FILL_BUFX2_571
timestamp 1516325494
transform 1 0 211 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_571
timestamp 1516325494
transform 1 0 219 0 -1 150
box 0 0 15 49
use AND2X2  AND2X2_527
timestamp 1516325494
transform 1 0 234 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_463
timestamp 1516325494
transform -1 0 272 0 -1 150
box 0 0 19 49
use BUFX2  BUFX2_888
timestamp 1516325494
transform 1 0 272 0 -1 150
box 0 0 15 49
use OR2X2  OR2X2_1301
timestamp 1516325494
transform -1 0 306 0 -1 150
box 0 0 19 49
use FILL  FILL_OR2X2_88
timestamp 1516325494
transform 1 0 306 0 -1 150
box 0 0 8 49
use OR2X2  OR2X2_88
timestamp 1516325494
transform 1 0 314 0 -1 150
box 0 0 19 49
use FILL  FILL_OR2X2_102
timestamp 1516325494
transform 1 0 333 0 -1 150
box 0 0 8 49
use OR2X2  OR2X2_102
timestamp 1516325494
transform 1 0 340 0 -1 150
box 0 0 19 49
use FILL  FILL_AND2X2_108
timestamp 1516325494
transform -1 0 367 0 -1 150
box 0 0 8 49
use AND2X2  AND2X2_108
timestamp 1516325494
transform -1 0 386 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1546
timestamp 1516325494
transform -1 0 405 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1523
timestamp 1516325494
transform -1 0 424 0 -1 150
box 0 0 19 49
use FILL  FILL_AND2X2_93
timestamp 1516325494
transform -1 0 432 0 -1 150
box 0 0 8 49
use AND2X2  AND2X2_93
timestamp 1516325494
transform -1 0 450 0 -1 150
box 0 0 19 49
use FILL  FILL_AND2X2_168
timestamp 1516325494
transform 1 0 450 0 -1 150
box 0 0 8 49
use AND2X2  AND2X2_168
timestamp 1516325494
transform 1 0 458 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1522
timestamp 1516325494
transform 1 0 477 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1431
timestamp 1516325494
transform -1 0 515 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1638
timestamp 1516325494
transform 1 0 515 0 -1 150
box 0 0 19 49
use FILL  FILL_OR2X2_158
timestamp 1516325494
transform 1 0 534 0 -1 150
box 0 0 8 49
use OR2X2  OR2X2_158
timestamp 1516325494
transform 1 0 542 0 -1 150
box 0 0 19 49
use FILL  FILL_AND2X2_167
timestamp 1516325494
transform -1 0 569 0 -1 150
box 0 0 8 49
use AND2X2  AND2X2_167
timestamp 1516325494
transform -1 0 587 0 -1 150
box 0 0 19 49
use FILL  FILL_AND2X2_33
timestamp 1516325494
transform 1 0 587 0 -1 150
box 0 0 8 49
use AND2X2  AND2X2_33
timestamp 1516325494
transform 1 0 595 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1636
timestamp 1516325494
transform 1 0 614 0 -1 150
box 0 0 19 49
use FILL  FILL_OR2X2_32
timestamp 1516325494
transform 1 0 633 0 -1 150
box 0 0 8 49
use OR2X2  OR2X2_32
timestamp 1516325494
transform 1 0 640 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_1293
timestamp 1516325494
transform -1 0 678 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_554
timestamp 1516325494
transform 1 0 678 0 -1 150
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_561
timestamp 1516325494
transform -1 0 785 0 -1 150
box 0 0 53 49
use OR2X2  OR2X2_1503
timestamp 1516325494
transform 1 0 785 0 -1 150
box 0 0 19 49
use NAND2X1  NAND2X1_458
timestamp 1516325494
transform 1 0 804 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_458
timestamp 1516325494
transform -1 0 849 0 -1 150
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_568
timestamp 1516325494
transform 1 0 849 0 -1 150
box 0 0 53 49
use AND2X2  AND2X2_1733
timestamp 1516325494
transform -1 0 922 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_1569
timestamp 1516325494
transform -1 0 941 0 -1 150
box 0 0 19 49
use MUX2X1  MUX2X1_472
timestamp 1516325494
transform 1 0 941 0 -1 150
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_696
timestamp 1516325494
transform 1 0 971 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_408
timestamp 1516325494
transform 1 0 1024 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_408
timestamp 1516325494
transform -1 0 1069 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_499
timestamp 1516325494
transform 1 0 1070 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_499
timestamp 1516325494
transform -1 0 1115 0 -1 150
box 0 0 30 49
use FILL  FILL_BUFX2_428
timestamp 1516325494
transform 1 0 1115 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_428
timestamp 1516325494
transform 1 0 1123 0 -1 150
box 0 0 15 49
use FILL  FILL_BUFX2_238
timestamp 1516325494
transform -1 0 1146 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_238
timestamp 1516325494
transform -1 0 1161 0 -1 150
box 0 0 15 49
use AND2X2  AND2X2_1430
timestamp 1516325494
transform -1 0 1180 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_1174
timestamp 1516325494
transform -1 0 1199 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_1173
timestamp 1516325494
transform -1 0 1218 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_678
timestamp 1516325494
transform 1 0 1218 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_294
timestamp 1516325494
transform 1 0 1271 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_294
timestamp 1516325494
transform -1 0 1316 0 -1 150
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_290
timestamp 1516325494
transform 1 0 1317 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_482
timestamp 1516325494
transform 1 0 1370 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_482
timestamp 1516325494
transform -1 0 1415 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_34
timestamp 1516325494
transform 1 0 1416 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_34
timestamp 1516325494
transform -1 0 1461 0 -1 150
box 0 0 30 49
use MUX2X1  MUX2X1_6
timestamp 1516325494
transform 1 0 1461 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_6
timestamp 1516325494
transform -1 0 1507 0 -1 150
box 0 0 15 49
use OR2X2  OR2X2_1171
timestamp 1516325494
transform 1 0 1507 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_550
timestamp 1516325494
transform 1 0 1526 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_454
timestamp 1516325494
transform 1 0 1579 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_454
timestamp 1516325494
transform -1 0 1624 0 -1 150
box 0 0 30 49
use FILL  FILL_BUFX2_444
timestamp 1516325494
transform 1 0 1625 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_444
timestamp 1516325494
transform 1 0 1632 0 -1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_300
timestamp 1516325494
transform 1 0 1647 0 -1 150
box 0 0 53 49
use OR2X2  OR2X2_1359
timestamp 1516325494
transform 1 0 1701 0 -1 150
box 0 0 19 49
use NAND2X1  NAND2X1_492
timestamp 1516325494
transform 1 0 1720 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_492
timestamp 1516325494
transform -1 0 1765 0 -1 150
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_44
timestamp 1516325494
transform 1 0 1765 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_428
timestamp 1516325494
transform 1 0 1818 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_428
timestamp 1516325494
transform -1 0 1864 0 -1 150
box 0 0 30 49
use OR2X2  OR2X2_1357
timestamp 1516325494
transform 1 0 1864 0 -1 150
box 0 0 19 49
use FILL  FILL_BUFX2_410
timestamp 1516325494
transform -1 0 1891 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_410
timestamp 1516325494
transform -1 0 1906 0 -1 150
box 0 0 15 49
use OR2X2  OR2X2_1356
timestamp 1516325494
transform -1 0 1925 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_620
timestamp 1516325494
transform 1 0 1925 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_890
timestamp 1516325494
transform 1 0 1978 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_835
timestamp 1516325494
transform -1 0 2023 0 -1 150
box 0 0 30 49
use FILL  FILL_BUFX2_20
timestamp 1516325494
transform 1 0 2024 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_20
timestamp 1516325494
transform 1 0 2031 0 -1 150
box 0 0 15 49
use AND2X2  AND2X2_1545
timestamp 1516325494
transform -1 0 2065 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_1323
timestamp 1516325494
transform -1 0 2084 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_1502
timestamp 1516325494
transform 1 0 2084 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_433
timestamp 1516325494
transform 1 0 2103 0 -1 150
box 0 0 53 49
use NAND2X1  NAND2X1_401
timestamp 1516325494
transform 1 0 2157 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_401
timestamp 1516325494
transform -1 0 2202 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_459
timestamp 1516325494
transform 1 0 2202 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_459
timestamp 1516325494
transform -1 0 2247 0 -1 150
box 0 0 30 49
use FILL  FILL_BUFX2_860
timestamp 1516325494
transform 1 0 2248 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_860
timestamp 1516325494
transform 1 0 2255 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_433
timestamp 1516325494
transform 1 0 2271 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_433
timestamp 1516325494
transform -1 0 2316 0 -1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_49
timestamp 1516325494
transform -1 0 2369 0 -1 150
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_61
timestamp 1516325494
transform 1 0 2369 0 -1 150
box 0 0 53 49
use MUX2X1  MUX2X1_445
timestamp 1516325494
transform 1 0 2423 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_445
timestamp 1516325494
transform 1 0 2453 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_490
timestamp 1516325494
transform 1 0 2468 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_490
timestamp 1516325494
transform -1 0 2514 0 -1 150
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_298
timestamp 1516325494
transform -1 0 2567 0 -1 150
box 0 0 53 49
use MUX2X1  MUX2X1_852
timestamp 1516325494
transform 1 0 2567 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_907
timestamp 1516325494
transform 1 0 2597 0 -1 150
box 0 0 15 49
use FILL  FILL_BUFX2_174
timestamp 1516325494
transform 1 0 2613 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_174
timestamp 1516325494
transform 1 0 2620 0 -1 150
box 0 0 15 49
use NAND2X1  NAND2X1_504
timestamp 1516325494
transform 1 0 2635 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_504
timestamp 1516325494
transform -1 0 2681 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_889
timestamp 1516325494
transform 1 0 2681 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_834
timestamp 1516325494
transform -1 0 2726 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_427
timestamp 1516325494
transform 1 0 2727 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_427
timestamp 1516325494
transform -1 0 2772 0 -1 150
box 0 0 30 49
use MUX2X1  MUX2X1_600
timestamp 1516325494
transform 1 0 2772 0 -1 150
box 0 0 30 49
use NAND2X1  NAND2X1_600
timestamp 1516325494
transform -1 0 2818 0 -1 150
box 0 0 15 49
use MUX2X1  MUX2X1_216
timestamp 1516325494
transform 1 0 2818 0 -1 150
box 0 0 30 49
use MUX2X1  MUX2X1_207
timestamp 1516325494
transform 1 0 2848 0 -1 150
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_267
timestamp 1516325494
transform -1 0 2932 0 -1 150
box 0 0 53 49
use XOR2X1  XOR2X1_69
timestamp 1516325494
transform -1 0 2966 0 -1 150
box 0 0 34 49
use AND2X2  AND2X2_1179
timestamp 1516325494
transform 1 0 2966 0 -1 150
box 0 0 19 49
use XOR2X1  XOR2X1_64
timestamp 1516325494
transform -1 0 3019 0 -1 150
box 0 0 34 49
use AND2X2  AND2X2_1159
timestamp 1516325494
transform 1 0 3019 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_755
timestamp 1516325494
transform -1 0 3091 0 -1 150
box 0 0 53 49
use FILL  FILL_BUFX2_199
timestamp 1516325494
transform -1 0 3099 0 -1 150
box 0 0 8 49
use BUFX2  BUFX2_199
timestamp 1516325494
transform -1 0 3114 0 -1 150
box 0 0 15 49
use INVX1  INVX1_260
timestamp 1516325494
transform 1 0 3114 0 -1 150
box 0 0 11 49
use DFFNEGX1  DFFNEGX1_5
timestamp 1516325494
transform 1 0 3126 0 -1 150
box 0 0 57 49
use AND2X2  AND2X2_1121
timestamp 1516325494
transform -1 0 3202 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1177
timestamp 1516325494
transform -1 0 3221 0 -1 150
box 0 0 19 49
use NOR2X1  NOR2X1_108
timestamp 1516325494
transform -1 0 3236 0 -1 150
box 0 0 15 49
use NAND2X1  NAND2X1_754
timestamp 1516325494
transform -1 0 3251 0 -1 150
box 0 0 15 49
use INVX1  INVX1_261
timestamp 1516325494
transform 1 0 3251 0 -1 150
box 0 0 11 49
use OR2X2  OR2X2_951
timestamp 1516325494
transform -1 0 3281 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1148
timestamp 1516325494
transform -1 0 3300 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_785
timestamp 1516325494
transform 1 0 3300 0 -1 150
box 0 0 53 49
use MUX2X1  MUX2X1_810
timestamp 1516325494
transform -1 0 3384 0 -1 150
box 0 0 30 49
use AND2X2  AND2X2_1157
timestamp 1516325494
transform 1 0 3384 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_941
timestamp 1516325494
transform 1 0 3403 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_932
timestamp 1516325494
transform 1 0 3422 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1145
timestamp 1516325494
transform -1 0 3460 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1152
timestamp 1516325494
transform 1 0 3460 0 -1 150
box 0 0 19 49
use INVX1  INVX1_254
timestamp 1516325494
transform 1 0 3479 0 -1 150
box 0 0 11 49
use AND2X2  AND2X2_1156
timestamp 1516325494
transform -1 0 3509 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_921
timestamp 1516325494
transform -1 0 3528 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1151
timestamp 1516325494
transform 1 0 3528 0 -1 150
box 0 0 19 49
use OR2X2  OR2X2_938
timestamp 1516325494
transform 1 0 3547 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1153
timestamp 1516325494
transform 1 0 3566 0 -1 150
box 0 0 19 49
use INVX1  INVX1_246
timestamp 1516325494
transform 1 0 3585 0 -1 150
box 0 0 11 49
use INVX1  INVX1_263
timestamp 1516325494
transform 1 0 3597 0 -1 150
box 0 0 11 49
use NOR3X1  NOR3X1_19
timestamp 1516325494
transform -1 0 3627 0 -1 150
box 0 0 19 49
use NOR3X1  NOR3X1_18
timestamp 1516325494
transform -1 0 3646 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1181
timestamp 1516325494
transform -1 0 3665 0 -1 150
box 0 0 19 49
use NOR3X1  NOR3X1_15
timestamp 1516325494
transform 1 0 3665 0 -1 150
box 0 0 19 49
use NOR3X1  NOR3X1_14
timestamp 1516325494
transform -1 0 3703 0 -1 150
box 0 0 19 49
use INVX1  INVX1_252
timestamp 1516325494
transform 1 0 3703 0 -1 150
box 0 0 11 49
use OR2X2  OR2X2_918
timestamp 1516325494
transform 1 0 3715 0 -1 150
box 0 0 19 49
use AND2X2  AND2X2_1130
timestamp 1516325494
transform 1 0 3734 0 -1 150
box 0 0 19 49
use NOR3X1  NOR3X1_23
timestamp 1516325494
transform -1 0 3772 0 -1 150
box 0 0 19 49
use INVX1  INVX1_251
timestamp 1516325494
transform -1 0 3783 0 -1 150
box 0 0 11 49
use INVX1  INVX1_250
timestamp 1516325494
transform 1 0 3783 0 -1 150
box 0 0 11 49
use OR2X2  OR2X2_919
timestamp 1516325494
transform 1 0 3794 0 -1 150
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_779
timestamp 1516325494
transform -1 0 3866 0 -1 150
box 0 0 53 49
use BUFX2  BUFX2_887
timestamp 1516325494
transform 1 0 2 0 1 51
box 0 0 15 49
use FILL  FILL_AND2X2_107
timestamp 1516325494
transform -1 0 25 0 1 51
box 0 0 8 49
use AND2X2  AND2X2_107
timestamp 1516325494
transform -1 0 44 0 1 51
box 0 0 19 49
use FILL  FILL_AND2X2_92
timestamp 1516325494
transform -1 0 52 0 1 51
box 0 0 8 49
use AND2X2  AND2X2_92
timestamp 1516325494
transform -1 0 70 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1331
timestamp 1516325494
transform -1 0 89 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1325
timestamp 1516325494
transform -1 0 108 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1544
timestamp 1516325494
transform -1 0 127 0 1 51
box 0 0 19 49
use FILL  FILL_AND2X2_95
timestamp 1516325494
transform -1 0 135 0 1 51
box 0 0 8 49
use AND2X2  AND2X2_95
timestamp 1516325494
transform -1 0 154 0 1 51
box 0 0 19 49
use FILL  FILL_OR2X2_89
timestamp 1516325494
transform 1 0 154 0 1 51
box 0 0 8 49
use OR2X2  OR2X2_89
timestamp 1516325494
transform 1 0 162 0 1 51
box 0 0 19 49
use FILL  FILL_AND2X2_94
timestamp 1516325494
transform -1 0 189 0 1 51
box 0 0 8 49
use AND2X2  AND2X2_94
timestamp 1516325494
transform -1 0 207 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1450
timestamp 1516325494
transform 1 0 207 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1527
timestamp 1516325494
transform 1 0 226 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1300
timestamp 1516325494
transform 1 0 245 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1525
timestamp 1516325494
transform -1 0 283 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1521
timestamp 1516325494
transform 1 0 283 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1295
timestamp 1516325494
transform -1 0 321 0 1 51
box 0 0 19 49
use FILL  FILL_AND2X2_32
timestamp 1516325494
transform -1 0 329 0 1 51
box 0 0 8 49
use AND2X2  AND2X2_32
timestamp 1516325494
transform -1 0 348 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1429
timestamp 1516325494
transform 1 0 348 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1175
timestamp 1516325494
transform -1 0 386 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1181
timestamp 1516325494
transform 1 0 386 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1637
timestamp 1516325494
transform 1 0 405 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1443
timestamp 1516325494
transform -1 0 443 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1444
timestamp 1516325494
transform -1 0 462 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1294
timestamp 1516325494
transform 1 0 462 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_682
timestamp 1516325494
transform 1 0 481 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_298
timestamp 1516325494
transform 1 0 534 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_298
timestamp 1516325494
transform -1 0 579 0 1 51
box 0 0 30 49
use BUFX2  BUFX2_882
timestamp 1516325494
transform 1 0 2 0 -1 51
box 0 0 15 49
use FILL  FILL_OR2X2_103
timestamp 1516325494
transform -1 0 25 0 -1 51
box 0 0 8 49
use OR2X2  OR2X2_103
timestamp 1516325494
transform -1 0 44 0 -1 51
box 0 0 19 49
use FILL  FILL_AND2X2_110
timestamp 1516325494
transform -1 0 52 0 -1 51
box 0 0 8 49
use AND2X2  AND2X2_110
timestamp 1516325494
transform -1 0 70 0 -1 51
box 0 0 19 49
use FILL  FILL_AND2X2_109
timestamp 1516325494
transform -1 0 78 0 -1 51
box 0 0 8 49
use AND2X2  AND2X2_109
timestamp 1516325494
transform -1 0 97 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1330
timestamp 1516325494
transform -1 0 116 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1550
timestamp 1516325494
transform -1 0 135 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1548
timestamp 1516325494
transform -1 0 154 0 -1 51
box 0 0 19 49
use FILL  FILL_AND2X2_169
timestamp 1516325494
transform -1 0 162 0 -1 51
box 0 0 8 49
use AND2X2  AND2X2_169
timestamp 1516325494
transform -1 0 181 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1640
timestamp 1516325494
transform 1 0 181 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1642
timestamp 1516325494
transform -1 0 219 0 -1 51
box 0 0 19 49
use FILL  FILL_AND2X2_170
timestamp 1516325494
transform 1 0 219 0 -1 51
box 0 0 8 49
use AND2X2  AND2X2_170
timestamp 1516325494
transform 1 0 226 0 -1 51
box 0 0 19 49
use FILL  FILL_OR2X2_159
timestamp 1516325494
transform 1 0 245 0 -1 51
box 0 0 8 49
use OR2X2  OR2X2_159
timestamp 1516325494
transform 1 0 253 0 -1 51
box 0 0 19 49
use FILL  FILL_AND2X2_35
timestamp 1516325494
transform -1 0 280 0 -1 51
box 0 0 8 49
use AND2X2  AND2X2_35
timestamp 1516325494
transform -1 0 298 0 -1 51
box 0 0 19 49
use FILL  FILL_OR2X2_33
timestamp 1516325494
transform 1 0 298 0 -1 51
box 0 0 8 49
use OR2X2  OR2X2_33
timestamp 1516325494
transform 1 0 306 0 -1 51
box 0 0 19 49
use FILL  FILL_AND2X2_34
timestamp 1516325494
transform -1 0 333 0 -1 51
box 0 0 8 49
use AND2X2  AND2X2_34
timestamp 1516325494
transform -1 0 352 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1435
timestamp 1516325494
transform 1 0 352 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1180
timestamp 1516325494
transform 1 0 371 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1433
timestamp 1516325494
transform -1 0 409 0 -1 51
box 0 0 19 49
use BUFX2  BUFX2_874
timestamp 1516325494
transform 1 0 409 0 -1 51
box 0 0 15 49
use AND2X2  AND2X2_1641
timestamp 1516325494
transform -1 0 443 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1448
timestamp 1516325494
transform -1 0 462 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1449
timestamp 1516325494
transform -1 0 481 0 -1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_655
timestamp 1516325494
transform 1 0 481 0 -1 51
box 0 0 53 49
use NAND2X1  NAND2X1_47
timestamp 1516325494
transform 1 0 534 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_47
timestamp 1516325494
transform -1 0 579 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_687
timestamp 1516325494
transform 1 0 580 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_303
timestamp 1516325494
transform 1 0 633 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_303
timestamp 1516325494
transform -1 0 678 0 1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_659
timestamp 1516325494
transform 1 0 678 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_559
timestamp 1516325494
transform 1 0 580 0 -1 51
box 0 0 53 49
use NAND2X1  NAND2X1_463
timestamp 1516325494
transform 1 0 633 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_463
timestamp 1516325494
transform -1 0 678 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_303
timestamp 1516325494
transform 1 0 678 0 -1 51
box 0 0 53 49
use OR2X2  OR2X2_1568
timestamp 1516325494
transform 1 0 732 0 1 51
box 0 0 19 49
use NAND2X1  NAND2X1_51
timestamp 1516325494
transform 1 0 751 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_51
timestamp 1516325494
transform -1 0 796 0 1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_586
timestamp 1516325494
transform 1 0 796 0 1 51
box 0 0 53 49
use MUX2X1  MUX2X1_10
timestamp 1516325494
transform 1 0 849 0 1 51
box 0 0 30 49
use FILL  FILL_BUFX2_69
timestamp 1516325494
transform -1 0 888 0 1 51
box 0 0 8 49
use BUFX2  BUFX2_69
timestamp 1516325494
transform -1 0 902 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_440
timestamp 1516325494
transform 1 0 903 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_307
timestamp 1516325494
transform 1 0 956 0 1 51
box 0 0 53 49
use OR2X2  OR2X2_1291
timestamp 1516325494
transform 1 0 1009 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1520
timestamp 1516325494
transform -1 0 1047 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1635
timestamp 1516325494
transform -1 0 1066 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1442
timestamp 1516325494
transform -1 0 1085 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1441
timestamp 1516325494
transform -1 0 1104 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_431
timestamp 1516325494
transform 1 0 1104 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_399
timestamp 1516325494
transform 1 0 1157 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_399
timestamp 1516325494
transform -1 0 1202 0 1 51
box 0 0 30 49
use MUX2X1  MUX2X1_15
timestamp 1516325494
transform 1 0 1203 0 1 51
box 0 0 30 49
use NAND2X1  NAND2X1_15
timestamp 1516325494
transform -1 0 1248 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_591
timestamp 1516325494
transform -1 0 1301 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_587
timestamp 1516325494
transform 1 0 1302 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_11
timestamp 1516325494
transform 1 0 1355 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_11
timestamp 1516325494
transform -1 0 1400 0 1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_642
timestamp 1516325494
transform 1 0 1400 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_496
timestamp 1516325494
transform -1 0 1469 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_582
timestamp 1516325494
transform -1 0 1522 0 1 51
box 0 0 53 49
use AND2X2  AND2X2_1428
timestamp 1516325494
transform -1 0 1541 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1479
timestamp 1516325494
transform 1 0 1541 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1662
timestamp 1516325494
transform -1 0 1579 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1477
timestamp 1516325494
transform -1 0 1598 0 1 51
box 0 0 19 49
use NAND2X1  NAND2X1_432
timestamp 1516325494
transform 1 0 1598 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_48
timestamp 1516325494
transform 1 0 1613 0 1 51
box 0 0 53 49
use MUX2X1  MUX2X1_432
timestamp 1516325494
transform -1 0 1696 0 1 51
box 0 0 30 49
use OR2X2  OR2X2_1172
timestamp 1516325494
transform -1 0 1716 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_422
timestamp 1516325494
transform 1 0 1716 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_390
timestamp 1516325494
transform 1 0 1769 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_390
timestamp 1516325494
transform -1 0 1814 0 1 51
box 0 0 30 49
use FILL  FILL_BUFX2_249
timestamp 1516325494
transform -1 0 1823 0 1 51
box 0 0 8 49
use BUFX2  BUFX2_249
timestamp 1516325494
transform -1 0 1837 0 1 51
box 0 0 15 49
use OR2X2  OR2X2_1476
timestamp 1516325494
transform -1 0 1856 0 1 51
box 0 0 19 49
use MUX2X1  MUX2X1_839
timestamp 1516325494
transform 1 0 1856 0 1 51
box 0 0 30 49
use NAND2X1  NAND2X1_495
timestamp 1516325494
transform 1 0 732 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_495
timestamp 1516325494
transform -1 0 777 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_299
timestamp 1516325494
transform 1 0 777 0 -1 51
box 0 0 53 49
use MUX2X1  MUX2X1_491
timestamp 1516325494
transform 1 0 830 0 -1 51
box 0 0 30 49
use NAND2X1  NAND2X1_491
timestamp 1516325494
transform -1 0 876 0 -1 51
box 0 0 15 49
use NAND2X1  NAND2X1_10
timestamp 1516325494
transform -1 0 891 0 -1 51
box 0 0 15 49
use OR2X2  OR2X2_1329
timestamp 1516325494
transform 1 0 891 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1549
timestamp 1516325494
transform -1 0 929 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1328
timestamp 1516325494
transform -1 0 948 0 -1 51
box 0 0 19 49
use FILL  FILL_BUFX2_177
timestamp 1516325494
transform 1 0 948 0 -1 51
box 0 0 8 49
use BUFX2  BUFX2_177
timestamp 1516325494
transform 1 0 956 0 -1 51
box 0 0 15 49
use NAND2X1  NAND2X1_43
timestamp 1516325494
transform 1 0 971 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_43
timestamp 1516325494
transform -1 0 1016 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_651
timestamp 1516325494
transform 1 0 1017 0 -1 51
box 0 0 53 49
use FILL  FILL_BUFX2_179
timestamp 1516325494
transform -1 0 1078 0 -1 51
box 0 0 8 49
use BUFX2  BUFX2_179
timestamp 1516325494
transform -1 0 1092 0 -1 51
box 0 0 15 49
use AND2X2  AND2X2_1543
timestamp 1516325494
transform -1 0 1112 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1321
timestamp 1516325494
transform -1 0 1131 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1322
timestamp 1516325494
transform -1 0 1150 0 -1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_427
timestamp 1516325494
transform 1 0 1150 0 -1 51
box 0 0 53 49
use NAND2X1  NAND2X1_395
timestamp 1516325494
transform 1 0 1203 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_395
timestamp 1516325494
transform -1 0 1248 0 -1 51
box 0 0 30 49
use OR2X2  OR2X2_1292
timestamp 1516325494
transform -1 0 1267 0 -1 51
box 0 0 19 49
use FILL  FILL_BUFX2_4
timestamp 1516325494
transform 1 0 1267 0 -1 51
box 0 0 8 49
use BUFX2  BUFX2_4
timestamp 1516325494
transform 1 0 1275 0 -1 51
box 0 0 15 49
use FILL  FILL_BUFX2_232
timestamp 1516325494
transform -1 0 1298 0 -1 51
box 0 0 8 49
use BUFX2  BUFX2_232
timestamp 1516325494
transform -1 0 1313 0 -1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_304
timestamp 1516325494
transform 1 0 1313 0 -1 51
box 0 0 53 49
use MUX2X1  MUX2X1_496
timestamp 1516325494
transform 1 0 1366 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_294
timestamp 1516325494
transform 1 0 1397 0 -1 51
box 0 0 53 49
use MUX2X1  MUX2X1_486
timestamp 1516325494
transform -1 0 1480 0 -1 51
box 0 0 30 49
use NAND2X1  NAND2X1_486
timestamp 1516325494
transform -1 0 1495 0 -1 51
box 0 0 15 49
use OR2X2  OR2X2_1179
timestamp 1516325494
transform 1 0 1495 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1434
timestamp 1516325494
transform -1 0 1533 0 -1 51
box 0 0 19 49
use NAND2X1  NAND2X1_394
timestamp 1516325494
transform 1 0 1533 0 -1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_426
timestamp 1516325494
transform 1 0 1549 0 -1 51
box 0 0 53 49
use MUX2X1  MUX2X1_394
timestamp 1516325494
transform -1 0 1632 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_618
timestamp 1516325494
transform -1 0 1685 0 -1 51
box 0 0 53 49
use AND2X2  AND2X2_1432
timestamp 1516325494
transform -1 0 1704 0 -1 51
box 0 0 19 49
use NAND2X1  NAND2X1_888
timestamp 1516325494
transform 1 0 1704 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_833
timestamp 1516325494
transform -1 0 1750 0 -1 51
box 0 0 30 49
use OR2X2  OR2X2_1178
timestamp 1516325494
transform -1 0 1769 0 -1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_646
timestamp 1516325494
transform 1 0 1769 0 -1 51
box 0 0 53 49
use OR2X2  OR2X2_1177
timestamp 1516325494
transform -1 0 1841 0 -1 51
box 0 0 19 49
use NAND2X1  NAND2X1_38
timestamp 1516325494
transform 1 0 1841 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_38
timestamp 1516325494
transform -1 0 1886 0 -1 51
box 0 0 30 49
use NAND2X1  NAND2X1_894
timestamp 1516325494
transform -1 0 1902 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_624
timestamp 1516325494
transform -1 0 1955 0 1 51
box 0 0 53 49
use OR2X2  OR2X2_1296
timestamp 1516325494
transform 1 0 1955 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1524
timestamp 1516325494
transform -1 0 1993 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_1176
timestamp 1516325494
transform -1 0 2012 0 1 51
box 0 0 19 49
use NAND2X1  NAND2X1_884
timestamp 1516325494
transform 1 0 2012 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_614
timestamp 1516325494
transform 1 0 2027 0 1 51
box 0 0 53 49
use MUX2X1  MUX2X1_829
timestamp 1516325494
transform -1 0 2111 0 1 51
box 0 0 30 49
use OR2X2  OR2X2_1297
timestamp 1516325494
transform -1 0 2130 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_555
timestamp 1516325494
transform 1 0 2130 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_42
timestamp 1516325494
transform 1 0 2183 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_426
timestamp 1516325494
transform 1 0 2236 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_38
timestamp 1516325494
transform 1 0 1887 0 -1 51
box 0 0 53 49
use NAND2X1  NAND2X1_422
timestamp 1516325494
transform 1 0 1940 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_422
timestamp 1516325494
transform -1 0 1985 0 -1 51
box 0 0 30 49
use MUX2X1  MUX2X1_42
timestamp 1516325494
transform 1 0 1986 0 -1 51
box 0 0 30 49
use NAND2X1  NAND2X1_42
timestamp 1516325494
transform -1 0 2031 0 -1 51
box 0 0 15 49
use AND2X2  AND2X2_1639
timestamp 1516325494
transform -1 0 2050 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1447
timestamp 1516325494
transform -1 0 2069 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1547
timestamp 1516325494
transform -1 0 2088 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1327
timestamp 1516325494
transform -1 0 2107 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1446
timestamp 1516325494
transform -1 0 2126 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_1326
timestamp 1516325494
transform -1 0 2145 0 -1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_47
timestamp 1516325494
transform 1 0 2145 0 -1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_623
timestamp 1516325494
transform 1 0 2198 0 -1 51
box 0 0 53 49
use MUX2X1  MUX2X1_426
timestamp 1516325494
transform -1 0 2282 0 1 51
box 0 0 30 49
use MUX2X1  MUX2X1_838
timestamp 1516325494
transform -1 0 2312 0 1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_625
timestamp 1516325494
transform 1 0 2312 0 1 51
box 0 0 53 49
use NAND2X1  NAND2X1_431
timestamp 1516325494
transform 1 0 2252 0 -1 51
box 0 0 15 49
use NAND2X1  NAND2X1_893
timestamp 1516325494
transform 1 0 2267 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_431
timestamp 1516325494
transform -1 0 2312 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_175
timestamp 1516325494
transform 1 0 2312 0 -1 51
box 0 0 53 49
use NAND2X1  NAND2X1_895
timestamp 1516325494
transform 1 0 2366 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_840
timestamp 1516325494
transform -1 0 2411 0 1 51
box 0 0 30 49
use OR2X2  OR2X2_1298
timestamp 1516325494
transform 1 0 2411 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1526
timestamp 1516325494
transform -1 0 2449 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_650
timestamp 1516325494
transform -1 0 2502 0 1 51
box 0 0 53 49
use OR2X2  OR2X2_1299
timestamp 1516325494
transform -1 0 2521 0 1 51
box 0 0 19 49
use FILL  FILL_BUFX2_68
timestamp 1516325494
transform -1 0 2529 0 1 51
box 0 0 8 49
use BUFX2  BUFX2_68
timestamp 1516325494
transform -1 0 2544 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_637
timestamp 1516325494
transform -1 0 2597 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_619
timestamp 1516325494
transform 1 0 2597 0 1 51
box 0 0 53 49
use FILL  FILL_BUFX2_252
timestamp 1516325494
transform -1 0 2659 0 1 51
box 0 0 8 49
use BUFX2  BUFX2_252
timestamp 1516325494
transform -1 0 2673 0 1 51
box 0 0 15 49
use FILL  FILL_BUFX2_246
timestamp 1516325494
transform -1 0 2681 0 1 51
box 0 0 8 49
use BUFX2  BUFX2_246
timestamp 1516325494
transform -1 0 2696 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_43
timestamp 1516325494
transform 1 0 2696 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_280
timestamp 1516325494
transform 1 0 2749 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_715
timestamp 1516325494
transform 1 0 2803 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_239
timestamp 1516325494
transform -1 0 2909 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_783
timestamp 1516325494
transform 1 0 2909 0 1 51
box 0 0 53 49
use XOR2X1  XOR2X1_68
timestamp 1516325494
transform 1 0 2962 0 1 51
box 0 0 34 49
use AOI21X1  AOI21X1_40
timestamp 1516325494
transform 1 0 2996 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1150
timestamp 1516325494
transform 1 0 3015 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_754
timestamp 1516325494
transform -1 0 3087 0 1 51
box 0 0 53 49
use INVX1  INVX1_232
timestamp 1516325494
transform 1 0 3088 0 1 51
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_775
timestamp 1516325494
transform 1 0 3099 0 1 51
box 0 0 53 49
use NOR2X1  NOR2X1_129
timestamp 1516325494
transform -1 0 3167 0 1 51
box 0 0 15 49
use AND2X2  AND2X2_1158
timestamp 1516325494
transform -1 0 3186 0 1 51
box 0 0 19 49
use FILL  FILL_BUFX2_224
timestamp 1516325494
transform 1 0 3186 0 1 51
box 0 0 8 49
use BUFX2  BUFX2_224
timestamp 1516325494
transform 1 0 3194 0 1 51
box 0 0 15 49
use NOR2X1  NOR2X1_127
timestamp 1516325494
transform 1 0 3209 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_773
timestamp 1516325494
transform -1 0 3277 0 1 51
box 0 0 53 49
use OR2X2  OR2X2_936
timestamp 1516325494
transform -1 0 3297 0 1 51
box 0 0 19 49
use NOR2X1  NOR2X1_161
timestamp 1516325494
transform -1 0 3312 0 1 51
box 0 0 15 49
use MUX2X1  MUX2X1_812
timestamp 1516325494
transform -1 0 3342 0 1 51
box 0 0 30 49
use NOR2X1  NOR2X1_167
timestamp 1516325494
transform -1 0 3357 0 1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_710
timestamp 1516325494
transform -1 0 3410 0 1 51
box 0 0 53 49
use OR2X2  OR2X2_942
timestamp 1516325494
transform -1 0 3430 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1146
timestamp 1516325494
transform -1 0 3449 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_931
timestamp 1516325494
transform -1 0 3468 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_940
timestamp 1516325494
transform -1 0 3487 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_939
timestamp 1516325494
transform -1 0 3506 0 1 51
box 0 0 19 49
use NOR2X1  NOR2X1_126
timestamp 1516325494
transform 1 0 3506 0 1 51
box 0 0 15 49
use NOR2X1  NOR2X1_131
timestamp 1516325494
transform 1 0 3521 0 1 51
box 0 0 15 49
use OR2X2  OR2X2_953
timestamp 1516325494
transform 1 0 3536 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_751
timestamp 1516325494
transform -1 0 3608 0 1 51
box 0 0 53 49
use NOR2X1  NOR2X1_119
timestamp 1516325494
transform 1 0 3608 0 1 51
box 0 0 15 49
use OR2X2  OR2X2_922
timestamp 1516325494
transform 1 0 3623 0 1 51
box 0 0 19 49
use AND2X2  AND2X2_1131
timestamp 1516325494
transform 1 0 3642 0 1 51
box 0 0 19 49
use OR2X2  OR2X2_923
timestamp 1516325494
transform 1 0 3661 0 1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_781
timestamp 1516325494
transform -1 0 3733 0 1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_153
timestamp 1516325494
transform 1 0 3734 0 1 51
box 0 0 53 49
use BUFX2  BUFX2_907
timestamp 1516325494
transform -1 0 3802 0 1 51
box 0 0 15 49
use BUFX2  BUFX2_878
timestamp 1516325494
transform -1 0 3817 0 1 51
box 0 0 15 49
use INVX1  INVX1_309
timestamp 1516325494
transform 1 0 3817 0 1 51
box 0 0 11 49
use BUFX2  BUFX2_908
timestamp 1516325494
transform -1 0 3844 0 1 51
box 0 0 15 49
use NAND2X1  NAND2X1_262
timestamp 1516325494
transform -1 0 3859 0 1 51
box 0 0 15 49
use FILL  FILL_2_1
timestamp 1516325494
transform 1 0 3859 0 1 51
box 0 0 8 49
use MUX2X1  MUX2X1_239
timestamp 1516325494
transform 1 0 2366 0 -1 51
box 0 0 30 49
use NAND2X1  NAND2X1_239
timestamp 1516325494
transform -1 0 2411 0 -1 51
box 0 0 15 49
use DFFNEGX1  DFFNEGX1_3
timestamp 1516325494
transform 1 0 2411 0 -1 51
box 0 0 57 49
use DFFNEGX1  DFFNEGX1_2
timestamp 1516325494
transform 1 0 2468 0 -1 51
box 0 0 57 49
use AND2X2  AND2X2_1118
timestamp 1516325494
transform -1 0 2544 0 -1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_782
timestamp 1516325494
transform 1 0 2544 0 -1 51
box 0 0 53 49
use AND2X2  AND2X2_1119
timestamp 1516325494
transform -1 0 2616 0 -1 51
box 0 0 19 49
use DFFNEGX1  DFFNEGX1_4
timestamp 1516325494
transform 1 0 2616 0 -1 51
box 0 0 57 49
use AND2X2  AND2X2_1120
timestamp 1516325494
transform -1 0 2692 0 -1 51
box 0 0 19 49
use DFFPOSX1  DFFPOSX1_784
timestamp 1516325494
transform 1 0 2692 0 -1 51
box 0 0 53 49
use INVX1  INVX1_259
timestamp 1516325494
transform -1 0 2757 0 -1 51
box 0 0 11 49
use NOR3X1  NOR3X1_28
timestamp 1516325494
transform -1 0 2776 0 -1 51
box 0 0 19 49
use NOR2X1  NOR2X1_107
timestamp 1516325494
transform -1 0 2791 0 -1 51
box 0 0 15 49
use NOR2X1  NOR2X1_109
timestamp 1516325494
transform -1 0 2806 0 -1 51
box 0 0 15 49
use INVX1  INVX1_258
timestamp 1516325494
transform 1 0 2806 0 -1 51
box 0 0 11 49
use OR2X2  OR2X2_937
timestamp 1516325494
transform -1 0 2837 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_934
timestamp 1516325494
transform -1 0 2856 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1149
timestamp 1516325494
transform 1 0 2856 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_1147
timestamp 1516325494
transform -1 0 2894 0 -1 51
box 0 0 19 49
use NAND2X1  NAND2X1_764
timestamp 1516325494
transform -1 0 2909 0 -1 51
box 0 0 15 49
use NAND2X1  NAND2X1_763
timestamp 1516325494
transform -1 0 2924 0 -1 51
box 0 0 15 49
use OR2X2  OR2X2_933
timestamp 1516325494
transform -1 0 2943 0 -1 51
box 0 0 19 49
use NOR3X1  NOR3X1_26
timestamp 1516325494
transform -1 0 2962 0 -1 51
box 0 0 19 49
use INVX1  INVX1_234
timestamp 1516325494
transform -1 0 2973 0 -1 51
box 0 0 11 49
use NOR3X1  NOR3X1_27
timestamp 1516325494
transform -1 0 2993 0 -1 51
box 0 0 19 49
use NAND2X1  NAND2X1_765
timestamp 1516325494
transform 1 0 2993 0 -1 51
box 0 0 15 49
use INVX1  INVX1_233
timestamp 1516325494
transform -1 0 3019 0 -1 51
box 0 0 11 49
use NAND3X1  NAND3X1_80
timestamp 1516325494
transform 1 0 3019 0 -1 51
box 0 0 19 49
use INVX1  INVX1_307
timestamp 1516325494
transform 1 0 3038 0 -1 51
box 0 0 11 49
use NOR2X1  NOR2X1_162
timestamp 1516325494
transform -1 0 3065 0 -1 51
box 0 0 15 49
use INVX1  INVX1_308
timestamp 1516325494
transform -1 0 3076 0 -1 51
box 0 0 11 49
use NOR2X1  NOR2X1_165
timestamp 1516325494
transform 1 0 3076 0 -1 51
box 0 0 15 49
use INVX1  INVX1_311
timestamp 1516325494
transform -1 0 3102 0 -1 51
box 0 0 11 49
use BUFX2  BUFX2_872
timestamp 1516325494
transform -1 0 3118 0 -1 51
box 0 0 15 49
use INVX1  INVX1_313
timestamp 1516325494
transform 1 0 3118 0 -1 51
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_822
timestamp 1516325494
transform -1 0 3182 0 -1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_798
timestamp 1516325494
transform 1 0 3183 0 -1 51
box 0 0 53 49
use AND2X2  AND2X2_1187
timestamp 1516325494
transform 1 0 3236 0 -1 51
box 0 0 19 49
use BUFX2  BUFX2_905
timestamp 1516325494
transform -1 0 3270 0 -1 51
box 0 0 15 49
use BUFX2  BUFX2_877
timestamp 1516325494
transform -1 0 3285 0 -1 51
box 0 0 15 49
use FILL  FILL_BUFX2_201
timestamp 1516325494
transform 1 0 3285 0 -1 51
box 0 0 8 49
use BUFX2  BUFX2_201
timestamp 1516325494
transform 1 0 3293 0 -1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_795
timestamp 1516325494
transform 1 0 3308 0 -1 51
box 0 0 53 49
use INVX1  INVX1_306
timestamp 1516325494
transform -1 0 3372 0 -1 51
box 0 0 11 49
use NAND2X1  NAND2X1_258
timestamp 1516325494
transform 1 0 3373 0 -1 51
box 0 0 15 49
use NOR2X1  NOR2X1_163
timestamp 1516325494
transform -1 0 3403 0 -1 51
box 0 0 15 49
use INVX1  INVX1_305
timestamp 1516325494
transform -1 0 3414 0 -1 51
box 0 0 11 49
use DFFPOSX1  DFFPOSX1_334
timestamp 1516325494
transform -1 0 3467 0 -1 51
box 0 0 53 49
use DFFPOSX1  DFFPOSX1_322
timestamp 1516325494
transform -1 0 3521 0 -1 51
box 0 0 53 49
use BUFX2  BUFX2_915
timestamp 1516325494
transform -1 0 3536 0 -1 51
box 0 0 15 49
use FILL  FILL_BUFX2_191
timestamp 1516325494
transform -1 0 3544 0 -1 51
box 0 0 8 49
use BUFX2  BUFX2_191
timestamp 1516325494
transform -1 0 3559 0 -1 51
box 0 0 15 49
use DFFPOSX1  DFFPOSX1_130
timestamp 1516325494
transform 1 0 3559 0 -1 51
box 0 0 53 49
use MUX2X1  MUX2X1_258
timestamp 1516325494
transform -1 0 3642 0 -1 51
box 0 0 30 49
use DFFPOSX1  DFFPOSX1_134
timestamp 1516325494
transform -1 0 3695 0 -1 51
box 0 0 53 49
use AND2X2  AND2X2_314
timestamp 1516325494
transform 1 0 3696 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_296
timestamp 1516325494
transform -1 0 3734 0 -1 51
box 0 0 19 49
use OR2X2  OR2X2_295
timestamp 1516325494
transform -1 0 3753 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_316
timestamp 1516325494
transform -1 0 3772 0 -1 51
box 0 0 19 49
use AND2X2  AND2X2_315
timestamp 1516325494
transform 1 0 3772 0 -1 51
box 0 0 19 49
use MUX2X1  MUX2X1_377
timestamp 1516325494
transform 1 0 3791 0 -1 51
box 0 0 30 49
use NAND2X1  NAND2X1_377
timestamp 1516325494
transform 1 0 3821 0 -1 51
box 0 0 15 49
use MUX2X1  MUX2X1_281
timestamp 1516325494
transform 1 0 3836 0 -1 51
box 0 0 30 49
<< labels >>
flabel space 3914 1227 3914 1227 3 FreeSans 48 0 0 0 IDATA_CORE_out<0>
port 0 nsew
flabel space 3914 509 3914 509 3 FreeSans 48 0 0 0 IDATA_CORE_out<1>
port 1 nsew
flabel space 3914 768 3914 768 3 FreeSans 48 0 0 0 IDATA_CORE_out<2>
port 2 nsew
flabel space 3914 42 3914 42 3 FreeSans 48 270 0 0 IDATA_CORE_out<3>
port 3 nsew
flabel space 3044 -38 3044 -38 7 FreeSans 48 270 0 0 IDATA_CORE_out<4>
port 4 nsew
flabel space 3097 -38 3097 -38 7 FreeSans 48 270 0 0 IDATA_CORE_out<5>
port 5 nsew
flabel space 3914 95 3914 95 3 FreeSans 48 0 0 0 IDATA_CORE_out<6>
port 6 nsew
flabel space 3914 1068 3914 1068 3 FreeSans 48 0 0 0 IDATA_CORE_out<7>
port 7 nsew
flabel space 3146 -38 3146 -38 7 FreeSans 48 270 0 0 IDATA_CORE_out<8>
port 8 nsew
flabel space 3914 2546 3914 2546 3 FreeSans 48 0 0 0 IDATA_CORE_out<9>
port 9 nsew
flabel space 3249 -38 3249 -38 7 FreeSans 48 270 0 0 IDATA_CORE_out<10>
port 10 nsew
flabel space 3914 1642 3914 1642 3 FreeSans 48 0 0 0 IDATA_CORE_out<11>
port 11 nsew
flabel space 3914 1455 3914 1455 3 FreeSans 48 0 0 0 IDATA_CORE_out<12>
port 12 nsew
flabel space 3914 559 3914 559 3 FreeSans 48 0 0 0 IDATA_CORE_out<13>
port 13 nsew
flabel space 3914 2117 3914 2117 3 FreeSans 48 0 0 0 IDATA_CORE_out<14>
port 14 nsew
flabel space 3914 2630 3914 2630 3 FreeSans 48 90 0 0 IDATA_CORE_out<15>
port 15 nsew
flabel space 3914 456 3914 456 3 FreeSans 48 0 0 0 IDATA_CORE_out<16>
port 16 nsew
flabel space 3914 1288 3914 1288 3 FreeSans 48 0 0 0 IDATA_CORE_out<17>
port 17 nsew
flabel space -38 1129 -38 1129 7 FreeSans 48 0 0 0 IDATA_CORE_out<18>
port 18 nsew
flabel space -38 95 -38 95 7 FreeSans 48 0 0 0 IDATA_CORE_out<19>
port 19 nsew
flabel space 1106 2709 1106 2709 3 FreeSans 48 90 0 0 IDATA_CORE_out<20>
port 20 nsew
flabel space 885 -38 885 -38 7 FreeSans 48 270 0 0 IDATA_CORE_out<21>
port 21 nsew
flabel space 1224 2709 1224 2709 3 FreeSans 48 90 0 0 IDATA_CORE_out<22>
port 22 nsew
flabel space 2930 2709 2930 2709 3 FreeSans 48 90 0 0 IDATA_CORE_out<23>
port 23 nsew
flabel space 1668 2709 1668 2709 3 FreeSans 48 90 0 0 IDATA_CORE_out<24>
port 24 nsew
flabel space 3914 2402 3914 2402 3 FreeSans 48 0 0 0 IDATA_CORE_out<25>
port 25 nsew
flabel space 217 -38 217 -38 7 FreeSans 48 270 0 0 IDATA_CORE_out<26>
port 26 nsew
flabel space 323 2709 323 2709 3 FreeSans 48 90 0 0 IDATA_CORE_out<27>
port 27 nsew
flabel space -38 2709 -38 2709 7 FreeSans 48 90 0 0 IDATA_CORE_out<28>
port 28 nsew
flabel space 3914 1163 3914 1163 3 FreeSans 48 0 0 0 IDATA_CORE_out<29>
port 29 nsew
flabel space 3652 2709 3652 2709 3 FreeSans 48 90 0 0 IDATA_CORE_out<30>
port 30 nsew
flabel space -38 148 -38 148 7 FreeSans 48 0 0 0 IDATA_CORE_out<31>
port 31 nsew
flabel space 1718 2709 1718 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<0>
port 32 nsew
flabel space 2310 2709 2310 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<1>
port 33 nsew
flabel space 2823 2709 2823 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<2>
port 34 nsew
flabel space 2721 2709 2721 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<3>
port 35 nsew
flabel space 2516 2709 2516 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<4>
port 36 nsew
flabel space 2671 2709 2671 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<5>
port 37 nsew
flabel space 2413 2709 2413 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<6>
port 38 nsew
flabel space 2360 2709 2360 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<7>
port 39 nsew
flabel space 1976 2709 1976 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<8>
port 40 nsew
flabel space 1505 -38 1505 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<9>
port 41 nsew
flabel space 1402 -38 1402 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<10>
port 42 nsew
flabel space 1566 -38 1566 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<11>
port 43 nsew
flabel space 2774 2709 2774 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<12>
port 44 nsew
flabel space 1425 2709 1425 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<13>
port 45 nsew
flabel space 935 -38 935 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<14>
port 46 nsew
flabel space 832 -38 832 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<15>
port 47 nsew
flabel space 988 -38 988 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<16>
port 48 nsew
flabel space 2569 2709 2569 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<17>
port 49 nsew
flabel space 1512 2709 1512 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<18>
port 50 nsew
flabel space 1873 2709 1873 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<19>
port 51 nsew
flabel space 1360 2709 1360 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<20>
port 52 nsew
flabel space 1927 2709 1927 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<21>
port 53 nsew
flabel space 2618 2709 2618 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<22>
port 54 nsew
flabel space 1455 -38 1455 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<23>
port 55 nsew
flabel space 1619 -38 1619 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<24>
port 56 nsew
flabel space 1771 2709 1771 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<25>
port 57 nsew
flabel space 2257 2709 2257 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<26>
port 58 nsew
flabel space 1820 2709 1820 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<27>
port 59 nsew
flabel space 1037 -38 1037 -38 7 FreeSans 48 270 0 0 DDATA_CORE_out<28>
port 60 nsew
flabel space 2204 2709 2204 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<29>
port 61 nsew
flabel space 2462 2709 2462 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<30>
port 62 nsew
flabel space 2155 2709 2155 2709 3 FreeSans 48 90 0 0 DDATA_CORE_out<31>
port 63 nsew
flabel space -38 1068 -38 1068 7 FreeSans 48 0 0 0 CORE_ctrl<0>
port 64 nsew
flabel space 3291 2709 3291 2709 3 FreeSans 48 90 0 0 CORE_ctrl<1>
port 65 nsew
flabel space 1300 -38 1300 -38 7 FreeSans 48 270 0 0 CORE_ctrl<2>
port 66 nsew
flabel space 3914 2037 3914 2037 3 FreeSans 48 0 0 0 INTERRUPT_ch<0>
port 67 nsew
flabel space 3238 2709 3238 2709 3 FreeSans 48 90 0 0 INTERRUPT_ch<1>
port 68 nsew
flabel space 3914 2166 3914 2166 3 FreeSans 48 0 0 0 INTERRUPT_ch<2>
port 69 nsew
flabel space 3857 2709 3857 2709 3 FreeSans 48 90 0 0 INTERRUPT_ch<3>
port 70 nsew
flabel space 3032 2709 3032 2709 3 FreeSans 48 90 0 0 INTERRUPT_ch<4>
port 71 nsew
flabel space 3914 2352 3914 2352 3 FreeSans 48 0 0 0 INTERRUPT_ch<5>
port 72 nsew
flabel space 3184 2709 3184 2709 3 FreeSans 48 90 0 0 INTERRUPT_ch<6>
port 73 nsew
flabel space 3135 2709 3135 2709 3 FreeSans 48 90 0 0 INTERRUPT_ch<7>
port 74 nsew
flabel space 1615 2709 1615 2709 3 FreeSans 48 90 0 0 INTERRUPT_flag
port 75 nsew
flabel space 1353 -38 1353 -38 7 FreeSans 48 270 0 0 clk
port 76 nsew
flabel space 3914 1015 3914 1015 3 FreeSans 48 0 0 0 rst
port 77 nsew
flabel space 3914 198 3914 198 3 FreeSans 48 0 0 0 IDATA_CORE_addr<0>
port 78 nsew
flabel space 3914 251 3914 251 3 FreeSans 48 0 0 0 IDATA_CORE_addr<1>
port 79 nsew
flabel space 3914 1406 3914 1406 3 FreeSans 48 0 0 0 IDATA_CORE_addr<2>
port 80 nsew
flabel space 3599 2709 3599 2709 3 FreeSans 48 90 0 0 IDATA_CORE_addr<3>
port 81 nsew
flabel space 3340 2709 3340 2709 3 FreeSans 48 90 0 0 IDATA_CORE_addr<4>
port 82 nsew
flabel space 3914 1695 3914 1695 3 FreeSans 48 0 0 0 IDATA_CORE_addr<5>
port 83 nsew
flabel space 3082 2709 3082 2709 3 FreeSans 48 90 0 0 IDATA_CORE_addr<6>
port 84 nsew
flabel space 2979 2709 2979 2709 3 FreeSans 48 90 0 0 IDATA_CORE_addr<7>
port 85 nsew
flabel space 3914 612 3914 612 3 FreeSans 48 0 0 0 IDATA_CORE_clk
port 86 nsew
flabel space 3443 2709 3443 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<0>
port 87 nsew
flabel space 3701 2709 3701 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<1>
port 88 nsew
flabel space 3804 2709 3804 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<2>
port 89 nsew
flabel space 3496 2709 3496 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<3>
port 90 nsew
flabel space 3754 2709 3754 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<4>
port 91 nsew
flabel space 3393 2709 3393 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<5>
port 92 nsew
flabel space 3549 2709 3549 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<6>
port 93 nsew
flabel space 3910 2709 3910 2709 3 FreeSans 48 90 0 0 DDATA_CORE_addr<7>
port 94 nsew
flabel space 1167 -38 1167 -38 7 FreeSans 48 270 0 0 DDATA_CORE_in<0>
port 95 nsew
flabel space 410 -38 410 -38 7 FreeSans 48 270 0 0 DDATA_CORE_in<1>
port 96 nsew
flabel space 3914 1562 3914 1562 3 FreeSans 48 0 0 0 DDATA_CORE_in<2>
port 97 nsew
flabel space 3914 2299 3914 2299 3 FreeSans 48 0 0 0 DDATA_CORE_in<3>
port 98 nsew
flabel space 3914 300 3914 300 3 FreeSans 48 0 0 0 DDATA_CORE_in<4>
port 99 nsew
flabel space 3914 148 3914 148 3 FreeSans 48 0 0 0 DDATA_CORE_in<5>
port 100 nsew
flabel space 2877 2709 2877 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<6>
port 101 nsew
flabel space 950 2709 950 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<7>
port 102 nsew
flabel space -38 1562 -38 1562 7 FreeSans 48 0 0 0 DDATA_CORE_in<8>
port 103 nsew
flabel space -38 42 -38 42 7 FreeSans 48 270 0 0 DDATA_CORE_in<9>
port 104 nsew
flabel space 1566 2709 1566 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<10>
port 105 nsew
flabel space 1003 2709 1003 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<11>
port 106 nsew
flabel space -38 2649 -38 2649 7 FreeSans 48 90 0 0 DDATA_CORE_in<12>
port 107 nsew
flabel space -38 1858 -38 1858 7 FreeSans 48 0 0 0 DDATA_CORE_in<13>
port 108 nsew
flabel space -38 198 -38 198 7 FreeSans 48 0 0 0 DDATA_CORE_in<14>
port 109 nsew
flabel space 277 -38 277 -38 7 FreeSans 48 270 0 0 DDATA_CORE_in<15>
port 110 nsew
flabel space 901 2709 901 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<16>
port 111 nsew
flabel space 642 2709 642 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<17>
port 112 nsew
flabel space 486 2709 486 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<18>
port 113 nsew
flabel space 1170 2709 1170 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<19>
port 114 nsew
flabel space 1056 2709 1056 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<20>
port 115 nsew
flabel space 798 2709 798 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<21>
port 116 nsew
flabel space 540 2709 540 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<22>
port 117 nsew
flabel space -38 2253 -38 2253 7 FreeSans 48 0 0 0 DDATA_CORE_in<23>
port 118 nsew
flabel space 692 2709 692 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<24>
port 119 nsew
flabel space 84 2709 84 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<25>
port 120 nsew
flabel space 426 2709 426 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<26>
port 121 nsew
flabel space 255 2709 255 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<27>
port 122 nsew
flabel space 745 2709 745 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<28>
port 123 nsew
flabel space 372 2709 372 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<29>
port 124 nsew
flabel space 847 2709 847 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<30>
port 125 nsew
flabel space 589 2709 589 2709 3 FreeSans 48 90 0 0 DDATA_CORE_in<31>
port 126 nsew
flabel space 3914 353 3914 353 3 FreeSans 48 0 0 0 DDATA_CORE_load
port 127 nsew
flabel space 3914 2683 3914 2683 3 FreeSans 48 90 0 0 DDATA_CORE_write
port 128 nsew
flabel space 3865 -38 3865 -38 3 FreeSans 48 270 0 0 DDATA_CORE_ctrl<0>
port 129 nsew
flabel space 3914 407 3914 407 3 FreeSans 48 0 0 0 DDATA_CORE_ctrl<1>
port 130 nsew
flabel space 3200 -38 3200 -38 7 FreeSans 48 270 0 0 DDATA_CORE_ctrl<2>
port 131 nsew
<< end >>
