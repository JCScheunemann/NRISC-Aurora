magic
tech scmos
magscale 1 4
timestamp 1513729314
<< metal1 >>
rect 93 2297 104 2303
rect 445 2297 456 2303
rect 141 2277 195 2283
rect 445 2283 451 2297
rect 509 2297 531 2303
rect 509 2283 515 2297
rect 653 2303 659 2323
rect 621 2297 659 2303
rect 877 2303 883 2323
rect 1816 2317 1832 2323
rect 845 2297 883 2303
rect 1357 2297 1384 2303
rect 1725 2297 1736 2303
rect 2008 2297 2019 2303
rect 2349 2297 2360 2303
rect 2600 2297 2611 2303
rect 2941 2303 2947 2323
rect 2792 2297 2803 2303
rect 2909 2297 2947 2303
rect 3117 2297 3128 2303
rect 429 2277 451 2283
rect 493 2277 515 2283
rect 776 2277 819 2283
rect 1565 2277 1576 2283
rect 1896 2277 1907 2283
rect 2269 2277 2296 2283
rect 3080 2277 3091 2283
rect 696 2157 707 2163
rect 2717 2157 2739 2163
rect 2877 2148 2883 2163
rect 152 2137 163 2143
rect 157 2123 163 2137
rect 232 2137 259 2143
rect 333 2137 360 2143
rect 376 2137 387 2143
rect 461 2137 488 2143
rect 669 2137 680 2143
rect 749 2137 819 2143
rect 973 2137 1000 2143
rect 1021 2137 1059 2143
rect 157 2117 179 2123
rect 540 2117 568 2123
rect 540 2116 548 2117
rect 824 2117 835 2123
rect 845 2117 884 2123
rect 876 2112 884 2117
rect 1261 2117 1272 2123
rect 1320 2117 1347 2123
rect 1373 2117 1384 2123
rect 1373 2097 1379 2117
rect 1565 2117 1576 2123
rect 1624 2117 1667 2123
rect 1741 2117 1859 2123
rect 2013 2117 2051 2123
rect 1704 2097 1715 2103
rect 2045 2097 2051 2117
rect 2173 2123 2179 2143
rect 2797 2137 2840 2143
rect 2888 2137 2899 2143
rect 3021 2143 3027 2152
rect 3021 2137 3043 2143
rect 3405 2137 3427 2143
rect 3469 2137 3491 2143
rect 2157 2117 2179 2123
rect 2301 2117 2328 2123
rect 2765 2117 2776 2123
rect 2824 2117 2867 2123
rect 2909 2117 2947 2123
rect 2941 2097 2947 2117
rect 3053 2117 3091 2123
rect 3085 2097 3091 2117
rect 3208 2117 3219 2123
rect 3421 2123 3427 2137
rect 3421 2117 3432 2123
rect 3485 2123 3491 2137
rect 3485 2117 3507 2123
rect 888 2077 915 2083
rect 1901 2077 1912 2083
rect 717 1937 728 1943
rect 1133 1917 1144 1923
rect 1832 1917 1859 1923
rect 2840 1917 2883 1923
rect 61 1897 72 1903
rect 253 1897 275 1903
rect 109 1877 136 1883
rect 269 1883 275 1897
rect 557 1897 579 1903
rect 941 1897 995 1903
rect 1005 1897 1016 1903
rect 1368 1897 1395 1903
rect 2413 1897 2435 1903
rect 2653 1897 2664 1903
rect 2749 1897 2787 1903
rect 2957 1903 2963 1923
rect 2925 1897 2963 1903
rect 2989 1897 3000 1903
rect 3069 1903 3075 1923
rect 3256 1916 3260 1924
rect 3277 1917 3288 1923
rect 3037 1897 3075 1903
rect 3208 1897 3251 1903
rect 3325 1897 3336 1903
rect 152 1877 163 1883
rect 269 1877 291 1883
rect 413 1877 451 1883
rect 1256 1877 1299 1883
rect 1597 1877 1635 1883
rect 1885 1877 1907 1883
rect 2360 1877 2371 1883
rect 2397 1877 2424 1883
rect 2461 1877 2499 1883
rect 2589 1877 2616 1883
rect 3389 1883 3395 1923
rect 3533 1897 3544 1903
rect 3597 1903 3603 1923
rect 3565 1897 3603 1903
rect 3389 1877 3427 1883
rect 1224 1857 1235 1863
rect 1805 1857 1832 1863
rect 2664 1857 2684 1863
rect 141 1737 163 1743
rect 157 1723 163 1737
rect 349 1737 360 1743
rect 589 1737 616 1743
rect 989 1743 995 1763
rect 1032 1757 1052 1763
rect 2749 1757 2771 1763
rect 957 1737 995 1743
rect 1453 1737 1491 1743
rect 1832 1737 1859 1743
rect 157 1717 179 1723
rect 269 1717 280 1723
rect 1021 1717 1032 1723
rect 1144 1717 1155 1723
rect 1245 1717 1272 1723
rect 1517 1717 1555 1723
rect 260 1696 264 1704
rect 324 1696 328 1704
rect 1517 1697 1523 1717
rect 1773 1717 1832 1723
rect 1928 1717 1971 1723
rect 2189 1723 2195 1743
rect 2557 1737 2568 1743
rect 2589 1737 2616 1743
rect 2701 1737 2712 1743
rect 3421 1737 3432 1743
rect 2125 1717 2195 1723
rect 2285 1717 2296 1723
rect 2632 1717 2643 1723
rect 2813 1717 2840 1723
rect 2968 1717 2979 1723
rect 3261 1717 3272 1723
rect 3432 1717 3459 1723
rect 3597 1717 3624 1723
rect 1837 1697 1843 1712
rect 285 1537 312 1543
rect 796 1537 824 1543
rect 796 1532 804 1537
rect 1053 1517 1064 1523
rect 140 1497 152 1503
rect 140 1492 148 1497
rect 237 1497 248 1503
rect 1208 1497 1219 1503
rect 1384 1497 1395 1503
rect 1592 1497 1619 1503
rect 1736 1497 1763 1503
rect 1800 1497 1859 1503
rect 1896 1497 1907 1503
rect 2077 1503 2083 1523
rect 2077 1497 2115 1503
rect 2253 1497 2275 1503
rect 2509 1503 2515 1523
rect 2477 1497 2515 1503
rect 2541 1497 2595 1503
rect 3069 1497 3123 1503
rect 173 1477 211 1483
rect 749 1477 760 1483
rect 749 1457 755 1477
rect 989 1477 1027 1483
rect 1357 1477 1368 1483
rect 1501 1477 1528 1483
rect 2733 1477 2776 1483
rect 2813 1457 2824 1463
rect 2877 1457 2915 1463
rect 3565 1457 3587 1463
rect 824 1437 851 1443
rect 1053 1437 1080 1443
rect 2621 1357 2643 1363
rect 157 1337 195 1343
rect 269 1337 307 1343
rect 360 1337 371 1343
rect 1213 1337 1224 1343
rect 1832 1337 1843 1343
rect 1944 1337 1971 1343
rect 1981 1337 2019 1343
rect 2056 1337 2083 1343
rect 2093 1337 2120 1343
rect 2173 1337 2184 1343
rect 2856 1337 2867 1343
rect 3016 1337 3027 1343
rect 3197 1337 3235 1343
rect 3336 1337 3347 1343
rect 301 1317 323 1323
rect 333 1317 387 1323
rect 397 1317 435 1323
rect 221 1297 243 1303
rect 429 1297 435 1317
rect 1053 1317 1091 1323
rect 1112 1317 1139 1323
rect 1224 1317 1251 1323
rect 2189 1317 2200 1323
rect 2312 1317 2323 1323
rect 2408 1317 2419 1323
rect 2669 1317 2712 1323
rect 2733 1317 2787 1323
rect 2989 1317 3027 1323
rect 749 1297 803 1303
rect 1800 1297 1843 1303
rect 2456 1297 2467 1303
rect 3021 1297 3027 1317
rect 3101 1317 3155 1323
rect 3373 1317 3411 1323
rect 3581 1317 3619 1323
rect 3485 1297 3523 1303
rect 808 1277 835 1283
rect 2984 1277 2995 1283
rect 445 1117 467 1123
rect 484 1116 488 1124
rect 173 1097 195 1103
rect 493 1097 504 1103
rect 685 1103 691 1123
rect 1037 1108 1043 1123
rect 2184 1117 2195 1123
rect 685 1097 723 1103
rect 733 1097 744 1103
rect 1021 1097 1032 1103
rect 1149 1097 1171 1103
rect 1693 1097 1720 1103
rect 1869 1097 1907 1103
rect 1976 1097 2019 1103
rect 2200 1097 2211 1103
rect 2221 1097 2259 1103
rect 3197 1097 3235 1103
rect 3325 1097 3352 1103
rect 3501 1097 3512 1103
rect 3597 1097 3608 1103
rect 621 1077 632 1083
rect 1197 1077 1224 1083
rect 1272 1077 1299 1083
rect 1517 1077 1544 1083
rect 1629 1077 1656 1083
rect 1773 1077 1843 1083
rect 1880 1077 1891 1083
rect 2120 1077 2131 1083
rect 2477 1077 2531 1083
rect 2968 1077 2979 1083
rect 1101 1057 1123 1063
rect 1160 1057 1171 1063
rect 1645 1057 1672 1063
rect 2696 1037 2707 1043
rect 541 977 552 983
rect 1821 977 1848 983
rect 1501 957 1512 963
rect 3277 957 3299 963
rect 781 937 792 943
rect 301 917 323 923
rect 781 923 787 937
rect 824 937 851 943
rect 888 937 915 943
rect 1117 937 1139 943
rect 1485 943 1491 952
rect 1469 937 1491 943
rect 2301 937 2323 943
rect 781 917 835 923
rect 893 917 904 923
rect 2157 917 2168 923
rect 2232 917 2243 923
rect 2317 923 2323 937
rect 2776 937 2787 943
rect 3165 937 3203 943
rect 3629 937 3656 943
rect 2317 917 2344 923
rect 2365 917 2404 923
rect 2396 912 2404 917
rect 2493 917 2531 923
rect 232 896 236 904
rect 957 897 968 903
rect 1821 897 1832 903
rect 1864 897 1875 903
rect 2493 897 2499 917
rect 2568 917 2579 923
rect 2589 917 2627 923
rect 2621 897 2627 917
rect 2941 917 2979 923
rect 3053 917 3091 923
rect 2765 897 2776 903
rect 3085 897 3091 917
rect 3304 917 3315 923
rect 541 877 584 883
rect 940 883 948 888
rect 940 877 979 883
rect 973 857 979 877
rect 1645 737 1656 743
rect 477 717 499 723
rect 989 717 1011 723
rect 1165 717 1187 723
rect 1325 717 1347 723
rect 157 697 195 703
rect 189 677 195 697
rect 296 697 323 703
rect 541 697 563 703
rect 1528 697 1539 703
rect 1560 697 1587 703
rect 1832 697 1859 703
rect 1917 697 1928 703
rect 2173 697 2184 703
rect 2285 697 2296 703
rect 568 677 579 683
rect 1037 677 1048 683
rect 1245 677 1288 683
rect 2285 683 2291 697
rect 2701 697 2712 703
rect 2765 697 2787 703
rect 3432 697 3443 703
rect 2136 677 2163 683
rect 2269 677 2291 683
rect 2333 677 2371 683
rect 2365 657 2371 677
rect 2424 677 2451 683
rect 2461 677 2499 683
rect 2461 657 2467 677
rect 2648 677 2675 683
rect 3293 677 3304 683
rect 3608 677 3619 683
rect 2045 637 2056 643
rect 125 577 136 583
rect 2093 557 2124 563
rect 461 537 499 543
rect 573 537 584 543
rect 669 537 680 543
rect 749 537 776 543
rect 1848 537 1859 543
rect 2253 537 2275 543
rect 360 517 371 523
rect 605 517 616 523
rect 760 517 819 523
rect 968 517 995 523
rect 1224 517 1251 523
rect 1789 517 1848 523
rect 2269 523 2275 537
rect 2653 537 2680 543
rect 2824 537 2867 543
rect 3021 537 3064 543
rect 3277 537 3331 543
rect 3405 537 3448 543
rect 3533 537 3544 543
rect 3645 537 3656 543
rect 2269 517 2308 523
rect 2300 516 2308 517
rect 2813 523 2819 532
rect 2797 517 2819 523
rect 3101 517 3112 523
rect 3240 517 3251 523
rect 3496 517 3507 523
rect 157 497 168 503
rect 1188 496 1192 504
rect 1444 496 1448 504
rect 3597 337 3656 343
rect 1021 317 1043 323
rect 1149 317 1171 323
rect 1332 316 1336 324
rect 1480 317 1491 323
rect 61 297 72 303
rect 221 297 232 303
rect 296 297 307 303
rect 525 297 536 303
rect 600 297 627 303
rect 712 297 723 303
rect 808 297 819 303
rect 1341 297 1368 303
rect 1437 297 1459 303
rect 1933 297 1944 303
rect 2205 297 2216 303
rect 2413 297 2435 303
rect 120 277 131 283
rect 312 277 323 283
rect 349 277 387 283
rect 957 277 984 283
rect 1629 277 1656 283
rect 2125 277 2179 283
rect 2413 283 2419 297
rect 2664 297 2675 303
rect 2776 297 2787 303
rect 2861 297 2883 303
rect 2280 277 2291 283
rect 2397 277 2419 283
rect 2461 277 2488 283
rect 2504 277 2515 283
rect 2701 277 2712 283
rect 2861 283 2867 297
rect 2989 297 3011 303
rect 2989 283 2995 297
rect 3064 297 3075 303
rect 3117 297 3139 303
rect 3181 297 3203 303
rect 3117 288 3123 297
rect 2813 277 2867 283
rect 2973 277 2995 283
rect 3101 277 3112 283
rect 3181 283 3187 297
rect 3437 297 3448 303
rect 3165 277 3187 283
rect 3293 277 3347 283
rect 1832 257 1843 263
rect 1805 177 1832 183
rect 77 137 88 143
rect 77 123 83 137
rect 61 117 83 123
rect 205 103 211 128
rect 456 117 467 123
rect 685 117 696 123
rect 760 117 792 123
rect 909 123 915 143
rect 2952 137 2963 143
rect 909 117 931 123
rect 1160 117 1187 123
rect 1320 117 1336 123
rect 1357 117 1379 123
rect 1517 117 1571 123
rect 1581 117 1603 123
rect 1997 117 2019 123
rect 2525 117 2536 123
rect 2957 123 2963 137
rect 3133 137 3155 143
rect 2957 117 2968 123
rect 3133 123 3139 137
rect 3389 137 3411 143
rect 3128 117 3139 123
rect 3192 117 3203 123
rect 3389 123 3395 137
rect 3464 137 3475 143
rect 3453 123 3459 132
rect 3373 117 3395 123
rect 3437 117 3459 123
rect 200 97 211 103
rect 1101 97 1123 103
rect 1236 96 1240 104
rect 1716 96 1720 104
rect 1832 97 1859 103
rect 157 77 200 83
<< m2contact >>
rect 765 2402 801 2418
rect 2813 2402 2849 2418
rect 312 2372 328 2388
rect 3272 2372 3288 2388
rect 3368 2372 3384 2388
rect 3480 2372 3496 2388
rect 8 2332 24 2348
rect 552 2312 568 2328
rect 632 2312 648 2328
rect 40 2292 56 2308
rect 104 2292 120 2308
rect 216 2292 248 2308
rect 280 2292 296 2308
rect 328 2292 344 2308
rect 392 2292 408 2308
rect 56 2272 72 2288
rect 264 2272 280 2288
rect 456 2292 472 2308
rect 600 2292 616 2308
rect 856 2312 872 2328
rect 680 2292 696 2308
rect 744 2292 760 2308
rect 824 2292 840 2308
rect 1160 2312 1176 2328
rect 1224 2312 1240 2328
rect 1272 2312 1288 2328
rect 1320 2312 1336 2328
rect 1384 2312 1400 2328
rect 1464 2312 1480 2328
rect 1528 2312 1544 2328
rect 1608 2312 1640 2328
rect 1800 2312 1816 2328
rect 1832 2312 1848 2328
rect 2920 2312 2936 2328
rect 904 2292 920 2308
rect 968 2292 984 2308
rect 1128 2292 1144 2308
rect 1192 2292 1208 2308
rect 1384 2292 1400 2308
rect 1448 2292 1464 2308
rect 1496 2292 1528 2308
rect 1736 2292 1752 2308
rect 1928 2292 1944 2308
rect 1992 2292 2008 2308
rect 2072 2292 2088 2308
rect 2136 2292 2152 2308
rect 2200 2292 2232 2308
rect 2264 2292 2280 2308
rect 2360 2292 2376 2308
rect 2424 2292 2440 2308
rect 2472 2292 2488 2308
rect 2536 2292 2552 2308
rect 2584 2292 2600 2308
rect 2664 2292 2680 2308
rect 2728 2292 2744 2308
rect 2776 2292 2792 2308
rect 3160 2312 3176 2328
rect 3512 2312 3528 2328
rect 3592 2312 3608 2328
rect 2968 2292 2984 2308
rect 3000 2292 3016 2308
rect 3128 2292 3144 2308
rect 3192 2292 3208 2308
rect 3240 2292 3256 2308
rect 3288 2292 3304 2308
rect 3336 2292 3352 2308
rect 3432 2292 3464 2308
rect 3544 2292 3576 2308
rect 1048 2288 1064 2292
rect 584 2272 600 2288
rect 696 2272 712 2288
rect 760 2272 776 2288
rect 888 2272 904 2288
rect 920 2272 936 2288
rect 984 2272 1000 2288
rect 1016 2276 1064 2288
rect 1016 2272 1048 2276
rect 1144 2272 1160 2288
rect 1176 2272 1192 2288
rect 1208 2272 1224 2288
rect 1256 2272 1272 2288
rect 1304 2272 1320 2288
rect 1336 2272 1352 2288
rect 1368 2272 1384 2288
rect 1416 2272 1432 2288
rect 1576 2272 1592 2288
rect 1656 2272 1672 2288
rect 1864 2272 1896 2288
rect 1960 2272 1976 2288
rect 2296 2272 2312 2288
rect 2888 2272 2904 2288
rect 2984 2272 3000 2288
rect 3032 2272 3080 2288
rect 3224 2272 3240 2288
rect 3320 2272 3336 2288
rect 1240 2252 1256 2268
rect 1688 2252 1704 2268
rect 2104 2252 2120 2268
rect 2456 2252 2472 2268
rect 136 2232 152 2248
rect 360 2232 376 2248
rect 424 2232 440 2248
rect 488 2232 504 2248
rect 648 2232 664 2248
rect 712 2232 728 2248
rect 936 2232 952 2248
rect 1000 2232 1016 2248
rect 1080 2232 1112 2248
rect 1288 2232 1304 2248
rect 1384 2232 1400 2248
rect 1528 2232 1544 2248
rect 1608 2232 1640 2248
rect 1768 2232 1784 2248
rect 1848 2232 1864 2248
rect 2040 2232 2056 2248
rect 2168 2232 2184 2248
rect 2312 2232 2328 2248
rect 2392 2232 2408 2248
rect 2440 2232 2456 2248
rect 2504 2232 2520 2248
rect 2568 2232 2584 2248
rect 2632 2232 2648 2248
rect 2696 2232 2712 2248
rect 2760 2232 2776 2248
rect 2824 2232 2840 2248
rect 2936 2232 2952 2248
rect 3400 2232 3416 2248
rect 1789 2202 1825 2218
rect 328 2172 344 2188
rect 456 2172 472 2188
rect 1160 2172 1176 2188
rect 1304 2172 1320 2188
rect 1928 2172 1944 2188
rect 2216 2172 2232 2188
rect 2376 2172 2392 2188
rect 3400 2172 3416 2188
rect 264 2154 280 2170
rect 680 2152 696 2168
rect 712 2152 744 2168
rect 936 2152 952 2168
rect 1000 2152 1016 2168
rect 1544 2152 1560 2168
rect 1768 2152 1784 2168
rect 1912 2152 1928 2168
rect 2808 2152 2824 2168
rect 3016 2152 3032 2168
rect 8 2132 24 2148
rect 56 2132 72 2148
rect 136 2132 152 2148
rect 40 2112 56 2128
rect 88 2112 120 2128
rect 200 2132 232 2148
rect 360 2132 376 2148
rect 488 2132 504 2148
rect 552 2132 584 2148
rect 680 2132 696 2148
rect 1000 2132 1016 2148
rect 1112 2132 1128 2148
rect 1272 2132 1288 2148
rect 1320 2132 1336 2148
rect 1480 2132 1496 2148
rect 1528 2132 1544 2148
rect 1576 2132 1592 2148
rect 1624 2132 1656 2148
rect 1672 2132 1688 2148
rect 1752 2132 1768 2148
rect 1832 2132 1848 2148
rect 1976 2132 2008 2148
rect 2088 2132 2120 2148
rect 280 2112 312 2128
rect 408 2112 440 2128
rect 568 2112 584 2128
rect 680 2112 696 2128
rect 760 2112 776 2128
rect 808 2112 824 2128
rect 888 2112 904 2128
rect 952 2112 968 2128
rect 984 2112 1000 2128
rect 1032 2112 1048 2128
rect 1064 2112 1080 2128
rect 1128 2112 1144 2128
rect 1192 2112 1208 2128
rect 1240 2112 1256 2128
rect 1272 2112 1288 2128
rect 1304 2112 1320 2128
rect 856 2092 872 2108
rect 1076 2092 1092 2108
rect 1096 2092 1112 2108
rect 1160 2092 1176 2108
rect 1304 2092 1320 2108
rect 1348 2092 1364 2108
rect 1384 2112 1416 2128
rect 1448 2112 1480 2128
rect 1512 2112 1528 2128
rect 1576 2112 1592 2128
rect 1608 2112 1624 2128
rect 1864 2112 1880 2128
rect 1960 2112 1976 2128
rect 1480 2092 1496 2108
rect 1576 2092 1592 2108
rect 1688 2092 1704 2108
rect 1724 2092 1740 2108
rect 1880 2092 1896 2108
rect 1928 2092 1944 2108
rect 2024 2092 2040 2108
rect 2056 2112 2088 2128
rect 2120 2112 2136 2128
rect 2392 2132 2424 2148
rect 2536 2132 2552 2148
rect 2600 2132 2616 2148
rect 2648 2132 2664 2148
rect 2680 2132 2696 2148
rect 2776 2132 2792 2148
rect 2840 2132 2856 2148
rect 2872 2132 2888 2148
rect 2984 2132 3000 2148
rect 3128 2132 3144 2148
rect 3240 2132 3256 2148
rect 2184 2112 2200 2128
rect 2232 2112 2264 2128
rect 2328 2112 2344 2128
rect 2456 2112 2472 2128
rect 2520 2112 2536 2128
rect 2552 2112 2568 2128
rect 2632 2112 2648 2128
rect 2664 2112 2680 2128
rect 2776 2112 2792 2128
rect 2808 2112 2824 2128
rect 2216 2092 2232 2108
rect 2564 2092 2580 2108
rect 2584 2092 2616 2108
rect 2728 2092 2744 2108
rect 2920 2092 2936 2108
rect 2952 2112 2984 2128
rect 3064 2092 3080 2108
rect 3096 2112 3128 2128
rect 3192 2112 3208 2128
rect 3272 2112 3304 2128
rect 3336 2112 3352 2128
rect 3368 2112 3384 2128
rect 3432 2112 3448 2128
rect 3560 2112 3576 2128
rect 872 2072 888 2088
rect 1912 2072 1928 2088
rect 3160 2052 3176 2068
rect 536 2032 552 2048
rect 616 2032 632 2048
rect 888 2032 904 2048
rect 1208 2032 1224 2048
rect 1416 2032 1432 2048
rect 2280 2032 2296 2048
rect 2424 2032 2440 2048
rect 2488 2032 2504 2048
rect 2712 2032 2728 2048
rect 3000 2032 3016 2048
rect 3304 2032 3320 2048
rect 3400 2032 3416 2048
rect 3464 2032 3480 2048
rect 3528 2032 3544 2048
rect 3592 2032 3608 2048
rect 765 2002 801 2018
rect 2813 2002 2849 2018
rect 872 1972 888 1988
rect 936 1972 952 1988
rect 2040 1972 2056 1988
rect 2296 1972 2312 1988
rect 2392 1972 2408 1988
rect 3496 1972 3512 1988
rect 1544 1952 1560 1968
rect 728 1932 744 1948
rect 888 1932 920 1948
rect 1464 1932 1480 1948
rect 1672 1932 1688 1948
rect 2072 1932 2088 1948
rect 2312 1932 2328 1948
rect 24 1912 40 1928
rect 216 1912 232 1928
rect 280 1912 296 1928
rect 376 1912 392 1928
rect 488 1912 504 1928
rect 680 1912 712 1928
rect 744 1912 760 1928
rect 968 1912 984 1928
rect 1064 1912 1080 1928
rect 1144 1912 1160 1928
rect 1336 1912 1352 1928
rect 1448 1912 1464 1928
rect 1496 1912 1528 1928
rect 1736 1912 1752 1928
rect 1816 1912 1832 1928
rect 1896 1912 1912 1928
rect 1992 1912 2024 1928
rect 2216 1912 2232 1928
rect 2280 1912 2296 1928
rect 2664 1912 2680 1928
rect 2760 1912 2776 1928
rect 2824 1912 2840 1928
rect 2888 1912 2904 1928
rect 2936 1912 2952 1928
rect 72 1892 88 1908
rect 184 1892 200 1908
rect 136 1872 152 1888
rect 312 1892 328 1908
rect 392 1892 408 1908
rect 456 1892 472 1908
rect 504 1892 520 1908
rect 632 1892 648 1908
rect 712 1892 728 1908
rect 840 1892 856 1908
rect 1016 1892 1032 1908
rect 1096 1892 1112 1908
rect 1208 1892 1224 1908
rect 1272 1892 1288 1908
rect 1320 1892 1336 1908
rect 1352 1892 1368 1908
rect 1416 1892 1432 1908
rect 1480 1892 1496 1908
rect 1544 1892 1560 1908
rect 1576 1892 1608 1908
rect 1928 1892 1944 1908
rect 2040 1892 2056 1908
rect 2120 1892 2152 1908
rect 2184 1892 2200 1908
rect 2232 1892 2264 1908
rect 2296 1892 2312 1908
rect 2344 1892 2360 1908
rect 2472 1892 2488 1908
rect 2568 1892 2584 1908
rect 2600 1892 2616 1908
rect 2664 1892 2680 1908
rect 2728 1892 2744 1908
rect 2792 1892 2808 1908
rect 3048 1912 3064 1928
rect 3000 1892 3016 1908
rect 3084 1912 3100 1928
rect 3240 1912 3256 1928
rect 3288 1912 3304 1928
rect 3096 1892 3112 1908
rect 3128 1892 3160 1908
rect 3192 1892 3208 1908
rect 3336 1892 3352 1908
rect 344 1888 360 1892
rect 328 1876 360 1888
rect 328 1872 344 1876
rect 520 1872 536 1888
rect 584 1872 600 1888
rect 616 1872 632 1888
rect 648 1872 664 1888
rect 856 1872 872 1888
rect 952 1872 968 1888
rect 1016 1872 1048 1888
rect 1080 1872 1096 1888
rect 1224 1872 1256 1888
rect 1368 1872 1384 1888
rect 1432 1872 1448 1888
rect 1560 1872 1576 1888
rect 1720 1872 1736 1888
rect 1768 1872 1784 1888
rect 1944 1872 1976 1888
rect 2056 1872 2072 1888
rect 2104 1872 2120 1888
rect 2264 1872 2280 1888
rect 2344 1872 2360 1888
rect 2424 1872 2440 1888
rect 2520 1872 2536 1888
rect 2616 1872 2648 1888
rect 2696 1872 2712 1888
rect 2808 1872 2824 1888
rect 2856 1872 2872 1888
rect 2904 1872 2920 1888
rect 2952 1872 2968 1888
rect 3000 1872 3032 1888
rect 3112 1872 3128 1888
rect 3224 1872 3240 1888
rect 3336 1872 3384 1888
rect 3576 1912 3592 1928
rect 3416 1892 3432 1908
rect 3464 1892 3496 1908
rect 3544 1892 3560 1908
rect 3624 1892 3640 1908
rect 3544 1872 3560 1888
rect 3640 1872 3656 1888
rect 424 1852 440 1868
rect 552 1852 568 1868
rect 664 1852 680 1868
rect 808 1852 824 1868
rect 1208 1852 1224 1868
rect 1320 1852 1336 1868
rect 1352 1852 1368 1868
rect 1608 1852 1624 1868
rect 1784 1852 1800 1868
rect 1832 1852 1848 1868
rect 1864 1852 1880 1868
rect 2088 1852 2104 1868
rect 2152 1852 2168 1868
rect 2424 1852 2440 1868
rect 2536 1852 2568 1868
rect 2616 1852 2632 1868
rect 2648 1852 2664 1868
rect 2712 1852 2728 1868
rect 104 1832 120 1848
rect 488 1832 504 1848
rect 600 1832 616 1848
rect 1048 1832 1064 1848
rect 1128 1832 1144 1848
rect 1224 1832 1240 1848
rect 1416 1832 1432 1848
rect 1752 1832 1768 1848
rect 1992 1832 2008 1848
rect 3160 1832 3176 1848
rect 3288 1832 3304 1848
rect 3592 1832 3608 1848
rect 1789 1802 1825 1818
rect 136 1772 152 1788
rect 200 1772 216 1788
rect 408 1772 424 1788
rect 744 1772 760 1788
rect 888 1772 904 1788
rect 1176 1772 1192 1788
rect 2008 1772 2024 1788
rect 2296 1772 2312 1788
rect 2456 1772 2472 1788
rect 3176 1772 3192 1788
rect 552 1752 568 1768
rect 664 1752 680 1768
rect 840 1752 856 1768
rect 8 1732 24 1748
rect 56 1732 72 1748
rect 40 1712 56 1728
rect 88 1712 120 1728
rect 280 1732 296 1748
rect 360 1732 376 1748
rect 440 1732 456 1748
rect 472 1732 488 1748
rect 616 1732 648 1748
rect 776 1732 792 1748
rect 824 1732 840 1748
rect 872 1732 888 1748
rect 1016 1752 1032 1768
rect 1496 1752 1512 1768
rect 1576 1752 1592 1768
rect 1992 1752 2008 1768
rect 2072 1752 2088 1768
rect 2664 1752 2680 1768
rect 2728 1752 2744 1768
rect 3048 1752 3064 1768
rect 3224 1752 3256 1768
rect 1064 1732 1080 1748
rect 1256 1732 1288 1748
rect 1336 1732 1352 1748
rect 1400 1732 1416 1748
rect 1560 1732 1576 1748
rect 1624 1732 1640 1748
rect 1688 1732 1704 1748
rect 1816 1732 1832 1748
rect 1864 1732 1896 1748
rect 1928 1732 1960 1748
rect 2056 1732 2072 1748
rect 2104 1732 2120 1748
rect 2168 1732 2184 1748
rect 280 1712 296 1728
rect 328 1712 344 1728
rect 376 1712 392 1728
rect 456 1712 472 1728
rect 488 1712 520 1728
rect 600 1712 632 1728
rect 648 1712 664 1728
rect 696 1712 712 1728
rect 920 1712 936 1728
rect 1000 1712 1016 1728
rect 1032 1712 1048 1728
rect 1080 1712 1096 1728
rect 1128 1712 1144 1728
rect 1224 1712 1240 1728
rect 1272 1712 1336 1728
rect 1384 1712 1400 1728
rect 1416 1712 1432 1728
rect 232 1692 248 1708
rect 264 1692 280 1708
rect 296 1692 312 1708
rect 328 1692 344 1708
rect 424 1692 440 1708
rect 680 1692 696 1708
rect 744 1692 760 1708
rect 904 1692 920 1708
rect 1032 1692 1048 1708
rect 1208 1692 1224 1708
rect 1352 1692 1368 1708
rect 1372 1692 1388 1708
rect 1608 1712 1624 1728
rect 1656 1712 1688 1728
rect 1704 1712 1736 1728
rect 1832 1712 1848 1728
rect 1912 1712 1928 1728
rect 2040 1712 2056 1728
rect 2328 1732 2344 1748
rect 2408 1732 2424 1748
rect 2504 1732 2520 1748
rect 2568 1732 2584 1748
rect 2616 1732 2632 1748
rect 2648 1732 2664 1748
rect 2712 1732 2728 1748
rect 2776 1732 2808 1748
rect 3096 1732 3112 1748
rect 3272 1732 3288 1748
rect 3320 1732 3336 1748
rect 3368 1732 3384 1748
rect 3432 1732 3448 1748
rect 2232 1712 2264 1728
rect 2296 1712 2312 1728
rect 2344 1712 2360 1728
rect 2616 1712 2632 1728
rect 2712 1712 2728 1728
rect 2840 1712 2888 1728
rect 2920 1712 2936 1728
rect 2952 1712 2968 1728
rect 3016 1712 3048 1728
rect 3080 1712 3096 1728
rect 3160 1712 3176 1728
rect 3272 1712 3288 1728
rect 3336 1712 3352 1728
rect 3416 1712 3432 1728
rect 3496 1712 3560 1728
rect 3624 1712 3640 1728
rect 1528 1692 1544 1708
rect 1576 1692 1592 1708
rect 1640 1692 1656 1708
rect 1880 1692 1896 1708
rect 1992 1692 2024 1708
rect 2072 1692 2088 1708
rect 2216 1692 2232 1708
rect 2296 1692 2312 1708
rect 2536 1692 2552 1708
rect 3128 1692 3160 1708
rect 3304 1692 3320 1708
rect 3368 1692 3384 1708
rect 520 1672 536 1688
rect 712 1672 728 1688
rect 856 1672 872 1688
rect 1736 1672 1752 1688
rect 2136 1672 2152 1688
rect 2600 1672 2632 1688
rect 3176 1672 3192 1688
rect 3384 1672 3416 1688
rect 552 1652 568 1668
rect 504 1632 520 1648
rect 696 1632 712 1648
rect 952 1632 968 1648
rect 1112 1632 1128 1648
rect 1176 1632 1192 1648
rect 1448 1632 1464 1648
rect 2200 1632 2216 1648
rect 2376 1632 2392 1648
rect 2664 1632 2680 1648
rect 2904 1632 2920 1648
rect 2984 1632 3000 1648
rect 3080 1632 3096 1648
rect 3112 1632 3128 1648
rect 3160 1632 3176 1648
rect 3208 1632 3224 1648
rect 3288 1632 3304 1648
rect 3464 1632 3480 1648
rect 3576 1632 3592 1648
rect 765 1602 801 1618
rect 2813 1602 2849 1618
rect 24 1572 40 1588
rect 296 1572 312 1588
rect 328 1572 344 1588
rect 376 1572 408 1588
rect 2344 1572 2360 1588
rect 3352 1572 3368 1588
rect 312 1532 328 1548
rect 520 1532 536 1548
rect 824 1532 856 1548
rect 1656 1532 1672 1548
rect 1752 1532 1768 1548
rect 248 1512 264 1528
rect 312 1512 328 1528
rect 488 1512 504 1528
rect 552 1512 568 1528
rect 952 1512 968 1528
rect 1064 1512 1080 1528
rect 1192 1512 1208 1528
rect 1288 1512 1320 1528
rect 1400 1512 1416 1528
rect 1624 1512 1640 1528
rect 1720 1512 1736 1528
rect 1784 1512 1800 1528
rect 1880 1512 1896 1528
rect 2008 1512 2024 1528
rect 88 1492 104 1508
rect 152 1492 168 1508
rect 184 1492 200 1508
rect 216 1492 232 1508
rect 248 1492 264 1508
rect 280 1492 296 1508
rect 536 1492 552 1508
rect 616 1492 632 1508
rect 680 1492 696 1508
rect 1000 1492 1016 1508
rect 1128 1492 1144 1508
rect 1192 1492 1208 1508
rect 1224 1492 1240 1508
rect 1336 1492 1352 1508
rect 1368 1492 1384 1508
rect 1432 1492 1464 1508
rect 1512 1492 1528 1508
rect 1576 1492 1592 1508
rect 1688 1492 1704 1508
rect 1720 1492 1736 1508
rect 1784 1492 1800 1508
rect 1880 1492 1896 1508
rect 1944 1492 1960 1508
rect 1976 1492 1992 1508
rect 2040 1492 2072 1508
rect 2088 1512 2104 1528
rect 2488 1512 2504 1528
rect 2136 1492 2152 1508
rect 2184 1492 2200 1508
rect 2328 1492 2360 1508
rect 2424 1492 2440 1508
rect 2568 1512 2584 1528
rect 2588 1512 2604 1528
rect 2648 1512 2664 1528
rect 3016 1512 3048 1528
rect 3096 1512 3112 1528
rect 3320 1512 3336 1528
rect 3368 1512 3400 1528
rect 3448 1512 3464 1528
rect 3468 1512 3484 1528
rect 3576 1512 3592 1528
rect 2600 1492 2616 1508
rect 2632 1492 2648 1508
rect 2664 1492 2696 1508
rect 2712 1492 2728 1508
rect 2744 1492 2776 1508
rect 2888 1492 2904 1508
rect 2952 1492 2968 1508
rect 2984 1492 3000 1508
rect 3048 1492 3064 1508
rect 3128 1492 3144 1508
rect 3288 1492 3320 1508
rect 3416 1492 3432 1508
rect 3480 1492 3496 1508
rect 3512 1492 3528 1508
rect 3608 1492 3624 1508
rect 72 1472 88 1488
rect 120 1476 136 1492
rect 344 1472 360 1488
rect 424 1472 440 1488
rect 456 1472 472 1488
rect 600 1472 616 1488
rect 664 1472 680 1488
rect 728 1472 744 1488
rect 152 1452 168 1468
rect 360 1452 376 1468
rect 440 1452 456 1468
rect 568 1452 584 1468
rect 632 1452 648 1468
rect 760 1472 776 1488
rect 872 1472 904 1488
rect 920 1472 936 1488
rect 1144 1472 1160 1488
rect 1240 1472 1272 1488
rect 1304 1472 1320 1488
rect 1368 1472 1384 1488
rect 1528 1472 1544 1488
rect 1560 1472 1576 1488
rect 1592 1472 1608 1488
rect 1672 1472 1688 1488
rect 1704 1472 1720 1488
rect 1736 1472 1752 1488
rect 1832 1472 1848 1488
rect 1928 1472 1944 1488
rect 1960 1472 1976 1488
rect 1992 1472 2008 1488
rect 2024 1472 2040 1488
rect 2120 1472 2136 1488
rect 2152 1472 2168 1488
rect 2216 1472 2232 1488
rect 2280 1472 2296 1488
rect 2312 1472 2328 1488
rect 2440 1472 2472 1488
rect 2552 1472 2568 1488
rect 2616 1472 2632 1488
rect 2696 1472 2712 1488
rect 2776 1472 2792 1488
rect 2936 1472 2952 1488
rect 2968 1472 2984 1488
rect 3000 1472 3016 1488
rect 3080 1472 3096 1488
rect 3144 1472 3176 1488
rect 3256 1472 3288 1488
rect 3336 1472 3352 1488
rect 3432 1472 3448 1488
rect 3496 1472 3512 1488
rect 3528 1472 3544 1488
rect 3624 1472 3640 1488
rect 968 1452 984 1468
rect 1160 1452 1176 1468
rect 1464 1452 1496 1468
rect 1528 1452 1544 1468
rect 1640 1452 1656 1468
rect 1896 1452 1912 1468
rect 2184 1452 2216 1468
rect 2296 1452 2312 1468
rect 2376 1452 2392 1468
rect 2664 1452 2680 1468
rect 2824 1452 2840 1468
rect 2856 1452 2872 1468
rect 3544 1452 3560 1468
rect 328 1432 344 1448
rect 488 1432 504 1448
rect 520 1432 536 1448
rect 584 1432 600 1448
rect 648 1432 664 1448
rect 696 1432 712 1448
rect 792 1432 824 1448
rect 904 1432 920 1448
rect 936 1432 952 1448
rect 1080 1432 1096 1448
rect 1144 1432 1160 1448
rect 1272 1432 1288 1448
rect 1416 1432 1432 1448
rect 1544 1432 1560 1448
rect 1880 1432 1896 1448
rect 2392 1432 2408 1448
rect 2504 1432 2520 1448
rect 2792 1432 2808 1448
rect 2920 1432 2936 1448
rect 3208 1432 3224 1448
rect 3384 1432 3400 1448
rect 1789 1402 1825 1418
rect 88 1372 104 1388
rect 216 1372 232 1388
rect 568 1372 584 1388
rect 744 1372 760 1388
rect 872 1372 888 1388
rect 1000 1372 1016 1388
rect 1288 1372 1304 1388
rect 1352 1372 1368 1388
rect 1640 1372 1656 1388
rect 1752 1372 1768 1388
rect 1928 1372 1944 1388
rect 2152 1372 2168 1388
rect 2248 1372 2264 1388
rect 2328 1372 2344 1388
rect 2440 1372 2456 1388
rect 2536 1372 2552 1388
rect 3176 1372 3192 1388
rect 3304 1372 3320 1388
rect 3560 1372 3576 1388
rect 168 1352 184 1368
rect 280 1352 296 1368
rect 328 1352 360 1368
rect 488 1352 504 1368
rect 552 1352 568 1368
rect 648 1352 664 1368
rect 1096 1352 1112 1368
rect 1992 1352 2008 1368
rect 2056 1352 2072 1368
rect 3240 1352 3256 1368
rect 3320 1352 3336 1368
rect 3416 1352 3432 1368
rect 3544 1352 3560 1368
rect 344 1332 360 1348
rect 440 1332 456 1348
rect 472 1332 488 1348
rect 536 1332 552 1348
rect 584 1332 600 1348
rect 728 1332 744 1348
rect 856 1332 872 1348
rect 968 1332 984 1348
rect 1064 1332 1080 1348
rect 1112 1332 1128 1348
rect 1224 1332 1240 1348
rect 1256 1332 1272 1348
rect 1336 1332 1352 1348
rect 1400 1332 1432 1348
rect 1464 1332 1480 1348
rect 1544 1332 1560 1348
rect 1608 1332 1624 1348
rect 1784 1332 1800 1348
rect 1816 1332 1832 1348
rect 1880 1332 1912 1348
rect 1928 1332 1944 1348
rect 2024 1332 2056 1348
rect 2120 1332 2152 1348
rect 2184 1332 2200 1348
rect 2392 1332 2408 1348
rect 2504 1332 2520 1348
rect 2552 1332 2568 1348
rect 2584 1332 2600 1348
rect 2680 1332 2712 1348
rect 2760 1332 2776 1348
rect 2840 1332 2856 1348
rect 2968 1332 2984 1348
rect 3000 1332 3016 1348
rect 3064 1332 3080 1348
rect 3112 1332 3144 1348
rect 3288 1332 3304 1348
rect 3320 1332 3336 1348
rect 3384 1332 3400 1348
rect 3432 1332 3448 1348
rect 3496 1332 3512 1348
rect 3624 1332 3640 1348
rect 56 1312 72 1328
rect 120 1312 152 1328
rect 248 1312 264 1328
rect 152 1292 168 1308
rect 408 1292 424 1308
rect 456 1312 472 1328
rect 520 1312 536 1328
rect 600 1312 632 1328
rect 696 1312 712 1328
rect 808 1312 824 1328
rect 936 1312 952 1328
rect 1096 1312 1112 1328
rect 1192 1312 1224 1328
rect 1320 1312 1336 1328
rect 1352 1312 1368 1328
rect 1384 1312 1400 1328
rect 1432 1312 1448 1328
rect 1480 1312 1496 1328
rect 1560 1312 1576 1328
rect 1672 1312 1688 1328
rect 1720 1312 1752 1328
rect 1864 1312 1880 1328
rect 2040 1312 2056 1328
rect 2104 1312 2136 1328
rect 2200 1312 2232 1328
rect 2264 1312 2312 1328
rect 2360 1312 2408 1328
rect 2472 1312 2504 1328
rect 2568 1312 2584 1328
rect 2600 1312 2616 1328
rect 2712 1312 2728 1328
rect 2792 1312 2808 1328
rect 2920 1312 2936 1328
rect 488 1292 504 1308
rect 632 1292 648 1308
rect 680 1292 696 1308
rect 712 1292 728 1308
rect 888 1292 904 1308
rect 952 1292 968 1308
rect 1000 1292 1032 1308
rect 1036 1292 1052 1308
rect 1144 1292 1176 1308
rect 1224 1292 1240 1308
rect 1464 1292 1480 1308
rect 1592 1292 1608 1308
rect 1640 1292 1656 1308
rect 1752 1292 1768 1308
rect 1784 1292 1800 1308
rect 1928 1292 1960 1308
rect 2232 1292 2248 1308
rect 2440 1292 2456 1308
rect 2520 1292 2536 1308
rect 2632 1292 2648 1308
rect 2744 1292 2760 1308
rect 2808 1292 2824 1308
rect 2872 1292 2920 1308
rect 3000 1292 3016 1308
rect 3048 1312 3064 1328
rect 3176 1312 3192 1328
rect 3208 1312 3224 1328
rect 3448 1312 3464 1328
rect 3080 1292 3096 1308
rect 3256 1292 3288 1308
rect 3336 1292 3352 1308
rect 3460 1292 3476 1308
rect 3528 1292 3544 1308
rect 3592 1292 3608 1308
rect 216 1272 232 1288
rect 792 1272 808 1288
rect 920 1272 936 1288
rect 1512 1272 1528 1288
rect 2936 1272 2952 1288
rect 2968 1272 2984 1288
rect 2920 1252 2936 1268
rect 24 1232 40 1248
rect 296 1232 312 1248
rect 696 1232 712 1248
rect 808 1232 824 1248
rect 936 1232 952 1248
rect 1192 1232 1208 1248
rect 1560 1232 1576 1248
rect 1688 1232 1704 1248
rect 765 1202 801 1218
rect 2813 1202 2849 1218
rect 168 1172 184 1188
rect 584 1172 600 1188
rect 1144 1172 1160 1188
rect 1352 1172 1368 1188
rect 1448 1172 1464 1188
rect 1896 1172 1912 1188
rect 1960 1172 1976 1188
rect 2328 1172 2344 1188
rect 2408 1172 2424 1188
rect 2920 1172 2936 1188
rect 3112 1172 3128 1188
rect 3384 1172 3400 1188
rect 1432 1132 1448 1148
rect 2392 1132 2408 1148
rect 2584 1132 2616 1148
rect 2696 1132 2712 1148
rect 3560 1132 3576 1148
rect 244 1112 260 1128
rect 264 1112 280 1128
rect 488 1112 504 1128
rect 520 1112 536 1128
rect 72 1092 104 1108
rect 120 1092 136 1108
rect 232 1092 248 1108
rect 312 1092 328 1108
rect 376 1092 408 1108
rect 504 1092 520 1108
rect 536 1092 568 1108
rect 696 1112 712 1128
rect 792 1112 808 1128
rect 840 1112 856 1128
rect 1464 1112 1480 1128
rect 1720 1112 1736 1128
rect 1912 1112 1944 1128
rect 2040 1112 2072 1128
rect 2168 1112 2184 1128
rect 2424 1112 2440 1128
rect 2504 1112 2520 1128
rect 2552 1112 2568 1128
rect 2616 1112 2648 1128
rect 2664 1112 2680 1128
rect 2792 1112 2808 1128
rect 3000 1112 3016 1128
rect 3032 1112 3064 1128
rect 3160 1112 3176 1128
rect 3288 1112 3304 1128
rect 744 1092 760 1108
rect 872 1092 888 1108
rect 952 1092 984 1108
rect 1032 1092 1048 1108
rect 1224 1092 1240 1108
rect 1320 1092 1336 1108
rect 1448 1092 1464 1108
rect 1480 1092 1496 1108
rect 1608 1092 1624 1108
rect 1672 1092 1688 1108
rect 1720 1092 1736 1108
rect 1752 1092 1768 1108
rect 1960 1092 1976 1108
rect 2072 1092 2104 1108
rect 2136 1092 2152 1108
rect 2184 1092 2200 1108
rect 2280 1092 2312 1108
rect 2344 1092 2360 1108
rect 2408 1092 2424 1108
rect 2488 1092 2504 1108
rect 2568 1092 2584 1108
rect 2680 1092 2696 1108
rect 2776 1092 2792 1108
rect 2872 1092 2904 1108
rect 2936 1092 2952 1108
rect 3064 1092 3096 1108
rect 3128 1092 3160 1108
rect 3176 1092 3192 1108
rect 3304 1092 3320 1108
rect 3352 1092 3384 1108
rect 3400 1092 3416 1108
rect 3432 1092 3464 1108
rect 3512 1092 3560 1108
rect 3608 1092 3624 1108
rect 24 1072 40 1088
rect 216 1072 232 1088
rect 296 1072 312 1088
rect 328 1072 344 1088
rect 360 1072 376 1088
rect 392 1072 424 1088
rect 504 1072 520 1088
rect 568 1072 584 1088
rect 632 1072 664 1088
rect 744 1072 776 1088
rect 856 1072 872 1088
rect 888 1072 904 1088
rect 936 1072 952 1088
rect 1000 1072 1016 1088
rect 1064 1072 1080 1088
rect 1224 1072 1272 1088
rect 1400 1072 1416 1088
rect 1544 1072 1560 1088
rect 1656 1072 1672 1088
rect 1720 1072 1736 1088
rect 1848 1072 1880 1088
rect 1976 1072 2008 1088
rect 2104 1072 2120 1088
rect 2168 1072 2184 1088
rect 2232 1072 2248 1088
rect 2536 1072 2552 1088
rect 2648 1072 2664 1088
rect 2760 1072 2776 1088
rect 2824 1072 2840 1088
rect 2952 1072 2968 1088
rect 3016 1072 3032 1088
rect 3208 1072 3224 1088
rect 3256 1072 3272 1088
rect 3352 1072 3368 1088
rect 3416 1072 3432 1088
rect 3496 1072 3512 1088
rect 8 1052 24 1068
rect 56 1052 72 1068
rect 136 1052 152 1068
rect 200 1052 216 1068
rect 280 1052 296 1068
rect 440 1052 456 1068
rect 632 1052 648 1068
rect 904 1052 920 1068
rect 968 1052 984 1068
rect 1080 1052 1096 1068
rect 1144 1052 1160 1068
rect 1208 1052 1224 1068
rect 1256 1052 1272 1068
rect 1624 1052 1640 1068
rect 1672 1052 1688 1068
rect 1704 1052 1720 1068
rect 1816 1052 1832 1068
rect 2040 1052 2056 1068
rect 2264 1052 2280 1068
rect 2440 1052 2472 1068
rect 2520 1052 2536 1068
rect 2728 1052 2744 1068
rect 3240 1052 3256 1068
rect 3336 1052 3352 1068
rect 360 1032 376 1048
rect 680 1032 696 1048
rect 792 1032 808 1048
rect 920 1032 936 1048
rect 1032 1032 1048 1048
rect 1096 1032 1112 1048
rect 1592 1032 1608 1048
rect 2680 1032 2696 1048
rect 2744 1032 2760 1048
rect 2792 1032 2808 1048
rect 2984 1032 3000 1048
rect 3096 1032 3112 1048
rect 3160 1032 3176 1048
rect 3272 1032 3288 1048
rect 1789 1002 1825 1018
rect 120 972 136 988
rect 392 972 408 988
rect 552 972 568 988
rect 632 972 648 988
rect 936 972 952 988
rect 1320 972 1336 988
rect 1608 972 1624 988
rect 1640 972 1672 988
rect 1752 972 1768 988
rect 1848 972 1864 988
rect 1944 972 1960 988
rect 1976 972 1992 988
rect 2056 972 2072 988
rect 2488 972 2504 988
rect 3000 972 3016 988
rect 3352 972 3368 988
rect 3528 972 3544 988
rect 264 952 280 968
rect 328 952 360 968
rect 664 952 680 968
rect 1032 952 1064 968
rect 1144 952 1160 968
rect 1368 952 1384 968
rect 1480 952 1496 968
rect 1512 952 1528 968
rect 1768 952 1784 968
rect 2040 952 2056 968
rect 2136 952 2152 968
rect 2504 952 2520 968
rect 2664 952 2696 968
rect 2856 952 2872 968
rect 2920 952 2936 968
rect 3176 952 3192 968
rect 3256 952 3272 968
rect 3512 952 3528 968
rect 72 944 88 948
rect 72 932 104 944
rect 136 932 152 948
rect 184 932 216 948
rect 440 944 472 948
rect 440 932 488 944
rect 584 932 600 948
rect 760 932 776 948
rect 88 928 104 932
rect 472 928 488 932
rect 56 912 72 928
rect 152 912 168 928
rect 216 912 232 928
rect 552 912 568 928
rect 600 912 616 928
rect 696 912 712 928
rect 792 932 824 948
rect 872 932 888 948
rect 1064 932 1080 948
rect 1176 932 1192 948
rect 1272 932 1288 948
rect 1560 932 1576 948
rect 1624 932 1640 948
rect 1704 932 1720 948
rect 1736 932 1752 948
rect 1784 932 1800 948
rect 1880 932 1896 948
rect 1912 932 1944 948
rect 2024 932 2040 948
rect 2088 932 2104 948
rect 2184 932 2200 948
rect 2216 932 2232 948
rect 904 912 920 928
rect 968 912 984 928
rect 1016 912 1032 928
rect 1096 912 1112 928
rect 1192 912 1208 928
rect 1240 912 1272 928
rect 1304 912 1320 928
rect 1384 912 1400 928
rect 1432 912 1464 928
rect 1544 912 1560 928
rect 1576 912 1592 928
rect 1688 912 1704 928
rect 1720 912 1736 928
rect 1896 912 1912 928
rect 2008 912 2024 928
rect 2072 912 2088 928
rect 2168 912 2184 928
rect 2200 912 2232 928
rect 2248 912 2264 928
rect 2296 912 2312 928
rect 2328 932 2344 948
rect 2456 932 2472 948
rect 2552 932 2568 948
rect 2632 932 2664 948
rect 2696 932 2712 948
rect 2728 932 2744 948
rect 2760 932 2776 948
rect 2872 932 2888 948
rect 2952 932 2968 948
rect 3016 932 3032 948
rect 3128 932 3144 948
rect 3224 932 3240 948
rect 3368 932 3384 948
rect 3480 932 3496 948
rect 3576 932 3592 948
rect 3656 932 3672 948
rect 2344 912 2360 928
rect 2408 912 2424 928
rect 184 892 200 908
rect 216 892 232 908
rect 248 892 264 908
rect 504 892 520 908
rect 568 892 584 908
rect 680 892 696 908
rect 712 892 728 908
rect 744 892 760 908
rect 936 892 952 908
rect 968 892 984 908
rect 1064 892 1080 908
rect 1176 892 1192 908
rect 1208 892 1240 908
rect 1288 892 1304 908
rect 1400 892 1432 908
rect 1608 892 1624 908
rect 1656 892 1672 908
rect 1832 892 1864 908
rect 1960 892 1992 908
rect 2104 892 2136 908
rect 2168 892 2184 908
rect 2376 892 2392 908
rect 2536 912 2568 928
rect 2600 892 2616 908
rect 2712 912 2728 928
rect 3032 912 3048 928
rect 2776 892 2792 908
rect 2808 892 2824 908
rect 3000 892 3016 908
rect 3064 892 3080 908
rect 3096 912 3128 928
rect 3144 912 3160 928
rect 3208 912 3224 928
rect 3288 912 3304 928
rect 3320 912 3336 928
rect 3384 912 3400 928
rect 3448 912 3464 928
rect 3544 912 3560 928
rect 3592 912 3608 928
rect 3240 892 3256 908
rect 3272 892 3288 908
rect 3336 892 3352 908
rect 296 872 312 888
rect 584 872 600 888
rect 984 872 1000 888
rect 1320 872 1336 888
rect 1368 872 1384 888
rect 2424 872 2440 888
rect 2536 872 2552 888
rect 24 832 40 848
rect 360 832 376 848
rect 648 832 664 848
rect 728 832 744 848
rect 840 832 856 848
rect 920 832 936 848
rect 1544 832 1560 848
rect 2440 832 2456 848
rect 2744 832 2760 848
rect 2792 832 2808 848
rect 2904 832 2920 848
rect 3416 832 3432 848
rect 3480 832 3496 848
rect 765 802 801 818
rect 2813 802 2849 818
rect 24 772 40 788
rect 88 772 104 788
rect 280 772 296 788
rect 696 772 712 788
rect 824 772 840 788
rect 1240 772 1256 788
rect 1576 772 1592 788
rect 1688 772 1704 788
rect 1768 772 1784 788
rect 1896 772 1912 788
rect 1944 772 1960 788
rect 1992 772 2008 788
rect 2952 772 2968 788
rect 3032 772 3048 788
rect 3512 772 3528 788
rect 648 752 664 768
rect 520 732 536 748
rect 632 732 648 748
rect 840 732 856 748
rect 904 732 920 748
rect 1656 732 1672 748
rect 2040 732 2056 748
rect 2120 732 2136 748
rect 3576 732 3592 748
rect 232 712 248 728
rect 324 712 340 728
rect 344 712 360 728
rect 392 712 408 728
rect 664 712 680 728
rect 744 712 760 728
rect 872 712 888 728
rect 936 712 952 728
rect 1096 712 1112 728
rect 1256 712 1272 728
rect 1448 712 1464 728
rect 1512 712 1528 728
rect 1608 712 1640 728
rect 1976 712 1992 728
rect 2072 712 2088 728
rect 2328 712 2344 728
rect 2488 712 2504 728
rect 2632 712 2648 728
rect 3256 712 3272 728
rect 56 692 72 708
rect 120 692 136 708
rect 168 672 184 688
rect 200 692 232 708
rect 280 692 296 708
rect 504 692 520 708
rect 648 692 664 708
rect 776 692 792 708
rect 856 692 872 708
rect 920 692 936 708
rect 1048 692 1064 708
rect 1112 692 1128 708
rect 1272 692 1288 708
rect 1352 692 1384 708
rect 1400 692 1416 708
rect 1480 692 1496 708
rect 1512 692 1528 708
rect 1544 692 1560 708
rect 1704 692 1752 708
rect 1784 692 1800 708
rect 1816 692 1832 708
rect 1864 692 1880 708
rect 1928 692 1944 708
rect 2056 692 2072 708
rect 2184 692 2200 708
rect 2216 692 2248 708
rect 296 672 312 688
rect 360 672 376 688
rect 424 672 456 688
rect 552 672 568 688
rect 712 672 728 688
rect 952 672 968 688
rect 1048 672 1080 688
rect 1128 672 1144 688
rect 1208 672 1240 688
rect 1288 672 1304 688
rect 1384 672 1400 688
rect 1416 672 1432 688
rect 1464 672 1480 688
rect 1512 672 1528 688
rect 1560 672 1576 688
rect 1656 672 1672 688
rect 2008 672 2024 688
rect 2088 672 2104 688
rect 2120 672 2136 688
rect 2296 692 2312 708
rect 2408 692 2440 708
rect 2520 692 2568 708
rect 2712 692 2744 708
rect 2872 692 2888 708
rect 2984 692 3016 708
rect 3064 692 3080 708
rect 3176 692 3208 708
rect 3352 692 3368 708
rect 3416 692 3432 708
rect 3480 692 3496 708
rect 3544 692 3560 708
rect 3640 692 3656 708
rect 248 652 264 668
rect 376 652 392 668
rect 456 652 472 668
rect 600 652 616 668
rect 904 652 920 668
rect 1000 652 1016 668
rect 1160 652 1176 668
rect 1320 652 1336 668
rect 1448 652 1464 668
rect 1544 652 1560 668
rect 1672 652 1688 668
rect 1960 652 1976 668
rect 2136 652 2152 668
rect 2184 652 2200 668
rect 2392 672 2424 688
rect 2600 672 2616 688
rect 2632 672 2648 688
rect 2680 672 2696 688
rect 2904 672 2920 688
rect 3096 672 3112 688
rect 3224 672 3240 688
rect 3304 672 3336 688
rect 3384 672 3400 688
rect 3464 672 3480 688
rect 3592 672 3608 688
rect 2648 652 2664 668
rect 3144 652 3160 668
rect 24 632 40 648
rect 152 632 168 648
rect 584 632 600 648
rect 984 632 1000 648
rect 1096 632 1112 648
rect 1192 632 1208 648
rect 2056 632 2072 648
rect 2104 632 2120 648
rect 2200 632 2216 648
rect 2376 632 2392 648
rect 2584 632 2600 648
rect 2632 632 2648 648
rect 2760 632 2776 648
rect 2808 632 2824 648
rect 2952 632 2968 648
rect 3256 632 3272 648
rect 1789 602 1825 618
rect 56 572 72 588
rect 136 572 152 588
rect 200 572 216 588
rect 888 572 904 588
rect 936 572 952 588
rect 1144 572 1160 588
rect 1496 572 1512 588
rect 1544 572 1560 588
rect 1624 572 1640 588
rect 2472 572 2488 588
rect 2632 572 2648 588
rect 2760 572 2776 588
rect 296 552 312 568
rect 392 552 408 568
rect 424 552 440 568
rect 504 552 520 568
rect 632 552 648 568
rect 904 552 936 568
rect 1352 552 1368 568
rect 1704 552 1720 568
rect 1736 552 1752 568
rect 2536 552 2552 568
rect 2616 552 2632 568
rect 8 532 24 548
rect 168 532 184 548
rect 344 532 360 548
rect 408 532 424 548
rect 584 532 600 548
rect 680 532 696 548
rect 776 532 808 548
rect 840 532 856 548
rect 872 532 888 548
rect 968 532 984 548
rect 1000 532 1016 548
rect 1032 532 1048 548
rect 1080 532 1112 548
rect 1208 532 1240 548
rect 1336 532 1352 548
rect 1384 532 1400 548
rect 1464 532 1480 548
rect 1592 532 1624 548
rect 1800 532 1816 548
rect 1832 532 1848 548
rect 2136 532 2152 548
rect 2200 532 2216 548
rect 72 512 88 528
rect 136 512 152 528
rect 248 512 264 528
rect 312 512 328 528
rect 344 512 360 528
rect 392 512 408 528
rect 440 512 456 528
rect 472 512 488 528
rect 520 512 536 528
rect 552 512 568 528
rect 616 512 632 528
rect 648 512 664 528
rect 680 512 696 528
rect 728 512 760 528
rect 856 512 872 528
rect 952 512 968 528
rect 1048 512 1064 528
rect 1112 512 1128 528
rect 1192 512 1224 528
rect 1304 512 1336 528
rect 1368 512 1384 528
rect 1400 512 1416 528
rect 1448 512 1464 528
rect 1512 512 1528 528
rect 1576 512 1592 528
rect 1656 512 1672 528
rect 1848 512 1864 528
rect 1960 512 1992 528
rect 2024 512 2040 528
rect 2056 512 2072 528
rect 2168 512 2200 528
rect 2216 512 2232 528
rect 2280 532 2296 548
rect 2424 532 2440 548
rect 2680 532 2696 548
rect 2808 532 2824 548
rect 2904 532 2920 548
rect 2952 532 2968 548
rect 3064 532 3080 548
rect 3144 532 3160 548
rect 3448 532 3464 548
rect 3544 532 3560 548
rect 3656 532 3672 548
rect 2376 512 2392 528
rect 2408 512 2424 528
rect 2504 512 2536 528
rect 2568 512 2584 528
rect 2664 512 2680 528
rect 2728 512 2744 528
rect 2888 512 2904 528
rect 2984 512 3000 528
rect 3112 512 3128 528
rect 3224 512 3240 528
rect 3352 512 3384 528
rect 3480 512 3496 528
rect 3608 512 3624 528
rect 88 492 104 508
rect 168 492 184 508
rect 200 492 216 508
rect 264 492 280 508
rect 328 492 344 508
rect 616 492 632 508
rect 696 492 712 508
rect 716 492 732 508
rect 840 492 856 508
rect 1016 492 1032 508
rect 1080 492 1096 508
rect 1144 492 1176 508
rect 1192 492 1208 508
rect 1252 492 1268 508
rect 1272 492 1304 508
rect 1416 492 1432 508
rect 1448 492 1464 508
rect 1528 492 1560 508
rect 1640 492 1656 508
rect 1768 492 1784 508
rect 1944 492 1960 508
rect 2040 492 2056 508
rect 2072 492 2088 508
rect 2104 492 2120 508
rect 2152 492 2168 508
rect 2600 492 2616 508
rect 24 472 40 488
rect 56 472 72 488
rect 120 472 136 488
rect 232 472 248 488
rect 296 472 312 488
rect 1496 472 1512 488
rect 1672 472 1688 488
rect 2008 472 2024 488
rect 2376 472 2392 488
rect 2568 472 2584 488
rect 3192 472 3208 488
rect 3272 472 3288 488
rect 248 452 264 468
rect 1656 452 1672 468
rect 1720 452 1736 468
rect 2024 452 2040 468
rect 1624 432 1640 448
rect 1752 432 1768 448
rect 1896 432 1912 448
rect 1960 432 1976 448
rect 2328 432 2344 448
rect 2392 432 2408 448
rect 2584 432 2600 448
rect 2696 432 2712 448
rect 2760 432 2776 448
rect 2856 432 2872 448
rect 3560 432 3576 448
rect 765 402 801 418
rect 2813 402 2849 418
rect 344 372 360 388
rect 488 372 504 388
rect 680 372 696 388
rect 904 372 920 388
rect 1064 372 1080 388
rect 1192 372 1208 388
rect 1384 372 1400 388
rect 1592 372 1608 388
rect 1720 372 1736 388
rect 2696 372 2712 388
rect 2808 372 2824 388
rect 2904 372 2920 388
rect 3288 372 3304 388
rect 3480 372 3496 388
rect 568 352 584 368
rect 104 332 120 348
rect 440 332 456 348
rect 1960 332 1976 348
rect 3656 332 3672 348
rect 280 312 296 328
rect 408 312 424 328
rect 1304 312 1320 328
rect 1336 312 1352 328
rect 1464 312 1480 328
rect 1688 312 1704 328
rect 1752 312 1768 328
rect 1944 312 1960 328
rect 2024 312 2040 328
rect 24 292 40 308
rect 72 292 88 308
rect 104 292 120 308
rect 152 292 168 308
rect 184 292 200 308
rect 232 292 264 308
rect 280 292 296 308
rect 360 292 376 308
rect 424 292 440 308
rect 456 292 472 308
rect 536 292 552 308
rect 584 292 600 308
rect 632 292 664 308
rect 696 292 712 308
rect 792 292 808 308
rect 872 292 888 308
rect 968 292 984 308
rect 1064 292 1080 308
rect 1096 292 1112 308
rect 1192 292 1208 308
rect 1368 292 1384 308
rect 1416 292 1432 308
rect 1496 292 1528 308
rect 1560 292 1576 308
rect 1640 292 1656 308
rect 1720 292 1736 308
rect 1848 292 1864 308
rect 1880 292 1896 308
rect 1912 292 1928 308
rect 1944 292 1960 308
rect 2056 292 2072 308
rect 2088 292 2104 308
rect 2216 292 2232 308
rect 2360 292 2376 308
rect 8 272 24 288
rect 104 272 120 288
rect 168 272 184 288
rect 200 272 216 288
rect 232 272 248 288
rect 296 272 312 288
rect 840 272 856 288
rect 984 272 1000 288
rect 1080 272 1096 288
rect 1112 272 1128 288
rect 1208 272 1224 288
rect 1288 272 1304 288
rect 1352 272 1368 288
rect 1528 272 1560 288
rect 1656 272 1672 288
rect 1704 272 1720 288
rect 1768 272 1784 288
rect 1864 272 1880 288
rect 1896 272 1912 288
rect 1992 272 2008 288
rect 2040 272 2056 288
rect 2072 272 2088 288
rect 2264 272 2280 288
rect 2536 292 2552 308
rect 2568 292 2600 308
rect 2648 292 2664 308
rect 2760 292 2776 308
rect 2488 272 2504 288
rect 2712 272 2728 288
rect 2936 292 2952 308
rect 3048 292 3064 308
rect 3112 272 3128 288
rect 3256 292 3272 308
rect 3368 292 3384 308
rect 3448 292 3464 308
rect 3512 292 3528 308
rect 3560 292 3576 308
rect 3544 272 3560 288
rect 72 252 88 268
rect 280 252 296 268
rect 392 252 408 268
rect 600 252 616 268
rect 744 252 760 268
rect 936 252 952 268
rect 1016 252 1032 268
rect 1144 252 1160 268
rect 1368 252 1384 268
rect 1400 252 1416 268
rect 1464 252 1480 268
rect 1608 252 1624 268
rect 1688 252 1704 268
rect 1816 252 1832 268
rect 1976 252 1992 268
rect 2552 252 2568 268
rect 136 232 152 248
rect 680 232 696 248
rect 1272 232 1288 248
rect 1784 232 1800 248
rect 2008 232 2024 248
rect 2120 232 2136 248
rect 2248 232 2264 248
rect 2328 232 2344 248
rect 2392 232 2408 248
rect 2616 232 2632 248
rect 2728 232 2744 248
rect 2968 232 2984 248
rect 3032 232 3048 248
rect 3160 232 3176 248
rect 3224 232 3240 248
rect 3400 232 3416 248
rect 3480 232 3496 248
rect 1789 202 1825 218
rect 248 172 264 188
rect 296 172 312 188
rect 360 172 376 188
rect 488 172 504 188
rect 616 172 632 188
rect 648 172 664 188
rect 712 172 728 188
rect 920 172 936 188
rect 1272 172 1288 188
rect 1560 172 1576 188
rect 1624 172 1640 188
rect 1832 172 1848 188
rect 1960 172 1976 188
rect 2024 172 2040 188
rect 2488 172 2504 188
rect 2568 172 2584 188
rect 3080 172 3096 188
rect 3400 172 3416 188
rect 824 152 840 168
rect 1096 152 1112 168
rect 1192 152 1208 168
rect 1336 152 1352 168
rect 1400 152 1416 168
rect 1432 152 1448 168
rect 1544 152 1560 168
rect 1608 152 1624 168
rect 1976 152 1992 168
rect 2040 152 2056 168
rect 24 132 40 148
rect 88 132 104 148
rect 584 132 600 148
rect 120 112 136 128
rect 168 112 184 128
rect 184 92 200 108
rect 216 112 232 128
rect 280 112 296 128
rect 328 112 344 128
rect 440 112 456 128
rect 520 112 536 128
rect 696 112 712 128
rect 744 112 760 128
rect 792 112 808 128
rect 888 112 904 128
rect 968 132 984 148
rect 1000 132 1016 148
rect 1032 132 1048 148
rect 1064 132 1080 148
rect 1128 132 1144 148
rect 1160 132 1176 148
rect 1256 132 1272 148
rect 1320 132 1336 148
rect 1384 132 1400 148
rect 1528 132 1544 148
rect 1672 132 1688 148
rect 1736 132 1768 148
rect 1896 132 1928 148
rect 2088 132 2104 148
rect 2152 132 2168 148
rect 2248 132 2264 148
rect 2312 132 2328 148
rect 2408 132 2424 148
rect 2616 132 2632 148
rect 2744 132 2760 148
rect 2792 132 2808 148
rect 2936 132 2952 148
rect 952 112 968 128
rect 1016 112 1032 128
rect 1048 112 1064 128
rect 1144 112 1160 128
rect 1240 112 1256 128
rect 1304 112 1320 128
rect 1336 112 1352 128
rect 1464 112 1480 128
rect 1656 112 1672 128
rect 1720 112 1736 128
rect 1768 112 1784 128
rect 1864 112 1896 128
rect 1928 112 1944 128
rect 2056 112 2072 128
rect 2120 112 2136 128
rect 2168 112 2184 128
rect 2216 112 2232 128
rect 2280 112 2296 128
rect 2328 112 2344 128
rect 2376 112 2392 128
rect 2424 112 2440 128
rect 2536 112 2552 128
rect 2648 112 2664 128
rect 2696 112 2728 128
rect 2760 112 2776 128
rect 2856 112 2872 128
rect 2904 112 2920 128
rect 3000 132 3016 148
rect 2968 112 2984 128
rect 3016 112 3032 128
rect 3112 112 3128 128
rect 3224 132 3240 148
rect 3336 132 3352 148
rect 3176 112 3192 128
rect 3240 112 3256 128
rect 3288 112 3304 128
rect 3448 132 3464 148
rect 3576 132 3592 148
rect 3496 112 3544 128
rect 3576 112 3592 128
rect 264 92 280 108
rect 408 92 424 108
rect 856 92 872 108
rect 984 92 1000 108
rect 1208 92 1224 108
rect 1240 92 1256 108
rect 1272 92 1288 108
rect 1480 92 1496 108
rect 1624 92 1640 108
rect 1688 92 1704 108
rect 1720 92 1736 108
rect 1816 92 1832 108
rect 200 72 216 88
rect 296 72 312 88
rect 552 72 568 88
rect 616 72 632 88
rect 1512 72 1528 88
rect 168 52 184 68
rect 888 52 904 68
rect 2200 32 2216 48
rect 2360 32 2376 48
rect 2456 32 2472 48
rect 2664 32 2680 48
rect 2888 32 2904 48
rect 3048 32 3064 48
rect 3272 32 3288 48
rect 3320 32 3336 48
rect 765 2 801 18
rect 2813 2 2849 18
<< metal2 >>
rect 317 2388 323 2463
rect 13 2328 19 2332
rect 557 2308 563 2312
rect 685 2308 691 2463
rect 813 2428 819 2463
rect 56 2297 67 2303
rect 61 2288 67 2297
rect 269 2297 280 2303
rect 109 2148 115 2292
rect 141 2148 147 2232
rect 221 2148 227 2292
rect 269 2288 275 2297
rect 333 2188 339 2292
rect 280 2157 291 2163
rect 13 2128 19 2132
rect 61 2123 67 2132
rect 109 2128 115 2132
rect 285 2128 291 2157
rect 365 2148 371 2232
rect 365 2128 371 2132
rect 429 2128 435 2232
rect 461 2188 467 2292
rect 493 2148 499 2232
rect 557 2148 563 2252
rect 605 2156 611 2292
rect 685 2268 691 2292
rect 701 2288 707 2332
rect 733 2297 744 2303
rect 664 2237 675 2243
rect 573 2148 579 2152
rect 56 2117 67 2123
rect 29 1908 35 1912
rect 93 1908 99 2112
rect 13 1728 19 1732
rect 29 1588 35 1892
rect 141 1888 147 1892
rect 61 1723 67 1732
rect 93 1728 99 1812
rect 109 1728 115 1832
rect 141 1788 147 1872
rect 205 1788 211 1892
rect 56 1717 67 1723
rect 93 1523 99 1712
rect 237 1688 243 1692
rect 93 1517 115 1523
rect 61 1328 67 1432
rect 45 1317 56 1323
rect 29 1203 35 1232
rect 45 1203 51 1317
rect 77 1208 83 1472
rect 109 1383 115 1517
rect 125 1468 131 1476
rect 104 1377 115 1383
rect 109 1323 115 1377
rect 173 1368 179 1512
rect 189 1368 195 1492
rect 237 1488 243 1672
rect 253 1528 259 1952
rect 317 1928 323 2112
rect 317 1908 323 1912
rect 285 1748 291 1872
rect 349 1848 355 1876
rect 333 1748 339 1772
rect 333 1728 339 1732
rect 285 1563 291 1712
rect 333 1588 339 1612
rect 349 1563 355 1832
rect 365 1748 371 2072
rect 429 1908 435 2112
rect 493 1928 499 1952
rect 461 1908 467 1912
rect 408 1897 419 1903
rect 397 1888 403 1892
rect 381 1728 387 1732
rect 397 1588 403 1792
rect 413 1788 419 1897
rect 429 1848 435 1852
rect 461 1728 467 1772
rect 285 1557 307 1563
rect 141 1328 147 1332
rect 109 1317 120 1323
rect 29 1197 51 1203
rect 13 1068 19 1152
rect 45 1043 51 1197
rect 77 1108 83 1152
rect 93 1088 99 1092
rect 45 1037 67 1043
rect 61 928 67 1037
rect 77 948 83 972
rect 29 788 35 832
rect 61 708 67 912
rect 109 783 115 1317
rect 125 1088 131 1092
rect 141 1068 147 1312
rect 157 988 163 1292
rect 173 1188 179 1212
rect 221 1108 227 1272
rect 269 1128 275 1472
rect 285 1348 291 1352
rect 301 1348 307 1557
rect 333 1557 355 1563
rect 317 1408 323 1512
rect 333 1468 339 1557
rect 429 1488 435 1552
rect 333 1383 339 1432
rect 349 1428 355 1472
rect 477 1468 483 1732
rect 493 1728 499 1832
rect 509 1808 515 1892
rect 509 1728 515 1752
rect 525 1668 531 1672
rect 493 1508 499 1512
rect 333 1377 355 1383
rect 349 1368 355 1377
rect 285 1308 291 1332
rect 269 1103 275 1112
rect 253 1097 275 1103
rect 205 1008 211 1052
rect 125 968 131 972
rect 141 948 147 972
rect 205 948 211 952
rect 141 888 147 932
rect 157 928 163 932
rect 237 928 243 1092
rect 253 908 259 1097
rect 285 1068 291 1072
rect 317 1068 323 1092
rect 333 1088 339 1112
rect 349 1108 355 1332
rect 365 1088 371 1452
rect 445 1368 451 1452
rect 477 1443 483 1452
rect 509 1448 515 1632
rect 541 1568 547 2032
rect 557 1943 563 2132
rect 557 1937 579 1943
rect 557 1868 563 1912
rect 557 1748 563 1752
rect 573 1708 579 1937
rect 621 1888 627 2032
rect 637 1968 643 2092
rect 669 2068 675 2237
rect 717 2208 723 2232
rect 717 2168 723 2172
rect 733 2168 739 2297
rect 829 2288 835 2292
rect 765 2248 771 2272
rect 637 1908 643 1952
rect 589 1848 595 1872
rect 653 1868 659 1872
rect 685 1868 691 1912
rect 717 1908 723 2052
rect 733 2048 739 2152
rect 765 2128 771 2232
rect 813 2128 819 2192
rect 829 2148 835 2272
rect 733 1928 739 1932
rect 749 1928 755 1932
rect 845 1908 851 2412
rect 861 2268 867 2312
rect 941 2308 947 2463
rect 989 2288 995 2412
rect 1021 2348 1027 2392
rect 1021 2288 1027 2332
rect 1053 2292 1059 2312
rect 1133 2308 1139 2463
rect 1277 2408 1283 2463
rect 904 2277 915 2283
rect 877 1988 883 2072
rect 893 1948 899 1952
rect 909 1948 915 2277
rect 1005 2188 1011 2232
rect 941 1988 947 2152
rect 989 2028 995 2112
rect 1005 2048 1011 2132
rect 605 1828 611 1832
rect 621 1748 627 1852
rect 669 1848 675 1852
rect 669 1768 675 1772
rect 621 1663 627 1712
rect 637 1708 643 1732
rect 701 1728 707 1732
rect 717 1708 723 1832
rect 749 1788 755 1792
rect 829 1748 835 1872
rect 845 1808 851 1892
rect 893 1788 899 1912
rect 957 1828 963 1872
rect 605 1657 627 1663
rect 605 1588 611 1657
rect 525 1508 531 1532
rect 621 1508 627 1632
rect 637 1528 643 1692
rect 717 1688 723 1692
rect 541 1488 547 1492
rect 685 1488 691 1492
rect 733 1488 739 1512
rect 461 1437 483 1443
rect 461 1388 467 1437
rect 477 1348 483 1412
rect 493 1388 499 1432
rect 461 1308 467 1312
rect 493 1308 499 1332
rect 525 1328 531 1372
rect 541 1348 547 1452
rect 573 1388 579 1392
rect 589 1363 595 1432
rect 605 1428 611 1472
rect 573 1357 595 1363
rect 413 1288 419 1292
rect 397 1108 403 1132
rect 269 908 275 952
rect 104 777 115 783
rect 45 697 56 703
rect 45 643 51 697
rect 109 703 115 777
rect 237 728 243 892
rect 221 708 227 712
rect 109 697 120 703
rect 184 677 195 683
rect 157 648 163 672
rect 40 637 51 643
rect 13 528 19 532
rect 13 288 19 512
rect 13 268 19 272
rect 29 128 35 132
rect 45 128 51 637
rect 61 588 67 592
rect 77 508 83 512
rect 93 488 99 492
rect 141 488 147 512
rect 157 508 163 632
rect 173 528 179 532
rect 189 508 195 677
rect 205 668 211 692
rect 205 588 211 652
rect 237 588 243 712
rect 253 708 259 892
rect 285 788 291 992
rect 333 968 339 972
rect 365 968 371 1032
rect 301 888 307 892
rect 333 788 339 952
rect 285 748 291 772
rect 285 668 291 692
rect 264 657 275 663
rect 269 508 275 657
rect 349 608 355 712
rect 365 688 371 772
rect 381 688 387 1092
rect 413 1088 419 1112
rect 461 1088 467 1292
rect 493 1108 499 1112
rect 509 1108 515 1112
rect 525 1108 531 1112
rect 541 1108 547 1192
rect 456 1057 467 1063
rect 397 988 403 992
rect 461 948 467 1057
rect 509 1008 515 1072
rect 445 928 451 932
rect 397 728 403 732
rect 461 708 467 932
rect 445 668 451 672
rect 301 548 307 552
rect 317 528 323 572
rect 413 548 419 652
rect 461 608 467 652
rect 493 568 499 692
rect 541 588 547 1092
rect 557 988 563 1092
rect 573 1088 579 1357
rect 589 1188 595 1332
rect 621 1328 627 1452
rect 669 1448 675 1472
rect 653 1383 659 1432
rect 701 1388 707 1432
rect 653 1377 675 1383
rect 605 1308 611 1312
rect 653 1263 659 1352
rect 637 1257 659 1263
rect 637 1128 643 1257
rect 637 1088 643 1112
rect 653 1088 659 1232
rect 648 1057 659 1063
rect 637 988 643 1032
rect 557 928 563 952
rect 557 668 563 672
rect 360 537 371 543
rect 61 468 67 472
rect 93 308 99 472
rect 125 468 131 472
rect 77 288 83 292
rect 93 283 99 292
rect 93 277 104 283
rect 125 148 131 452
rect 157 308 163 492
rect 205 488 211 492
rect 189 308 195 312
rect 253 308 259 332
rect 237 288 243 292
rect 248 277 259 283
rect 205 248 211 272
rect 93 128 99 132
rect 173 128 179 132
rect 189 -43 195 92
rect 205 88 211 232
rect 221 128 227 252
rect 253 188 259 277
rect 269 108 275 492
rect 285 328 291 472
rect 301 328 307 472
rect 333 468 339 492
rect 349 388 355 512
rect 365 488 371 537
rect 445 508 451 512
rect 477 348 483 512
rect 493 388 499 552
rect 509 548 515 552
rect 509 508 515 532
rect 365 228 371 292
rect 429 268 435 292
rect 397 208 403 252
rect 365 188 371 192
rect 397 188 403 192
rect 557 188 563 512
rect 573 368 579 892
rect 589 788 595 872
rect 605 728 611 912
rect 621 703 627 812
rect 637 748 643 932
rect 653 868 659 1057
rect 669 1028 675 1377
rect 701 1348 707 1372
rect 717 1323 723 1392
rect 749 1388 755 1632
rect 829 1548 835 1652
rect 845 1548 851 1692
rect 861 1628 867 1672
rect 877 1648 883 1732
rect 925 1728 931 1792
rect 973 1788 979 1912
rect 989 1908 995 2012
rect 1021 1908 1027 2192
rect 1037 2128 1043 2272
rect 1053 2168 1059 2276
rect 1085 2123 1091 2232
rect 1101 2143 1107 2232
rect 1165 2188 1171 2312
rect 1213 2288 1219 2332
rect 1277 2328 1283 2392
rect 1101 2137 1112 2143
rect 1101 2128 1107 2137
rect 1133 2128 1139 2132
rect 1080 2117 1091 2123
rect 1085 2068 1091 2092
rect 1069 1928 1075 1992
rect 1101 1948 1107 2092
rect 1021 1868 1027 1872
rect 909 1708 915 1712
rect 877 1608 883 1632
rect 957 1628 963 1632
rect 973 1588 979 1772
rect 1021 1768 1027 1772
rect 1037 1743 1043 1872
rect 1085 1828 1091 1872
rect 1021 1737 1043 1743
rect 765 1488 771 1532
rect 733 1348 739 1352
rect 712 1317 723 1323
rect 701 1228 707 1232
rect 701 1128 707 1132
rect 717 1103 723 1232
rect 749 1108 755 1332
rect 797 1288 803 1432
rect 813 1408 819 1432
rect 861 1348 867 1512
rect 877 1488 883 1492
rect 925 1488 931 1512
rect 957 1488 963 1512
rect 877 1388 883 1452
rect 813 1328 819 1332
rect 893 1328 899 1472
rect 973 1468 979 1532
rect 1021 1508 1027 1737
rect 1037 1708 1043 1712
rect 1053 1588 1059 1732
rect 1069 1628 1075 1732
rect 1085 1728 1091 1792
rect 1069 1528 1075 1592
rect 1005 1488 1011 1492
rect 909 1428 915 1432
rect 941 1368 947 1432
rect 1005 1388 1011 1392
rect 941 1328 947 1352
rect 973 1348 979 1352
rect 893 1288 899 1292
rect 797 1108 803 1112
rect 701 1097 723 1103
rect 669 968 675 972
rect 685 968 691 1032
rect 701 928 707 1097
rect 749 1068 755 1072
rect 717 908 723 1052
rect 749 908 755 952
rect 797 948 803 1032
rect 861 1023 867 1072
rect 877 1048 883 1092
rect 893 1088 899 1172
rect 909 1068 915 1312
rect 957 1308 963 1332
rect 1021 1308 1027 1312
rect 925 1288 931 1292
rect 1037 1268 1043 1292
rect 1037 1248 1043 1252
rect 941 1088 947 1232
rect 957 1117 995 1123
rect 957 1108 963 1117
rect 989 1108 995 1117
rect 1037 1088 1043 1092
rect 1069 1088 1075 1332
rect 1085 1168 1091 1432
rect 1101 1408 1107 1892
rect 1133 1888 1139 2112
rect 1165 1848 1171 2092
rect 1181 1928 1187 2272
rect 1261 2148 1267 2272
rect 1309 2268 1315 2272
rect 1325 2243 1331 2312
rect 1389 2308 1395 2312
rect 1453 2308 1459 2392
rect 1501 2308 1507 2463
rect 1565 2328 1571 2463
rect 1629 2348 1635 2463
rect 1693 2408 1699 2463
rect 1805 2428 1811 2463
rect 1613 2328 1619 2332
rect 1693 2328 1699 2392
rect 1805 2328 1811 2412
rect 1741 2308 1747 2312
rect 1309 2237 1331 2243
rect 1277 2128 1283 2132
rect 1213 1908 1219 2032
rect 1245 1968 1251 2112
rect 1277 1988 1283 2112
rect 1277 1908 1283 1912
rect 1213 1883 1219 1892
rect 1197 1877 1219 1883
rect 1133 1728 1139 1792
rect 1181 1788 1187 1852
rect 1197 1728 1203 1877
rect 1229 1868 1235 1872
rect 1229 1748 1235 1832
rect 1213 1648 1219 1692
rect 1117 1548 1123 1632
rect 1101 1348 1107 1352
rect 1117 1348 1123 1492
rect 1133 1488 1139 1492
rect 1149 1488 1155 1552
rect 1133 1468 1139 1472
rect 1165 1468 1171 1532
rect 1181 1528 1187 1632
rect 1197 1528 1203 1532
rect 1149 1368 1155 1432
rect 1165 1308 1171 1412
rect 1149 1288 1155 1292
rect 1181 1268 1187 1512
rect 1213 1428 1219 1632
rect 1245 1608 1251 1872
rect 1293 1788 1299 2232
rect 1309 2188 1315 2237
rect 1341 2208 1347 2272
rect 1421 2248 1427 2272
rect 1389 2128 1395 2232
rect 1453 2228 1459 2292
rect 1501 2288 1507 2292
rect 1533 2208 1539 2232
rect 1405 2128 1411 2152
rect 1453 2128 1459 2132
rect 1309 2108 1315 2112
rect 1469 2108 1475 2112
rect 1501 2103 1507 2192
rect 1517 2128 1523 2172
rect 1549 2168 1555 2272
rect 1581 2228 1587 2272
rect 1613 2208 1619 2232
rect 1629 2188 1635 2232
rect 1773 2228 1779 2232
rect 1533 2148 1539 2152
rect 1496 2097 1507 2103
rect 1309 2068 1315 2092
rect 1549 2088 1555 2152
rect 1597 2103 1603 2172
rect 1645 2148 1651 2152
rect 1677 2148 1683 2152
rect 1693 2108 1699 2192
rect 1741 2143 1747 2212
rect 1837 2188 1843 2312
rect 1869 2288 1875 2292
rect 1869 2268 1875 2272
rect 1773 2168 1779 2172
rect 1837 2148 1843 2152
rect 1741 2137 1752 2143
rect 1592 2097 1603 2103
rect 1740 2097 1747 2103
rect 1741 2088 1747 2097
rect 1421 2008 1427 2032
rect 1309 1883 1315 1932
rect 1357 1908 1363 1912
rect 1421 1908 1427 1992
rect 1469 1948 1475 1952
rect 1309 1877 1331 1883
rect 1325 1868 1331 1877
rect 1357 1868 1363 1892
rect 1373 1868 1379 1872
rect 1293 1668 1299 1712
rect 1325 1708 1331 1712
rect 1341 1708 1347 1732
rect 1357 1708 1363 1772
rect 1421 1728 1427 1792
rect 1437 1708 1443 1872
rect 1373 1668 1379 1692
rect 1357 1608 1363 1632
rect 1309 1528 1315 1552
rect 1373 1508 1379 1652
rect 1453 1568 1459 1632
rect 1469 1508 1475 1812
rect 1485 1548 1491 1892
rect 1501 1868 1507 1912
rect 1517 1688 1523 1912
rect 1533 1768 1539 1952
rect 1533 1708 1539 1752
rect 1565 1748 1571 1852
rect 1581 1828 1587 1892
rect 1565 1648 1571 1732
rect 1613 1728 1619 1852
rect 1629 1748 1635 1992
rect 1725 1923 1731 2072
rect 1741 2068 1747 2072
rect 1725 1917 1736 1923
rect 1757 1888 1763 2132
rect 1773 1888 1779 2132
rect 1837 2008 1843 2132
rect 1853 2008 1859 2232
rect 1917 2168 1923 2332
rect 2141 2328 2147 2463
rect 1933 2308 1939 2312
rect 1997 2308 2003 2312
rect 2077 2308 2083 2312
rect 2141 2308 2147 2312
rect 2221 2308 2227 2463
rect 2589 2308 2595 2463
rect 3277 2388 3283 2463
rect 3373 2388 3379 2463
rect 3485 2388 3491 2463
rect 1965 2288 1971 2292
rect 2221 2283 2227 2292
rect 2269 2288 2275 2292
rect 2429 2288 2435 2292
rect 2205 2277 2227 2283
rect 1965 2148 1971 2272
rect 1981 2148 1987 2252
rect 1997 2148 2003 2192
rect 2045 2168 2051 2232
rect 2045 2148 2051 2152
rect 2109 2148 2115 2232
rect 2125 2128 2131 2212
rect 1869 2108 1875 2112
rect 2029 2108 2035 2112
rect 1821 1908 1827 1912
rect 1661 1728 1667 1732
rect 1677 1728 1683 1832
rect 1693 1748 1699 1752
rect 1709 1728 1715 1732
rect 1757 1728 1763 1832
rect 1581 1688 1587 1692
rect 1645 1608 1651 1692
rect 1725 1668 1731 1712
rect 1821 1568 1827 1732
rect 1837 1728 1843 1732
rect 1229 1428 1235 1492
rect 1245 1488 1251 1492
rect 1341 1488 1347 1492
rect 1384 1477 1395 1483
rect 1197 1328 1203 1352
rect 1229 1348 1235 1352
rect 1261 1348 1267 1472
rect 1293 1388 1299 1392
rect 1293 1348 1299 1372
rect 1325 1368 1331 1392
rect 1357 1388 1363 1392
rect 1389 1368 1395 1477
rect 1437 1448 1443 1492
rect 1485 1483 1491 1532
rect 1565 1488 1571 1552
rect 1469 1477 1491 1483
rect 1469 1468 1475 1477
rect 1501 1463 1507 1472
rect 1496 1457 1507 1463
rect 1341 1348 1347 1352
rect 973 1068 979 1072
rect 861 1017 883 1023
rect 877 948 883 1017
rect 925 1008 931 1032
rect 1037 983 1043 1032
rect 1069 1028 1075 1072
rect 1021 977 1043 983
rect 813 908 819 932
rect 973 928 979 932
rect 1021 928 1027 977
rect 909 908 915 912
rect 1021 908 1027 912
rect 653 828 659 832
rect 669 728 675 732
rect 653 708 659 712
rect 669 708 675 712
rect 605 697 627 703
rect 605 668 611 697
rect 589 628 595 632
rect 589 548 595 592
rect 589 308 595 472
rect 621 388 627 492
rect 637 448 643 552
rect 685 548 691 832
rect 701 788 707 792
rect 717 608 723 672
rect 733 588 739 832
rect 845 788 851 832
rect 845 748 851 772
rect 877 728 883 812
rect 909 748 915 772
rect 925 748 931 832
rect 941 737 952 743
rect 941 728 947 737
rect 781 708 787 712
rect 696 537 707 543
rect 701 528 707 537
rect 749 528 755 612
rect 893 588 899 692
rect 957 668 963 672
rect 973 668 979 892
rect 989 888 995 892
rect 1085 888 1091 1052
rect 1101 968 1107 1032
rect 1053 708 1059 852
rect 1101 808 1107 912
rect 1101 728 1107 772
rect 1117 708 1123 1232
rect 1149 1188 1155 1212
rect 1261 1208 1267 1332
rect 1357 1328 1363 1352
rect 1405 1348 1411 1372
rect 1421 1363 1427 1432
rect 1533 1388 1539 1452
rect 1421 1357 1443 1363
rect 1437 1328 1443 1357
rect 1549 1348 1555 1432
rect 1597 1408 1603 1472
rect 1613 1348 1619 1432
rect 1629 1408 1635 1512
rect 1709 1503 1715 1532
rect 1725 1528 1731 1532
rect 1789 1528 1795 1532
rect 1709 1497 1720 1503
rect 1645 1448 1651 1452
rect 1645 1388 1651 1412
rect 1565 1328 1571 1332
rect 1325 1308 1331 1312
rect 1229 1108 1235 1132
rect 1229 1088 1235 1092
rect 1261 1088 1267 1192
rect 1325 1188 1331 1292
rect 1389 1188 1395 1312
rect 1485 1308 1491 1312
rect 1453 1297 1464 1303
rect 1453 1188 1459 1297
rect 1325 1108 1331 1172
rect 1069 688 1075 692
rect 1133 688 1139 832
rect 1149 788 1155 952
rect 1181 928 1187 932
rect 1197 928 1203 1032
rect 1229 908 1235 932
rect 1261 928 1267 1052
rect 1277 948 1283 992
rect 1245 903 1251 912
rect 1277 908 1283 932
rect 1245 897 1267 903
rect 1213 883 1219 892
rect 1261 883 1267 897
rect 1293 883 1299 892
rect 1213 877 1235 883
rect 1261 877 1299 883
rect 1213 688 1219 852
rect 1229 688 1235 877
rect 1357 883 1363 1152
rect 1421 1137 1432 1143
rect 1421 1048 1427 1137
rect 1469 1128 1475 1132
rect 1453 928 1459 1072
rect 1469 1008 1475 1112
rect 1485 1108 1491 1292
rect 1613 1283 1619 1332
rect 1597 1277 1619 1283
rect 1597 1148 1603 1277
rect 1613 1108 1619 1252
rect 1485 968 1491 1072
rect 1517 968 1523 1052
rect 1549 1028 1555 1072
rect 1629 1068 1635 1332
rect 1549 928 1555 1012
rect 1645 988 1651 1292
rect 1661 1088 1667 1472
rect 1693 1448 1699 1492
rect 1837 1488 1843 1492
rect 1709 1468 1715 1472
rect 1725 1328 1731 1392
rect 1757 1388 1763 1452
rect 1741 1328 1747 1332
rect 1789 1328 1795 1332
rect 1677 1248 1683 1312
rect 1693 1188 1699 1232
rect 1693 1103 1699 1172
rect 1688 1097 1699 1103
rect 1709 1068 1715 1272
rect 1757 1248 1763 1292
rect 1789 1208 1795 1292
rect 1789 1188 1795 1192
rect 1661 988 1667 992
rect 1565 948 1571 952
rect 1629 948 1635 952
rect 1581 908 1587 912
rect 1405 888 1411 892
rect 1357 877 1368 883
rect 1325 868 1331 872
rect 1261 708 1267 712
rect 1357 708 1363 772
rect 1229 668 1235 672
rect 797 548 803 572
rect 909 568 915 612
rect 925 548 931 552
rect 653 463 659 512
rect 685 488 691 512
rect 765 503 771 512
rect 732 497 771 503
rect 701 463 707 492
rect 781 488 787 532
rect 845 528 851 532
rect 989 528 995 632
rect 1005 548 1011 652
rect 1101 588 1107 632
rect 1165 583 1171 652
rect 1160 577 1171 583
rect 1037 548 1043 572
rect 1085 528 1091 532
rect 1197 528 1203 572
rect 1213 548 1219 632
rect 1277 608 1283 692
rect 1293 668 1299 672
rect 1325 588 1331 652
rect 1229 548 1235 572
rect 1341 548 1347 672
rect 1373 668 1379 692
rect 1389 688 1395 852
rect 1421 828 1427 892
rect 1613 868 1619 892
rect 1661 868 1667 892
rect 1464 717 1512 723
rect 1549 708 1555 832
rect 1501 697 1512 703
rect 1389 588 1395 672
rect 1357 568 1363 572
rect 829 503 835 512
rect 829 497 840 503
rect 653 457 707 463
rect 685 388 691 432
rect 605 268 611 332
rect 589 257 600 263
rect 589 148 595 257
rect 621 188 627 212
rect 333 68 339 112
rect 589 -43 595 132
rect 621 28 627 72
rect 637 28 643 292
rect 717 188 723 232
rect 797 128 803 292
rect 845 288 851 472
rect 861 468 867 512
rect 957 508 963 512
rect 1117 508 1123 512
rect 1165 508 1171 512
rect 1005 497 1016 503
rect 973 308 979 472
rect 925 257 936 263
rect 893 128 899 192
rect 925 188 931 257
rect 973 188 979 292
rect 989 288 995 292
rect 1005 148 1011 497
rect 1069 497 1080 503
rect 1021 268 1027 412
rect 1069 388 1075 497
rect 1213 503 1219 512
rect 1309 508 1315 512
rect 1208 497 1219 503
rect 1101 288 1107 292
rect 1117 288 1123 292
rect 1101 248 1107 272
rect 653 -43 659 12
rect 749 -37 755 112
rect 957 108 963 112
rect 1021 108 1027 112
rect 957 -37 963 92
rect 989 68 995 92
rect 1037 48 1043 132
rect 1053 128 1059 232
rect 1117 228 1123 272
rect 1101 168 1107 172
rect 1133 148 1139 452
rect 1149 448 1155 492
rect 1197 388 1203 392
rect 1261 388 1267 492
rect 1277 408 1283 492
rect 1293 468 1299 492
rect 1357 428 1363 552
rect 1389 528 1395 532
rect 1405 528 1411 692
rect 1485 688 1491 692
rect 1501 688 1507 697
rect 1453 568 1459 652
rect 1469 548 1475 672
rect 1549 668 1555 692
rect 1565 688 1571 792
rect 1581 788 1587 812
rect 1661 748 1667 852
rect 1677 828 1683 1052
rect 1757 988 1763 1072
rect 1821 1068 1827 1332
rect 1837 1208 1843 1472
rect 1853 1108 1859 1872
rect 1869 1848 1875 1852
rect 1869 1748 1875 1792
rect 1885 1788 1891 2092
rect 1901 1928 1907 1952
rect 1869 1548 1875 1732
rect 1917 1728 1923 2072
rect 2045 1988 2051 2092
rect 1949 1888 1955 1932
rect 1997 1928 2003 1932
rect 2061 1923 2067 2112
rect 2189 2108 2195 2112
rect 2077 1948 2083 2072
rect 2189 2068 2195 2092
rect 2061 1917 2083 1923
rect 1949 1868 1955 1872
rect 1965 1743 1971 1872
rect 1997 1828 2003 1832
rect 2045 1788 2051 1892
rect 1960 1737 1971 1743
rect 1981 1743 1987 1752
rect 2061 1748 2067 1872
rect 2077 1828 2083 1917
rect 2109 1888 2115 1952
rect 2205 1948 2211 2277
rect 2397 2248 2403 2252
rect 2221 2188 2227 2192
rect 2253 2128 2259 2132
rect 2317 2128 2323 2232
rect 2381 2168 2387 2172
rect 2397 2148 2403 2232
rect 2445 2148 2451 2232
rect 2221 2108 2227 2112
rect 2285 1948 2291 2032
rect 2301 1988 2307 2032
rect 2397 1988 2403 2072
rect 2413 1968 2419 2132
rect 2461 2128 2467 2152
rect 2429 2008 2435 2032
rect 2493 2008 2499 2032
rect 2493 1988 2499 1992
rect 2317 1928 2323 1932
rect 2125 1888 2131 1892
rect 2104 1857 2115 1863
rect 2109 1748 2115 1857
rect 2173 1748 2179 1752
rect 1981 1737 2019 1743
rect 1885 1708 1891 1712
rect 1997 1708 2003 1712
rect 2013 1708 2019 1737
rect 2109 1728 2115 1732
rect 2029 1703 2035 1712
rect 2221 1708 2227 1712
rect 2029 1697 2072 1703
rect 1885 1528 1891 1672
rect 1901 1548 1907 1612
rect 1885 1463 1891 1492
rect 1901 1468 1907 1532
rect 1869 1457 1891 1463
rect 1869 1368 1875 1457
rect 1885 1428 1891 1432
rect 1885 1348 1891 1352
rect 1901 1348 1907 1392
rect 1949 1383 1955 1492
rect 1965 1488 1971 1652
rect 2013 1528 2019 1652
rect 2141 1648 2147 1672
rect 1965 1408 1971 1472
rect 1981 1468 1987 1492
rect 2029 1488 2035 1632
rect 2045 1508 2051 1632
rect 2061 1508 2067 1552
rect 1997 1448 2003 1472
rect 1944 1377 1955 1383
rect 1997 1368 2003 1412
rect 1933 1308 1939 1312
rect 1949 1308 1955 1332
rect 1869 1208 1875 1212
rect 1837 1097 1848 1103
rect 1837 988 1843 1097
rect 1869 1088 1875 1192
rect 1853 988 1859 1012
rect 1725 928 1731 972
rect 1773 968 1779 972
rect 1789 948 1795 972
rect 1885 948 1891 1192
rect 1901 1188 1907 1232
rect 1965 1188 1971 1312
rect 1997 1208 2003 1352
rect 2029 1348 2035 1472
rect 2045 1368 2051 1492
rect 2093 1488 2099 1512
rect 2109 1368 2115 1512
rect 2125 1488 2131 1492
rect 2141 1488 2147 1492
rect 2157 1488 2163 1612
rect 2205 1528 2211 1632
rect 2237 1608 2243 1712
rect 2253 1668 2259 1712
rect 2200 1497 2243 1503
rect 2221 1468 2227 1472
rect 2237 1468 2243 1497
rect 2205 1448 2211 1452
rect 2029 1328 2035 1332
rect 1917 1128 1923 1132
rect 2029 1123 2035 1232
rect 2045 1148 2051 1312
rect 2061 1308 2067 1352
rect 2109 1328 2115 1352
rect 2125 1348 2131 1432
rect 2157 1388 2163 1412
rect 2125 1268 2131 1312
rect 2141 1308 2147 1332
rect 2029 1117 2040 1123
rect 1917 963 1923 1092
rect 1933 1028 1939 1112
rect 1949 988 1955 1012
rect 1965 963 1971 1092
rect 2061 1088 2067 1112
rect 2077 1108 2083 1232
rect 1997 1068 2003 1072
rect 2045 968 2051 1012
rect 2093 968 2099 1092
rect 2109 1088 2115 1212
rect 2141 988 2147 1092
rect 1917 957 1939 963
rect 1933 948 1939 957
rect 1949 957 1971 963
rect 1741 928 1747 932
rect 1917 928 1923 932
rect 1885 917 1896 923
rect 1693 908 1699 912
rect 1613 728 1619 732
rect 1613 688 1619 712
rect 1565 668 1571 672
rect 1629 663 1635 712
rect 1677 668 1683 752
rect 1709 708 1715 732
rect 1725 708 1731 852
rect 1821 788 1827 812
rect 1821 708 1827 772
rect 1613 657 1635 663
rect 1373 508 1379 512
rect 1149 268 1155 352
rect 1149 228 1155 252
rect 1165 168 1171 352
rect 1213 288 1219 352
rect 1293 288 1299 372
rect 1277 188 1283 192
rect 1165 148 1171 152
rect 1197 148 1203 152
rect 1325 148 1331 392
rect 1389 388 1395 512
rect 1405 368 1411 512
rect 1469 488 1475 532
rect 1517 388 1523 512
rect 1533 508 1539 612
rect 1549 588 1555 612
rect 1613 548 1619 657
rect 1629 588 1635 632
rect 1581 468 1587 512
rect 1597 388 1603 492
rect 1501 308 1507 312
rect 1565 308 1571 312
rect 1613 308 1619 532
rect 1661 528 1667 652
rect 1709 568 1715 572
rect 1725 548 1731 692
rect 1741 588 1747 692
rect 1837 588 1843 892
rect 1741 568 1747 572
rect 1677 488 1683 492
rect 1149 128 1155 132
rect 1245 128 1251 132
rect 1261 128 1267 132
rect 1213 88 1219 92
rect 749 -43 771 -37
rect 941 -43 963 -37
rect 1229 -43 1235 12
rect 1309 -43 1315 112
rect 1325 28 1331 132
rect 1341 128 1347 152
rect 1357 128 1363 272
rect 1373 268 1379 292
rect 1469 268 1475 292
rect 1533 288 1539 292
rect 1549 263 1555 272
rect 1629 268 1635 432
rect 1741 408 1747 552
rect 1757 368 1763 432
rect 1645 308 1651 332
rect 1661 288 1667 292
rect 1773 288 1779 492
rect 1533 257 1555 263
rect 1405 168 1411 192
rect 1437 168 1443 232
rect 1533 188 1539 257
rect 1549 168 1555 232
rect 1613 188 1619 252
rect 1469 128 1475 152
rect 1613 148 1619 152
rect 1677 148 1683 192
rect 1533 128 1539 132
rect 1661 128 1667 132
rect 1629 88 1635 92
rect 1373 -43 1379 12
rect 1469 -43 1475 12
rect 1533 -43 1539 12
rect 1661 -43 1667 112
rect 1677 28 1683 132
rect 1725 128 1731 172
rect 1757 148 1763 212
rect 1773 208 1779 272
rect 1821 268 1827 552
rect 1837 488 1843 532
rect 1853 528 1859 892
rect 1869 588 1875 692
rect 1885 648 1891 917
rect 1901 908 1907 912
rect 1901 788 1907 812
rect 1917 748 1923 852
rect 1949 788 1955 957
rect 2029 948 2035 952
rect 2013 908 2019 912
rect 1992 897 2003 903
rect 1933 708 1939 732
rect 1901 428 1907 432
rect 1837 188 1843 392
rect 1853 308 1859 312
rect 1869 288 1875 292
rect 1885 288 1891 292
rect 1901 288 1907 332
rect 1917 308 1923 332
rect 1933 228 1939 692
rect 1949 508 1955 692
rect 1965 668 1971 892
rect 1997 788 2003 897
rect 2045 748 2051 912
rect 2125 888 2131 892
rect 2157 868 2163 1372
rect 2173 1163 2179 1432
rect 2189 1348 2195 1412
rect 2253 1388 2259 1632
rect 2269 1628 2275 1872
rect 2301 1788 2307 1892
rect 2429 1848 2435 1852
rect 2509 1808 2515 2232
rect 2637 2228 2643 2232
rect 2669 2168 2675 2292
rect 2525 2128 2531 2152
rect 2685 2148 2691 2172
rect 2701 2168 2707 2232
rect 2765 2148 2771 2232
rect 2813 2168 2819 2172
rect 2781 2148 2787 2152
rect 2557 2128 2563 2132
rect 2637 2128 2643 2132
rect 2573 2083 2579 2092
rect 2557 2077 2579 2083
rect 2525 1848 2531 1872
rect 2557 1868 2563 2077
rect 2589 2028 2595 2092
rect 2653 2008 2659 2132
rect 2669 2128 2675 2132
rect 2669 2048 2675 2112
rect 2765 2108 2771 2132
rect 2792 2117 2808 2123
rect 2653 1948 2659 1992
rect 2621 1928 2627 1932
rect 2541 1848 2547 1852
rect 2605 1748 2611 1892
rect 2621 1888 2627 1912
rect 2680 1897 2691 1903
rect 2653 1748 2659 1852
rect 2669 1748 2675 1752
rect 2632 1737 2643 1743
rect 2333 1728 2339 1732
rect 2301 1648 2307 1692
rect 2317 1488 2323 1512
rect 2333 1508 2339 1712
rect 2349 1648 2355 1712
rect 2381 1628 2387 1632
rect 2349 1588 2355 1612
rect 2413 1568 2419 1732
rect 2525 1668 2531 1732
rect 2557 1703 2563 1732
rect 2605 1728 2611 1732
rect 2621 1703 2627 1712
rect 2557 1697 2627 1703
rect 2637 1683 2643 1737
rect 2632 1677 2643 1683
rect 2285 1468 2291 1472
rect 2349 1428 2355 1492
rect 2461 1488 2467 1552
rect 2605 1543 2611 1672
rect 2589 1537 2611 1543
rect 2589 1528 2595 1537
rect 2653 1528 2659 1712
rect 2493 1488 2499 1512
rect 2557 1488 2563 1512
rect 2573 1488 2579 1512
rect 2333 1388 2339 1412
rect 2397 1408 2403 1432
rect 2445 1388 2451 1472
rect 2541 1388 2547 1472
rect 2205 1328 2211 1332
rect 2221 1328 2227 1372
rect 2269 1308 2275 1312
rect 2301 1308 2307 1312
rect 2333 1188 2339 1292
rect 2173 1157 2195 1163
rect 2173 1128 2179 1132
rect 2189 1108 2195 1157
rect 2205 1068 2211 1132
rect 2349 1128 2355 1332
rect 2365 1328 2371 1372
rect 2397 1348 2403 1352
rect 2509 1328 2515 1332
rect 2397 1308 2403 1312
rect 2477 1308 2483 1312
rect 2493 1308 2499 1312
rect 2525 1308 2531 1352
rect 2557 1348 2563 1452
rect 2605 1448 2611 1492
rect 2621 1488 2627 1512
rect 2685 1508 2691 1897
rect 2701 1888 2707 2092
rect 2829 2048 2835 2232
rect 2893 2188 2899 2272
rect 2925 2188 2931 2312
rect 3565 2308 3571 2312
rect 3229 2297 3240 2303
rect 2973 2288 2979 2292
rect 3005 2208 3011 2292
rect 2845 2157 2899 2163
rect 2845 2148 2851 2157
rect 2893 2148 2899 2157
rect 2989 2148 2995 2172
rect 2973 2128 2979 2132
rect 2925 2068 2931 2092
rect 2717 1868 2723 2032
rect 2957 2028 2963 2112
rect 2765 1928 2771 2012
rect 2797 1888 2803 1892
rect 2893 1888 2899 1912
rect 2909 1888 2915 1952
rect 2749 1868 2755 1872
rect 2733 1768 2739 1852
rect 2717 1508 2723 1712
rect 2733 1568 2739 1752
rect 2557 1328 2563 1332
rect 2573 1328 2579 1412
rect 2589 1348 2595 1392
rect 2621 1388 2627 1472
rect 2669 1468 2675 1492
rect 2605 1308 2611 1312
rect 2445 1208 2451 1292
rect 2413 1188 2419 1192
rect 2237 1088 2243 1092
rect 2221 948 2227 1072
rect 2269 1068 2275 1092
rect 2285 1088 2291 1092
rect 2221 928 2227 932
rect 2253 928 2259 952
rect 2301 928 2307 1052
rect 2333 948 2339 1072
rect 2349 968 2355 1092
rect 1981 728 1987 732
rect 2029 688 2035 712
rect 2093 688 2099 832
rect 1981 528 1987 652
rect 2061 588 2067 632
rect 2109 628 2115 632
rect 2029 528 2035 552
rect 1965 503 1971 512
rect 2045 508 2051 512
rect 2061 508 2067 512
rect 1965 497 1987 503
rect 1965 368 1971 432
rect 1981 323 1987 497
rect 2029 468 2035 492
rect 2077 488 2083 492
rect 1965 317 1987 323
rect 1901 148 1907 212
rect 1965 188 1971 317
rect 2029 308 2035 312
rect 2045 303 2051 352
rect 2093 308 2099 412
rect 2045 297 2056 303
rect 2077 288 2083 292
rect 1981 208 1987 252
rect 1997 228 2003 272
rect 1981 188 1987 192
rect 2013 188 2019 232
rect 2029 188 2035 192
rect 2045 168 2051 172
rect 1741 128 1747 132
rect 1885 108 1891 112
rect 1725 -43 1731 12
rect 1789 -43 1795 32
rect 1853 -43 1859 92
rect 1901 -37 1907 132
rect 1981 108 1987 152
rect 2093 148 2099 292
rect 2109 288 2115 492
rect 2125 308 2131 672
rect 2141 668 2147 752
rect 2189 708 2195 852
rect 2221 788 2227 912
rect 2301 888 2307 912
rect 2381 908 2387 1152
rect 2397 1028 2403 1132
rect 2509 1128 2515 1132
rect 2557 1128 2563 1152
rect 2589 1128 2595 1132
rect 2493 1108 2499 1112
rect 2413 1068 2419 1092
rect 2445 1068 2451 1092
rect 2541 1088 2547 1092
rect 2573 1068 2579 1092
rect 2461 948 2467 1032
rect 2621 1028 2627 1112
rect 2653 1088 2659 1312
rect 2669 1228 2675 1452
rect 2685 1348 2691 1452
rect 2701 1368 2707 1472
rect 2701 1268 2707 1332
rect 2733 1308 2739 1552
rect 2749 1508 2755 1852
rect 2797 1728 2803 1732
rect 2765 1508 2771 1712
rect 2813 1708 2819 1872
rect 2861 1868 2867 1872
rect 2877 1728 2883 1852
rect 2925 1728 2931 1752
rect 2845 1708 2851 1712
rect 2861 1688 2867 1712
rect 2749 1428 2755 1492
rect 2829 1468 2835 1492
rect 2797 1368 2803 1432
rect 2845 1348 2851 1532
rect 2861 1468 2867 1632
rect 2909 1503 2915 1632
rect 2904 1497 2915 1503
rect 2781 1317 2792 1323
rect 2717 1163 2723 1252
rect 2701 1157 2723 1163
rect 2701 1148 2707 1157
rect 2749 1148 2755 1292
rect 2669 1008 2675 1112
rect 2685 1108 2691 1132
rect 2765 1088 2771 1292
rect 2781 1108 2787 1317
rect 2813 1308 2819 1332
rect 2893 1308 2899 1432
rect 2909 1408 2915 1497
rect 2941 1488 2947 1632
rect 2925 1348 2931 1432
rect 2957 1428 2963 1492
rect 2973 1488 2979 1932
rect 3005 1908 3011 2032
rect 3021 1888 3027 1912
rect 3005 1548 3011 1872
rect 3037 1748 3043 2092
rect 3053 1928 3059 2272
rect 3069 2108 3075 2272
rect 3133 2168 3139 2292
rect 3229 2288 3235 2297
rect 3325 2297 3336 2303
rect 3293 2288 3299 2292
rect 3325 2288 3331 2297
rect 3197 2128 3203 2152
rect 3293 2128 3299 2232
rect 3405 2188 3411 2232
rect 3101 2108 3107 2112
rect 3053 1888 3059 1912
rect 3069 1888 3075 2092
rect 3117 1888 3123 1932
rect 3149 1908 3155 2012
rect 3133 1888 3139 1892
rect 3085 1808 3091 1812
rect 3053 1768 3059 1792
rect 3037 1728 3043 1732
rect 3037 1528 3043 1552
rect 2989 1448 2995 1492
rect 2973 1348 2979 1372
rect 3069 1348 3075 1792
rect 3085 1728 3091 1792
rect 3133 1788 3139 1872
rect 3165 1728 3171 1812
rect 3181 1788 3187 2012
rect 3197 1908 3203 1912
rect 3277 1888 3283 2112
rect 3309 1928 3315 2032
rect 3293 1908 3299 1912
rect 3229 1768 3235 1852
rect 3293 1788 3299 1832
rect 3245 1748 3251 1752
rect 3325 1748 3331 2172
rect 3437 2128 3443 2292
rect 3341 2108 3347 2112
rect 3341 1908 3347 2092
rect 3373 2088 3379 2112
rect 3373 2048 3379 2072
rect 3501 1988 3507 2292
rect 3421 1908 3427 1912
rect 3549 1908 3555 2292
rect 3565 2028 3571 2112
rect 3597 2028 3603 2032
rect 3581 1928 3587 1932
rect 3469 1888 3475 1892
rect 3341 1828 3347 1872
rect 3357 1848 3363 1872
rect 3437 1748 3443 1832
rect 3133 1708 3139 1712
rect 3149 1648 3155 1692
rect 3085 1488 3091 1632
rect 3117 1528 3123 1632
rect 3165 1628 3171 1632
rect 3101 1428 3107 1512
rect 3213 1508 3219 1632
rect 3261 1488 3267 1652
rect 3293 1528 3299 1632
rect 3325 1568 3331 1732
rect 3421 1728 3427 1732
rect 3357 1697 3368 1703
rect 3357 1588 3363 1697
rect 3389 1543 3395 1672
rect 3389 1537 3411 1543
rect 3373 1528 3379 1532
rect 3325 1477 3336 1483
rect 3165 1463 3171 1472
rect 3149 1457 3171 1463
rect 3133 1348 3139 1452
rect 3005 1328 3011 1332
rect 2925 1308 2931 1312
rect 2893 1208 2899 1292
rect 2909 1288 2915 1292
rect 3005 1268 3011 1292
rect 3085 1288 3091 1292
rect 2941 1248 2947 1252
rect 2925 1188 2931 1192
rect 2829 1088 2835 1172
rect 2893 1108 2899 1152
rect 2925 1128 2931 1172
rect 2941 1108 2947 1232
rect 3005 1128 3011 1192
rect 3053 1128 3059 1132
rect 2493 988 2499 992
rect 2557 948 2563 952
rect 2653 948 2659 992
rect 2685 988 2691 1032
rect 2733 948 2739 952
rect 2749 943 2755 1032
rect 2749 937 2760 943
rect 2717 928 2723 932
rect 2413 848 2419 912
rect 2557 903 2563 912
rect 2781 908 2787 952
rect 2797 908 2803 1032
rect 2813 908 2819 992
rect 2861 968 2867 1052
rect 2925 968 2931 1032
rect 2877 928 2883 932
rect 2541 897 2563 903
rect 2429 888 2435 892
rect 2541 888 2547 897
rect 2989 903 2995 1032
rect 3005 988 3011 1032
rect 3021 1028 3027 1072
rect 3053 948 3059 1112
rect 3085 1108 3091 1272
rect 3117 1188 3123 1232
rect 3133 1108 3139 1272
rect 3149 1188 3155 1457
rect 3325 1448 3331 1477
rect 3181 1328 3187 1352
rect 3213 1348 3219 1432
rect 3245 1348 3251 1352
rect 3213 1288 3219 1312
rect 3293 1288 3299 1332
rect 3309 1328 3315 1372
rect 3325 1368 3331 1432
rect 3373 1368 3379 1512
rect 3389 1468 3395 1512
rect 3389 1408 3395 1432
rect 3325 1303 3331 1332
rect 3389 1328 3395 1332
rect 3309 1297 3331 1303
rect 3181 1108 3187 1172
rect 3245 1168 3251 1272
rect 3101 943 3107 1032
rect 3085 937 3107 943
rect 3069 908 3075 932
rect 2989 897 3000 903
rect 2237 708 2243 712
rect 2301 708 2307 712
rect 2413 708 2419 732
rect 2429 708 2435 792
rect 2397 688 2403 692
rect 2141 648 2147 652
rect 2189 648 2195 652
rect 2205 608 2211 632
rect 2189 528 2195 572
rect 2205 548 2211 572
rect 2381 528 2387 632
rect 2413 528 2419 672
rect 2445 668 2451 832
rect 2493 688 2499 712
rect 2525 708 2531 712
rect 2541 708 2547 772
rect 2557 708 2563 732
rect 2637 728 2643 752
rect 2749 708 2755 832
rect 2797 788 2803 832
rect 2989 708 2995 772
rect 3005 728 3011 792
rect 3037 788 3043 792
rect 3069 748 3075 892
rect 3085 888 3091 937
rect 3117 928 3123 972
rect 3133 948 3139 1072
rect 3149 1048 3155 1092
rect 3213 1088 3219 1112
rect 3245 1068 3251 1152
rect 3261 1088 3267 1112
rect 3309 1108 3315 1297
rect 3405 1183 3411 1537
rect 3421 1508 3427 1712
rect 3437 1588 3443 1732
rect 3469 1608 3475 1632
rect 3453 1528 3459 1572
rect 3485 1548 3491 1892
rect 3549 1868 3555 1872
rect 3501 1728 3507 1832
rect 3517 1728 3523 1812
rect 3629 1808 3635 1892
rect 3645 1888 3651 2132
rect 3533 1728 3539 1732
rect 3629 1728 3635 1792
rect 3645 1748 3651 1872
rect 3469 1528 3475 1532
rect 3517 1508 3523 1712
rect 3581 1548 3587 1632
rect 3485 1468 3491 1492
rect 3517 1488 3523 1492
rect 3501 1448 3507 1472
rect 3421 1288 3427 1352
rect 3437 1348 3443 1352
rect 3453 1328 3459 1372
rect 3421 1268 3427 1272
rect 3400 1177 3411 1183
rect 3405 1108 3411 1132
rect 3437 1108 3443 1292
rect 3261 1043 3267 1072
rect 3245 1037 3267 1043
rect 3101 868 3107 912
rect 3149 868 3155 912
rect 3165 768 3171 1032
rect 3245 908 3251 1037
rect 3261 968 3267 1012
rect 3277 1008 3283 1032
rect 3309 988 3315 1092
rect 3341 1068 3347 1092
rect 3357 1068 3363 1072
rect 3341 948 3347 1052
rect 3373 1043 3379 1092
rect 3421 1088 3427 1092
rect 3437 1088 3443 1092
rect 3453 1088 3459 1092
rect 3469 1088 3475 1292
rect 3501 1288 3507 1332
rect 3517 1308 3523 1472
rect 3533 1368 3539 1472
rect 3549 1368 3555 1412
rect 3565 1388 3571 1432
rect 3581 1428 3587 1512
rect 3533 1308 3539 1312
rect 3549 1283 3555 1352
rect 3597 1288 3603 1292
rect 3533 1277 3555 1283
rect 3517 1188 3523 1272
rect 3517 1108 3523 1172
rect 3533 1108 3539 1277
rect 3613 1203 3619 1492
rect 3597 1197 3619 1203
rect 3565 1128 3571 1132
rect 3501 1088 3507 1092
rect 3357 1037 3379 1043
rect 3357 988 3363 1037
rect 3517 968 3523 1072
rect 3533 1028 3539 1092
rect 3533 988 3539 992
rect 3597 968 3603 1197
rect 3261 728 3267 812
rect 3005 708 3011 712
rect 2605 688 2611 692
rect 2733 688 2739 692
rect 2877 688 2883 692
rect 3069 688 3075 692
rect 2637 668 2643 672
rect 2477 588 2483 592
rect 2429 548 2435 552
rect 2173 508 2179 512
rect 2157 388 2163 492
rect 2221 448 2227 512
rect 2381 468 2387 472
rect 2125 148 2131 232
rect 2221 148 2227 292
rect 2253 148 2259 232
rect 2333 188 2339 232
rect 2365 188 2371 292
rect 2397 268 2403 432
rect 2397 188 2403 232
rect 2493 188 2499 272
rect 2061 128 2067 132
rect 2125 128 2131 132
rect 2157 123 2163 132
rect 2221 128 2227 132
rect 2285 128 2291 172
rect 2157 117 2168 123
rect 2317 123 2323 132
rect 2317 117 2328 123
rect 2413 123 2419 132
rect 2509 128 2515 512
rect 2589 488 2595 632
rect 2605 508 2611 652
rect 2621 568 2627 632
rect 2669 528 2675 632
rect 2685 548 2691 632
rect 2765 588 2771 632
rect 2813 548 2819 632
rect 2877 608 2883 672
rect 3181 668 3187 692
rect 3197 688 3203 692
rect 3309 688 3315 932
rect 3453 928 3459 932
rect 3389 848 3395 912
rect 3485 788 3491 832
rect 3517 828 3523 952
rect 3485 708 3491 772
rect 3357 688 3363 692
rect 3421 688 3427 692
rect 2957 568 2963 632
rect 2701 448 2707 512
rect 2589 308 2595 432
rect 2701 388 2707 432
rect 2765 388 2771 432
rect 2861 388 2867 432
rect 2893 388 2899 512
rect 2909 508 2915 532
rect 2989 528 2995 532
rect 3117 528 3123 532
rect 3229 488 3235 512
rect 2765 308 2771 372
rect 3261 308 3267 472
rect 3293 388 3299 472
rect 2541 188 2547 292
rect 2541 128 2547 172
rect 2621 148 2627 232
rect 2653 148 2659 292
rect 2717 148 2723 272
rect 2653 128 2659 132
rect 2717 128 2723 132
rect 2733 128 2739 232
rect 2765 148 2771 152
rect 2941 148 2947 292
rect 2749 128 2755 132
rect 2765 128 2771 132
rect 2909 128 2915 132
rect 2973 128 2979 232
rect 3117 188 3123 272
rect 3165 188 3171 232
rect 3229 188 3235 232
rect 2413 117 2424 123
rect 3005 123 3011 132
rect 3117 128 3123 172
rect 3181 128 3187 172
rect 3309 148 3315 672
rect 3373 528 3379 532
rect 3485 528 3491 532
rect 3357 488 3363 512
rect 3373 308 3379 472
rect 3485 388 3491 392
rect 3453 248 3459 292
rect 3405 188 3411 232
rect 3453 148 3459 232
rect 3005 117 3016 123
rect 3229 123 3235 132
rect 3341 128 3347 132
rect 3501 128 3507 232
rect 3517 128 3523 132
rect 3533 128 3539 952
rect 3549 928 3555 932
rect 3581 923 3587 932
rect 3581 917 3592 923
rect 3581 728 3587 732
rect 3549 688 3555 692
rect 3597 688 3603 772
rect 3613 548 3619 1092
rect 3661 928 3667 932
rect 3645 708 3651 772
rect 3549 528 3555 532
rect 3565 408 3571 432
rect 3549 297 3560 303
rect 3549 288 3555 297
rect 3581 148 3587 532
rect 3661 528 3667 532
rect 3661 328 3667 332
rect 3229 117 3240 123
rect 1901 -43 1923 -37
rect 2205 -43 2211 32
rect 2365 -43 2371 32
rect 2461 -43 2467 32
rect 2669 -43 2675 32
rect 2893 28 2899 32
rect 3053 28 3059 32
rect 2861 -43 2867 12
rect 3021 -43 3027 12
rect 3277 -43 3283 32
rect 3325 -37 3331 32
rect 3325 -43 3347 -37
<< m3contact >>
rect 8 2312 24 2328
rect 632 2312 648 2328
rect 765 2402 801 2418
rect 808 2412 824 2428
rect 840 2412 856 2428
rect 696 2332 712 2348
rect 232 2292 248 2308
rect 328 2292 344 2308
rect 392 2292 408 2308
rect 456 2292 472 2308
rect 552 2292 568 2308
rect 104 2132 120 2148
rect 136 2132 152 2148
rect 200 2132 216 2148
rect 8 2112 24 2128
rect 584 2272 600 2288
rect 552 2252 568 2268
rect 568 2152 584 2168
rect 680 2252 696 2268
rect 296 2112 312 2128
rect 312 2112 328 2128
rect 360 2112 376 2128
rect 408 2112 424 2128
rect 248 1952 264 1968
rect 216 1912 232 1928
rect 24 1892 40 1908
rect 72 1892 88 1908
rect 88 1892 104 1908
rect 136 1892 152 1908
rect 184 1892 200 1908
rect 200 1892 216 1908
rect 8 1712 24 1728
rect 88 1812 104 1828
rect 232 1672 248 1688
rect 88 1492 104 1508
rect 56 1432 72 1448
rect 168 1512 184 1528
rect 152 1492 168 1508
rect 120 1452 136 1468
rect 152 1452 168 1468
rect 184 1492 200 1508
rect 200 1492 216 1508
rect 360 2072 376 2088
rect 280 1912 296 1928
rect 312 1912 328 1928
rect 280 1872 296 1888
rect 328 1872 344 1888
rect 344 1832 360 1848
rect 328 1772 344 1788
rect 328 1732 344 1748
rect 280 1712 296 1728
rect 264 1692 280 1708
rect 296 1692 312 1708
rect 328 1692 344 1708
rect 328 1612 344 1628
rect 312 1572 328 1588
rect 376 1912 392 1928
rect 488 1952 504 1968
rect 456 1912 472 1928
rect 392 1872 408 1888
rect 392 1792 408 1808
rect 376 1732 392 1748
rect 424 1892 440 1908
rect 424 1832 440 1848
rect 456 1772 472 1788
rect 440 1732 456 1748
rect 424 1692 440 1708
rect 376 1572 392 1588
rect 248 1492 264 1508
rect 280 1492 296 1508
rect 232 1472 248 1488
rect 264 1472 280 1488
rect 216 1372 232 1388
rect 184 1352 200 1368
rect 136 1332 152 1348
rect 8 1152 24 1168
rect 24 1072 40 1088
rect 72 1192 88 1208
rect 72 1152 88 1168
rect 88 1072 104 1088
rect 56 1052 72 1068
rect 72 972 88 988
rect 88 944 104 948
rect 88 932 104 944
rect 136 1312 152 1328
rect 248 1312 264 1328
rect 120 1072 136 1088
rect 168 1212 184 1228
rect 312 1532 328 1548
rect 424 1552 440 1568
rect 456 1472 472 1488
rect 328 1452 344 1468
rect 312 1392 328 1408
rect 520 1872 536 1888
rect 504 1792 520 1808
rect 504 1752 520 1768
rect 520 1652 536 1668
rect 488 1492 504 1508
rect 376 1452 392 1468
rect 472 1452 488 1468
rect 344 1412 360 1428
rect 328 1352 344 1368
rect 280 1332 312 1348
rect 344 1332 360 1348
rect 280 1292 296 1308
rect 296 1232 312 1248
rect 248 1112 260 1128
rect 260 1112 264 1128
rect 328 1112 344 1128
rect 216 1092 232 1108
rect 232 1092 248 1108
rect 216 1072 232 1088
rect 200 992 216 1008
rect 136 972 168 988
rect 120 952 136 968
rect 200 952 216 968
rect 152 932 168 948
rect 184 932 200 948
rect 152 912 168 928
rect 216 912 232 928
rect 232 912 248 928
rect 280 1072 296 1088
rect 296 1072 312 1088
rect 344 1092 360 1108
rect 568 2112 584 2128
rect 632 2092 648 2108
rect 552 1912 568 1928
rect 552 1732 568 1748
rect 712 2192 728 2208
rect 712 2172 728 2188
rect 824 2272 840 2288
rect 760 2232 776 2248
rect 680 2152 696 2168
rect 728 2152 744 2168
rect 680 2132 696 2148
rect 680 2112 696 2128
rect 664 2052 680 2068
rect 712 2052 728 2068
rect 632 1952 648 1968
rect 696 1912 712 1928
rect 808 2192 824 2208
rect 824 2132 840 2148
rect 728 2032 744 2048
rect 765 2002 801 2018
rect 744 1932 760 1948
rect 728 1912 744 1928
rect 856 2312 872 2328
rect 984 2412 1000 2428
rect 904 2292 920 2308
rect 936 2292 952 2308
rect 968 2292 984 2308
rect 1016 2392 1032 2408
rect 1016 2332 1032 2348
rect 1048 2312 1064 2328
rect 1272 2392 1288 2408
rect 1448 2392 1464 2408
rect 1208 2332 1224 2348
rect 1128 2292 1144 2308
rect 856 2252 872 2268
rect 888 2112 904 2128
rect 856 2092 872 2108
rect 888 2032 904 2048
rect 888 1952 904 1968
rect 920 2272 936 2288
rect 984 2272 1000 2288
rect 936 2232 952 2248
rect 1016 2192 1032 2208
rect 1000 2172 1016 2188
rect 1000 2152 1016 2168
rect 952 2112 968 2128
rect 1000 2032 1016 2048
rect 984 2012 1000 2028
rect 888 1912 904 1928
rect 824 1872 840 1888
rect 616 1852 632 1868
rect 648 1852 664 1868
rect 680 1852 696 1868
rect 808 1852 824 1868
rect 584 1832 600 1848
rect 600 1812 616 1828
rect 664 1832 680 1848
rect 712 1832 728 1848
rect 664 1772 680 1788
rect 696 1732 712 1748
rect 600 1712 616 1728
rect 568 1692 584 1708
rect 552 1652 568 1668
rect 648 1712 664 1728
rect 744 1792 760 1808
rect 856 1872 872 1888
rect 840 1792 856 1808
rect 952 1872 968 1888
rect 952 1812 968 1828
rect 920 1792 936 1808
rect 840 1752 856 1768
rect 792 1732 808 1748
rect 824 1732 840 1748
rect 632 1692 648 1708
rect 680 1692 696 1708
rect 712 1692 728 1708
rect 744 1692 760 1708
rect 840 1692 856 1708
rect 616 1632 632 1648
rect 600 1572 616 1588
rect 536 1552 552 1568
rect 552 1512 568 1528
rect 824 1652 840 1668
rect 696 1632 712 1648
rect 744 1632 760 1648
rect 632 1512 648 1528
rect 728 1512 744 1528
rect 520 1492 536 1508
rect 536 1472 552 1488
rect 680 1472 696 1488
rect 536 1452 552 1468
rect 568 1452 584 1468
rect 504 1432 520 1448
rect 520 1432 536 1448
rect 472 1412 488 1428
rect 456 1372 472 1388
rect 440 1352 456 1368
rect 488 1372 504 1388
rect 520 1372 536 1388
rect 488 1352 504 1368
rect 440 1332 456 1348
rect 488 1332 504 1348
rect 568 1392 584 1408
rect 552 1352 568 1368
rect 616 1452 632 1468
rect 632 1452 648 1468
rect 600 1412 616 1428
rect 536 1332 552 1348
rect 456 1292 472 1308
rect 408 1272 424 1288
rect 392 1132 408 1148
rect 408 1112 424 1128
rect 312 1052 328 1068
rect 280 992 296 1008
rect 184 892 200 908
rect 216 892 232 908
rect 232 892 248 908
rect 264 892 280 908
rect 136 872 152 888
rect 216 712 232 728
rect 152 672 168 688
rect 8 512 24 528
rect 24 472 40 488
rect 24 292 40 308
rect 8 252 24 268
rect 56 592 72 608
rect 136 572 152 588
rect 72 492 88 508
rect 168 512 184 528
rect 200 652 216 668
rect 328 972 344 988
rect 344 952 360 968
rect 360 952 376 968
rect 296 892 312 908
rect 360 832 376 848
rect 328 772 344 788
rect 360 772 376 788
rect 280 732 296 748
rect 328 712 340 728
rect 340 712 344 728
rect 248 692 264 708
rect 296 672 312 688
rect 232 572 248 588
rect 248 512 264 528
rect 280 652 296 668
rect 536 1192 552 1208
rect 504 1112 520 1128
rect 488 1092 504 1108
rect 520 1092 536 1108
rect 392 1072 408 1088
rect 456 1072 472 1088
rect 392 992 408 1008
rect 504 992 520 1008
rect 472 944 488 948
rect 472 932 488 944
rect 440 912 456 928
rect 392 732 408 748
rect 504 892 520 908
rect 520 732 536 748
rect 456 692 472 708
rect 488 692 504 708
rect 504 692 520 708
rect 376 672 392 688
rect 424 672 440 688
rect 376 652 392 668
rect 408 652 424 668
rect 440 652 456 668
rect 344 592 360 608
rect 312 572 328 588
rect 296 532 312 548
rect 392 552 408 568
rect 456 592 472 608
rect 664 1432 680 1448
rect 712 1392 728 1408
rect 648 1352 664 1368
rect 616 1312 632 1328
rect 600 1292 616 1308
rect 632 1292 648 1308
rect 648 1232 664 1248
rect 632 1112 648 1128
rect 632 1032 648 1048
rect 552 952 568 968
rect 584 932 600 948
rect 632 932 648 948
rect 552 652 568 668
rect 536 572 552 588
rect 424 552 440 568
rect 488 552 504 568
rect 152 492 168 508
rect 168 492 184 508
rect 184 492 200 508
rect 264 492 280 508
rect 56 472 72 488
rect 88 472 104 488
rect 136 472 152 488
rect 56 452 72 468
rect 120 452 136 468
rect 104 332 120 348
rect 88 292 104 308
rect 104 292 120 308
rect 72 272 88 288
rect 72 252 88 268
rect 200 472 216 488
rect 232 472 248 488
rect 248 452 264 468
rect 248 332 264 348
rect 184 312 200 328
rect 152 292 168 308
rect 248 292 264 308
rect 168 272 184 288
rect 200 272 216 288
rect 216 252 232 268
rect 136 232 152 248
rect 200 232 216 248
rect 120 132 136 148
rect 168 132 184 148
rect 24 112 56 128
rect 88 112 104 128
rect 120 112 136 128
rect 184 92 200 108
rect 168 52 184 68
rect 216 112 232 128
rect 280 472 296 488
rect 328 452 344 468
rect 408 512 424 528
rect 472 512 488 528
rect 440 492 456 508
rect 360 472 376 488
rect 504 532 520 548
rect 520 512 536 528
rect 504 492 520 508
rect 440 332 456 348
rect 472 332 488 348
rect 296 312 312 328
rect 408 312 424 328
rect 280 292 296 308
rect 456 292 472 308
rect 536 292 552 308
rect 296 272 312 288
rect 280 252 296 268
rect 424 252 440 268
rect 360 212 376 228
rect 360 192 376 208
rect 392 192 408 208
rect 584 772 600 788
rect 616 812 632 828
rect 600 712 616 728
rect 696 1372 712 1388
rect 696 1332 712 1348
rect 765 1602 801 1618
rect 1144 2272 1160 2288
rect 1048 2152 1064 2168
rect 1032 2112 1048 2128
rect 1192 2292 1208 2308
rect 1224 2312 1240 2328
rect 1384 2312 1400 2328
rect 1208 2272 1224 2288
rect 1128 2132 1144 2148
rect 1096 2112 1112 2128
rect 1096 2092 1112 2108
rect 1080 2052 1096 2068
rect 1064 1992 1080 2008
rect 1096 1932 1112 1948
rect 984 1892 1000 1908
rect 1016 1872 1032 1888
rect 1016 1852 1032 1868
rect 968 1772 984 1788
rect 1016 1772 1032 1788
rect 904 1712 920 1728
rect 872 1632 888 1648
rect 856 1612 872 1628
rect 952 1612 968 1628
rect 872 1592 888 1608
rect 1048 1832 1064 1848
rect 1080 1812 1096 1828
rect 1080 1792 1096 1808
rect 1000 1712 1016 1728
rect 968 1572 984 1588
rect 760 1532 776 1548
rect 968 1532 984 1548
rect 856 1512 872 1528
rect 920 1512 936 1528
rect 728 1352 744 1368
rect 744 1332 760 1348
rect 680 1292 696 1308
rect 712 1292 728 1308
rect 712 1232 728 1248
rect 696 1212 712 1228
rect 696 1132 712 1148
rect 808 1392 824 1408
rect 872 1492 888 1508
rect 952 1472 968 1488
rect 872 1452 888 1468
rect 808 1332 824 1348
rect 856 1332 872 1348
rect 1048 1732 1064 1748
rect 1032 1712 1048 1728
rect 1064 1612 1080 1628
rect 1064 1592 1080 1608
rect 1048 1572 1064 1588
rect 1016 1492 1032 1508
rect 1000 1472 1016 1488
rect 904 1412 920 1428
rect 1000 1392 1016 1408
rect 936 1352 952 1368
rect 968 1352 984 1368
rect 952 1332 968 1348
rect 888 1312 920 1328
rect 888 1272 904 1288
rect 808 1232 824 1248
rect 765 1202 801 1218
rect 888 1172 904 1188
rect 840 1112 856 1128
rect 664 1012 680 1028
rect 664 972 680 988
rect 680 952 696 968
rect 792 1092 808 1108
rect 760 1072 776 1088
rect 712 1052 728 1068
rect 744 1052 760 1068
rect 744 952 760 968
rect 888 1072 904 1088
rect 1016 1312 1032 1328
rect 920 1292 936 1308
rect 1000 1292 1016 1308
rect 1032 1252 1048 1268
rect 1032 1232 1048 1248
rect 968 1092 984 1108
rect 984 1092 1000 1108
rect 1144 1912 1160 1928
rect 1128 1872 1144 1888
rect 1240 2252 1256 2268
rect 1304 2252 1320 2268
rect 1464 2312 1480 2328
rect 1800 2412 1816 2428
rect 1688 2392 1704 2408
rect 1608 2332 1640 2348
rect 1912 2332 1928 2348
rect 1528 2312 1544 2328
rect 1560 2312 1576 2328
rect 1624 2312 1640 2328
rect 1688 2312 1704 2328
rect 1736 2312 1752 2328
rect 1512 2292 1528 2308
rect 1368 2272 1384 2288
rect 1256 2132 1272 2148
rect 1192 2112 1208 2128
rect 1176 1912 1192 1928
rect 1272 1972 1288 1988
rect 1240 1952 1256 1968
rect 1272 1912 1288 1928
rect 1176 1852 1192 1868
rect 1144 1832 1176 1848
rect 1128 1792 1144 1808
rect 1208 1852 1224 1868
rect 1224 1852 1240 1868
rect 1224 1732 1240 1748
rect 1192 1712 1208 1728
rect 1224 1712 1240 1728
rect 1208 1632 1224 1648
rect 1144 1552 1160 1568
rect 1112 1532 1128 1548
rect 1112 1492 1128 1508
rect 1096 1392 1112 1408
rect 1160 1532 1176 1548
rect 1128 1472 1144 1488
rect 1192 1532 1208 1548
rect 1176 1512 1192 1528
rect 1128 1452 1144 1468
rect 1160 1412 1176 1428
rect 1144 1352 1160 1368
rect 1096 1332 1112 1348
rect 1112 1332 1128 1348
rect 1096 1312 1112 1328
rect 1144 1272 1160 1288
rect 1192 1492 1208 1508
rect 1416 2232 1432 2248
rect 1336 2192 1352 2208
rect 1304 2132 1320 2148
rect 1496 2272 1512 2288
rect 1544 2272 1560 2288
rect 1656 2272 1672 2288
rect 1448 2212 1464 2228
rect 1496 2192 1512 2208
rect 1528 2192 1544 2208
rect 1400 2152 1416 2168
rect 1448 2132 1464 2148
rect 1480 2132 1496 2148
rect 1448 2112 1464 2128
rect 1352 2092 1364 2108
rect 1364 2092 1368 2108
rect 1464 2092 1480 2108
rect 1512 2172 1528 2188
rect 1688 2252 1704 2268
rect 1576 2212 1592 2228
rect 1608 2192 1624 2208
rect 1736 2212 1752 2228
rect 1768 2212 1784 2228
rect 1688 2192 1704 2208
rect 1592 2172 1608 2188
rect 1624 2172 1640 2188
rect 1528 2152 1544 2168
rect 1576 2132 1592 2148
rect 1576 2112 1592 2128
rect 1640 2152 1656 2168
rect 1672 2152 1688 2168
rect 1624 2132 1640 2148
rect 1608 2112 1624 2128
rect 1789 2202 1825 2218
rect 1864 2292 1880 2308
rect 1880 2272 1896 2288
rect 1864 2252 1880 2268
rect 1768 2172 1784 2188
rect 1832 2172 1848 2188
rect 1832 2152 1848 2168
rect 1768 2132 1784 2148
rect 1544 2072 1560 2088
rect 1720 2072 1752 2088
rect 1304 2052 1320 2068
rect 1416 1992 1432 2008
rect 1624 1992 1640 2008
rect 1304 1932 1320 1948
rect 1336 1912 1352 1928
rect 1352 1912 1368 1928
rect 1464 1952 1480 1968
rect 1528 1952 1544 1968
rect 1544 1952 1560 1968
rect 1448 1912 1464 1928
rect 1320 1892 1336 1908
rect 1368 1852 1384 1868
rect 1416 1832 1432 1848
rect 1416 1792 1432 1808
rect 1288 1772 1304 1788
rect 1352 1772 1368 1788
rect 1256 1732 1272 1748
rect 1288 1732 1304 1748
rect 1272 1712 1288 1728
rect 1304 1712 1320 1728
rect 1400 1732 1416 1748
rect 1368 1712 1384 1728
rect 1464 1812 1480 1828
rect 1320 1692 1352 1708
rect 1432 1692 1448 1708
rect 1288 1652 1304 1668
rect 1368 1652 1384 1668
rect 1352 1632 1368 1648
rect 1240 1592 1256 1608
rect 1352 1592 1368 1608
rect 1304 1552 1320 1568
rect 1288 1512 1304 1528
rect 1448 1552 1464 1568
rect 1400 1512 1416 1528
rect 1496 1852 1512 1868
rect 1496 1752 1512 1768
rect 1544 1892 1560 1908
rect 1592 1892 1608 1908
rect 1560 1872 1576 1888
rect 1560 1852 1576 1868
rect 1528 1752 1544 1768
rect 1608 1852 1624 1868
rect 1576 1812 1592 1828
rect 1576 1752 1592 1768
rect 1512 1672 1528 1688
rect 1672 1932 1688 1948
rect 1736 2052 1752 2068
rect 1928 2312 1944 2328
rect 1992 2312 2008 2328
rect 2072 2312 2088 2328
rect 2136 2312 2152 2328
rect 2813 2402 2849 2418
rect 2920 2312 2936 2328
rect 3160 2312 3176 2328
rect 3512 2312 3528 2328
rect 3560 2312 3576 2328
rect 3592 2312 3608 2328
rect 1960 2292 1976 2308
rect 2200 2292 2216 2308
rect 2360 2292 2376 2308
rect 2472 2292 2488 2308
rect 2536 2292 2552 2308
rect 2584 2292 2600 2308
rect 2664 2292 2680 2308
rect 2728 2292 2744 2308
rect 2776 2292 2792 2308
rect 1928 2172 1944 2188
rect 1976 2252 1992 2268
rect 2104 2252 2120 2268
rect 2104 2232 2120 2248
rect 2168 2232 2184 2248
rect 1992 2192 2008 2208
rect 2040 2152 2056 2168
rect 2120 2212 2136 2228
rect 1960 2132 1976 2148
rect 1976 2132 1992 2148
rect 2040 2132 2056 2148
rect 2088 2132 2104 2148
rect 1944 2112 1960 2128
rect 2024 2112 2040 2128
rect 2088 2112 2104 2128
rect 1864 2092 1880 2108
rect 1912 2092 1928 2108
rect 2040 2092 2056 2108
rect 1832 1992 1864 2008
rect 1816 1892 1832 1908
rect 1720 1872 1736 1888
rect 1752 1872 1768 1888
rect 1848 1872 1864 1888
rect 1784 1852 1800 1868
rect 1832 1852 1848 1868
rect 1672 1832 1688 1848
rect 1624 1732 1640 1748
rect 1656 1732 1672 1748
rect 1688 1752 1704 1768
rect 1704 1732 1720 1748
rect 1789 1802 1825 1818
rect 1832 1732 1848 1748
rect 1752 1712 1768 1728
rect 1576 1672 1592 1688
rect 1560 1632 1576 1648
rect 1736 1672 1752 1688
rect 1720 1652 1736 1668
rect 1640 1592 1656 1608
rect 1560 1552 1576 1568
rect 1816 1552 1832 1568
rect 1480 1532 1496 1548
rect 1240 1492 1256 1508
rect 1464 1492 1480 1508
rect 1288 1472 1304 1488
rect 1336 1472 1352 1488
rect 1208 1412 1240 1428
rect 1192 1352 1208 1368
rect 1224 1352 1240 1368
rect 1272 1432 1288 1448
rect 1288 1392 1304 1408
rect 1320 1392 1336 1408
rect 1352 1392 1368 1408
rect 1512 1492 1528 1508
rect 1656 1532 1672 1548
rect 1704 1532 1736 1548
rect 1752 1532 1768 1548
rect 1784 1532 1800 1548
rect 1576 1492 1592 1508
rect 1496 1472 1512 1488
rect 1528 1472 1544 1488
rect 1560 1472 1576 1488
rect 1432 1432 1448 1448
rect 1400 1372 1416 1388
rect 1320 1352 1368 1368
rect 1384 1352 1400 1368
rect 1288 1332 1304 1348
rect 1208 1312 1224 1328
rect 1240 1292 1256 1308
rect 1176 1252 1192 1268
rect 1112 1232 1128 1248
rect 1192 1232 1208 1248
rect 1080 1152 1096 1168
rect 968 1072 984 1088
rect 1016 1072 1048 1088
rect 872 1032 888 1048
rect 920 992 936 1008
rect 952 972 968 988
rect 1064 1012 1080 1028
rect 760 932 776 948
rect 968 932 984 948
rect 1032 952 1064 968
rect 1064 932 1080 948
rect 680 892 696 908
rect 744 892 760 908
rect 808 892 824 908
rect 904 892 920 908
rect 936 892 952 908
rect 984 892 1000 908
rect 1016 892 1032 908
rect 1064 892 1080 908
rect 648 852 664 868
rect 680 832 696 848
rect 648 812 664 828
rect 648 752 664 768
rect 632 732 648 748
rect 664 732 680 748
rect 648 712 664 728
rect 664 692 680 708
rect 584 612 600 628
rect 584 592 600 608
rect 584 532 600 548
rect 616 512 632 528
rect 584 472 600 488
rect 568 352 584 368
rect 696 792 712 808
rect 712 592 728 608
rect 765 802 801 818
rect 872 812 888 828
rect 824 772 840 788
rect 840 772 856 788
rect 904 772 920 788
rect 920 732 936 748
rect 952 732 968 748
rect 744 712 760 728
rect 776 712 792 728
rect 856 692 872 708
rect 888 692 904 708
rect 920 692 936 708
rect 744 612 760 628
rect 728 572 744 588
rect 1096 952 1112 968
rect 1080 872 1096 888
rect 1048 852 1064 868
rect 1096 792 1112 808
rect 1096 772 1112 788
rect 1144 1212 1160 1228
rect 1528 1372 1544 1388
rect 1416 1332 1432 1348
rect 1608 1432 1624 1448
rect 1592 1392 1608 1408
rect 1784 1492 1800 1508
rect 1832 1492 1848 1508
rect 1656 1472 1672 1488
rect 1640 1432 1656 1448
rect 1640 1412 1656 1428
rect 1624 1392 1640 1408
rect 1464 1332 1480 1348
rect 1560 1332 1576 1348
rect 1624 1332 1640 1348
rect 1320 1292 1336 1308
rect 1256 1192 1272 1208
rect 1224 1132 1240 1148
rect 1480 1292 1496 1308
rect 1576 1292 1592 1308
rect 1320 1172 1336 1188
rect 1352 1172 1368 1188
rect 1384 1172 1400 1188
rect 1352 1152 1368 1168
rect 1240 1072 1256 1088
rect 1144 1052 1160 1068
rect 1208 1052 1224 1068
rect 1256 1052 1272 1068
rect 1192 1032 1208 1048
rect 1128 832 1144 848
rect 1064 692 1080 708
rect 1224 932 1240 948
rect 1176 912 1192 928
rect 1272 992 1288 1008
rect 1336 972 1352 988
rect 1176 892 1192 908
rect 1208 892 1224 908
rect 1304 912 1320 928
rect 1272 892 1288 908
rect 1208 852 1224 868
rect 1144 772 1160 788
rect 1400 1072 1416 1088
rect 1464 1132 1480 1148
rect 1432 1092 1448 1108
rect 1448 1072 1464 1088
rect 1416 1032 1432 1048
rect 1384 952 1400 968
rect 1512 1272 1528 1288
rect 1576 1232 1592 1248
rect 1608 1252 1624 1268
rect 1592 1132 1608 1148
rect 1480 1072 1496 1088
rect 1464 992 1480 1008
rect 1512 1052 1528 1068
rect 1592 1032 1608 1048
rect 1544 1012 1560 1028
rect 1736 1472 1752 1488
rect 1704 1452 1720 1468
rect 1752 1452 1768 1468
rect 1688 1432 1704 1448
rect 1720 1392 1736 1408
rect 1789 1402 1825 1418
rect 1736 1332 1752 1348
rect 1784 1312 1800 1328
rect 1704 1272 1720 1288
rect 1672 1232 1688 1248
rect 1688 1172 1704 1188
rect 1752 1232 1768 1248
rect 1784 1192 1800 1208
rect 1784 1172 1800 1188
rect 1720 1112 1736 1128
rect 1720 1092 1736 1108
rect 1752 1092 1768 1108
rect 1736 1072 1768 1088
rect 1656 992 1672 1008
rect 1624 972 1640 988
rect 1640 972 1656 988
rect 1560 952 1576 968
rect 1624 952 1640 968
rect 1384 912 1400 928
rect 1432 912 1448 928
rect 1576 892 1592 908
rect 1400 872 1416 888
rect 1320 852 1336 868
rect 1384 852 1400 868
rect 1240 772 1256 788
rect 1352 772 1368 788
rect 1256 692 1272 708
rect 1048 672 1064 688
rect 1128 672 1144 688
rect 904 652 920 668
rect 952 652 984 668
rect 1224 652 1240 668
rect 904 612 920 628
rect 792 572 808 588
rect 936 572 952 588
rect 872 532 888 548
rect 920 532 936 548
rect 968 532 984 548
rect 696 512 712 528
rect 728 512 744 528
rect 760 512 776 528
rect 680 472 696 488
rect 1032 572 1048 588
rect 1096 572 1112 588
rect 1176 632 1192 648
rect 1208 632 1224 648
rect 1192 572 1208 588
rect 1096 532 1112 548
rect 1336 672 1352 688
rect 1288 652 1304 668
rect 1272 592 1288 608
rect 1224 572 1240 588
rect 1320 572 1336 588
rect 1608 852 1624 868
rect 1656 852 1672 868
rect 1416 812 1432 828
rect 1576 812 1592 828
rect 1560 792 1576 808
rect 1368 652 1384 668
rect 1352 572 1368 588
rect 1384 572 1400 588
rect 824 512 856 528
rect 984 512 1000 528
rect 1048 512 1064 528
rect 1080 512 1096 528
rect 1160 512 1176 528
rect 1320 512 1336 528
rect 776 472 792 488
rect 840 472 856 488
rect 632 432 648 448
rect 680 432 696 448
rect 765 402 801 418
rect 616 372 632 388
rect 600 332 616 348
rect 648 292 664 308
rect 696 292 712 308
rect 792 292 808 308
rect 296 172 312 188
rect 392 172 408 188
rect 488 172 504 188
rect 552 172 568 188
rect 616 212 632 228
rect 280 112 296 128
rect 328 112 344 128
rect 440 112 456 128
rect 520 112 536 128
rect 264 92 280 108
rect 200 72 216 88
rect 296 72 312 88
rect 408 92 424 108
rect 552 72 568 88
rect 328 52 344 68
rect 744 252 760 268
rect 680 232 696 248
rect 712 232 728 248
rect 648 172 664 188
rect 952 492 968 508
rect 968 472 984 488
rect 856 452 872 468
rect 920 372 936 388
rect 872 292 888 308
rect 984 292 1000 308
rect 840 272 856 288
rect 888 192 904 208
rect 824 152 840 168
rect 968 172 984 188
rect 1016 412 1032 428
rect 1112 492 1128 508
rect 1304 492 1320 508
rect 1128 452 1144 468
rect 1064 292 1080 308
rect 1112 292 1128 308
rect 1064 272 1080 288
rect 1096 272 1112 288
rect 1016 252 1032 268
rect 1048 232 1064 248
rect 1096 232 1112 248
rect 968 132 984 148
rect 1032 132 1048 148
rect 696 112 712 128
rect 744 112 760 128
rect 888 112 904 128
rect 616 12 664 28
rect 856 92 872 108
rect 952 92 968 108
rect 1016 92 1032 108
rect 888 52 904 68
rect 765 2 801 18
rect 984 52 1000 68
rect 1112 212 1128 228
rect 1096 172 1112 188
rect 1144 432 1160 448
rect 1192 392 1208 408
rect 1288 452 1304 468
rect 1416 672 1432 688
rect 1480 672 1512 688
rect 1528 672 1544 688
rect 1448 552 1464 568
rect 1832 1192 1848 1208
rect 1864 1832 1880 1848
rect 1864 1792 1880 1808
rect 1896 1952 1912 1968
rect 1880 1772 1896 1788
rect 1880 1732 1896 1748
rect 1944 1932 1960 1948
rect 1992 1932 2008 1948
rect 1928 1892 1944 1908
rect 2008 1912 2024 1928
rect 2184 2092 2200 2108
rect 2072 2072 2088 2088
rect 2184 2052 2200 2068
rect 2104 1952 2120 1968
rect 2040 1892 2056 1908
rect 1960 1872 1976 1888
rect 1944 1852 1960 1868
rect 1928 1732 1944 1748
rect 1992 1812 2008 1828
rect 2024 1772 2056 1788
rect 1976 1752 1992 1768
rect 1992 1752 2008 1768
rect 2264 2272 2280 2288
rect 2296 2272 2312 2288
rect 2424 2272 2440 2288
rect 2392 2252 2408 2268
rect 2456 2252 2472 2268
rect 2584 2232 2600 2248
rect 2216 2192 2232 2208
rect 2248 2132 2264 2148
rect 2376 2152 2392 2168
rect 2456 2152 2472 2168
rect 2440 2132 2456 2148
rect 2216 2112 2232 2128
rect 2232 2112 2248 2128
rect 2312 2112 2328 2128
rect 2328 2112 2344 2128
rect 2392 2072 2408 2088
rect 2296 2032 2312 2048
rect 2424 1992 2440 2008
rect 2488 1992 2504 2008
rect 2488 1972 2504 1988
rect 2408 1952 2424 1968
rect 2200 1932 2216 1948
rect 2280 1932 2296 1948
rect 2216 1912 2232 1928
rect 2280 1912 2296 1928
rect 2312 1912 2328 1928
rect 2152 1892 2168 1908
rect 2200 1892 2232 1908
rect 2264 1892 2280 1908
rect 2328 1892 2344 1908
rect 2472 1892 2488 1908
rect 2120 1872 2136 1888
rect 2072 1812 2088 1828
rect 2088 1752 2104 1768
rect 2152 1852 2168 1868
rect 2168 1752 2184 1768
rect 1880 1712 1896 1728
rect 1992 1712 2008 1728
rect 2056 1732 2072 1748
rect 2024 1712 2040 1728
rect 2056 1712 2072 1728
rect 2104 1712 2120 1728
rect 2216 1712 2232 1728
rect 1880 1672 1896 1688
rect 1864 1532 1880 1548
rect 1960 1652 1976 1668
rect 2008 1652 2024 1668
rect 1896 1612 1912 1628
rect 1896 1532 1912 1548
rect 1928 1472 1944 1488
rect 1880 1412 1896 1428
rect 1896 1392 1912 1408
rect 1864 1352 1896 1368
rect 2024 1632 2056 1648
rect 2136 1632 2152 1648
rect 2152 1612 2168 1628
rect 2056 1552 2072 1568
rect 2104 1512 2120 1528
rect 1976 1452 1992 1468
rect 1992 1432 2008 1448
rect 1992 1412 2008 1428
rect 1960 1392 1976 1408
rect 1928 1332 1944 1348
rect 1944 1332 1960 1348
rect 1864 1312 1880 1328
rect 1928 1312 1944 1328
rect 1960 1312 1976 1328
rect 1896 1232 1912 1248
rect 1864 1212 1880 1228
rect 1864 1192 1896 1208
rect 1789 1002 1825 1018
rect 1848 1092 1864 1108
rect 1848 1072 1864 1088
rect 1848 1012 1864 1028
rect 1720 972 1736 988
rect 1768 972 1800 988
rect 1832 972 1848 988
rect 1704 932 1720 948
rect 2088 1472 2104 1488
rect 2120 1492 2136 1508
rect 2248 1652 2264 1668
rect 2248 1632 2264 1648
rect 2232 1592 2248 1608
rect 2200 1512 2216 1528
rect 2136 1472 2152 1488
rect 2152 1472 2168 1488
rect 2184 1452 2200 1468
rect 2216 1452 2248 1468
rect 2120 1432 2136 1448
rect 2168 1432 2184 1448
rect 2200 1432 2216 1448
rect 2040 1352 2056 1368
rect 2104 1352 2120 1368
rect 2040 1332 2056 1348
rect 2024 1312 2040 1328
rect 2024 1232 2040 1248
rect 1992 1192 2008 1208
rect 1912 1132 1928 1148
rect 2152 1412 2168 1428
rect 2056 1292 2072 1308
rect 2136 1292 2152 1308
rect 2120 1252 2136 1268
rect 2072 1232 2088 1248
rect 2040 1132 2056 1148
rect 1912 1092 1928 1108
rect 1928 1012 1960 1028
rect 2104 1212 2120 1228
rect 1976 1072 1992 1088
rect 2056 1072 2072 1088
rect 1992 1052 2008 1068
rect 2040 1052 2056 1068
rect 2040 1012 2056 1028
rect 1976 972 1992 988
rect 2056 972 2072 988
rect 2136 972 2152 988
rect 1736 912 1752 928
rect 1688 892 1704 908
rect 1848 892 1864 908
rect 1720 852 1736 868
rect 1672 812 1688 828
rect 1688 772 1704 788
rect 1672 752 1688 768
rect 1608 732 1624 748
rect 1608 672 1624 688
rect 1560 652 1576 668
rect 1656 672 1672 688
rect 1704 732 1720 748
rect 1816 812 1832 828
rect 1784 772 1800 788
rect 1816 772 1832 788
rect 1720 692 1736 708
rect 1784 692 1800 708
rect 1528 612 1560 628
rect 1496 572 1512 588
rect 1384 512 1400 528
rect 1448 512 1464 528
rect 1368 492 1384 508
rect 1352 412 1368 428
rect 1272 392 1288 408
rect 1320 392 1336 408
rect 1256 372 1272 388
rect 1288 372 1304 388
rect 1144 352 1176 368
rect 1208 352 1224 368
rect 1144 212 1160 228
rect 1192 292 1208 308
rect 1304 312 1320 328
rect 1272 232 1288 248
rect 1272 192 1288 208
rect 1160 152 1176 168
rect 1416 492 1432 508
rect 1448 492 1464 508
rect 1464 472 1480 488
rect 1496 472 1512 488
rect 1656 652 1672 668
rect 1624 632 1640 648
rect 1576 532 1592 548
rect 1544 492 1560 508
rect 1592 492 1608 508
rect 1576 452 1592 468
rect 1512 372 1528 388
rect 1400 352 1416 368
rect 1336 312 1352 328
rect 1464 312 1480 328
rect 1496 312 1512 328
rect 1560 312 1576 328
rect 1704 572 1720 588
rect 1789 602 1825 618
rect 1736 572 1752 588
rect 1832 572 1848 588
rect 1816 552 1832 568
rect 1720 532 1736 548
rect 1640 492 1656 508
rect 1672 492 1688 508
rect 1656 452 1672 468
rect 1720 452 1736 468
rect 1368 292 1384 308
rect 1416 292 1432 308
rect 1464 292 1480 308
rect 1512 292 1528 308
rect 1528 292 1544 308
rect 1608 292 1624 308
rect 1064 132 1080 148
rect 1144 132 1160 148
rect 1192 132 1208 148
rect 1240 132 1256 148
rect 1256 112 1272 128
rect 1240 92 1256 108
rect 1272 92 1288 108
rect 1208 72 1224 88
rect 1032 32 1048 48
rect 1224 12 1240 28
rect 1400 252 1416 268
rect 1800 532 1816 548
rect 1752 432 1768 448
rect 1736 392 1752 408
rect 1720 372 1736 388
rect 1752 352 1768 368
rect 1640 332 1656 348
rect 1688 312 1704 328
rect 1752 312 1768 328
rect 1656 292 1672 308
rect 1720 292 1736 308
rect 1704 272 1720 288
rect 1432 232 1448 248
rect 1400 192 1416 208
rect 1624 252 1640 268
rect 1688 252 1704 268
rect 1544 232 1560 248
rect 1528 172 1544 188
rect 1752 212 1768 228
rect 1672 192 1688 208
rect 1560 172 1576 188
rect 1608 172 1624 188
rect 1640 172 1656 188
rect 1432 152 1448 168
rect 1464 152 1480 168
rect 1384 132 1400 148
rect 1720 172 1736 188
rect 1608 132 1624 148
rect 1656 132 1672 148
rect 1352 112 1368 128
rect 1528 112 1544 128
rect 1480 92 1496 108
rect 1512 72 1528 88
rect 1624 72 1640 88
rect 1320 12 1336 28
rect 1368 12 1384 28
rect 1464 12 1480 28
rect 1528 12 1544 28
rect 1912 912 1928 928
rect 1896 892 1912 908
rect 1912 852 1928 868
rect 1896 812 1912 828
rect 2024 952 2040 968
rect 2088 952 2104 968
rect 2120 952 2136 968
rect 2088 932 2104 948
rect 2040 912 2056 928
rect 2072 912 2088 928
rect 1912 732 1944 748
rect 1944 692 1960 708
rect 1880 632 1896 648
rect 1864 572 1880 588
rect 1832 472 1848 488
rect 1896 412 1912 428
rect 1832 392 1848 408
rect 1816 252 1832 268
rect 1784 232 1800 248
rect 1768 192 1784 208
rect 1789 202 1825 218
rect 1896 332 1928 348
rect 1848 312 1864 328
rect 1864 292 1880 308
rect 1912 292 1928 308
rect 1880 272 1896 288
rect 2008 892 2024 908
rect 2104 892 2120 908
rect 2120 872 2136 888
rect 2184 1412 2200 1428
rect 2344 1872 2360 1888
rect 2424 1872 2440 1888
rect 2424 1832 2440 1848
rect 2632 2212 2648 2228
rect 2680 2172 2696 2188
rect 2520 2152 2536 2168
rect 2664 2152 2680 2168
rect 2696 2152 2712 2168
rect 2808 2172 2824 2188
rect 2776 2152 2792 2168
rect 2536 2132 2552 2148
rect 2552 2132 2568 2148
rect 2600 2132 2616 2148
rect 2632 2132 2648 2148
rect 2664 2132 2680 2148
rect 2760 2132 2776 2148
rect 2600 2092 2616 2108
rect 2584 2012 2600 2028
rect 2808 2112 2824 2128
rect 2696 2092 2712 2108
rect 2728 2092 2744 2108
rect 2760 2092 2776 2108
rect 2664 2032 2680 2048
rect 2648 1992 2664 2008
rect 2616 1932 2632 1948
rect 2648 1932 2664 1948
rect 2616 1912 2632 1928
rect 2664 1912 2680 1928
rect 2568 1892 2584 1908
rect 2520 1832 2552 1848
rect 2504 1792 2520 1808
rect 2456 1772 2472 1788
rect 2632 1872 2648 1888
rect 2616 1852 2632 1868
rect 2520 1732 2536 1748
rect 2552 1732 2568 1748
rect 2568 1732 2584 1748
rect 2600 1732 2616 1748
rect 2296 1712 2312 1728
rect 2328 1712 2344 1728
rect 2296 1632 2312 1648
rect 2264 1612 2280 1628
rect 2312 1512 2328 1528
rect 2344 1632 2360 1648
rect 2344 1612 2360 1628
rect 2376 1612 2392 1628
rect 2536 1692 2552 1708
rect 2600 1712 2616 1728
rect 2664 1732 2680 1748
rect 2648 1712 2664 1728
rect 2520 1652 2536 1668
rect 2408 1552 2424 1568
rect 2456 1552 2472 1568
rect 2424 1492 2440 1508
rect 2280 1452 2296 1468
rect 2312 1452 2328 1468
rect 2664 1632 2680 1648
rect 2552 1512 2568 1528
rect 2616 1512 2632 1528
rect 2440 1472 2456 1488
rect 2488 1472 2504 1488
rect 2536 1472 2552 1488
rect 2568 1472 2584 1488
rect 2376 1452 2392 1468
rect 2328 1412 2360 1428
rect 2392 1392 2408 1408
rect 2504 1432 2520 1448
rect 2552 1452 2568 1468
rect 2216 1372 2232 1388
rect 2360 1372 2376 1388
rect 2200 1332 2216 1348
rect 2344 1332 2360 1348
rect 2280 1312 2296 1328
rect 2232 1292 2248 1308
rect 2264 1292 2280 1308
rect 2296 1292 2312 1308
rect 2328 1292 2344 1308
rect 2168 1132 2184 1148
rect 2200 1132 2216 1148
rect 2184 1072 2200 1088
rect 2392 1352 2408 1368
rect 2520 1352 2536 1368
rect 2376 1312 2392 1328
rect 2504 1312 2520 1328
rect 3000 2292 3016 2308
rect 3128 2292 3144 2308
rect 3192 2292 3208 2308
rect 2968 2272 2984 2288
rect 2984 2272 3000 2288
rect 2936 2232 2952 2248
rect 3032 2272 3048 2288
rect 3000 2192 3016 2208
rect 2888 2172 2904 2188
rect 2920 2172 2936 2188
rect 2984 2172 3000 2188
rect 3016 2152 3032 2168
rect 2872 2132 2888 2148
rect 2888 2132 2904 2148
rect 2968 2132 2984 2148
rect 2920 2052 2936 2068
rect 2824 2032 2840 2048
rect 2696 1872 2712 1888
rect 3032 2092 3048 2108
rect 2760 2012 2776 2028
rect 2813 2002 2849 2018
rect 2952 2012 2968 2028
rect 2904 1952 2920 1968
rect 2824 1912 2840 1928
rect 2744 1892 2760 1908
rect 2968 1932 2984 1948
rect 2936 1912 2952 1928
rect 2744 1872 2760 1888
rect 2792 1872 2808 1888
rect 2888 1872 2904 1888
rect 2952 1872 2968 1888
rect 2728 1852 2760 1868
rect 2712 1732 2728 1748
rect 2728 1552 2744 1568
rect 2632 1492 2648 1508
rect 2600 1432 2616 1448
rect 2568 1412 2584 1428
rect 2584 1392 2600 1408
rect 2680 1452 2696 1468
rect 2616 1372 2632 1388
rect 2552 1312 2568 1328
rect 2648 1312 2664 1328
rect 2392 1292 2408 1308
rect 2472 1292 2504 1308
rect 2600 1292 2616 1308
rect 2632 1292 2648 1308
rect 2408 1192 2424 1208
rect 2440 1192 2456 1208
rect 2376 1152 2392 1168
rect 2552 1152 2568 1168
rect 2344 1112 2360 1128
rect 2232 1092 2248 1108
rect 2264 1092 2280 1108
rect 2312 1092 2328 1108
rect 2216 1072 2232 1088
rect 2200 1052 2216 1068
rect 2280 1072 2296 1088
rect 2328 1072 2344 1088
rect 2296 1052 2312 1068
rect 2248 952 2264 968
rect 2184 932 2200 948
rect 2344 952 2360 968
rect 2168 912 2184 928
rect 2200 912 2216 928
rect 2344 912 2360 928
rect 2168 892 2184 908
rect 2152 852 2168 868
rect 2184 852 2200 868
rect 2088 832 2104 848
rect 1976 732 1992 748
rect 2024 712 2040 728
rect 2072 712 2088 728
rect 2040 692 2056 708
rect 2136 752 2152 768
rect 2120 732 2136 748
rect 2008 672 2024 688
rect 2024 672 2040 688
rect 1960 652 1976 668
rect 1976 652 1992 668
rect 2104 612 2120 628
rect 2056 572 2072 588
rect 2024 552 2040 568
rect 2024 512 2040 528
rect 2040 512 2056 528
rect 1960 352 1976 368
rect 1960 332 1976 348
rect 1944 312 1960 328
rect 2024 492 2040 508
rect 2056 492 2072 508
rect 2008 472 2024 488
rect 2072 472 2088 488
rect 2088 412 2104 428
rect 2040 352 2056 368
rect 1944 292 1960 308
rect 1896 212 1912 228
rect 1928 212 1944 228
rect 2024 292 2040 308
rect 2072 292 2088 308
rect 2040 272 2056 288
rect 1992 212 2008 228
rect 1976 192 1992 208
rect 2024 192 2040 208
rect 1976 172 1992 188
rect 2008 172 2024 188
rect 2040 172 2056 188
rect 1752 132 1768 148
rect 1912 132 1928 148
rect 1736 112 1752 128
rect 1768 112 1784 128
rect 1864 112 1880 128
rect 1688 92 1704 108
rect 1720 92 1736 108
rect 1816 92 1832 108
rect 1848 92 1864 108
rect 1880 92 1896 108
rect 1784 32 1800 48
rect 1672 12 1688 28
rect 1720 12 1736 28
rect 1928 112 1944 128
rect 2504 1132 2520 1148
rect 2600 1132 2616 1148
rect 2424 1112 2440 1128
rect 2488 1112 2504 1128
rect 2584 1112 2600 1128
rect 2632 1112 2648 1128
rect 2440 1092 2456 1108
rect 2536 1092 2552 1108
rect 2408 1052 2424 1068
rect 2472 1052 2488 1068
rect 2520 1052 2536 1068
rect 2568 1052 2584 1068
rect 2456 1032 2472 1048
rect 2392 1012 2408 1028
rect 2696 1352 2712 1368
rect 2712 1312 2728 1328
rect 2776 1732 2792 1748
rect 2760 1712 2776 1728
rect 2792 1712 2808 1728
rect 2856 1852 2888 1868
rect 2920 1752 2936 1768
rect 2936 1712 2952 1728
rect 2808 1692 2824 1708
rect 2840 1692 2856 1708
rect 2856 1672 2872 1688
rect 2856 1632 2872 1648
rect 2936 1632 2952 1648
rect 2813 1602 2849 1618
rect 2840 1532 2856 1548
rect 2824 1492 2840 1508
rect 2776 1472 2792 1488
rect 2744 1412 2760 1428
rect 2792 1352 2808 1368
rect 2856 1452 2872 1468
rect 2888 1432 2904 1448
rect 2760 1332 2776 1348
rect 2808 1332 2824 1348
rect 2728 1292 2744 1308
rect 2760 1292 2776 1308
rect 2696 1252 2728 1268
rect 2664 1212 2680 1228
rect 2680 1132 2696 1148
rect 2744 1132 2760 1148
rect 2648 1072 2664 1088
rect 2616 1012 2632 1028
rect 2904 1392 2920 1408
rect 3016 1912 3032 1928
rect 3000 1892 3016 1908
rect 2984 1632 3000 1648
rect 3432 2292 3464 2308
rect 3496 2292 3512 2308
rect 3288 2272 3304 2288
rect 3288 2232 3304 2248
rect 3128 2152 3144 2168
rect 3192 2152 3208 2168
rect 3128 2132 3144 2148
rect 3240 2132 3256 2148
rect 3320 2172 3336 2188
rect 3112 2112 3128 2128
rect 3096 2092 3112 2108
rect 3160 2052 3176 2068
rect 3144 2012 3160 2028
rect 3176 2012 3192 2028
rect 3112 1932 3128 1948
rect 3080 1912 3084 1928
rect 3084 1912 3096 1928
rect 3096 1892 3112 1908
rect 3048 1872 3080 1888
rect 3112 1872 3128 1888
rect 3128 1872 3144 1888
rect 3080 1812 3096 1828
rect 3048 1792 3096 1808
rect 3032 1732 3048 1748
rect 3016 1712 3032 1728
rect 3032 1552 3048 1568
rect 3000 1532 3016 1548
rect 3016 1512 3032 1528
rect 3048 1492 3064 1508
rect 3000 1472 3016 1488
rect 2984 1432 3000 1448
rect 2952 1412 2968 1428
rect 2968 1372 2984 1388
rect 3160 1832 3176 1848
rect 3160 1812 3176 1828
rect 3128 1772 3144 1788
rect 3096 1732 3112 1748
rect 3192 1912 3208 1928
rect 3240 1912 3256 1928
rect 3304 1912 3320 1928
rect 3288 1892 3304 1908
rect 3224 1872 3240 1888
rect 3272 1872 3288 1888
rect 3224 1852 3240 1868
rect 3288 1772 3304 1788
rect 3240 1752 3256 1768
rect 3336 2092 3352 2108
rect 3368 2072 3384 2088
rect 3368 2032 3384 2048
rect 3400 2032 3416 2048
rect 3464 2032 3480 2048
rect 3528 2032 3544 2048
rect 3416 1912 3432 1928
rect 3640 2132 3656 2148
rect 3560 2012 3576 2028
rect 3592 2012 3608 2028
rect 3576 1932 3592 1948
rect 3480 1892 3496 1908
rect 3544 1892 3560 1908
rect 3336 1872 3352 1888
rect 3384 1872 3400 1888
rect 3464 1872 3480 1888
rect 3352 1832 3368 1848
rect 3432 1832 3448 1848
rect 3336 1812 3352 1828
rect 3240 1732 3256 1748
rect 3272 1732 3288 1748
rect 3368 1732 3384 1748
rect 3416 1732 3432 1748
rect 3080 1712 3096 1728
rect 3128 1712 3144 1728
rect 3272 1712 3288 1728
rect 3288 1692 3304 1708
rect 3176 1672 3192 1688
rect 3256 1652 3272 1668
rect 3144 1632 3160 1648
rect 3160 1612 3176 1628
rect 3112 1512 3128 1528
rect 3128 1492 3144 1508
rect 3208 1492 3224 1508
rect 3336 1712 3352 1728
rect 3400 1672 3416 1688
rect 3320 1552 3336 1568
rect 3368 1532 3384 1548
rect 3288 1512 3304 1528
rect 3320 1512 3336 1528
rect 3384 1512 3400 1528
rect 3288 1492 3320 1508
rect 3144 1472 3160 1488
rect 3272 1472 3288 1488
rect 3128 1452 3144 1468
rect 3096 1412 3112 1428
rect 2920 1332 2936 1348
rect 3096 1332 3112 1348
rect 3000 1312 3016 1328
rect 3048 1312 3064 1328
rect 2872 1292 2888 1308
rect 2920 1292 2936 1308
rect 2813 1202 2849 1218
rect 2904 1272 2920 1288
rect 2936 1272 2952 1288
rect 2968 1272 2984 1288
rect 3080 1272 3096 1288
rect 3128 1272 3144 1288
rect 2920 1252 2936 1268
rect 2936 1252 2952 1268
rect 3000 1252 3016 1268
rect 2936 1232 2952 1248
rect 2888 1192 2904 1208
rect 2920 1192 2936 1208
rect 2824 1172 2840 1188
rect 2792 1112 2808 1128
rect 2888 1152 2904 1168
rect 2920 1112 2936 1128
rect 3000 1192 3016 1208
rect 3048 1132 3064 1148
rect 3032 1112 3048 1128
rect 2872 1092 2888 1108
rect 2952 1072 2968 1088
rect 2728 1052 2744 1068
rect 2856 1052 2872 1068
rect 2488 992 2504 1008
rect 2648 992 2680 1008
rect 2520 952 2536 968
rect 2552 952 2568 968
rect 2680 972 2696 988
rect 2664 952 2696 968
rect 2728 952 2744 968
rect 2632 932 2648 948
rect 2696 932 2712 948
rect 2712 932 2728 948
rect 2776 952 2792 968
rect 2536 912 2552 928
rect 2296 872 2312 888
rect 2424 892 2440 908
rect 2808 992 2824 1008
rect 2920 1032 2936 1048
rect 3000 1032 3016 1048
rect 2952 932 2968 948
rect 2872 912 2888 928
rect 2600 892 2616 908
rect 2792 892 2808 908
rect 3016 1012 3032 1028
rect 3112 1232 3128 1248
rect 3320 1432 3336 1448
rect 3160 1372 3176 1388
rect 3176 1352 3192 1368
rect 3304 1372 3320 1388
rect 3208 1332 3224 1348
rect 3240 1332 3256 1348
rect 3256 1292 3288 1308
rect 3384 1452 3400 1468
rect 3384 1392 3400 1408
rect 3368 1352 3384 1368
rect 3304 1312 3320 1328
rect 3384 1312 3400 1328
rect 3208 1272 3224 1288
rect 3240 1272 3256 1288
rect 3288 1272 3304 1288
rect 3144 1172 3160 1188
rect 3176 1172 3192 1188
rect 3160 1112 3176 1128
rect 3240 1152 3256 1168
rect 3208 1112 3224 1128
rect 3064 1092 3080 1108
rect 3128 1072 3144 1088
rect 3016 932 3032 948
rect 3048 932 3080 948
rect 3112 972 3128 988
rect 3032 912 3048 928
rect 2408 832 2424 848
rect 2904 832 2920 848
rect 2424 792 2440 808
rect 2216 772 2232 788
rect 2408 732 2424 748
rect 2232 712 2248 728
rect 2296 712 2312 728
rect 2328 712 2344 728
rect 2216 692 2232 708
rect 2392 692 2408 708
rect 2136 632 2152 648
rect 2184 632 2200 648
rect 2200 592 2216 608
rect 2184 572 2216 588
rect 2136 532 2152 548
rect 2280 532 2296 548
rect 2536 772 2552 788
rect 2488 712 2504 728
rect 2520 712 2536 728
rect 2632 752 2648 768
rect 2552 732 2568 748
rect 2813 802 2849 818
rect 3000 792 3016 808
rect 3032 792 3048 808
rect 2792 772 2808 788
rect 2952 772 2968 788
rect 2984 772 3000 788
rect 3256 1112 3272 1128
rect 3288 1112 3304 1128
rect 3336 1292 3352 1308
rect 3464 1592 3480 1608
rect 3432 1572 3464 1588
rect 3544 1852 3560 1868
rect 3496 1832 3512 1848
rect 3592 1832 3608 1848
rect 3512 1812 3528 1828
rect 3624 1792 3640 1808
rect 3528 1732 3544 1748
rect 3640 1732 3656 1748
rect 3544 1712 3560 1728
rect 3464 1532 3496 1548
rect 3576 1532 3592 1548
rect 3576 1512 3592 1528
rect 3432 1472 3448 1488
rect 3512 1472 3528 1488
rect 3480 1452 3496 1468
rect 3496 1432 3512 1448
rect 3448 1372 3464 1388
rect 3432 1352 3448 1368
rect 3432 1292 3448 1308
rect 3416 1272 3432 1288
rect 3416 1252 3432 1268
rect 3400 1132 3416 1148
rect 3336 1092 3352 1108
rect 3352 1092 3368 1108
rect 3416 1092 3432 1108
rect 3144 1032 3160 1048
rect 3128 932 3144 948
rect 3080 872 3096 888
rect 3096 852 3112 868
rect 3144 852 3160 868
rect 3176 952 3192 968
rect 3224 932 3240 948
rect 3208 912 3224 928
rect 3256 1012 3272 1028
rect 3272 992 3288 1008
rect 3352 1052 3368 1068
rect 3304 972 3320 988
rect 3256 952 3272 968
rect 3544 1452 3560 1468
rect 3560 1432 3576 1448
rect 3544 1412 3560 1428
rect 3608 1492 3624 1508
rect 3576 1412 3592 1428
rect 3528 1352 3544 1368
rect 3528 1312 3544 1328
rect 3512 1292 3528 1308
rect 3528 1292 3544 1308
rect 3496 1272 3528 1288
rect 3512 1172 3528 1188
rect 3592 1272 3608 1288
rect 3624 1472 3640 1488
rect 3624 1332 3640 1348
rect 3560 1112 3576 1128
rect 3496 1092 3512 1108
rect 3544 1092 3560 1108
rect 3432 1072 3480 1088
rect 3512 1072 3528 1088
rect 3528 1012 3544 1028
rect 3528 992 3544 1008
rect 3528 952 3544 968
rect 3592 952 3608 968
rect 3304 932 3320 948
rect 3336 932 3352 948
rect 3368 932 3384 948
rect 3448 932 3464 948
rect 3480 932 3496 948
rect 3288 912 3304 928
rect 3272 892 3288 908
rect 3256 812 3272 828
rect 3160 752 3176 768
rect 3064 732 3080 748
rect 3000 712 3016 728
rect 2536 692 2552 708
rect 2600 692 2616 708
rect 2712 692 2728 708
rect 2744 692 2760 708
rect 2488 672 2504 688
rect 2680 672 2696 688
rect 2728 672 2744 688
rect 2872 672 2888 688
rect 2904 672 2920 688
rect 3064 672 3080 688
rect 3096 672 3112 688
rect 2440 652 2456 668
rect 2600 652 2616 668
rect 2632 652 2648 668
rect 2648 652 2664 668
rect 2472 592 2488 608
rect 2424 552 2440 568
rect 2536 552 2552 568
rect 2168 512 2184 528
rect 2520 512 2536 528
rect 2568 512 2584 528
rect 2168 492 2184 508
rect 2376 452 2392 468
rect 2216 432 2232 448
rect 2328 432 2344 448
rect 2152 372 2168 388
rect 2120 292 2136 308
rect 2104 272 2120 288
rect 2264 272 2280 288
rect 2392 252 2408 268
rect 2280 172 2296 188
rect 2328 172 2344 188
rect 2360 172 2376 188
rect 2392 172 2408 188
rect 2488 172 2504 188
rect 2056 132 2072 148
rect 2088 132 2104 148
rect 2120 132 2136 148
rect 2216 132 2232 148
rect 2248 132 2264 148
rect 2360 112 2376 128
rect 2616 632 2632 648
rect 2632 632 2648 648
rect 2664 632 2696 648
rect 2632 572 2648 588
rect 3336 912 3352 928
rect 3336 892 3352 908
rect 3384 832 3416 848
rect 3512 812 3528 828
rect 3480 772 3496 788
rect 3512 772 3528 788
rect 3192 672 3208 688
rect 3224 672 3240 688
rect 3320 672 3336 688
rect 3352 672 3368 688
rect 3384 672 3400 688
rect 3416 672 3432 688
rect 3464 672 3480 688
rect 3144 652 3160 668
rect 3176 652 3192 668
rect 3256 632 3272 648
rect 2872 592 2888 608
rect 2952 552 2968 568
rect 2952 532 2968 548
rect 2984 532 3000 548
rect 3064 532 3080 548
rect 3112 532 3128 548
rect 3144 532 3160 548
rect 2696 512 2712 528
rect 2728 512 2744 528
rect 2568 472 2584 488
rect 2584 472 2600 488
rect 2696 432 2712 448
rect 2813 402 2849 418
rect 2904 492 2920 508
rect 3192 472 3208 488
rect 3224 472 3240 488
rect 3256 472 3272 488
rect 3272 472 3288 488
rect 3288 472 3304 488
rect 2760 372 2776 388
rect 2808 372 2824 388
rect 2856 372 2872 388
rect 2888 372 2904 388
rect 2904 372 2920 388
rect 2568 292 2584 308
rect 3048 292 3064 308
rect 2552 252 2568 268
rect 2536 172 2552 188
rect 2568 172 2584 188
rect 2616 132 2632 148
rect 2648 132 2664 148
rect 2712 132 2728 148
rect 2760 152 2776 168
rect 2968 232 2984 248
rect 3032 232 3048 248
rect 2760 132 2776 148
rect 2792 132 2808 148
rect 2904 132 2920 148
rect 2936 132 2952 148
rect 3080 172 3096 188
rect 3112 172 3128 188
rect 3160 172 3192 188
rect 3224 172 3240 188
rect 2504 112 2520 128
rect 2696 112 2712 128
rect 2728 112 2760 128
rect 2856 112 2872 128
rect 3368 532 3384 548
rect 3448 532 3464 548
rect 3480 532 3496 548
rect 3352 472 3384 488
rect 3480 392 3496 408
rect 3368 292 3384 308
rect 3512 292 3528 308
rect 3400 232 3416 248
rect 3448 232 3464 248
rect 3480 232 3496 248
rect 3496 232 3512 248
rect 3304 132 3320 148
rect 3512 132 3528 148
rect 3544 932 3560 948
rect 3592 772 3608 788
rect 3576 712 3592 728
rect 3544 672 3560 688
rect 3656 912 3672 928
rect 3640 772 3656 788
rect 3576 532 3592 548
rect 3608 532 3624 548
rect 3544 512 3560 528
rect 3560 392 3576 408
rect 3608 512 3624 528
rect 3656 512 3672 528
rect 3656 312 3672 328
rect 3288 112 3304 128
rect 3336 112 3352 128
rect 3592 112 3608 128
rect 1976 92 1992 108
rect 2813 2 2849 18
rect 2856 12 2872 28
rect 2888 12 2904 28
rect 3016 12 3032 28
rect 3048 12 3064 28
<< metal3 >>
rect 824 2417 840 2423
rect 1000 2417 1800 2423
rect 1032 2397 1272 2403
rect 1464 2397 1688 2403
rect 712 2337 1016 2343
rect 1224 2337 1608 2343
rect 1640 2337 1912 2343
rect -51 2317 8 2323
rect 648 2317 856 2323
rect 1064 2317 1224 2323
rect 1400 2317 1464 2323
rect 1544 2317 1560 2323
rect 1640 2317 1688 2323
rect 1752 2317 1928 2323
rect 1944 2317 1992 2323
rect 2008 2317 2072 2323
rect 2088 2317 2136 2323
rect 2936 2317 3160 2323
rect 3528 2317 3560 2323
rect 3576 2317 3592 2323
rect 248 2297 328 2303
rect 408 2297 456 2303
rect 472 2297 552 2303
rect 920 2297 936 2303
rect 952 2297 968 2303
rect 1144 2297 1192 2303
rect 1528 2297 1864 2303
rect 1976 2297 2200 2303
rect 2376 2297 2472 2303
rect 2488 2297 2536 2303
rect 2552 2297 2584 2303
rect 2680 2297 2728 2303
rect 2744 2297 2776 2303
rect 3016 2297 3128 2303
rect 3208 2297 3432 2303
rect 3464 2297 3496 2303
rect 472 2277 584 2283
rect 600 2277 824 2283
rect 936 2277 984 2283
rect 1160 2277 1208 2283
rect 1384 2277 1432 2283
rect 1512 2277 1544 2283
rect 1672 2277 1880 2283
rect 2088 2277 2264 2283
rect 2312 2277 2424 2283
rect 2440 2277 2968 2283
rect 3000 2277 3032 2283
rect 568 2257 680 2263
rect 872 2257 1064 2263
rect 1256 2257 1288 2263
rect 1320 2257 1688 2263
rect 1704 2257 1848 2263
rect 1880 2257 1976 2263
rect 1992 2257 2104 2263
rect 2408 2257 2456 2263
rect 776 2237 936 2243
rect 1432 2237 1843 2243
rect 600 2217 1448 2223
rect 1592 2217 1736 2223
rect 1752 2217 1768 2223
rect 1837 2223 1843 2237
rect 1880 2237 2104 2243
rect 2120 2237 2168 2243
rect 2952 2237 3288 2243
rect 728 2197 808 2203
rect 1032 2197 1336 2203
rect 1512 2197 1528 2203
rect 1624 2197 1688 2203
rect 1837 2217 2120 2223
rect 2136 2217 2616 2223
rect 1864 2197 1880 2203
rect 1896 2197 1992 2203
rect 2232 2197 3000 2203
rect 728 2177 1000 2183
rect 1016 2177 1512 2183
rect 1528 2177 1576 2183
rect 1608 2177 1624 2183
rect 1640 2177 1752 2183
rect 1784 2177 1832 2183
rect 1944 2177 2680 2183
rect 2696 2177 2808 2183
rect 2824 2177 2888 2183
rect 2936 2177 2984 2183
rect 3000 2177 3320 2183
rect 584 2157 680 2163
rect 744 2157 1000 2163
rect 1016 2157 1048 2163
rect 1416 2157 1523 2163
rect 120 2137 136 2143
rect 152 2137 200 2143
rect 696 2137 728 2143
rect 840 2137 1128 2143
rect 1272 2137 1304 2143
rect 1464 2137 1480 2143
rect 1517 2143 1523 2157
rect 1544 2157 1640 2163
rect 1848 2157 2040 2163
rect 2392 2157 2456 2163
rect 2472 2157 2520 2163
rect 2536 2157 2664 2163
rect 2712 2157 2760 2163
rect 2808 2157 3016 2163
rect 3144 2157 3192 2163
rect 1517 2137 1576 2143
rect 1640 2137 1768 2143
rect 1784 2137 1960 2143
rect 2056 2137 2088 2143
rect 2456 2137 2536 2143
rect 2568 2137 2600 2143
rect 2680 2137 2760 2143
rect 2792 2137 2872 2143
rect 2904 2137 2968 2143
rect 3144 2137 3240 2143
rect 3256 2137 3640 2143
rect -51 2117 8 2123
rect 328 2117 360 2123
rect 376 2117 408 2123
rect 584 2117 680 2123
rect 904 2117 952 2123
rect 1048 2117 1096 2123
rect 1208 2117 1448 2123
rect 1592 2117 1608 2123
rect 1976 2117 2024 2123
rect 2072 2117 2088 2123
rect 2248 2117 2264 2123
rect 2280 2117 2312 2123
rect 2344 2117 2792 2123
rect 2824 2117 3112 2123
rect 1869 2108 1875 2112
rect 2221 2108 2227 2112
rect 648 2097 856 2103
rect 872 2097 952 2103
rect 968 2097 1096 2103
rect 1320 2097 1352 2103
rect 1480 2097 1608 2103
rect 2056 2097 2184 2103
rect 2616 2097 2696 2103
rect 2712 2097 2728 2103
rect 2776 2097 3032 2103
rect 3112 2097 3336 2103
rect 376 2077 1544 2083
rect 1560 2077 1720 2083
rect 1752 2077 2072 2083
rect 2408 2077 3368 2083
rect 680 2057 712 2063
rect 1320 2057 1736 2063
rect 2200 2057 2504 2063
rect 2936 2057 3160 2063
rect 3176 2057 3304 2063
rect 568 2037 728 2043
rect 872 2037 888 2043
rect 1016 2037 2296 2043
rect 2344 2037 2664 2043
rect 2840 2037 3016 2043
rect 3416 2037 3464 2043
rect 3480 2037 3528 2043
rect 1000 2017 2584 2023
rect 2600 2017 2696 2023
rect 2712 2017 2760 2023
rect 1080 1997 1416 2003
rect 1640 1997 1832 2003
rect 1864 1997 1960 2003
rect 2376 1997 2424 2003
rect 2504 1997 2648 2003
rect 2968 2017 3144 2023
rect 3192 2017 3560 2023
rect 3576 2017 3592 2023
rect 1288 1977 1736 1983
rect 1752 1977 2488 1983
rect 264 1957 488 1963
rect 504 1957 632 1963
rect 904 1957 1224 1963
rect 1256 1957 1464 1963
rect 1480 1957 1528 1963
rect 1560 1957 1896 1963
rect 2120 1957 2216 1963
rect 2232 1957 2408 1963
rect 2584 1957 2904 1963
rect 760 1937 1048 1943
rect 1112 1937 1304 1943
rect 1320 1937 1336 1943
rect 1688 1937 1848 1943
rect 1960 1937 1992 1943
rect 2008 1937 2200 1943
rect 2296 1937 2616 1943
rect 2664 1937 2968 1943
rect 3128 1937 3240 1943
rect 3256 1937 3576 1943
rect 232 1917 280 1923
rect 296 1917 312 1923
rect 392 1917 456 1923
rect 568 1917 696 1923
rect 744 1917 888 1923
rect 1160 1917 1176 1923
rect 1288 1917 1336 1923
rect 1368 1917 1448 1923
rect 1512 1917 2008 1923
rect 2232 1917 2280 1923
rect 2632 1917 2664 1923
rect 2696 1917 2824 1923
rect 2920 1917 2936 1923
rect 2952 1917 3016 1923
rect 3096 1917 3192 1923
rect 3224 1917 3240 1923
rect 3320 1917 3416 1923
rect 40 1897 72 1903
rect 104 1897 136 1903
rect 152 1897 184 1903
rect 312 1897 424 1903
rect 632 1897 984 1903
rect 1336 1897 1528 1903
rect 1560 1897 1592 1903
rect 1944 1897 2040 1903
rect 2488 1897 2568 1903
rect 2728 1897 2744 1903
rect 3016 1897 3096 1903
rect 3224 1897 3288 1903
rect 3304 1897 3480 1903
rect 3512 1897 3544 1903
rect 296 1877 328 1883
rect 344 1877 392 1883
rect 536 1877 632 1883
rect 664 1877 824 1883
rect 840 1877 856 1883
rect 888 1877 952 1883
rect 1032 1877 1096 1883
rect 1144 1877 1560 1883
rect 1592 1877 1720 1883
rect 1768 1877 1848 1883
rect 1864 1877 1960 1883
rect 2136 1877 2232 1883
rect 2296 1877 2344 1883
rect 2440 1877 2600 1883
rect 2648 1877 2696 1883
rect 2712 1877 2744 1883
rect 2808 1877 2888 1883
rect 2904 1877 2952 1883
rect 3080 1877 3112 1883
rect 3144 1877 3224 1883
rect 3240 1877 3272 1883
rect 3288 1877 3336 1883
rect 3368 1877 3384 1883
rect 653 1868 659 1872
rect 440 1857 616 1863
rect 824 1857 1016 1863
rect 1192 1857 1208 1863
rect 1256 1857 1368 1863
rect 1512 1857 1560 1863
rect 1624 1857 1784 1863
rect 1848 1857 1944 1863
rect 1965 1857 2019 1863
rect 360 1837 424 1843
rect 440 1837 552 1843
rect 600 1837 664 1843
rect 728 1837 1048 1843
rect 1176 1837 1192 1843
rect 1432 1837 1672 1843
rect 1965 1843 1971 1857
rect 1880 1837 1971 1843
rect 2013 1843 2019 1857
rect 2040 1857 2152 1863
rect 2712 1857 2728 1863
rect 2760 1857 2856 1863
rect 2888 1857 3224 1863
rect 3240 1857 3544 1863
rect 2541 1848 2547 1852
rect 2013 1837 2424 1843
rect 2568 1837 3160 1843
rect 3368 1837 3432 1843
rect 3512 1837 3592 1843
rect 1997 1828 2003 1832
rect 104 1817 600 1823
rect 616 1817 888 1823
rect 968 1817 1080 1823
rect 1448 1817 1464 1823
rect 1480 1817 1576 1823
rect 408 1797 504 1803
rect 525 1797 744 1803
rect -51 1777 328 1783
rect 525 1783 531 1797
rect 856 1797 920 1803
rect 936 1797 1080 1803
rect 1096 1797 1128 1803
rect 1144 1797 1416 1803
rect 2088 1817 3080 1823
rect 3112 1817 3160 1823
rect 3352 1817 3512 1823
rect 1880 1797 2264 1803
rect 2488 1797 2504 1803
rect 2520 1797 3048 1803
rect 3096 1797 3624 1803
rect 472 1777 531 1783
rect 680 1777 936 1783
rect 984 1777 1016 1783
rect 1304 1777 1352 1783
rect 1864 1777 1880 1783
rect 2013 1777 2024 1783
rect 2056 1777 2088 1783
rect 2472 1777 3128 1783
rect 3208 1777 3288 1783
rect 520 1757 840 1763
rect 1048 1757 1496 1763
rect 1544 1757 1576 1763
rect 1704 1757 1720 1763
rect 1960 1757 1976 1763
rect 2120 1757 2168 1763
rect 2184 1757 2328 1763
rect 2360 1757 2920 1763
rect 2936 1757 3240 1763
rect 344 1737 376 1743
rect 456 1737 552 1743
rect 712 1737 792 1743
rect 840 1737 1048 1743
rect 1240 1737 1256 1743
rect 1368 1737 1400 1743
rect 1416 1737 1624 1743
rect 1848 1737 1880 1743
rect 1912 1737 1928 1743
rect 1944 1737 2056 1743
rect 2584 1737 2600 1743
rect 2648 1737 2664 1743
rect 2728 1737 2776 1743
rect 3048 1737 3096 1743
rect 3256 1737 3272 1743
rect 3384 1737 3416 1743
rect 3560 1737 3640 1743
rect -51 1717 8 1723
rect 296 1717 456 1723
rect 616 1717 648 1723
rect 920 1717 1000 1723
rect 1048 1717 1192 1723
rect 1288 1717 1304 1723
rect 1661 1723 1667 1732
rect 1661 1717 1672 1723
rect 1709 1717 1715 1732
rect 1768 1717 1880 1723
rect 1896 1717 1944 1723
rect 1976 1717 1992 1723
rect 2120 1717 2216 1723
rect 2344 1717 2600 1723
rect 2616 1717 2648 1723
rect 2664 1717 2760 1723
rect 2776 1717 2792 1723
rect 2952 1717 2963 1723
rect 3032 1717 3080 1723
rect 3144 1717 3272 1723
rect 3288 1717 3336 1723
rect 280 1697 296 1703
rect 344 1697 424 1703
rect 584 1697 632 1703
rect 648 1697 680 1703
rect 728 1697 744 1703
rect 856 1697 1304 1703
rect 1352 1697 1432 1703
rect 1448 1697 2536 1703
rect 2552 1697 2808 1703
rect 2856 1697 2920 1703
rect 248 1677 1512 1683
rect 1560 1677 1576 1683
rect 1688 1677 1736 1683
rect 1896 1677 1960 1683
rect 2280 1677 2856 1683
rect 3192 1677 3400 1683
rect 536 1657 552 1663
rect 840 1657 1288 1663
rect 1384 1657 1720 1663
rect 2024 1657 2248 1663
rect 2536 1657 3256 1663
rect 632 1637 696 1643
rect 760 1637 872 1643
rect 1224 1637 1352 1643
rect 1576 1637 2024 1643
rect 2056 1637 2136 1643
rect 2264 1637 2296 1643
rect 2360 1637 2376 1643
rect 2680 1637 2808 1643
rect 2840 1637 2856 1643
rect 2952 1637 2984 1643
rect 2381 1628 2387 1632
rect 344 1617 744 1623
rect 872 1617 936 1623
rect 968 1617 1064 1623
rect 1080 1617 1896 1623
rect 2104 1617 2152 1623
rect 2280 1617 2344 1623
rect 888 1597 1064 1603
rect 1080 1597 1240 1603
rect 1368 1597 1592 1603
rect 1608 1597 1640 1603
rect 1672 1597 2232 1603
rect 3336 1597 3464 1603
rect 392 1577 600 1583
rect 776 1577 968 1583
rect 1064 1577 3256 1583
rect 3272 1577 3432 1583
rect 440 1557 536 1563
rect 552 1557 616 1563
rect 632 1557 1144 1563
rect 1160 1557 1240 1563
rect 1256 1557 1304 1563
rect 1576 1557 1816 1563
rect 1944 1557 2056 1563
rect 2269 1557 2408 1563
rect 328 1537 728 1543
rect 776 1537 968 1543
rect 984 1537 1112 1543
rect 1128 1537 1160 1543
rect 1176 1537 1192 1543
rect 1304 1537 1480 1543
rect 1672 1537 1704 1543
rect 1736 1537 1752 1543
rect 1800 1537 1864 1543
rect 2269 1543 2275 1557
rect 2424 1557 2456 1563
rect 2744 1557 3032 1563
rect 3304 1557 3320 1563
rect 1912 1537 2275 1543
rect 2376 1537 2840 1543
rect 3320 1537 3368 1543
rect 184 1517 552 1523
rect 568 1517 632 1523
rect 648 1517 728 1523
rect 744 1517 856 1523
rect 936 1517 1176 1523
rect 1304 1517 1400 1523
rect 1421 1517 2104 1523
rect 104 1497 120 1503
rect 168 1497 184 1503
rect 216 1497 227 1503
rect 264 1497 280 1503
rect 504 1497 520 1503
rect 536 1497 824 1503
rect 888 1497 1016 1503
rect 1032 1497 1112 1503
rect 1256 1497 1320 1503
rect 1421 1503 1427 1517
rect 2216 1517 2312 1523
rect 2456 1517 2552 1523
rect 2568 1517 2600 1523
rect 3032 1517 3112 1523
rect 3304 1517 3320 1523
rect 3485 1523 3491 1532
rect 3400 1517 3576 1523
rect 1336 1497 1427 1503
rect 1528 1497 1576 1503
rect 1672 1497 1784 1503
rect 1864 1497 1923 1503
rect 248 1477 264 1483
rect 472 1477 536 1483
rect 552 1477 632 1483
rect 696 1477 936 1483
rect 968 1477 1000 1483
rect 1016 1477 1128 1483
rect 1304 1477 1320 1483
rect 1352 1477 1496 1483
rect 1544 1477 1560 1483
rect 1672 1477 1688 1483
rect 1752 1477 1896 1483
rect 1917 1483 1923 1497
rect 1944 1497 2120 1503
rect 2136 1497 2392 1503
rect 2440 1497 2632 1503
rect 2840 1497 3048 1503
rect 3144 1497 3208 1503
rect 3224 1497 3288 1503
rect 3320 1497 3608 1503
rect 1917 1477 1928 1483
rect 2024 1477 2088 1483
rect 2104 1477 2136 1483
rect 2168 1477 2435 1483
rect 136 1457 152 1463
rect 168 1457 328 1463
rect 488 1457 536 1463
rect 584 1457 616 1463
rect 888 1457 1112 1463
rect 1144 1457 1704 1463
rect 1768 1457 1848 1463
rect 1880 1457 1976 1463
rect 2088 1457 2184 1463
rect 2248 1457 2280 1463
rect 2301 1457 2312 1463
rect 2344 1457 2376 1463
rect 2429 1463 2435 1477
rect 2456 1477 2488 1483
rect 2552 1477 2568 1483
rect 2792 1477 3000 1483
rect 3032 1477 3144 1483
rect 3448 1477 3512 1483
rect 3528 1477 3624 1483
rect 2429 1457 2552 1463
rect 2696 1457 2856 1463
rect 3144 1457 3384 1463
rect 3496 1457 3544 1463
rect 72 1437 504 1443
rect 536 1437 664 1443
rect 840 1437 1272 1443
rect 1448 1437 1560 1443
rect 1624 1437 1640 1443
rect 1704 1437 1992 1443
rect 2136 1437 2168 1443
rect 2184 1437 2200 1443
rect 2360 1437 2504 1443
rect 2520 1437 2536 1443
rect 2904 1437 2984 1443
rect 3000 1437 3320 1443
rect 3512 1437 3560 1443
rect 360 1417 472 1423
rect 488 1417 584 1423
rect 616 1417 888 1423
rect 920 1417 1160 1423
rect 1176 1417 1208 1423
rect 1240 1417 1640 1423
rect 328 1397 568 1403
rect 728 1397 808 1403
rect 1016 1397 1096 1403
rect 1336 1397 1352 1403
rect 1640 1397 1720 1403
rect 1864 1417 1880 1423
rect 1976 1417 1992 1423
rect 2200 1417 2328 1423
rect 2440 1417 2568 1423
rect 2584 1417 2744 1423
rect 2760 1417 2952 1423
rect 2968 1417 3096 1423
rect 3560 1417 3576 1423
rect 2072 1397 2392 1403
rect 2600 1397 2904 1403
rect 232 1377 456 1383
rect 504 1377 520 1383
rect 712 1377 1272 1383
rect 1288 1377 1400 1383
rect 1416 1377 1528 1383
rect 1544 1377 2072 1383
rect 2168 1377 2216 1383
rect 2232 1377 2360 1383
rect 2376 1377 2499 1383
rect 200 1357 328 1363
rect 504 1357 552 1363
rect 632 1357 648 1363
rect 669 1357 728 1363
rect 152 1337 280 1343
rect 312 1337 344 1343
rect 456 1337 488 1343
rect 669 1343 675 1357
rect 744 1357 872 1363
rect 952 1357 968 1363
rect 1160 1357 1192 1363
rect 1240 1357 1320 1363
rect 1400 1357 1864 1363
rect 1896 1357 1928 1363
rect 1976 1357 2040 1363
rect 2120 1357 2392 1363
rect 2408 1357 2472 1363
rect 2493 1363 2499 1377
rect 2520 1377 2616 1383
rect 2632 1377 2968 1383
rect 2984 1377 3000 1383
rect 3320 1377 3448 1383
rect 2493 1357 2520 1363
rect 2584 1357 2696 1363
rect 2728 1357 2792 1363
rect 3240 1357 3368 1363
rect 3384 1357 3432 1363
rect 1101 1348 1107 1352
rect 1341 1348 1347 1352
rect 552 1337 675 1343
rect 712 1337 744 1343
rect 872 1337 952 1343
rect 1128 1337 1288 1343
rect 1352 1337 1416 1343
rect 1480 1337 1560 1343
rect 1768 1337 1928 1343
rect 1960 1337 2040 1343
rect 2216 1337 2328 1343
rect 2360 1337 2520 1343
rect 2536 1337 2760 1343
rect 2824 1337 2920 1343
rect 3112 1337 3208 1343
rect 3224 1337 3240 1343
rect 3256 1337 3624 1343
rect -51 1317 136 1323
rect 264 1317 616 1323
rect 632 1317 888 1323
rect 1032 1317 1096 1323
rect 1117 1317 1208 1323
rect 296 1297 456 1303
rect 648 1297 680 1303
rect 728 1297 760 1303
rect 936 1297 1000 1303
rect 1117 1303 1123 1317
rect 1288 1317 1768 1323
rect 1880 1317 1928 1323
rect 1944 1317 1960 1323
rect 2040 1317 2280 1323
rect 2296 1317 2360 1323
rect 2392 1317 2456 1323
rect 2568 1317 2648 1323
rect 2728 1317 3000 1323
rect 3064 1317 3304 1323
rect 3368 1317 3384 1323
rect 3400 1317 3528 1323
rect 2477 1308 2483 1312
rect 2493 1308 2499 1312
rect 1016 1297 1123 1303
rect 1336 1297 1480 1303
rect 1624 1297 2056 1303
rect 2072 1297 2136 1303
rect 2184 1297 2232 1303
rect 2280 1297 2296 1303
rect 2312 1297 2328 1303
rect 2344 1297 2392 1303
rect 2536 1297 2600 1303
rect 2648 1297 2728 1303
rect 2744 1297 2760 1303
rect 2888 1297 2920 1303
rect 3288 1297 3336 1303
rect 3448 1297 3512 1303
rect 893 1288 899 1292
rect 1149 1288 1155 1292
rect 424 1277 616 1283
rect 1528 1277 1704 1283
rect 1720 1277 2632 1283
rect 2648 1277 2904 1283
rect 2952 1277 2968 1283
rect 3000 1277 3080 1283
rect 3144 1277 3208 1283
rect 3256 1277 3288 1283
rect 3432 1277 3496 1283
rect 3528 1277 3592 1283
rect 456 1257 1032 1263
rect 1192 1257 1608 1263
rect 1624 1257 2120 1263
rect 2136 1257 2696 1263
rect 2728 1257 2920 1263
rect 2952 1257 3000 1263
rect 3016 1257 3416 1263
rect 312 1237 648 1243
rect 728 1237 808 1243
rect 1048 1237 1112 1243
rect 1208 1237 1224 1243
rect 1688 1237 1752 1243
rect 1912 1237 2024 1243
rect 2088 1237 2936 1243
rect 3128 1237 3464 1243
rect 184 1217 424 1223
rect 88 1197 536 1203
rect 1112 1217 1144 1223
rect 1160 1217 1608 1223
rect 1880 1217 2104 1223
rect 2152 1217 2648 1223
rect 1272 1197 1784 1203
rect 1848 1197 1864 1203
rect 1896 1197 1960 1203
rect 2008 1197 2328 1203
rect 2424 1197 2440 1203
rect 2872 1197 2888 1203
rect 3016 1197 3288 1203
rect 360 1177 696 1183
rect 712 1177 888 1183
rect 1336 1177 1352 1183
rect 1400 1177 1688 1183
rect 1800 1177 2824 1183
rect 2840 1177 3144 1183
rect 3192 1177 3512 1183
rect -51 1157 8 1163
rect 24 1157 72 1163
rect 88 1157 600 1163
rect 1096 1157 1352 1163
rect 1448 1157 2376 1163
rect 2392 1157 2552 1163
rect 2573 1157 2888 1163
rect 408 1137 696 1143
rect 712 1137 904 1143
rect 1240 1137 1272 1143
rect 1480 1137 1592 1143
rect 1848 1137 1912 1143
rect 1928 1137 1992 1143
rect 2216 1137 2504 1143
rect 2573 1143 2579 1157
rect 2904 1157 3240 1163
rect 2520 1137 2579 1143
rect 2616 1137 2680 1143
rect 2696 1137 2744 1143
rect 264 1117 328 1123
rect 424 1117 504 1123
rect 648 1117 840 1123
rect 856 1117 1720 1123
rect 1736 1117 2344 1123
rect 2504 1117 2584 1123
rect 2600 1117 2632 1123
rect 2808 1117 2920 1123
rect 3048 1117 3160 1123
rect 3224 1117 3240 1123
rect 3304 1117 3560 1123
rect 248 1097 344 1103
rect 504 1097 520 1103
rect 808 1097 968 1103
rect 1000 1097 1416 1103
rect 1736 1097 1752 1103
rect 1864 1097 1912 1103
rect 1960 1097 2232 1103
rect 2296 1097 2312 1103
rect 2344 1097 2440 1103
rect 2552 1097 2760 1103
rect 2776 1097 2872 1103
rect 3080 1097 3096 1103
rect 3112 1097 3336 1103
rect 3368 1097 3416 1103
rect 3512 1097 3544 1103
rect -51 1077 24 1083
rect 40 1077 88 1083
rect 136 1077 216 1083
rect 232 1077 280 1083
rect 312 1077 392 1083
rect 472 1077 760 1083
rect 904 1077 968 1083
rect 1048 1077 1240 1083
rect 1416 1077 1432 1083
rect 1496 1077 1512 1083
rect 1720 1077 1736 1083
rect 1768 1077 1848 1083
rect 1912 1077 1976 1083
rect 2173 1077 2184 1083
rect 2232 1077 2280 1083
rect 2344 1077 2648 1083
rect 2680 1077 2952 1083
rect 3144 1077 3432 1083
rect 3480 1077 3512 1083
rect 72 1057 312 1063
rect 760 1057 1144 1063
rect 1224 1057 1240 1063
rect 1272 1057 1352 1063
rect 1528 1057 1864 1063
rect 1896 1057 1992 1063
rect 2056 1057 2200 1063
rect 2312 1057 2408 1063
rect 2536 1057 2568 1063
rect 2600 1057 2728 1063
rect 2760 1057 2856 1063
rect 2872 1057 3224 1063
rect 888 1037 1192 1043
rect 1208 1037 1416 1043
rect 1432 1037 1592 1043
rect 1773 1037 2456 1043
rect 680 1017 1016 1023
rect 1080 1017 1544 1023
rect 1773 1023 1779 1037
rect 2632 1037 2904 1043
rect 3016 1037 3144 1043
rect 1560 1017 1779 1023
rect 216 997 280 1003
rect 344 997 392 1003
rect 520 997 728 1003
rect 936 997 1224 1003
rect 1288 997 1464 1003
rect 1864 1017 1912 1023
rect 1992 1017 2040 1023
rect 2056 1017 2392 1023
rect 2424 1017 2616 1023
rect 2632 1017 3016 1023
rect 3272 1017 3528 1023
rect 1944 997 2488 1003
rect 2504 997 2568 1003
rect 2824 997 3272 1003
rect 3533 988 3539 992
rect -51 977 72 983
rect 88 977 136 983
rect 168 977 328 983
rect 680 977 867 983
rect 136 957 200 963
rect 216 957 344 963
rect 376 957 552 963
rect 696 957 744 963
rect 861 963 867 977
rect 1325 977 1336 983
rect 1656 977 1720 983
rect 1736 977 1752 983
rect 1800 977 1832 983
rect 2184 977 2680 983
rect 3128 977 3304 983
rect 861 957 888 963
rect 904 957 1032 963
rect 1064 957 1096 963
rect 1576 957 1624 963
rect 1640 957 1944 963
rect 1960 957 2024 963
rect 2136 957 2248 963
rect 2141 948 2147 957
rect 2264 957 2344 963
rect 2568 957 2632 963
rect 2696 957 2728 963
rect 2792 957 3171 963
rect 104 937 152 943
rect 200 937 472 943
rect 600 937 632 943
rect 648 937 760 943
rect 1080 937 1224 943
rect 1368 937 1704 943
rect 1720 937 2088 943
rect 2200 937 2408 943
rect 2648 937 2696 943
rect 2968 937 3016 943
rect 3032 937 3048 943
rect 3080 937 3128 943
rect 3165 943 3171 957
rect 3192 957 3256 963
rect 3544 957 3592 963
rect 3165 937 3224 943
rect 3320 937 3336 943
rect 3352 937 3368 943
rect 3464 937 3480 943
rect 3496 937 3544 943
rect 973 928 979 932
rect -51 917 152 923
rect 456 917 920 923
rect 1192 917 1304 923
rect 1400 917 1432 923
rect 1464 917 1736 923
rect 1752 917 1864 923
rect 1896 917 1912 923
rect 1960 917 2040 923
rect 2088 917 2168 923
rect 2184 917 2200 923
rect 2360 917 2536 923
rect 2552 917 2872 923
rect 2888 917 3032 923
rect 3224 917 3288 923
rect 3672 917 3715 923
rect 200 897 216 903
rect 248 897 264 903
rect 520 897 680 903
rect 760 897 808 903
rect 920 897 936 903
rect 1000 897 1016 903
rect 1048 897 1064 903
rect 1096 897 1176 903
rect 1224 897 1272 903
rect 1592 897 1640 903
rect 1912 897 2008 903
rect 2120 897 2168 903
rect 2440 897 2600 903
rect 2616 897 2792 903
rect 3288 897 3336 903
rect 1405 888 1411 892
rect 152 877 1080 883
rect 1096 877 1384 883
rect 1512 877 2120 883
rect 2136 877 2296 883
rect 2328 877 3080 883
rect 664 857 1048 863
rect 1064 857 1176 863
rect 1400 857 1576 863
rect 1624 857 1656 863
rect 1736 857 1880 863
rect 1928 857 2152 863
rect 2200 857 3096 863
rect 3112 857 3144 863
rect 376 837 680 843
rect 1144 837 2088 843
rect 2104 837 2408 843
rect 2424 837 2664 843
rect 2728 837 2904 843
rect 2920 837 3352 843
rect 3416 837 3427 843
rect 632 817 648 823
rect 888 817 1288 823
rect 1432 817 1576 823
rect 1688 817 1816 823
rect 1912 817 2008 823
rect 1112 797 1560 803
rect 1640 797 2424 803
rect 2440 797 2792 803
rect 3272 817 3512 823
rect 3016 797 3032 803
rect 3048 797 3496 803
rect 701 788 707 792
rect 344 777 360 783
rect 600 777 680 783
rect 728 777 824 783
rect 856 777 904 783
rect 920 777 1096 783
rect 1160 777 1240 783
rect 1384 777 1688 783
rect 1832 777 2216 783
rect 2552 777 2792 783
rect 2968 777 2984 783
rect 3000 777 3144 783
rect 3160 777 3480 783
rect 3496 777 3512 783
rect 3528 777 3592 783
rect 3608 777 3640 783
rect 664 757 1672 763
rect 1688 757 2136 763
rect 2168 757 2632 763
rect 2648 757 3160 763
rect 296 737 392 743
rect 536 737 632 743
rect 680 737 920 743
rect 1208 737 1608 743
rect 1720 737 1912 743
rect 1944 737 1976 743
rect 2136 737 2344 743
rect 2376 737 2408 743
rect 2424 737 2552 743
rect 2616 737 3064 743
rect 344 717 600 723
rect 616 717 648 723
rect 760 717 776 723
rect 792 717 856 723
rect 872 717 2024 723
rect 2088 717 2168 723
rect 2248 717 2296 723
rect 2312 717 2328 723
rect 2344 717 2376 723
rect 2504 717 2520 723
rect 2536 717 3000 723
rect 3592 717 3715 723
rect 221 708 227 712
rect 472 697 488 703
rect 520 697 664 703
rect 872 697 888 703
rect 904 697 920 703
rect 936 697 1064 703
rect 1272 697 1720 703
rect 1848 697 1944 703
rect 2232 697 2312 703
rect 2408 697 2536 703
rect 2728 697 2744 703
rect 168 677 296 683
rect 392 677 424 683
rect 440 677 1048 683
rect 1064 677 1128 683
rect 1352 677 1368 683
rect 1432 677 1480 683
rect 1672 677 1896 683
rect 1912 677 2008 683
rect 2040 677 2488 683
rect 2520 677 2680 683
rect 2696 677 2728 683
rect 2888 677 2904 683
rect 2920 677 3064 683
rect 3080 677 3096 683
rect 3112 677 3192 683
rect 3208 677 3224 683
rect 3240 677 3320 683
rect 3336 677 3352 683
rect 3368 677 3384 683
rect 3400 677 3416 683
rect 3480 677 3544 683
rect 1565 668 1571 672
rect 216 657 280 663
rect 392 657 408 663
rect 424 657 440 663
rect 456 657 552 663
rect 920 657 952 663
rect 1304 657 1368 663
rect 1384 657 1544 663
rect 1784 657 1960 663
rect 1992 657 2440 663
rect 2616 657 2632 663
rect 2664 657 3144 663
rect 3160 657 3176 663
rect 3192 657 3384 663
rect 936 637 1027 643
rect 600 617 744 623
rect 920 617 984 623
rect 1021 623 1027 637
rect 1224 637 1592 643
rect 1640 637 1880 643
rect 2152 637 2184 643
rect 2200 637 2616 643
rect 2648 637 2664 643
rect 2696 637 3256 643
rect 1021 617 1528 623
rect 72 597 344 603
rect 360 597 456 603
rect 472 597 584 603
rect 920 597 1272 603
rect 1288 597 1528 603
rect 1848 617 2104 623
rect 1864 597 2200 603
rect 2488 597 2872 603
rect 152 577 232 583
rect 248 577 312 583
rect 552 577 696 583
rect 744 577 792 583
rect 1112 577 1192 583
rect 1336 577 1352 583
rect 1512 577 1704 583
rect 1752 577 1832 583
rect 1848 577 1864 583
rect 2072 577 2184 583
rect 2216 577 2632 583
rect 408 557 424 563
rect 504 557 1448 563
rect 1464 557 1816 563
rect 2040 557 2424 563
rect 2552 557 2952 563
rect 312 537 504 543
rect 600 537 872 543
rect 952 537 968 543
rect 984 537 1096 543
rect 1117 537 1475 543
rect -51 517 8 523
rect 24 517 168 523
rect 184 517 248 523
rect 488 517 520 523
rect 632 517 680 523
rect 712 517 728 523
rect 776 517 824 523
rect 1000 517 1048 523
rect 1117 523 1123 537
rect 1096 517 1123 523
rect 1400 517 1448 523
rect 1469 523 1475 537
rect 1592 537 1603 543
rect 1736 537 1800 543
rect 1832 537 2136 543
rect 2152 537 2280 543
rect 2968 537 2984 543
rect 3000 537 3064 543
rect 3080 537 3112 543
rect 3128 537 3144 543
rect 3160 537 3368 543
rect 3384 537 3448 543
rect 3464 537 3480 543
rect 3592 537 3608 543
rect 1469 517 2024 523
rect 2056 517 2168 523
rect 2536 517 2568 523
rect 2712 517 2728 523
rect 3560 517 3608 523
rect 3672 517 3715 523
rect 88 497 152 503
rect 200 497 264 503
rect 456 497 488 503
rect 520 497 952 503
rect 968 497 1112 503
rect 1165 503 1171 512
rect 1309 508 1315 512
rect 1160 497 1171 503
rect 1384 497 1416 503
rect 1464 497 1544 503
rect 1608 497 1640 503
rect 1688 497 1832 503
rect 2040 497 2056 503
rect 2184 497 2904 503
rect 40 477 56 483
rect 104 477 136 483
rect 152 477 200 483
rect 216 477 232 483
rect 248 477 280 483
rect 376 477 584 483
rect 696 477 712 483
rect 760 477 776 483
rect 792 477 840 483
rect 984 477 1464 483
rect 1512 477 1832 483
rect 1912 477 2008 483
rect 2088 477 2568 483
rect 2600 477 3192 483
rect 3208 477 3224 483
rect 3240 477 3256 483
rect 3304 477 3352 483
rect 72 457 120 463
rect 264 457 328 463
rect 344 457 856 463
rect 1144 457 1288 463
rect 1592 457 1656 463
rect 1736 457 2376 463
rect 648 437 680 443
rect 1768 437 2120 443
rect 2232 437 2328 443
rect 2344 437 2696 443
rect 1032 417 1048 423
rect 1064 417 1352 423
rect 1912 417 2088 423
rect 1208 397 1272 403
rect 1336 397 1736 403
rect 1848 397 2056 403
rect 3496 397 3560 403
rect 1272 377 1288 383
rect 1304 377 1512 383
rect 1736 377 2152 383
rect 2776 377 2808 383
rect 2824 377 2856 383
rect 2872 377 2888 383
rect 584 357 1144 363
rect 1176 357 1208 363
rect 1224 357 1400 363
rect 1448 357 1752 363
rect 1976 357 2040 363
rect 120 337 248 343
rect 456 337 472 343
rect 616 337 1448 343
rect 1544 337 1640 343
rect 1656 337 1896 343
rect 1928 337 1960 343
rect 200 317 296 323
rect 312 317 408 323
rect 936 317 1304 323
rect 1352 317 1464 323
rect 1512 317 1560 323
rect 1704 317 1752 323
rect 1864 317 1944 323
rect 3672 317 3715 323
rect -51 297 24 303
rect 40 297 88 303
rect 120 297 152 303
rect 264 297 280 303
rect 472 297 536 303
rect 552 297 648 303
rect 664 297 696 303
rect 808 297 872 303
rect 1000 297 1064 303
rect 1128 297 1192 303
rect 1384 297 1416 303
rect 1480 297 1512 303
rect 1560 297 1608 303
rect 1672 297 1720 303
rect 1880 297 1912 303
rect 1960 297 2024 303
rect 2088 297 2120 303
rect 2584 297 3048 303
rect 3384 297 3512 303
rect 88 277 168 283
rect 216 277 296 283
rect 856 277 1064 283
rect 1080 277 1091 283
rect 1112 277 1384 283
rect 1400 277 1704 283
rect 1736 277 1880 283
rect 2056 277 2104 283
rect 2120 277 2264 283
rect 24 257 72 263
rect 88 257 216 263
rect 296 257 424 263
rect 760 257 1016 263
rect 1416 257 1624 263
rect 1704 257 1816 263
rect 2408 257 2552 263
rect 152 237 200 243
rect 744 237 1048 243
rect 1064 237 1096 243
rect 1288 237 1432 243
rect 1560 237 1640 243
rect 1656 237 1784 243
rect 2984 237 3032 243
rect 3416 237 3448 243
rect 3464 237 3480 243
rect 376 217 616 223
rect 632 217 1112 223
rect 1160 217 1320 223
rect 1336 217 1752 223
rect 264 197 360 203
rect 408 197 888 203
rect 1160 197 1272 203
rect 1416 197 1432 203
rect 1688 197 1768 203
rect 1912 217 1928 223
rect 1944 217 1992 223
rect 1992 197 2024 203
rect 248 177 296 183
rect 312 177 392 183
rect 504 177 552 183
rect 568 177 632 183
rect 664 177 680 183
rect 696 177 968 183
rect 1000 177 1096 183
rect 1112 177 1400 183
rect 1416 177 1528 183
rect 1576 177 1608 183
rect 1629 177 1640 183
rect 1736 177 1976 183
rect 2024 177 2040 183
rect 2056 177 2088 183
rect 2296 177 2328 183
rect 2344 177 2360 183
rect 2376 177 2392 183
rect 2408 177 2488 183
rect 2504 177 2536 183
rect 2552 177 2568 183
rect 3096 177 3112 183
rect 3128 177 3160 183
rect 3192 177 3224 183
rect 840 157 968 163
rect 984 157 1160 163
rect 1448 157 1464 163
rect 1480 157 2760 163
rect 136 137 168 143
rect 984 137 1032 143
rect 1080 137 1144 143
rect 1208 137 1240 143
rect 1256 137 1384 143
rect 1624 137 1656 143
rect 1768 137 1912 143
rect 2072 137 2088 143
rect 2104 137 2120 143
rect 2136 137 2216 143
rect 2232 137 2248 143
rect 2632 137 2648 143
rect 2664 137 2712 143
rect 2776 137 2792 143
rect 2808 137 2904 143
rect 2920 137 2936 143
rect 3320 137 3512 143
rect 56 117 88 123
rect 104 117 120 123
rect 136 117 200 123
rect 232 117 280 123
rect 344 117 440 123
rect 456 117 520 123
rect 712 117 744 123
rect 904 117 1256 123
rect 1272 117 1352 123
rect 1368 117 1528 123
rect 1544 117 1560 123
rect 1576 117 1736 123
rect 1880 117 1928 123
rect 2376 117 2504 123
rect 2712 117 2728 123
rect 2760 117 2856 123
rect 3304 117 3336 123
rect 200 97 264 103
rect 424 97 616 103
rect 632 97 856 103
rect 872 97 936 103
rect 968 97 1016 103
rect 1256 97 1272 103
rect 1368 97 1480 103
rect 1544 97 1608 103
rect 1624 97 1688 103
rect 1736 97 1816 103
rect 1864 97 1880 103
rect 1896 97 1976 103
rect 216 77 296 83
rect 568 77 1032 83
rect 1048 77 1208 83
rect 1528 77 1624 83
rect 184 57 328 63
rect 904 57 984 63
rect 1048 37 1768 43
rect 1336 17 1368 23
rect 1688 17 1720 23
rect 2872 17 2888 23
rect 3032 17 3048 23
<< m4contact >>
rect 766 2402 794 2418
rect 2814 2402 2842 2418
rect 1512 2312 1528 2328
rect 456 2272 472 2288
rect 1432 2272 1448 2288
rect 1896 2272 1912 2288
rect 2072 2272 2088 2288
rect 3272 2272 3288 2288
rect 1064 2252 1080 2268
rect 1288 2252 1304 2268
rect 1848 2252 1864 2268
rect 584 2212 600 2228
rect 1864 2232 1880 2248
rect 2568 2232 2584 2248
rect 1790 2202 1818 2218
rect 2616 2212 2632 2228
rect 1848 2192 1864 2208
rect 1880 2192 1896 2208
rect 1576 2172 1592 2188
rect 1752 2172 1768 2188
rect 728 2132 744 2148
rect 1320 2132 1336 2148
rect 1656 2152 1672 2168
rect 1672 2152 1688 2168
rect 2760 2152 2776 2168
rect 2792 2152 2808 2168
rect 1624 2132 1640 2148
rect 1976 2132 1992 2148
rect 2248 2132 2264 2148
rect 2648 2132 2664 2148
rect 2776 2132 2792 2148
rect 2888 2132 2904 2148
rect 1864 2112 1880 2128
rect 1960 2112 1976 2128
rect 2056 2112 2072 2128
rect 2264 2112 2280 2128
rect 2328 2112 2344 2128
rect 2792 2112 2808 2128
rect 952 2092 968 2108
rect 1304 2092 1320 2108
rect 1608 2092 1624 2108
rect 1928 2092 1944 2108
rect 2216 2092 2232 2108
rect 1096 2052 1112 2068
rect 2504 2052 2520 2068
rect 3304 2052 3320 2068
rect 552 2032 568 2048
rect 856 2032 872 2048
rect 2328 2032 2344 2048
rect 3016 2032 3032 2048
rect 3384 2032 3400 2048
rect 766 2002 794 2018
rect 2696 2012 2712 2028
rect 1960 1992 1976 2008
rect 2360 1992 2376 2008
rect 2814 2002 2842 2018
rect 1736 1972 1752 1988
rect 1224 1952 1240 1968
rect 2216 1952 2232 1968
rect 2568 1952 2584 1968
rect 1048 1932 1064 1948
rect 1336 1932 1352 1948
rect 1848 1932 1864 1948
rect 3240 1932 3256 1948
rect 328 1912 344 1928
rect 1496 1912 1512 1928
rect 2200 1912 2216 1928
rect 2296 1912 2312 1928
rect 2680 1912 2696 1928
rect 2904 1912 2920 1928
rect 3208 1912 3224 1928
rect 296 1892 312 1908
rect 616 1892 632 1908
rect 1528 1892 1544 1908
rect 1816 1892 1832 1908
rect 2136 1892 2152 1908
rect 2184 1892 2200 1908
rect 2232 1892 2264 1908
rect 2344 1892 2360 1908
rect 2712 1892 2728 1908
rect 3208 1892 3224 1908
rect 3496 1892 3512 1908
rect 632 1872 664 1888
rect 872 1872 888 1888
rect 1096 1872 1112 1888
rect 1576 1872 1592 1888
rect 2120 1872 2136 1888
rect 2232 1872 2248 1888
rect 2280 1872 2296 1888
rect 2600 1872 2616 1888
rect 3048 1872 3064 1888
rect 3352 1872 3368 1888
rect 3464 1872 3480 1888
rect 424 1852 440 1868
rect 616 1852 632 1868
rect 696 1852 712 1868
rect 1240 1852 1256 1868
rect 552 1832 568 1848
rect 1128 1832 1144 1848
rect 1192 1832 1208 1848
rect 1992 1832 2008 1848
rect 2024 1852 2040 1868
rect 2536 1852 2552 1868
rect 2600 1852 2616 1868
rect 2696 1852 2712 1868
rect 2872 1852 2888 1868
rect 2520 1832 2536 1848
rect 2552 1832 2568 1848
rect 888 1812 904 1828
rect 1432 1812 1448 1828
rect 1790 1802 1818 1818
rect 3096 1812 3112 1828
rect 2264 1792 2280 1808
rect 2472 1792 2488 1808
rect 936 1772 952 1788
rect 1848 1772 1864 1788
rect 2024 1772 2040 1788
rect 2088 1772 2104 1788
rect 3192 1772 3208 1788
rect 1032 1752 1048 1768
rect 1720 1752 1736 1768
rect 1944 1752 1960 1768
rect 2008 1752 2024 1768
rect 2072 1752 2088 1768
rect 2104 1752 2120 1768
rect 2328 1752 2360 1768
rect 792 1732 808 1748
rect 1272 1732 1288 1748
rect 1352 1732 1368 1748
rect 1704 1732 1720 1748
rect 1896 1732 1912 1748
rect 2504 1732 2520 1748
rect 2552 1732 2568 1748
rect 2632 1732 2648 1748
rect 3544 1732 3560 1748
rect 456 1712 472 1728
rect 1208 1712 1224 1728
rect 1384 1712 1400 1728
rect 1672 1712 1688 1728
rect 1944 1712 1976 1728
rect 2008 1712 2024 1728
rect 2040 1712 2056 1728
rect 2312 1712 2328 1728
rect 2936 1712 2952 1728
rect 3528 1712 3544 1728
rect 1304 1692 1320 1708
rect 1336 1692 1352 1708
rect 2824 1692 2840 1708
rect 2920 1692 2936 1708
rect 3304 1692 3320 1708
rect 1544 1672 1560 1688
rect 1672 1672 1688 1688
rect 1960 1672 1976 1688
rect 2264 1672 2280 1688
rect 1304 1652 1320 1668
rect 1976 1652 2008 1668
rect 2376 1632 2392 1648
rect 2808 1632 2840 1648
rect 3128 1632 3144 1648
rect 744 1612 760 1628
rect 766 1602 794 1618
rect 936 1612 952 1628
rect 2088 1612 2104 1628
rect 1592 1592 1608 1608
rect 1656 1592 1672 1608
rect 2814 1602 2842 1618
rect 3144 1612 3160 1628
rect 3320 1592 3336 1608
rect 296 1572 312 1588
rect 760 1572 776 1588
rect 3256 1572 3272 1588
rect 616 1552 632 1568
rect 1240 1552 1256 1568
rect 1432 1552 1448 1568
rect 1928 1552 1944 1568
rect 728 1532 744 1548
rect 1288 1532 1304 1548
rect 1768 1532 1784 1548
rect 3288 1552 3304 1568
rect 2360 1532 2376 1548
rect 3000 1532 3016 1548
rect 3304 1532 3320 1548
rect 3448 1532 3464 1548
rect 3576 1532 3592 1548
rect 120 1492 136 1508
rect 200 1492 216 1508
rect 824 1492 840 1508
rect 1176 1492 1192 1508
rect 1320 1492 1336 1508
rect 2440 1512 2456 1528
rect 2600 1512 2616 1528
rect 2616 1512 2632 1528
rect 1448 1492 1464 1508
rect 1656 1492 1672 1508
rect 1832 1492 1848 1508
rect 1848 1492 1864 1508
rect 632 1472 648 1488
rect 936 1472 952 1488
rect 1320 1472 1336 1488
rect 1688 1472 1704 1488
rect 1896 1472 1912 1488
rect 1928 1492 1944 1508
rect 2392 1492 2408 1508
rect 2632 1492 2648 1508
rect 2008 1472 2024 1488
rect 344 1452 376 1468
rect 1112 1452 1128 1468
rect 1848 1452 1880 1468
rect 2072 1452 2088 1468
rect 2216 1452 2232 1468
rect 2312 1452 2328 1468
rect 2328 1452 2344 1468
rect 3016 1472 3032 1488
rect 3288 1472 3304 1488
rect 2568 1452 2584 1468
rect 824 1432 840 1448
rect 1560 1432 1576 1448
rect 1672 1432 1688 1448
rect 2344 1432 2360 1448
rect 2536 1432 2552 1448
rect 2616 1432 2632 1448
rect 584 1412 600 1428
rect 888 1412 904 1428
rect 1640 1412 1656 1428
rect 1288 1392 1304 1408
rect 1608 1392 1624 1408
rect 1720 1392 1736 1408
rect 1790 1402 1818 1418
rect 1848 1412 1864 1428
rect 1960 1412 1976 1428
rect 2136 1412 2152 1428
rect 2424 1412 2440 1428
rect 1912 1392 1928 1408
rect 1944 1392 1960 1408
rect 2056 1392 2072 1408
rect 3400 1392 3416 1408
rect 1272 1372 1288 1388
rect 2072 1372 2088 1388
rect 2152 1372 2168 1388
rect 440 1352 456 1368
rect 616 1352 632 1368
rect 872 1352 888 1368
rect 1096 1352 1112 1368
rect 1368 1352 1384 1368
rect 1928 1352 1944 1368
rect 1960 1352 1976 1368
rect 2472 1352 2488 1368
rect 2504 1372 2520 1388
rect 3000 1372 3016 1388
rect 3176 1372 3192 1388
rect 2568 1352 2584 1368
rect 2712 1352 2728 1368
rect 3192 1352 3208 1368
rect 3224 1352 3240 1368
rect 3528 1352 3544 1368
rect 808 1332 824 1348
rect 968 1332 984 1348
rect 1336 1332 1352 1348
rect 1624 1332 1640 1348
rect 1736 1332 1752 1348
rect 1752 1332 1768 1348
rect 2328 1332 2344 1348
rect 2520 1332 2536 1348
rect 3096 1332 3112 1348
rect 616 1292 632 1308
rect 760 1292 776 1308
rect 888 1292 904 1308
rect 1272 1312 1288 1328
rect 1768 1312 1784 1328
rect 2360 1312 2376 1328
rect 2456 1312 2504 1328
rect 2520 1312 2536 1328
rect 3352 1312 3368 1328
rect 1144 1292 1160 1308
rect 1224 1292 1240 1308
rect 1592 1292 1624 1308
rect 2168 1292 2184 1308
rect 2392 1292 2408 1308
rect 2520 1292 2536 1308
rect 3240 1292 3256 1308
rect 3544 1292 3560 1308
rect 616 1272 632 1288
rect 2632 1272 2648 1288
rect 2984 1272 3000 1288
rect 440 1252 456 1268
rect 1224 1232 1240 1248
rect 1560 1232 1576 1248
rect 1672 1232 1688 1248
rect 3464 1232 3480 1248
rect 424 1212 440 1228
rect 712 1212 728 1228
rect 766 1202 794 1218
rect 1096 1212 1112 1228
rect 1608 1212 1624 1228
rect 2136 1212 2152 1228
rect 2648 1212 2664 1228
rect 1960 1192 1976 1208
rect 2328 1192 2344 1208
rect 2814 1202 2842 1218
rect 2856 1192 2872 1208
rect 2920 1192 2936 1208
rect 3288 1192 3304 1208
rect 344 1172 360 1188
rect 696 1172 712 1188
rect 600 1152 616 1168
rect 1432 1152 1448 1168
rect 904 1132 920 1148
rect 1272 1132 1288 1148
rect 1832 1132 1848 1148
rect 1992 1132 2008 1148
rect 2040 1132 2056 1148
rect 2184 1132 2200 1148
rect 3048 1132 3064 1148
rect 3400 1132 3416 1148
rect 2408 1112 2424 1128
rect 3240 1112 3256 1128
rect 3256 1112 3272 1128
rect 216 1092 232 1108
rect 1416 1092 1432 1108
rect 1448 1092 1464 1108
rect 1944 1092 1960 1108
rect 2280 1092 2296 1108
rect 2328 1092 2344 1108
rect 2440 1092 2456 1108
rect 2760 1092 2776 1108
rect 3096 1092 3112 1108
rect 1000 1072 1016 1088
rect 1432 1072 1448 1088
rect 1512 1072 1528 1088
rect 1704 1072 1720 1088
rect 1896 1072 1912 1088
rect 2056 1072 2072 1088
rect 2184 1072 2200 1088
rect 2664 1072 2680 1088
rect 712 1052 728 1068
rect 1240 1052 1256 1068
rect 1352 1052 1368 1068
rect 1864 1052 1896 1068
rect 2456 1052 2472 1068
rect 2584 1052 2600 1068
rect 2744 1052 2760 1068
rect 3224 1052 3240 1068
rect 3352 1052 3368 1068
rect 648 1032 664 1048
rect 1016 1012 1032 1028
rect 2616 1032 2632 1048
rect 2904 1032 2920 1048
rect 328 992 344 1008
rect 728 992 744 1008
rect 1224 992 1240 1008
rect 1672 992 1688 1008
rect 1790 1002 1818 1018
rect 1912 1012 1928 1028
rect 1960 1012 1992 1028
rect 2408 1012 2424 1028
rect 1928 992 1944 1008
rect 2568 992 2584 1008
rect 2648 992 2680 1008
rect 936 972 952 988
rect 1336 972 1352 988
rect 1608 972 1624 988
rect 1752 972 1768 988
rect 1768 972 1784 988
rect 1992 972 2008 988
rect 2040 972 2056 988
rect 2120 972 2136 988
rect 2168 972 2184 988
rect 3528 972 3544 988
rect 888 952 904 968
rect 1368 952 1384 968
rect 1944 952 1960 968
rect 2088 952 2104 968
rect 2504 952 2520 968
rect 2632 952 2664 968
rect 1352 932 1368 948
rect 2136 932 2152 948
rect 2408 932 2424 948
rect 2712 932 2728 948
rect 232 912 248 928
rect 920 912 936 928
rect 968 912 984 928
rect 1448 912 1464 928
rect 1864 912 1896 928
rect 1944 912 1960 928
rect 3320 912 3336 928
rect 312 892 328 908
rect 1032 892 1048 908
rect 1064 892 1080 908
rect 1080 892 1096 908
rect 1400 892 1416 908
rect 1640 892 1656 908
rect 1704 892 1720 908
rect 1848 892 1864 908
rect 1384 872 1400 888
rect 1496 872 1512 888
rect 2312 872 2328 888
rect 1176 852 1192 868
rect 1208 852 1224 868
rect 1320 852 1336 868
rect 1576 852 1592 868
rect 1880 852 1896 868
rect 2664 832 2680 848
rect 2712 832 2728 848
rect 3352 832 3368 848
rect 3400 832 3416 848
rect 766 802 794 818
rect 1288 812 1304 828
rect 2008 812 2024 828
rect 1624 792 1640 808
rect 2792 792 2808 808
rect 2814 802 2842 818
rect 3496 792 3512 808
rect 680 772 728 788
rect 1352 772 1368 788
rect 1368 772 1384 788
rect 1768 772 1784 788
rect 3144 772 3160 788
rect 2152 752 2168 768
rect 936 732 952 748
rect 1192 732 1208 748
rect 2344 732 2376 748
rect 2600 732 2616 748
rect 856 712 872 728
rect 2168 712 2184 728
rect 2376 712 2392 728
rect 216 692 232 708
rect 248 692 264 708
rect 1240 692 1256 708
rect 1768 692 1784 708
rect 1832 692 1848 708
rect 2056 692 2072 708
rect 2312 692 2328 708
rect 2600 692 2616 708
rect 1368 672 1384 688
rect 1512 672 1528 688
rect 1560 672 1576 688
rect 1608 672 1624 688
rect 1896 672 1912 688
rect 2504 672 2520 688
rect 968 652 984 668
rect 1240 652 1256 668
rect 1544 652 1560 668
rect 1656 652 1672 668
rect 1768 652 1784 668
rect 3384 652 3400 668
rect 920 632 936 648
rect 984 612 1000 628
rect 1192 632 1208 648
rect 1592 632 1608 648
rect 712 592 728 608
rect 904 592 920 608
rect 1528 592 1544 608
rect 1790 602 1818 618
rect 1832 612 1848 628
rect 1848 592 1864 608
rect 696 572 712 588
rect 952 572 968 588
rect 1016 572 1032 588
rect 1224 572 1240 588
rect 1384 572 1400 588
rect 936 532 952 548
rect 392 512 408 528
rect 680 512 696 528
rect 856 512 872 528
rect 1304 512 1320 528
rect 1336 512 1352 528
rect 1576 532 1592 548
rect 1816 532 1832 548
rect 488 492 504 508
rect 1144 492 1160 508
rect 1832 492 1848 508
rect 680 472 696 488
rect 712 472 728 488
rect 744 472 760 488
rect 1480 472 1496 488
rect 1896 472 1912 488
rect 1144 432 1160 448
rect 2120 432 2136 448
rect 766 402 794 418
rect 1048 412 1064 428
rect 2056 392 2072 408
rect 2814 402 2842 418
rect 616 372 632 388
rect 904 372 920 388
rect 1432 352 1448 368
rect 1448 332 1464 348
rect 1528 332 1544 348
rect 920 312 936 328
rect 1464 292 1480 308
rect 1544 292 1560 308
rect 1064 272 1080 288
rect 1384 272 1400 288
rect 1720 272 1736 288
rect 696 232 712 248
rect 728 232 744 248
rect 1640 232 1656 248
rect 1320 212 1336 228
rect 248 192 264 208
rect 1144 192 1160 208
rect 1432 192 1448 208
rect 1790 202 1818 218
rect 232 172 248 188
rect 632 172 648 188
rect 680 172 696 188
rect 984 172 1000 188
rect 1400 172 1416 188
rect 1640 172 1656 188
rect 2088 172 2104 188
rect 968 152 984 168
rect 200 112 216 128
rect 1560 112 1576 128
rect 1752 112 1768 128
rect 2360 112 2376 128
rect 3576 112 3592 128
rect 616 92 632 108
rect 936 92 952 108
rect 1352 92 1368 108
rect 1528 92 1544 108
rect 1608 92 1624 108
rect 1032 72 1048 88
rect 1768 32 1784 48
rect 766 2 794 18
rect 1240 12 1256 28
rect 1464 12 1480 28
rect 1544 12 1560 28
rect 2814 2 2842 18
<< metal4 >>
rect 794 2406 800 2414
rect 2842 2406 2848 2414
rect 301 1588 307 1892
rect 220 1503 228 1504
rect 216 1497 228 1503
rect 220 1496 228 1497
rect 301 1244 307 1572
rect 300 1236 308 1244
rect 221 708 227 1092
rect 333 1008 339 1912
rect 349 1188 355 1452
rect 365 1344 371 1452
rect 364 1336 372 1344
rect 429 1228 435 1852
rect 461 1728 467 2272
rect 557 1848 563 2032
rect 589 1428 595 2212
rect 733 1924 739 2132
rect 794 2006 800 2014
rect 732 1916 740 1924
rect 636 1896 644 1904
rect 621 1868 627 1892
rect 637 1888 643 1896
rect 621 1368 627 1552
rect 636 1496 644 1504
rect 637 1488 643 1496
rect 445 1268 451 1352
rect 604 1303 612 1304
rect 604 1297 616 1303
rect 604 1296 612 1297
rect 605 1144 611 1152
rect 604 1136 612 1144
rect 237 188 243 912
rect 300 903 308 904
rect 300 897 312 903
rect 300 896 308 897
rect 253 324 259 692
rect 396 556 404 564
rect 397 528 403 556
rect 621 388 627 1272
rect 653 1048 659 1872
rect 684 1863 692 1864
rect 684 1857 696 1863
rect 684 1856 692 1857
rect 733 1583 739 1916
rect 780 1743 788 1744
rect 780 1737 792 1743
rect 780 1736 788 1737
rect 748 1676 756 1684
rect 749 1628 755 1676
rect 794 1606 800 1614
rect 733 1577 755 1583
rect 701 788 707 1172
rect 717 1068 723 1212
rect 684 536 692 544
rect 685 528 691 536
rect 717 488 723 592
rect 252 316 260 324
rect 253 208 259 316
rect 621 108 627 372
rect 685 188 691 472
rect 733 248 739 992
rect 749 488 755 1577
rect 765 1308 771 1572
rect 829 1448 835 1492
rect 812 1396 820 1404
rect 813 1348 819 1396
rect 794 1206 800 1214
rect 794 806 800 814
rect 861 728 867 2032
rect 877 1368 883 1872
rect 893 1604 899 1812
rect 892 1596 900 1604
rect 941 1524 947 1612
rect 940 1516 948 1524
rect 892 1456 900 1464
rect 893 1428 899 1456
rect 893 968 899 1292
rect 940 1176 948 1184
rect 909 608 915 1132
rect 941 988 947 1176
rect 925 648 931 912
rect 844 523 852 524
rect 844 517 856 523
rect 844 516 852 517
rect 794 406 800 414
rect 909 388 915 592
rect 957 588 963 2092
rect 1037 1744 1043 1752
rect 1036 1736 1044 1744
rect 973 1124 979 1332
rect 1004 1216 1012 1224
rect 972 1116 980 1124
rect 973 928 979 1116
rect 1005 1088 1011 1216
rect 988 676 996 684
rect 924 543 932 544
rect 924 537 936 543
rect 924 536 932 537
rect 637 104 643 172
rect 973 168 979 652
rect 989 628 995 676
rect 1021 588 1027 1012
rect 988 236 996 244
rect 989 188 995 236
rect 636 96 644 104
rect 941 84 947 92
rect 1037 88 1043 892
rect 1053 428 1059 1932
rect 1069 908 1075 2252
rect 1084 2063 1092 2064
rect 1084 2057 1096 2063
rect 1084 2056 1092 2057
rect 1229 1944 1235 1952
rect 1228 1936 1236 1944
rect 1101 1644 1107 1872
rect 1116 1836 1124 1844
rect 1100 1636 1108 1644
rect 1117 1468 1123 1836
rect 1133 1744 1139 1832
rect 1132 1736 1140 1744
rect 1101 1228 1107 1352
rect 1149 1264 1155 1292
rect 1148 1256 1156 1264
rect 1180 876 1188 884
rect 1181 868 1187 876
rect 1197 748 1203 1832
rect 1213 868 1219 1712
rect 1245 1568 1251 1852
rect 1277 1388 1283 1732
rect 1309 1708 1315 2092
rect 1309 1564 1315 1652
rect 1308 1556 1316 1564
rect 1293 1408 1299 1532
rect 1325 1508 1331 2132
rect 1341 1884 1347 1932
rect 1340 1876 1348 1884
rect 1437 1828 1443 2272
rect 1517 2124 1523 2312
rect 1756 2236 1764 2244
rect 1757 2188 1763 2236
rect 1818 2206 1824 2214
rect 1853 2208 1859 2252
rect 1676 2176 1684 2184
rect 1581 2144 1587 2172
rect 1677 2168 1683 2176
rect 1644 2163 1652 2164
rect 1644 2157 1656 2163
rect 1644 2156 1652 2157
rect 1869 2164 1875 2232
rect 1836 2156 1844 2164
rect 1868 2156 1876 2164
rect 1580 2136 1588 2144
rect 1516 2116 1524 2124
rect 1308 1483 1316 1484
rect 1308 1477 1320 1483
rect 1308 1476 1316 1477
rect 1341 1348 1347 1692
rect 1228 1316 1236 1324
rect 1229 1308 1235 1316
rect 1229 1104 1235 1232
rect 1277 1148 1283 1312
rect 1292 1276 1300 1284
rect 1228 1096 1236 1104
rect 1197 544 1203 632
rect 1229 588 1235 992
rect 1245 708 1251 1052
rect 1293 828 1299 1276
rect 1357 1068 1363 1732
rect 1389 1684 1395 1712
rect 1388 1676 1396 1684
rect 1372 1496 1380 1504
rect 1373 1368 1379 1496
rect 1373 1324 1379 1352
rect 1372 1316 1380 1324
rect 1437 1168 1443 1552
rect 1453 1384 1459 1492
rect 1452 1376 1460 1384
rect 1421 1084 1427 1092
rect 1437 1088 1443 1152
rect 1452 1116 1460 1124
rect 1453 1108 1459 1116
rect 1517 1088 1523 2116
rect 1532 1916 1540 1924
rect 1533 1908 1539 1916
rect 1420 1076 1428 1084
rect 1324 983 1332 984
rect 1324 977 1336 983
rect 1324 976 1332 977
rect 1357 948 1363 1052
rect 1373 944 1379 952
rect 1372 936 1380 944
rect 1388 896 1396 904
rect 1389 888 1395 896
rect 1196 536 1204 544
rect 1164 503 1172 504
rect 1160 497 1172 503
rect 1164 496 1172 497
rect 1084 283 1092 284
rect 1080 277 1092 283
rect 1084 276 1092 277
rect 1149 208 1155 432
rect 940 76 948 84
rect 1245 28 1251 652
rect 1309 484 1315 512
rect 1308 476 1316 484
rect 1325 228 1331 852
rect 1357 764 1363 772
rect 1356 756 1364 764
rect 1373 688 1379 772
rect 1340 536 1348 544
rect 1341 528 1347 536
rect 1389 288 1395 572
rect 1405 188 1411 892
rect 1437 208 1443 352
rect 1453 348 1459 912
rect 1500 896 1508 904
rect 1501 888 1507 896
rect 1516 696 1524 704
rect 1517 688 1523 696
rect 1549 668 1555 1672
rect 1565 924 1571 1232
rect 1564 916 1572 924
rect 1581 868 1587 1872
rect 1597 1308 1603 1592
rect 1613 1408 1619 2092
rect 1613 1364 1619 1392
rect 1612 1356 1620 1364
rect 1629 1348 1635 2132
rect 1661 1717 1672 1723
rect 1661 1704 1667 1717
rect 1709 1724 1715 1732
rect 1708 1716 1716 1724
rect 1725 1704 1731 1752
rect 1660 1696 1668 1704
rect 1724 1696 1732 1704
rect 1661 1523 1667 1592
rect 1645 1517 1667 1523
rect 1645 1428 1651 1517
rect 1677 1504 1683 1672
rect 1676 1496 1684 1504
rect 1661 1403 1667 1492
rect 1676 1483 1684 1484
rect 1676 1477 1688 1483
rect 1676 1476 1684 1477
rect 1692 1443 1700 1444
rect 1688 1437 1700 1443
rect 1692 1436 1700 1437
rect 1724 1436 1732 1444
rect 1725 1408 1731 1436
rect 1645 1397 1667 1403
rect 1613 1228 1619 1292
rect 1628 1236 1636 1244
rect 1612 1036 1620 1044
rect 1613 988 1619 1036
rect 1596 836 1604 844
rect 1533 348 1539 592
rect 1357 84 1363 92
rect 1356 76 1364 84
rect 1469 28 1475 292
rect 1549 28 1555 292
rect 1565 128 1571 672
rect 1597 648 1603 836
rect 1629 808 1635 1236
rect 1645 908 1651 1397
rect 1741 1348 1747 1972
rect 1820 1916 1828 1924
rect 1821 1908 1827 1916
rect 1818 1806 1824 1814
rect 1756 1396 1764 1404
rect 1757 1348 1763 1396
rect 1773 1328 1779 1532
rect 1837 1508 1843 2156
rect 1869 2104 1875 2112
rect 1868 2096 1876 2104
rect 1853 1924 1859 1932
rect 1852 1916 1860 1924
rect 1853 1764 1859 1772
rect 1852 1756 1860 1764
rect 1853 1468 1859 1492
rect 1852 1436 1860 1444
rect 1853 1428 1859 1436
rect 1818 1406 1824 1414
rect 1660 1316 1668 1324
rect 1596 543 1604 544
rect 1592 537 1604 543
rect 1596 536 1604 537
rect 1613 108 1619 672
rect 1645 248 1651 892
rect 1661 668 1667 1316
rect 1852 1236 1860 1244
rect 1677 1008 1683 1232
rect 1836 1096 1844 1104
rect 1724 1083 1732 1084
rect 1720 1077 1732 1083
rect 1724 1076 1732 1077
rect 1772 1076 1780 1084
rect 1756 1056 1764 1064
rect 1757 988 1763 1056
rect 1773 988 1779 1076
rect 1818 1006 1824 1014
rect 1772 796 1780 804
rect 1773 788 1779 796
rect 1837 708 1843 1096
rect 1853 908 1859 1236
rect 1869 1068 1875 1452
rect 1885 1068 1891 2192
rect 1901 1748 1907 2272
rect 1932 2236 1940 2244
rect 1933 2108 1939 2236
rect 1964 2136 1972 2144
rect 1965 2128 1971 2136
rect 1901 1488 1907 1732
rect 1949 1728 1955 1752
rect 1965 1728 1971 1992
rect 1965 1688 1971 1712
rect 1981 1668 1987 2132
rect 2077 2124 2083 2272
rect 2220 2256 2228 2264
rect 2076 2123 2084 2124
rect 2072 2117 2084 2123
rect 2076 2116 2084 2117
rect 2221 2108 2227 2256
rect 2252 2176 2260 2184
rect 2253 2148 2259 2176
rect 2253 2124 2259 2132
rect 2252 2116 2260 2124
rect 1997 1668 2003 1832
rect 2012 1783 2020 1784
rect 2012 1777 2024 1783
rect 2012 1776 2020 1777
rect 2013 1704 2019 1712
rect 2012 1696 2020 1704
rect 2045 1684 2051 1712
rect 2044 1676 2052 1684
rect 1964 1636 1972 1644
rect 1901 1088 1907 1472
rect 1916 1416 1924 1424
rect 1917 1408 1923 1416
rect 1917 1364 1923 1392
rect 1933 1384 1939 1492
rect 1965 1428 1971 1636
rect 1932 1376 1940 1384
rect 1933 1368 1939 1376
rect 1916 1356 1924 1364
rect 1949 1108 1955 1392
rect 1965 1208 1971 1352
rect 1964 1136 1972 1144
rect 1868 956 1876 964
rect 1869 928 1875 956
rect 1885 928 1891 1052
rect 1885 868 1891 912
rect 1773 668 1779 692
rect 1901 688 1907 1072
rect 1917 1004 1923 1012
rect 1916 996 1924 1004
rect 1628 183 1636 184
rect 1628 177 1640 183
rect 1628 176 1636 177
rect 1756 176 1764 184
rect 1757 128 1763 176
rect 1773 48 1779 652
rect 1818 606 1824 614
rect 1821 524 1827 532
rect 1820 516 1828 524
rect 1837 508 1843 612
rect 1853 544 1859 592
rect 1900 576 1908 584
rect 1852 536 1860 544
rect 1901 488 1907 576
rect 1933 564 1939 992
rect 1949 968 1955 1092
rect 1965 1028 1971 1136
rect 1997 1104 2003 1132
rect 1996 1096 2004 1104
rect 1980 1056 1988 1064
rect 1981 1028 1987 1056
rect 1996 1016 2004 1024
rect 1997 988 2003 1016
rect 2013 828 2019 1472
rect 2077 1468 2083 1752
rect 2093 1628 2099 1772
rect 2109 1724 2115 1752
rect 2108 1716 2116 1724
rect 2061 1344 2067 1392
rect 2077 1388 2083 1452
rect 2060 1336 2068 1344
rect 2125 1184 2131 1872
rect 2141 1428 2147 1892
rect 2189 1864 2195 1892
rect 2188 1856 2196 1864
rect 2205 1844 2211 1912
rect 2204 1836 2212 1844
rect 2221 1484 2227 1952
rect 2236 1936 2244 1944
rect 2252 1936 2260 1944
rect 2237 1908 2243 1936
rect 2253 1908 2259 1936
rect 2237 1844 2243 1872
rect 2236 1836 2244 1844
rect 2269 1808 2275 2112
rect 2333 2104 2339 2112
rect 2332 2096 2340 2104
rect 2284 1916 2292 1924
rect 2285 1888 2291 1916
rect 2316 1923 2324 1924
rect 2312 1917 2324 1923
rect 2316 1916 2324 1917
rect 2269 1688 2275 1792
rect 2333 1768 2339 2032
rect 2349 1884 2355 1892
rect 2348 1876 2356 1884
rect 2365 1548 2371 1992
rect 2381 1604 2387 1632
rect 2380 1596 2388 1604
rect 2220 1476 2228 1484
rect 2221 1468 2227 1476
rect 2300 1463 2308 1464
rect 2300 1457 2312 1463
rect 2300 1456 2308 1457
rect 2221 1404 2227 1452
rect 2220 1396 2228 1404
rect 2124 1176 2132 1184
rect 2045 988 2051 1132
rect 2141 1124 2147 1212
rect 2140 1116 2148 1124
rect 2061 1004 2067 1072
rect 2060 996 2068 1004
rect 2093 904 2099 952
rect 2092 896 2100 904
rect 1932 556 1940 564
rect 2061 408 2067 692
rect 1818 206 1824 214
rect 2093 188 2099 896
rect 2125 448 2131 972
rect 2140 956 2148 964
rect 2141 948 2147 956
rect 2157 804 2163 1372
rect 2333 1348 2339 1452
rect 2173 1264 2179 1292
rect 2172 1256 2180 1264
rect 2172 1143 2180 1144
rect 2172 1137 2184 1143
rect 2172 1136 2180 1137
rect 2333 1108 2339 1192
rect 2300 1103 2308 1104
rect 2296 1097 2308 1103
rect 2300 1096 2308 1097
rect 2172 1083 2180 1084
rect 2172 1077 2184 1083
rect 2172 1076 2180 1077
rect 2156 796 2164 804
rect 2157 744 2163 752
rect 2156 736 2164 744
rect 2173 728 2179 972
rect 2317 708 2323 872
rect 2349 748 2355 1432
rect 2365 1328 2371 1532
rect 2364 756 2372 764
rect 2365 748 2371 756
rect 2381 728 2387 1596
rect 2412 1396 2420 1404
rect 2396 1316 2404 1324
rect 2397 1308 2403 1316
rect 2413 1128 2419 1396
rect 2429 1224 2435 1412
rect 2428 1216 2436 1224
rect 2445 1108 2451 1512
rect 2477 1368 2483 1792
rect 2509 1748 2515 2052
rect 2573 1968 2579 2232
rect 2556 1856 2564 1864
rect 2460 1356 2468 1364
rect 2461 1328 2467 1356
rect 2477 1284 2483 1312
rect 2476 1276 2484 1284
rect 2493 1124 2499 1312
rect 2492 1116 2500 1124
rect 2509 1064 2515 1372
rect 2525 1348 2531 1832
rect 2541 1448 2547 1852
rect 2557 1848 2563 1856
rect 2556 1796 2564 1804
rect 2557 1748 2563 1796
rect 2573 1468 2579 1952
rect 2605 1528 2611 1852
rect 2621 1528 2627 2212
rect 2701 1868 2707 2012
rect 2732 1903 2740 1904
rect 2728 1897 2740 1903
rect 2732 1896 2740 1897
rect 2508 1056 2516 1064
rect 2413 948 2419 1012
rect 2461 884 2467 1052
rect 2509 968 2515 1056
rect 2573 1008 2579 1352
rect 2589 984 2595 1052
rect 2621 1048 2627 1432
rect 2637 1288 2643 1492
rect 2765 1424 2771 2152
rect 2781 2124 2787 2132
rect 2797 2128 2803 2152
rect 2780 2116 2788 2124
rect 3100 2056 3108 2064
rect 2842 2006 2848 2014
rect 2877 1784 2883 1852
rect 2876 1776 2884 1784
rect 2829 1648 2835 1692
rect 2842 1606 2848 1614
rect 2764 1416 2772 1424
rect 2621 1024 2627 1032
rect 2620 1016 2628 1024
rect 2588 976 2596 984
rect 2637 968 2643 1272
rect 2653 1008 2659 1212
rect 2653 944 2659 952
rect 2652 936 2660 944
rect 2460 876 2468 884
rect 2669 848 2675 992
rect 2717 948 2723 1352
rect 2748 1116 2756 1124
rect 2749 1068 2755 1116
rect 2765 1108 2771 1416
rect 2842 1206 2848 1214
rect 2861 1044 2867 1192
rect 2909 1048 2915 1912
rect 2956 1723 2964 1724
rect 2952 1717 2964 1723
rect 2956 1716 2964 1717
rect 2925 1208 2931 1692
rect 3005 1388 3011 1532
rect 3021 1504 3027 2032
rect 3020 1496 3028 1504
rect 3021 1488 3027 1496
rect 3053 1148 3059 1872
rect 3101 1828 3107 2056
rect 3212 1936 3220 1944
rect 3213 1928 3219 1936
rect 3213 1844 3219 1892
rect 3212 1836 3220 1844
rect 3148 1643 3156 1644
rect 3144 1637 3156 1643
rect 3148 1636 3156 1637
rect 3116 1343 3124 1344
rect 3112 1337 3124 1343
rect 3116 1336 3124 1337
rect 3101 1108 3107 1332
rect 2860 1036 2868 1044
rect 2796 836 2804 844
rect 2797 808 2803 836
rect 2842 806 2848 814
rect 3149 788 3155 1612
rect 3180 1516 3188 1524
rect 3181 1388 3187 1516
rect 3197 1368 3203 1772
rect 3229 1068 3235 1352
rect 3245 1308 3251 1932
rect 3245 1128 3251 1292
rect 3261 1128 3267 1572
rect 3277 844 3283 2272
rect 3309 1708 3315 2052
rect 3372 1883 3380 1884
rect 3368 1877 3380 1883
rect 3372 1876 3380 1877
rect 3293 1488 3299 1552
rect 3309 1548 3315 1692
rect 3293 1208 3299 1472
rect 3325 928 3331 1592
rect 3356 1356 3364 1364
rect 3357 1328 3363 1356
rect 3357 848 3363 1052
rect 3276 836 3284 844
rect 2605 708 2611 732
rect 2508 696 2516 704
rect 2509 688 2515 696
rect 2605 684 2611 692
rect 2604 676 2612 684
rect 3389 668 3395 2032
rect 3405 1148 3411 1392
rect 3469 1248 3475 1872
rect 3420 843 3428 844
rect 3416 837 3428 843
rect 3420 836 3428 837
rect 3501 808 3507 1892
rect 3533 988 3539 1352
rect 3549 1308 3555 1732
rect 2842 406 2848 414
rect 3581 128 3587 1532
rect 2380 123 2388 124
rect 2376 117 2388 123
rect 2380 116 2388 117
rect 794 6 800 14
rect 2842 6 2848 14
use BUFX2  BUFX2_36
timestamp 1513729314
transform -1 0 56 0 1 2210
box 0 0 48 200
use BUFX2  BUFX2_17
timestamp 1513729314
transform -1 0 104 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_18
timestamp 1513729314
transform 1 0 104 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_35
timestamp 1513729314
transform -1 0 232 0 1 2210
box 0 0 64 200
use BUFX2  BUFX2_10
timestamp 1513729314
transform 1 0 232 0 1 2210
box 0 0 48 200
use BUFX2  BUFX2_29
timestamp 1513729314
transform 1 0 280 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_9
timestamp 1513729314
transform 1 0 328 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_88
timestamp 1513729314
transform 1 0 392 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_4
timestamp 1513729314
transform 1 0 456 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_96
timestamp 1513729314
transform 1 0 520 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_45
timestamp 1513729314
transform 1 0 584 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_48
timestamp 1513729314
transform -1 0 712 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_10
timestamp 1513729314
transform -1 0 776 0 1 2210
box 0 0 64 200
use FILL  FILL_11_0_0
timestamp 1513729314
transform 1 0 776 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1513729314
transform 1 0 792 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_75
timestamp 1513729314
transform 1 0 808 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_79
timestamp 1513729314
transform -1 0 936 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_15
timestamp 1513729314
transform -1 0 1000 0 1 2210
box 0 0 64 200
use INVX2  INVX2_10
timestamp 1513729314
transform -1 0 1032 0 1 2210
box 0 0 32 200
use AND2X2  AND2X2_14
timestamp 1513729314
transform 1 0 1032 0 1 2210
box 0 0 64 200
use AND2X2  AND2X2_13
timestamp 1513729314
transform -1 0 1160 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_66
timestamp 1513729314
transform -1 0 1224 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_55
timestamp 1513729314
transform -1 0 1272 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_61
timestamp 1513729314
transform -1 0 1320 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_103
timestamp 1513729314
transform -1 0 1384 0 1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_31
timestamp 1513729314
transform -1 0 1432 0 1 2210
box 0 0 48 200
use MUX2X1  MUX2X1_22
timestamp 1513729314
transform -1 0 1528 0 1 2210
box 0 0 96 200
use NAND2X1  NAND2X1_52
timestamp 1513729314
transform -1 0 1576 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_11
timestamp 1513729314
transform 1 0 1576 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_7
timestamp 1513729314
transform -1 0 1672 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_130
timestamp 1513729314
transform -1 0 1736 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_128
timestamp 1513729314
transform 1 0 1736 0 1 2210
box 0 0 64 200
use FILL  FILL_11_1_0
timestamp 1513729314
transform -1 0 1816 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1513729314
transform -1 0 1832 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_4
timestamp 1513729314
transform -1 0 1880 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_126
timestamp 1513729314
transform -1 0 1944 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_113
timestamp 1513729314
transform -1 0 2008 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_36
timestamp 1513729314
transform 1 0 2008 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_127
timestamp 1513729314
transform 1 0 2072 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_132
timestamp 1513729314
transform 1 0 2136 0 1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_4
timestamp 1513729314
transform 1 0 2200 0 1 2210
box 0 0 96 200
use BUFX4  BUFX4_121
timestamp 1513729314
transform -1 0 2360 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_123
timestamp 1513729314
transform 1 0 2360 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_46
timestamp 1513729314
transform -1 0 2472 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_120
timestamp 1513729314
transform 1 0 2472 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_125
timestamp 1513729314
transform 1 0 2536 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_119
timestamp 1513729314
transform 1 0 2600 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_34
timestamp 1513729314
transform 1 0 2664 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_37
timestamp 1513729314
transform 1 0 2728 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_31
timestamp 1513729314
transform 1 0 2792 0 1 2210
box 0 0 64 200
use FILL  FILL_11_2_0
timestamp 1513729314
transform 1 0 2856 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1513729314
transform 1 0 2872 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_9
timestamp 1513729314
transform 1 0 2888 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_137
timestamp 1513729314
transform -1 0 3000 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_114
timestamp 1513729314
transform 1 0 3000 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_116
timestamp 1513729314
transform -1 0 3128 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_112
timestamp 1513729314
transform 1 0 3128 0 1 2210
box 0 0 64 200
use BUFX2  BUFX2_2
timestamp 1513729314
transform 1 0 3192 0 1 2210
box 0 0 48 200
use BUFX2  BUFX2_21
timestamp 1513729314
transform 1 0 3240 0 1 2210
box 0 0 48 200
use BUFX2  BUFX2_5
timestamp 1513729314
transform 1 0 3288 0 1 2210
box 0 0 48 200
use BUFX2  BUFX2_24
timestamp 1513729314
transform 1 0 3336 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_91
timestamp 1513729314
transform -1 0 3448 0 1 2210
box 0 0 64 200
use BUFX2  BUFX2_27
timestamp 1513729314
transform 1 0 3448 0 1 2210
box 0 0 48 200
use BUFX4  BUFX4_69
timestamp 1513729314
transform -1 0 3560 0 1 2210
box 0 0 64 200
use BUFX4  BUFX4_7
timestamp 1513729314
transform 1 0 3560 0 1 2210
box 0 0 64 200
use FILL  FILL_12_1
timestamp 1513729314
transform 1 0 3624 0 1 2210
box 0 0 16 200
use FILL  FILL_12_2
timestamp 1513729314
transform 1 0 3640 0 1 2210
box 0 0 16 200
use BUFX2  BUFX2_33
timestamp 1513729314
transform -1 0 56 0 -1 2210
box 0 0 48 200
use BUFX2  BUFX2_14
timestamp 1513729314
transform -1 0 104 0 -1 2210
box 0 0 48 200
use BUFX4  BUFX4_83
timestamp 1513729314
transform 1 0 104 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_51
timestamp 1513729314
transform 1 0 168 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_65
timestamp 1513729314
transform -1 0 296 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_117
timestamp 1513729314
transform 1 0 296 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_44
timestamp 1513729314
transform -1 0 424 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_98
timestamp 1513729314
transform 1 0 424 0 -1 2210
box 0 0 64 200
use INVX8  INVX8_1
timestamp 1513729314
transform -1 0 568 0 -1 2210
box 0 0 80 200
use XNOR2X1  XNOR2X1_4
timestamp 1513729314
transform 1 0 568 0 -1 2210
box 0 0 112 200
use NOR2X1  NOR2X1_37
timestamp 1513729314
transform -1 0 728 0 -1 2210
box 0 0 48 200
use NOR2X1  NOR2X1_45
timestamp 1513729314
transform 1 0 728 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_0_0
timestamp 1513729314
transform 1 0 776 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1513729314
transform 1 0 792 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_135
timestamp 1513729314
transform 1 0 808 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_29
timestamp 1513729314
transform 1 0 872 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_16
timestamp 1513729314
transform -1 0 1000 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_12
timestamp 1513729314
transform 1 0 1000 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_70
timestamp 1513729314
transform 1 0 1048 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_65
timestamp 1513729314
transform 1 0 1112 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_27
timestamp 1513729314
transform -1 0 1272 0 -1 2210
box 0 0 96 200
use NAND2X1  NAND2X1_99
timestamp 1513729314
transform 1 0 1272 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_61
timestamp 1513729314
transform 1 0 1320 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_3
timestamp 1513729314
transform -1 0 1480 0 -1 2210
box 0 0 96 200
use OAI21X1  OAI21X1_44
timestamp 1513729314
transform -1 0 1544 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_32
timestamp 1513729314
transform 1 0 1544 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_57
timestamp 1513729314
transform -1 0 1640 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_138
timestamp 1513729314
transform 1 0 1640 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_35
timestamp 1513729314
transform -1 0 1768 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_27
timestamp 1513729314
transform 1 0 1768 0 -1 2210
box 0 0 32 200
use FILL  FILL_10_1_0
timestamp 1513729314
transform 1 0 1800 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1513729314
transform 1 0 1816 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_139
timestamp 1513729314
transform 1 0 1832 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_4
timestamp 1513729314
transform -1 0 1928 0 -1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_136
timestamp 1513729314
transform -1 0 1992 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_74
timestamp 1513729314
transform 1 0 1992 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_123
timestamp 1513729314
transform -1 0 2104 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_5
timestamp 1513729314
transform 1 0 2104 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_113
timestamp 1513729314
transform 1 0 2168 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_19
timestamp 1513729314
transform 1 0 2232 0 -1 2210
box 0 0 96 200
use INVX8  INVX8_5
timestamp 1513729314
transform -1 0 2408 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_32
timestamp 1513729314
transform -1 0 2472 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_38
timestamp 1513729314
transform -1 0 2536 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_16
timestamp 1513729314
transform 1 0 2536 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_14
timestamp 1513729314
transform -1 0 2664 0 -1 2210
box 0 0 64 200
use AOI21X1  AOI21X1_31
timestamp 1513729314
transform 1 0 2664 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_33
timestamp 1513729314
transform -1 0 2792 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_36
timestamp 1513729314
transform -1 0 2824 0 -1 2210
box 0 0 32 200
use FILL  FILL_10_2_0
timestamp 1513729314
transform -1 0 2840 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1513729314
transform -1 0 2856 0 -1 2210
box 0 0 16 200
use INVX1  INVX1_34
timestamp 1513729314
transform -1 0 2888 0 -1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_45
timestamp 1513729314
transform 1 0 2888 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_140
timestamp 1513729314
transform -1 0 3000 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_19
timestamp 1513729314
transform -1 0 3032 0 -1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_14
timestamp 1513729314
transform 1 0 3032 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_141
timestamp 1513729314
transform -1 0 3144 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_111
timestamp 1513729314
transform -1 0 3208 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_109
timestamp 1513729314
transform 1 0 3208 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_14
timestamp 1513729314
transform 1 0 3272 0 -1 2210
box 0 0 96 200
use BUFX4  BUFX4_27
timestamp 1513729314
transform 1 0 3368 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_61
timestamp 1513729314
transform 1 0 3432 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_33
timestamp 1513729314
transform 1 0 3496 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_118
timestamp 1513729314
transform 1 0 3560 0 -1 2210
box 0 0 64 200
use FILL  FILL_11_1
timestamp 1513729314
transform -1 0 3640 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_2
timestamp 1513729314
transform -1 0 3656 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_97
timestamp 1513729314
transform -1 0 72 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_48
timestamp 1513729314
transform 1 0 72 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_59
timestamp 1513729314
transform -1 0 200 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_71
timestamp 1513729314
transform -1 0 264 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_53
timestamp 1513729314
transform -1 0 328 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_11
timestamp 1513729314
transform 1 0 328 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_40
timestamp 1513729314
transform -1 0 440 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_59
timestamp 1513729314
transform 1 0 440 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_32
timestamp 1513729314
transform 1 0 504 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_5
timestamp 1513729314
transform -1 0 648 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_49
timestamp 1513729314
transform 1 0 648 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_25
timestamp 1513729314
transform -1 0 760 0 1 1810
box 0 0 64 200
use FILL  FILL_9_0_0
timestamp 1513729314
transform -1 0 776 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1513729314
transform -1 0 792 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_39
timestamp 1513729314
transform -1 0 856 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_93
timestamp 1513729314
transform 1 0 856 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_11
timestamp 1513729314
transform -1 0 968 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_118
timestamp 1513729314
transform -1 0 1032 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_77
timestamp 1513729314
transform 1 0 1032 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_69
timestamp 1513729314
transform 1 0 1080 0 1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_3
timestamp 1513729314
transform -1 0 1272 0 1 1810
box 0 0 128 200
use AOI21X1  AOI21X1_27
timestamp 1513729314
transform 1 0 1272 0 1 1810
box 0 0 64 200
use INVX1  INVX1_39
timestamp 1513729314
transform -1 0 1368 0 1 1810
box 0 0 32 200
use OAI22X1  OAI22X1_4
timestamp 1513729314
transform 1 0 1368 0 1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_22
timestamp 1513729314
transform -1 0 1512 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_17
timestamp 1513729314
transform -1 0 1576 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_26
timestamp 1513729314
transform -1 0 1624 0 1 1810
box 0 0 48 200
use XNOR2X1  XNOR2X1_3
timestamp 1513729314
transform 1 0 1624 0 1 1810
box 0 0 112 200
use NAND2X1  NAND2X1_89
timestamp 1513729314
transform -1 0 1784 0 1 1810
box 0 0 48 200
use INVX1  INVX1_37
timestamp 1513729314
transform -1 0 1816 0 1 1810
box 0 0 32 200
use FILL  FILL_9_1_0
timestamp 1513729314
transform -1 0 1832 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1513729314
transform -1 0 1848 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_29
timestamp 1513729314
transform -1 0 1896 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_18
timestamp 1513729314
transform -1 0 1960 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_10
timestamp 1513729314
transform 1 0 1960 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_95
timestamp 1513729314
transform -1 0 2072 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_46
timestamp 1513729314
transform -1 0 2120 0 1 1810
box 0 0 48 200
use MUX2X1  MUX2X1_24
timestamp 1513729314
transform 1 0 2120 0 1 1810
box 0 0 96 200
use OAI21X1  OAI21X1_74
timestamp 1513729314
transform -1 0 2280 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_27
timestamp 1513729314
transform 1 0 2280 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_3
timestamp 1513729314
transform 1 0 2344 0 1 1810
box 0 0 80 200
use AOI21X1  AOI21X1_28
timestamp 1513729314
transform -1 0 2488 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_3
timestamp 1513729314
transform -1 0 2552 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_26
timestamp 1513729314
transform -1 0 2616 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_41
timestamp 1513729314
transform 1 0 2616 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_66
timestamp 1513729314
transform -1 0 2712 0 1 1810
box 0 0 48 200
use NOR2X1  NOR2X1_33
timestamp 1513729314
transform 1 0 2712 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_43
timestamp 1513729314
transform -1 0 2824 0 1 1810
box 0 0 64 200
use FILL  FILL_9_2_0
timestamp 1513729314
transform 1 0 2824 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1513729314
transform 1 0 2840 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_94
timestamp 1513729314
transform 1 0 2856 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_51
timestamp 1513729314
transform 1 0 2904 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_42
timestamp 1513729314
transform -1 0 3016 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_47
timestamp 1513729314
transform 1 0 3016 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_115
timestamp 1513729314
transform -1 0 3128 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_23
timestamp 1513729314
transform 1 0 3128 0 1 1810
box 0 0 96 200
use OAI21X1  OAI21X1_72
timestamp 1513729314
transform 1 0 3224 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_52
timestamp 1513729314
transform -1 0 3352 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_21
timestamp 1513729314
transform 1 0 3352 0 1 1810
box 0 0 48 200
use MUX2X1  MUX2X1_17
timestamp 1513729314
transform -1 0 3496 0 1 1810
box 0 0 96 200
use BUFX2  BUFX2_8
timestamp 1513729314
transform -1 0 3544 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_30
timestamp 1513729314
transform 1 0 3544 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_28
timestamp 1513729314
transform -1 0 3656 0 1 1810
box 0 0 64 200
use BUFX2  BUFX2_23
timestamp 1513729314
transform -1 0 56 0 -1 1810
box 0 0 48 200
use BUFX2  BUFX2_4
timestamp 1513729314
transform -1 0 104 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_14
timestamp 1513729314
transform 1 0 104 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_80
timestamp 1513729314
transform 1 0 168 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_53
timestamp 1513729314
transform -1 0 296 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_54
timestamp 1513729314
transform -1 0 360 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_9
timestamp 1513729314
transform 1 0 360 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_58
timestamp 1513729314
transform -1 0 488 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1513729314
transform 1 0 488 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_37
timestamp 1513729314
transform -1 0 616 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_36
timestamp 1513729314
transform 1 0 616 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_40
timestamp 1513729314
transform 1 0 680 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_78
timestamp 1513729314
transform -1 0 792 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_0_0
timestamp 1513729314
transform 1 0 792 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1513729314
transform 1 0 808 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_65
timestamp 1513729314
transform 1 0 824 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_53
timestamp 1513729314
transform 1 0 872 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_106
timestamp 1513729314
transform 1 0 920 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_35
timestamp 1513729314
transform 1 0 984 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_97
timestamp 1513729314
transform -1 0 1080 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_102
timestamp 1513729314
transform 1 0 1080 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_105
timestamp 1513729314
transform 1 0 1144 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_92
timestamp 1513729314
transform -1 0 1272 0 -1 1810
box 0 0 64 200
use OAI22X1  OAI22X1_6
timestamp 1513729314
transform 1 0 1272 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_2
timestamp 1513729314
transform -1 0 1416 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_103
timestamp 1513729314
transform 1 0 1416 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_76
timestamp 1513729314
transform 1 0 1480 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_69
timestamp 1513729314
transform -1 0 1576 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_20
timestamp 1513729314
transform -1 0 1640 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_82
timestamp 1513729314
transform -1 0 1704 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_5
timestamp 1513729314
transform 1 0 1704 0 -1 1810
box 0 0 96 200
use FILL  FILL_8_1_0
timestamp 1513729314
transform -1 0 1816 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1513729314
transform -1 0 1832 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_22
timestamp 1513729314
transform -1 0 1880 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_68
timestamp 1513729314
transform -1 0 1944 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_125
timestamp 1513729314
transform 1 0 1944 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_124
timestamp 1513729314
transform -1 0 2072 0 -1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_44
timestamp 1513729314
transform -1 0 2136 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_34
timestamp 1513729314
transform -1 0 2184 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_24
timestamp 1513729314
transform 1 0 2184 0 -1 1810
box 0 0 48 200
use AND2X2  AND2X2_3
timestamp 1513729314
transform 1 0 2232 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_96
timestamp 1513729314
transform -1 0 2344 0 -1 1810
box 0 0 48 200
use BUFX4  BUFX4_86
timestamp 1513729314
transform 1 0 2344 0 -1 1810
box 0 0 64 200
use XNOR2X1  XNOR2X1_2
timestamp 1513729314
transform -1 0 2520 0 -1 1810
box 0 0 112 200
use INVX4  INVX4_4
timestamp 1513729314
transform -1 0 2568 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_67
timestamp 1513729314
transform 1 0 2568 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_68
timestamp 1513729314
transform -1 0 2664 0 -1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_4
timestamp 1513729314
transform -1 0 2728 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_3
timestamp 1513729314
transform 1 0 2728 0 -1 1810
box 0 0 32 200
use AOI21X1  AOI21X1_39
timestamp 1513729314
transform -1 0 2824 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_2_0
timestamp 1513729314
transform 1 0 2824 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1513729314
transform 1 0 2840 0 -1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_13
timestamp 1513729314
transform 1 0 2856 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_11
timestamp 1513729314
transform -1 0 3048 0 -1 1810
box 0 0 96 200
use NOR2X1  NOR2X1_34
timestamp 1513729314
transform 1 0 3048 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_39
timestamp 1513729314
transform 1 0 3096 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_26
timestamp 1513729314
transform 1 0 3144 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_41
timestamp 1513729314
transform -1 0 3240 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_42
timestamp 1513729314
transform 1 0 3240 0 -1 1810
box 0 0 32 200
use NAND2X1  NAND2X1_15
timestamp 1513729314
transform 1 0 3272 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_29
timestamp 1513729314
transform 1 0 3320 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_80
timestamp 1513729314
transform -1 0 3432 0 -1 1810
box 0 0 48 200
use MUX2X1  MUX2X1_20
timestamp 1513729314
transform -1 0 3528 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_1
timestamp 1513729314
transform 1 0 3528 0 -1 1810
box 0 0 96 200
use FILL  FILL_9_1
timestamp 1513729314
transform -1 0 3640 0 -1 1810
box 0 0 16 200
use FILL  FILL_9_2
timestamp 1513729314
transform -1 0 3656 0 -1 1810
box 0 0 16 200
use INVX8  INVX8_11
timestamp 1513729314
transform -1 0 88 0 1 1410
box 0 0 80 200
use AND2X2  AND2X2_8
timestamp 1513729314
transform -1 0 152 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_38
timestamp 1513729314
transform 1 0 152 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_46
timestamp 1513729314
transform 1 0 200 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_34
timestamp 1513729314
transform -1 0 328 0 1 1410
box 0 0 64 200
use INVX2  INVX2_4
timestamp 1513729314
transform -1 0 360 0 1 1410
box 0 0 32 200
use INVX1  INVX1_2
timestamp 1513729314
transform 1 0 360 0 1 1410
box 0 0 32 200
use OR2X2  OR2X2_4
timestamp 1513729314
transform -1 0 456 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_63
timestamp 1513729314
transform 1 0 456 0 1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_23
timestamp 1513729314
transform -1 0 568 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_11
timestamp 1513729314
transform -1 0 632 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1513729314
transform -1 0 696 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_2
timestamp 1513729314
transform -1 0 760 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_20
timestamp 1513729314
transform 1 0 760 0 1 1410
box 0 0 48 200
use FILL  FILL_7_0_0
timestamp 1513729314
transform -1 0 824 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1513729314
transform -1 0 840 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_2
timestamp 1513729314
transform -1 0 888 0 1 1410
box 0 0 48 200
use INVX2  INVX2_2
timestamp 1513729314
transform 1 0 888 0 1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_84
timestamp 1513729314
transform 1 0 920 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_8
timestamp 1513729314
transform 1 0 968 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_41
timestamp 1513729314
transform 1 0 1016 0 1 1410
box 0 0 48 200
use NOR3X1  NOR3X1_2
timestamp 1513729314
transform -1 0 1192 0 1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_133
timestamp 1513729314
transform -1 0 1256 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_62
timestamp 1513729314
transform 1 0 1256 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_104
timestamp 1513729314
transform -1 0 1368 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_2
timestamp 1513729314
transform -1 0 1464 0 1 1410
box 0 0 96 200
use AOI21X1  AOI21X1_2
timestamp 1513729314
transform -1 0 1528 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_41
timestamp 1513729314
transform -1 0 1592 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_48
timestamp 1513729314
transform 1 0 1592 0 1 1410
box 0 0 48 200
use INVX1  INVX1_9
timestamp 1513729314
transform 1 0 1640 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_91
timestamp 1513729314
transform 1 0 1672 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_76
timestamp 1513729314
transform 1 0 1736 0 1 1410
box 0 0 64 200
use FILL  FILL_7_1_0
timestamp 1513729314
transform 1 0 1800 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1513729314
transform 1 0 1816 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_47
timestamp 1513729314
transform 1 0 1832 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_49
timestamp 1513729314
transform -1 0 1960 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_108
timestamp 1513729314
transform 1 0 1960 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_85
timestamp 1513729314
transform 1 0 2024 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_44
timestamp 1513729314
transform -1 0 2136 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_10
timestamp 1513729314
transform 1 0 2136 0 1 1410
box 0 0 64 200
use OR2X2  OR2X2_7
timestamp 1513729314
transform 1 0 2200 0 1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_8
timestamp 1513729314
transform 1 0 2264 0 1 1410
box 0 0 80 200
use NOR2X1  NOR2X1_43
timestamp 1513729314
transform -1 0 2392 0 1 1410
box 0 0 48 200
use AND2X2  AND2X2_4
timestamp 1513729314
transform -1 0 2456 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_25
timestamp 1513729314
transform 1 0 2456 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_12
timestamp 1513729314
transform -1 0 2568 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1513729314
transform -1 0 2632 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_20
timestamp 1513729314
transform -1 0 2680 0 1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_6
timestamp 1513729314
transform 1 0 2680 0 1 1410
box 0 0 80 200
use AOI21X1  AOI21X1_29
timestamp 1513729314
transform 1 0 2760 0 1 1410
box 0 0 64 200
use FILL  FILL_7_2_0
timestamp 1513729314
transform 1 0 2824 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1513729314
transform 1 0 2840 0 1 1410
box 0 0 16 200
use NOR2X1  NOR2X1_22
timestamp 1513729314
transform 1 0 2856 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_24
timestamp 1513729314
transform -1 0 2968 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_37
timestamp 1513729314
transform 1 0 2968 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_62
timestamp 1513729314
transform -1 0 3096 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_40
timestamp 1513729314
transform -1 0 3160 0 1 1410
box 0 0 64 200
use XNOR2X1  XNOR2X1_1
timestamp 1513729314
transform -1 0 3272 0 1 1410
box 0 0 112 200
use OAI21X1  OAI21X1_126
timestamp 1513729314
transform 1 0 3272 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_32
timestamp 1513729314
transform 1 0 3336 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_63
timestamp 1513729314
transform -1 0 3448 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_50
timestamp 1513729314
transform -1 0 3512 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_33
timestamp 1513729314
transform 1 0 3512 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_49
timestamp 1513729314
transform -1 0 3640 0 1 1410
box 0 0 64 200
use FILL  FILL_8_1
timestamp 1513729314
transform 1 0 3640 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_67
timestamp 1513729314
transform -1 0 72 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_77
timestamp 1513729314
transform -1 0 136 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_24
timestamp 1513729314
transform -1 0 184 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_27
timestamp 1513729314
transform 1 0 184 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_26
timestamp 1513729314
transform -1 0 280 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_46
timestamp 1513729314
transform 1 0 280 0 -1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_16
timestamp 1513729314
transform -1 0 360 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_100
timestamp 1513729314
transform 1 0 360 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_111
timestamp 1513729314
transform -1 0 488 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_24
timestamp 1513729314
transform -1 0 552 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_35
timestamp 1513729314
transform -1 0 616 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_36
timestamp 1513729314
transform -1 0 664 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_30
timestamp 1513729314
transform -1 0 728 0 -1 1410
box 0 0 64 200
use INVX2  INVX2_1
timestamp 1513729314
transform 1 0 728 0 -1 1410
box 0 0 32 200
use FILL  FILL_6_0_0
timestamp 1513729314
transform 1 0 760 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1513729314
transform 1 0 776 0 -1 1410
box 0 0 16 200
use NAND3X1  NAND3X1_39
timestamp 1513729314
transform 1 0 792 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_90
timestamp 1513729314
transform 1 0 856 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_1
timestamp 1513729314
transform -1 0 968 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_88
timestamp 1513729314
transform 1 0 968 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_5
timestamp 1513729314
transform -1 0 1080 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_45
timestamp 1513729314
transform -1 0 1112 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_50
timestamp 1513729314
transform 1 0 1112 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_120
timestamp 1513729314
transform -1 0 1224 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_86
timestamp 1513729314
transform -1 0 1272 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_1
timestamp 1513729314
transform -1 0 1336 0 -1 1410
box 0 0 64 200
use OAI22X1  OAI22X1_5
timestamp 1513729314
transform -1 0 1416 0 -1 1410
box 0 0 80 200
use OAI21X1  OAI21X1_19
timestamp 1513729314
transform 1 0 1416 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_138
timestamp 1513729314
transform 1 0 1480 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_89
timestamp 1513729314
transform 1 0 1544 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_37
timestamp 1513729314
transform 1 0 1608 0 -1 1410
box 0 0 48 200
use MUX2X1  MUX2X1_6
timestamp 1513729314
transform -1 0 1752 0 -1 1410
box 0 0 96 200
use NAND2X1  NAND2X1_42
timestamp 1513729314
transform -1 0 1800 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_1_0
timestamp 1513729314
transform -1 0 1816 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1513729314
transform -1 0 1832 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_129
timestamp 1513729314
transform -1 0 1896 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_28
timestamp 1513729314
transform 1 0 1896 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_81
timestamp 1513729314
transform -1 0 1992 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_19
timestamp 1513729314
transform -1 0 2056 0 -1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_18
timestamp 1513729314
transform -1 0 2120 0 -1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_4
timestamp 1513729314
transform 1 0 2120 0 -1 1410
box 0 0 80 200
use MUX2X1  MUX2X1_26
timestamp 1513729314
transform -1 0 2296 0 -1 1410
box 0 0 96 200
use MUX2X1  MUX2X1_15
timestamp 1513729314
transform -1 0 2392 0 -1 1410
box 0 0 96 200
use OAI21X1  OAI21X1_10
timestamp 1513729314
transform 1 0 2392 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_142
timestamp 1513729314
transform -1 0 2520 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_23
timestamp 1513729314
transform -1 0 2568 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_8
timestamp 1513729314
transform 1 0 2568 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_78
timestamp 1513729314
transform -1 0 2696 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_77
timestamp 1513729314
transform 1 0 2696 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_96
timestamp 1513729314
transform 1 0 2760 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_2_0
timestamp 1513729314
transform 1 0 2824 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1513729314
transform 1 0 2840 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_3
timestamp 1513729314
transform 1 0 2856 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_4
timestamp 1513729314
transform 1 0 2904 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_70
timestamp 1513729314
transform 1 0 2968 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_64
timestamp 1513729314
transform -1 0 3080 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_64
timestamp 1513729314
transform -1 0 3128 0 -1 1410
box 0 0 48 200
use OAI22X1  OAI22X1_2
timestamp 1513729314
transform 1 0 3128 0 -1 1410
box 0 0 80 200
use NOR2X1  NOR2X1_39
timestamp 1513729314
transform -1 0 3256 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_33
timestamp 1513729314
transform -1 0 3304 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_29
timestamp 1513729314
transform -1 0 3336 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_31
timestamp 1513729314
transform -1 0 3400 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_43
timestamp 1513729314
transform -1 0 3432 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_38
timestamp 1513729314
transform 1 0 3432 0 -1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_72
timestamp 1513729314
transform 1 0 3496 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_4
timestamp 1513729314
transform 1 0 3544 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_60
timestamp 1513729314
transform -1 0 3640 0 -1 1410
box 0 0 48 200
use FILL  FILL_7_1
timestamp 1513729314
transform -1 0 3656 0 -1 1410
box 0 0 16 200
use OR2X2  OR2X2_8
timestamp 1513729314
transform 1 0 8 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_21
timestamp 1513729314
transform 1 0 72 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_19
timestamp 1513729314
transform 1 0 136 0 1 1010
box 0 0 48 200
use INVX1  INVX1_24
timestamp 1513729314
transform -1 0 216 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_116
timestamp 1513729314
transform 1 0 216 0 1 1010
box 0 0 64 200
use INVX1  INVX1_22
timestamp 1513729314
transform 1 0 280 0 1 1010
box 0 0 32 200
use AOI22X1  AOI22X1_9
timestamp 1513729314
transform 1 0 312 0 1 1010
box 0 0 80 200
use AOI21X1  AOI21X1_13
timestamp 1513729314
transform 1 0 392 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_117
timestamp 1513729314
transform -1 0 520 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_121
timestamp 1513729314
transform -1 0 584 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_5
timestamp 1513729314
transform -1 0 648 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_98
timestamp 1513729314
transform 1 0 648 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_67
timestamp 1513729314
transform -1 0 760 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_85
timestamp 1513729314
transform 1 0 760 0 1 1010
box 0 0 48 200
use FILL  FILL_5_0_0
timestamp 1513729314
transform -1 0 824 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1513729314
transform -1 0 840 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_132
timestamp 1513729314
transform -1 0 904 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_46
timestamp 1513729314
transform -1 0 968 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_22
timestamp 1513729314
transform -1 0 1032 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_75
timestamp 1513729314
transform -1 0 1080 0 1 1010
box 0 0 48 200
use INVX1  INVX1_44
timestamp 1513729314
transform 1 0 1080 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_32
timestamp 1513729314
transform 1 0 1112 0 1 1010
box 0 0 48 200
use OR2X2  OR2X2_1
timestamp 1513729314
transform -1 0 1224 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_21
timestamp 1513729314
transform -1 0 1272 0 1 1010
box 0 0 48 200
use BUFX4  BUFX4_137
timestamp 1513729314
transform -1 0 1336 0 1 1010
box 0 0 64 200
use INVX8  INVX8_4
timestamp 1513729314
transform -1 0 1416 0 1 1010
box 0 0 80 200
use NAND3X1  NAND3X1_32
timestamp 1513729314
transform -1 0 1480 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_25
timestamp 1513729314
transform 1 0 1480 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1513729314
transform -1 0 1672 0 1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_1
timestamp 1513729314
transform -1 0 1720 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_73
timestamp 1513729314
transform -1 0 1784 0 1 1010
box 0 0 64 200
use FILL  FILL_5_1_0
timestamp 1513729314
transform -1 0 1800 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1513729314
transform -1 0 1816 0 1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_38
timestamp 1513729314
transform -1 0 1880 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_56
timestamp 1513729314
transform 1 0 1880 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_101
timestamp 1513729314
transform -1 0 1992 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_127
timestamp 1513729314
transform 1 0 1992 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_25
timestamp 1513729314
transform -1 0 2120 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_4
timestamp 1513729314
transform 1 0 2120 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_114
timestamp 1513729314
transform -1 0 2248 0 1 1010
box 0 0 64 200
use INVX1  INVX1_21
timestamp 1513729314
transform -1 0 2280 0 1 1010
box 0 0 32 200
use MUX2X1  MUX2X1_16
timestamp 1513729314
transform 1 0 2280 0 1 1010
box 0 0 96 200
use NAND3X1  NAND3X1_20
timestamp 1513729314
transform -1 0 2440 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_34
timestamp 1513729314
transform -1 0 2504 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_95
timestamp 1513729314
transform -1 0 2552 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_13
timestamp 1513729314
transform 1 0 2552 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_59
timestamp 1513729314
transform -1 0 2664 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_16
timestamp 1513729314
transform 1 0 2664 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_25
timestamp 1513729314
transform -1 0 2792 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_35
timestamp 1513729314
transform -1 0 2840 0 1 1010
box 0 0 48 200
use FILL  FILL_5_2_0
timestamp 1513729314
transform 1 0 2840 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1513729314
transform 1 0 2856 0 1 1010
box 0 0 16 200
use MUX2X1  MUX2X1_21
timestamp 1513729314
transform 1 0 2872 0 1 1010
box 0 0 96 200
use NAND2X1  NAND2X1_19
timestamp 1513729314
transform 1 0 2968 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_87
timestamp 1513729314
transform 1 0 3016 0 1 1010
box 0 0 48 200
use MUX2X1  MUX2X1_7
timestamp 1513729314
transform 1 0 3064 0 1 1010
box 0 0 96 200
use OAI21X1  OAI21X1_131
timestamp 1513729314
transform -1 0 3224 0 1 1010
box 0 0 64 200
use INVX1  INVX1_23
timestamp 1513729314
transform -1 0 3256 0 1 1010
box 0 0 32 200
use NAND2X1  NAND2X1_83
timestamp 1513729314
transform 1 0 3256 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_42
timestamp 1513729314
transform -1 0 3352 0 1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_3
timestamp 1513729314
transform 1 0 3352 0 1 1010
box 0 0 80 200
use MUX2X1  MUX2X1_9
timestamp 1513729314
transform 1 0 3432 0 1 1010
box 0 0 96 200
use MUX2X1  MUX2X1_10
timestamp 1513729314
transform 1 0 3528 0 1 1010
box 0 0 96 200
use FILL  FILL_6_1
timestamp 1513729314
transform 1 0 3624 0 1 1010
box 0 0 16 200
use FILL  FILL_6_2
timestamp 1513729314
transform 1 0 3640 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_110
timestamp 1513729314
transform -1 0 72 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_1
timestamp 1513729314
transform 1 0 72 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_41
timestamp 1513729314
transform 1 0 136 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_13
timestamp 1513729314
transform 1 0 200 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_25
timestamp 1513729314
transform 1 0 264 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_31
timestamp 1513729314
transform -1 0 344 0 -1 1010
box 0 0 32 200
use INVX1  INVX1_20
timestamp 1513729314
transform 1 0 344 0 -1 1010
box 0 0 32 200
use INVX8  INVX8_7
timestamp 1513729314
transform -1 0 456 0 -1 1010
box 0 0 80 200
use AND2X2  AND2X2_12
timestamp 1513729314
transform 1 0 456 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_2
timestamp 1513729314
transform -1 0 584 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_6
timestamp 1513729314
transform 1 0 584 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_38
timestamp 1513729314
transform -1 0 680 0 -1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_3
timestamp 1513729314
transform 1 0 680 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_58
timestamp 1513729314
transform -1 0 792 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_0_0
timestamp 1513729314
transform -1 0 808 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1513729314
transform -1 0 824 0 -1 1010
box 0 0 16 200
use AOI22X1  AOI22X1_7
timestamp 1513729314
transform -1 0 904 0 -1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_91
timestamp 1513729314
transform 1 0 904 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_11
timestamp 1513729314
transform 1 0 952 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_23
timestamp 1513729314
transform -1 0 1064 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_102
timestamp 1513729314
transform -1 0 1128 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_30
timestamp 1513729314
transform -1 0 1160 0 -1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_18
timestamp 1513729314
transform -1 0 1224 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_128
timestamp 1513729314
transform -1 0 1288 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_28
timestamp 1513729314
transform 1 0 1288 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_24
timestamp 1513729314
transform -1 0 1416 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_119
timestamp 1513729314
transform -1 0 1480 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_13
timestamp 1513729314
transform 1 0 1480 0 -1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_27
timestamp 1513729314
transform 1 0 1512 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_134
timestamp 1513729314
transform 1 0 1560 0 -1 1010
box 0 0 64 200
use INVX2  INVX2_9
timestamp 1513729314
transform 1 0 1624 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_90
timestamp 1513729314
transform -1 0 1720 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_14
timestamp 1513729314
transform 1 0 1720 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_57
timestamp 1513729314
transform 1 0 1784 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_1_0
timestamp 1513729314
transform -1 0 1848 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1513729314
transform -1 0 1864 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_81
timestamp 1513729314
transform -1 0 1928 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_17
timestamp 1513729314
transform 1 0 1928 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_143
timestamp 1513729314
transform -1 0 2040 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_44
timestamp 1513729314
transform 1 0 2040 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_73
timestamp 1513729314
transform 1 0 2088 0 -1 1010
box 0 0 48 200
use INVX1  INVX1_26
timestamp 1513729314
transform 1 0 2136 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_130
timestamp 1513729314
transform -1 0 2232 0 -1 1010
box 0 0 64 200
use MUX2X1  MUX2X1_12
timestamp 1513729314
transform 1 0 2232 0 -1 1010
box 0 0 96 200
use OAI21X1  OAI21X1_3
timestamp 1513729314
transform 1 0 2328 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_37
timestamp 1513729314
transform 1 0 2392 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_82
timestamp 1513729314
transform 1 0 2456 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_31
timestamp 1513729314
transform 1 0 2504 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_36
timestamp 1513729314
transform 1 0 2552 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_36
timestamp 1513729314
transform -1 0 2664 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_30
timestamp 1513729314
transform -1 0 2728 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_43
timestamp 1513729314
transform 1 0 2728 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_92
timestamp 1513729314
transform 1 0 2776 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_2_0
timestamp 1513729314
transform 1 0 2824 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1513729314
transform 1 0 2840 0 -1 1010
box 0 0 16 200
use OR2X2  OR2X2_6
timestamp 1513729314
transform 1 0 2856 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_28
timestamp 1513729314
transform 1 0 2920 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_7
timestamp 1513729314
transform 1 0 2952 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_30
timestamp 1513729314
transform 1 0 3016 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_32
timestamp 1513729314
transform -1 0 3144 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_30
timestamp 1513729314
transform -1 0 3192 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_34
timestamp 1513729314
transform 1 0 3192 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_40
timestamp 1513729314
transform 1 0 3256 0 -1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_29
timestamp 1513729314
transform 1 0 3288 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_79
timestamp 1513729314
transform -1 0 3384 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_66
timestamp 1513729314
transform 1 0 3384 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_6
timestamp 1513729314
transform 1 0 3448 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_47
timestamp 1513729314
transform 1 0 3512 0 -1 1010
box 0 0 32 200
use BUFX2  BUFX2_7
timestamp 1513729314
transform 1 0 3544 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_26
timestamp 1513729314
transform 1 0 3592 0 -1 1010
box 0 0 48 200
use FILL  FILL_5_1
timestamp 1513729314
transform -1 0 3656 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_107
timestamp 1513729314
transform -1 0 72 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_42
timestamp 1513729314
transform -1 0 136 0 1 610
box 0 0 64 200
use INVX4  INVX4_2
timestamp 1513729314
transform -1 0 184 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_21
timestamp 1513729314
transform 1 0 184 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_6
timestamp 1513729314
transform 1 0 248 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_51
timestamp 1513729314
transform 1 0 296 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_5
timestamp 1513729314
transform 1 0 360 0 1 610
box 0 0 48 200
use INVX4  INVX4_1
timestamp 1513729314
transform -1 0 456 0 1 610
box 0 0 48 200
use INVX1  INVX1_8
timestamp 1513729314
transform 1 0 456 0 1 610
box 0 0 32 200
use NAND3X1  NAND3X1_14
timestamp 1513729314
transform 1 0 488 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_17
timestamp 1513729314
transform 1 0 552 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_31
timestamp 1513729314
transform -1 0 680 0 1 610
box 0 0 64 200
use INVX4  INVX4_3
timestamp 1513729314
transform -1 0 728 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_129
timestamp 1513729314
transform -1 0 792 0 1 610
box 0 0 64 200
use FILL  FILL_3_0_0
timestamp 1513729314
transform -1 0 808 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1513729314
transform -1 0 824 0 1 610
box 0 0 16 200
use NAND3X1  NAND3X1_42
timestamp 1513729314
transform -1 0 888 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_38
timestamp 1513729314
transform -1 0 952 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_8
timestamp 1513729314
transform 1 0 952 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_7
timestamp 1513729314
transform -1 0 1064 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_1
timestamp 1513729314
transform 1 0 1064 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_45
timestamp 1513729314
transform 1 0 1112 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_13
timestamp 1513729314
transform -1 0 1224 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_54
timestamp 1513729314
transform 1 0 1224 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_6
timestamp 1513729314
transform 1 0 1272 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_55
timestamp 1513729314
transform -1 0 1400 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_48
timestamp 1513729314
transform 1 0 1400 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1513729314
transform 1 0 1464 0 1 610
box 0 0 64 200
use INVX1  INVX1_33
timestamp 1513729314
transform -1 0 1560 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_105
timestamp 1513729314
transform 1 0 1560 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_101
timestamp 1513729314
transform -1 0 1672 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_9
timestamp 1513729314
transform 1 0 1672 0 1 610
box 0 0 48 200
use MUX2X1  MUX2X1_18
timestamp 1513729314
transform 1 0 1720 0 1 610
box 0 0 96 200
use FILL  FILL_3_1_0
timestamp 1513729314
transform 1 0 1816 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1513729314
transform 1 0 1832 0 1 610
box 0 0 16 200
use MUX2X1  MUX2X1_8
timestamp 1513729314
transform 1 0 1848 0 1 610
box 0 0 96 200
use INVX1  INVX1_15
timestamp 1513729314
transform -1 0 1976 0 1 610
box 0 0 32 200
use NAND2X1  NAND2X1_16
timestamp 1513729314
transform -1 0 2024 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_33
timestamp 1513729314
transform -1 0 2088 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_18
timestamp 1513729314
transform 1 0 2088 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_5
timestamp 1513729314
transform 1 0 2136 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_2
timestamp 1513729314
transform 1 0 2184 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_3
timestamp 1513729314
transform 1 0 2232 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_85
timestamp 1513729314
transform 1 0 2296 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_21
timestamp 1513729314
transform -1 0 2424 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_11
timestamp 1513729314
transform -1 0 2472 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_92
timestamp 1513729314
transform -1 0 2536 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_7
timestamp 1513729314
transform 1 0 2536 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_100
timestamp 1513729314
transform 1 0 2600 0 1 610
box 0 0 48 200
use AOI21X1  AOI21X1_43
timestamp 1513729314
transform -1 0 2712 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_2
timestamp 1513729314
transform 1 0 2712 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_2
timestamp 1513729314
transform 1 0 2776 0 1 610
box 0 0 64 200
use FILL  FILL_3_2_0
timestamp 1513729314
transform 1 0 2840 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1513729314
transform 1 0 2856 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_13
timestamp 1513729314
transform 1 0 2872 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_90
timestamp 1513729314
transform -1 0 3000 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_134
timestamp 1513729314
transform 1 0 3000 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_47
timestamp 1513729314
transform 1 0 3064 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_63
timestamp 1513729314
transform -1 0 3192 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_58
timestamp 1513729314
transform 1 0 3192 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_102
timestamp 1513729314
transform -1 0 3304 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_95
timestamp 1513729314
transform -1 0 3368 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_79
timestamp 1513729314
transform -1 0 3432 0 1 610
box 0 0 64 200
use BUFX2  BUFX2_13
timestamp 1513729314
transform 1 0 3432 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_122
timestamp 1513729314
transform 1 0 3480 0 1 610
box 0 0 64 200
use BUFX2  BUFX2_32
timestamp 1513729314
transform 1 0 3544 0 1 610
box 0 0 48 200
use BUFX4  BUFX4_68
timestamp 1513729314
transform -1 0 3656 0 1 610
box 0 0 64 200
use INVX2  INVX2_6
timestamp 1513729314
transform 1 0 8 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_21
timestamp 1513729314
transform -1 0 104 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_17
timestamp 1513729314
transform -1 0 168 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_71
timestamp 1513729314
transform 1 0 168 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_41
timestamp 1513729314
transform -1 0 280 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_19
timestamp 1513729314
transform -1 0 344 0 -1 610
box 0 0 64 200
use OAI22X1  OAI22X1_1
timestamp 1513729314
transform 1 0 344 0 -1 610
box 0 0 80 200
use AOI21X1  AOI21X1_15
timestamp 1513729314
transform -1 0 488 0 -1 610
box 0 0 64 200
use INVX1  INVX1_1
timestamp 1513729314
transform -1 0 520 0 -1 610
box 0 0 32 200
use AND2X2  AND2X2_18
timestamp 1513729314
transform -1 0 584 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_6
timestamp 1513729314
transform 1 0 584 0 -1 610
box 0 0 48 200
use AOI21X1  AOI21X1_20
timestamp 1513729314
transform -1 0 696 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_122
timestamp 1513729314
transform -1 0 760 0 -1 610
box 0 0 64 200
use FILL  FILL_2_0_0
timestamp 1513729314
transform 1 0 760 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1513729314
transform 1 0 776 0 -1 610
box 0 0 16 200
use OAI21X1  OAI21X1_60
timestamp 1513729314
transform 1 0 792 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_5
timestamp 1513729314
transform 1 0 856 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_28
timestamp 1513729314
transform 1 0 920 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_109
timestamp 1513729314
transform 1 0 968 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_112
timestamp 1513729314
transform 1 0 1032 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_97
timestamp 1513729314
transform 1 0 1096 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_6
timestamp 1513729314
transform -1 0 1224 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_22
timestamp 1513729314
transform 1 0 1224 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_99
timestamp 1513729314
transform -1 0 1352 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_12
timestamp 1513729314
transform -1 0 1416 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_87
timestamp 1513729314
transform -1 0 1480 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1513729314
transform -1 0 1544 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_88
timestamp 1513729314
transform -1 0 1608 0 -1 610
box 0 0 64 200
use INVX2  INVX2_3
timestamp 1513729314
transform 1 0 1608 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_35
timestamp 1513729314
transform 1 0 1640 0 -1 610
box 0 0 64 200
use INVX1  INVX1_25
timestamp 1513729314
transform 1 0 1704 0 -1 610
box 0 0 32 200
use INVX1  INVX1_35
timestamp 1513729314
transform 1 0 1736 0 -1 610
box 0 0 32 200
use NAND2X1  NAND2X1_12
timestamp 1513729314
transform -1 0 1816 0 -1 610
box 0 0 48 200
use FILL  FILL_2_1_0
timestamp 1513729314
transform 1 0 1816 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1513729314
transform 1 0 1832 0 -1 610
box 0 0 16 200
use INVX8  INVX8_9
timestamp 1513729314
transform 1 0 1848 0 -1 610
box 0 0 80 200
use NAND3X1  NAND3X1_12
timestamp 1513729314
transform -1 0 1992 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1513729314
transform -1 0 2056 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_15
timestamp 1513729314
transform -1 0 2104 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_38
timestamp 1513729314
transform -1 0 2152 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_80
timestamp 1513729314
transform -1 0 2216 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_28
timestamp 1513729314
transform 1 0 2216 0 -1 610
box 0 0 64 200
use INVX8  INVX8_3
timestamp 1513729314
transform 1 0 2280 0 -1 610
box 0 0 80 200
use NAND3X1  NAND3X1_7
timestamp 1513729314
transform -1 0 2424 0 -1 610
box 0 0 64 200
use INVX8  INVX8_10
timestamp 1513729314
transform 1 0 2424 0 -1 610
box 0 0 80 200
use NOR2X1  NOR2X1_13
timestamp 1513729314
transform -1 0 2552 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_10
timestamp 1513729314
transform -1 0 2616 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_40
timestamp 1513729314
transform -1 0 2680 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_100
timestamp 1513729314
transform -1 0 2744 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_74
timestamp 1513729314
transform -1 0 2808 0 -1 610
box 0 0 64 200
use FILL  FILL_2_2_0
timestamp 1513729314
transform -1 0 2824 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1513729314
transform -1 0 2840 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_115
timestamp 1513729314
transform -1 0 2904 0 -1 610
box 0 0 64 200
use INVX8  INVX8_6
timestamp 1513729314
transform 1 0 2904 0 -1 610
box 0 0 80 200
use BUFX4  BUFX4_29
timestamp 1513729314
transform 1 0 2984 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_40
timestamp 1513729314
transform -1 0 3112 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_70
timestamp 1513729314
transform 1 0 3112 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_101
timestamp 1513729314
transform -1 0 3240 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_64
timestamp 1513729314
transform 1 0 3240 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_52
timestamp 1513729314
transform -1 0 3368 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_93
timestamp 1513729314
transform 1 0 3368 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_8
timestamp 1513729314
transform -1 0 3496 0 -1 610
box 0 0 64 200
use BUFX2  BUFX2_9
timestamp 1513729314
transform 1 0 3496 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_104
timestamp 1513729314
transform -1 0 3608 0 -1 610
box 0 0 64 200
use BUFX2  BUFX2_28
timestamp 1513729314
transform 1 0 3608 0 -1 610
box 0 0 48 200
use AND2X2  AND2X2_23
timestamp 1513729314
transform 1 0 8 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_18
timestamp 1513729314
transform 1 0 72 0 1 210
box 0 0 48 200
use INVX2  INVX2_8
timestamp 1513729314
transform 1 0 120 0 1 210
box 0 0 32 200
use AOI22X1  AOI22X1_2
timestamp 1513729314
transform -1 0 232 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_86
timestamp 1513729314
transform 1 0 232 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_1
timestamp 1513729314
transform 1 0 296 0 1 210
box 0 0 80 200
use INVX1  INVX1_11
timestamp 1513729314
transform -1 0 408 0 1 210
box 0 0 32 200
use NAND3X1  NAND3X1_6
timestamp 1513729314
transform 1 0 408 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_30
timestamp 1513729314
transform -1 0 536 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_139
timestamp 1513729314
transform 1 0 536 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_14
timestamp 1513729314
transform 1 0 600 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_15
timestamp 1513729314
transform 1 0 648 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_12
timestamp 1513729314
transform 1 0 712 0 1 210
box 0 0 64 200
use FILL  FILL_1_0_0
timestamp 1513729314
transform 1 0 776 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1513729314
transform 1 0 792 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_124
timestamp 1513729314
transform 1 0 808 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_136
timestamp 1513729314
transform 1 0 872 0 1 210
box 0 0 64 200
use INVX1  INVX1_18
timestamp 1513729314
transform 1 0 936 0 1 210
box 0 0 32 200
use AOI21X1  AOI21X1_9
timestamp 1513729314
transform 1 0 968 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_110
timestamp 1513729314
transform -1 0 1096 0 1 210
box 0 0 64 200
use AOI21X1  AOI21X1_1
timestamp 1513729314
transform 1 0 1096 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_1
timestamp 1513729314
transform -1 0 1224 0 1 210
box 0 0 64 200
use INVX8  INVX8_2
timestamp 1513729314
transform -1 0 1304 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_83
timestamp 1513729314
transform -1 0 1368 0 1 210
box 0 0 64 200
use INVX1  INVX1_10
timestamp 1513729314
transform 1 0 1368 0 1 210
box 0 0 32 200
use NOR2X1  NOR2X1_3
timestamp 1513729314
transform 1 0 1400 0 1 210
box 0 0 48 200
use INVX1  INVX1_7
timestamp 1513729314
transform -1 0 1480 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_84
timestamp 1513729314
transform -1 0 1544 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_17
timestamp 1513729314
transform 1 0 1544 0 1 210
box 0 0 64 200
use INVX1  INVX1_6
timestamp 1513729314
transform 1 0 1608 0 1 210
box 0 0 32 200
use AOI21X1  AOI21X1_42
timestamp 1513729314
transform 1 0 1640 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_71
timestamp 1513729314
transform 1 0 1704 0 1 210
box 0 0 64 200
use INVX2  INVX2_7
timestamp 1513729314
transform 1 0 1768 0 1 210
box 0 0 32 200
use FILL  FILL_1_1_0
timestamp 1513729314
transform -1 0 1816 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1513729314
transform -1 0 1832 0 1 210
box 0 0 16 200
use AOI21X1  AOI21X1_23
timestamp 1513729314
transform -1 0 1896 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_39
timestamp 1513729314
transform 1 0 1896 0 1 210
box 0 0 64 200
use INVX1  INVX1_14
timestamp 1513729314
transform -1 0 1992 0 1 210
box 0 0 32 200
use INVX2  INVX2_5
timestamp 1513729314
transform 1 0 1992 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_56
timestamp 1513729314
transform -1 0 2088 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_94
timestamp 1513729314
transform 1 0 2088 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_11
timestamp 1513729314
transform -1 0 2216 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_76
timestamp 1513729314
transform 1 0 2216 0 1 210
box 0 0 64 200
use INVX8  INVX8_8
timestamp 1513729314
transform 1 0 2280 0 1 210
box 0 0 80 200
use BUFX4  BUFX4_72
timestamp 1513729314
transform 1 0 2360 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_45
timestamp 1513729314
transform 1 0 2424 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_56
timestamp 1513729314
transform -1 0 2552 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_17
timestamp 1513729314
transform 1 0 2552 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_82
timestamp 1513729314
transform -1 0 2664 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_50
timestamp 1513729314
transform 1 0 2664 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_3
timestamp 1513729314
transform -1 0 2776 0 1 210
box 0 0 48 200
use BUFX4  BUFX4_41
timestamp 1513729314
transform 1 0 2776 0 1 210
box 0 0 64 200
use FILL  FILL_1_2_0
timestamp 1513729314
transform 1 0 2840 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1513729314
transform 1 0 2856 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_73
timestamp 1513729314
transform 1 0 2872 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_81
timestamp 1513729314
transform 1 0 2936 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_60
timestamp 1513729314
transform 1 0 3000 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_78
timestamp 1513729314
transform 1 0 3064 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_19
timestamp 1513729314
transform 1 0 3128 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_54
timestamp 1513729314
transform 1 0 3192 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_131
timestamp 1513729314
transform 1 0 3256 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_26
timestamp 1513729314
transform -1 0 3384 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_62
timestamp 1513729314
transform -1 0 3448 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_87
timestamp 1513729314
transform 1 0 3448 0 1 210
box 0 0 64 200
use BUFX2  BUFX2_1
timestamp 1513729314
transform 1 0 3512 0 1 210
box 0 0 48 200
use BUFX2  BUFX2_20
timestamp 1513729314
transform 1 0 3560 0 1 210
box 0 0 48 200
use FILL  FILL_2_1
timestamp 1513729314
transform 1 0 3608 0 1 210
box 0 0 16 200
use FILL  FILL_2_2
timestamp 1513729314
transform 1 0 3624 0 1 210
box 0 0 16 200
use FILL  FILL_2_3
timestamp 1513729314
transform 1 0 3640 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_5
timestamp 1513729314
transform -1 0 72 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_89
timestamp 1513729314
transform -1 0 136 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_36
timestamp 1513729314
transform -1 0 200 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_22
timestamp 1513729314
transform 1 0 200 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_15
timestamp 1513729314
transform 1 0 264 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_21
timestamp 1513729314
transform 1 0 328 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_24
timestamp 1513729314
transform -1 0 456 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_22
timestamp 1513729314
transform 1 0 456 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_23
timestamp 1513729314
transform 1 0 520 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_40
timestamp 1513729314
transform 1 0 584 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_108
timestamp 1513729314
transform -1 0 696 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_133
timestamp 1513729314
transform -1 0 760 0 -1 210
box 0 0 64 200
use FILL  FILL_0_0_0
timestamp 1513729314
transform 1 0 760 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1513729314
transform 1 0 776 0 -1 210
box 0 0 16 200
use BUFX4  BUFX4_135
timestamp 1513729314
transform 1 0 792 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_106
timestamp 1513729314
transform -1 0 920 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_20
timestamp 1513729314
transform -1 0 984 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_107
timestamp 1513729314
transform -1 0 1048 0 -1 210
box 0 0 64 200
use AOI21X1  AOI21X1_47
timestamp 1513729314
transform 1 0 1048 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_98
timestamp 1513729314
transform -1 0 1176 0 -1 210
box 0 0 64 200
use INVX1  INVX1_17
timestamp 1513729314
transform -1 0 1208 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_93
timestamp 1513729314
transform -1 0 1272 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_94
timestamp 1513729314
transform -1 0 1336 0 -1 210
box 0 0 64 200
use INVX1  INVX1_16
timestamp 1513729314
transform 1 0 1336 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_10
timestamp 1513729314
transform -1 0 1416 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_99
timestamp 1513729314
transform -1 0 1480 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_8
timestamp 1513729314
transform -1 0 1544 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_47
timestamp 1513729314
transform 1 0 1544 0 -1 210
box 0 0 48 200
use INVX1  INVX1_5
timestamp 1513729314
transform -1 0 1624 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_23
timestamp 1513729314
transform -1 0 1688 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_15
timestamp 1513729314
transform -1 0 1752 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_16
timestamp 1513729314
transform 1 0 1752 0 -1 210
box 0 0 64 200
use FILL  FILL_0_1_0
timestamp 1513729314
transform -1 0 1832 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1513729314
transform -1 0 1848 0 -1 210
box 0 0 16 200
use OAI21X1  OAI21X1_27
timestamp 1513729314
transform -1 0 1912 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_19
timestamp 1513729314
transform 1 0 1912 0 -1 210
box 0 0 64 200
use INVX1  INVX1_12
timestamp 1513729314
transform 1 0 1976 0 -1 210
box 0 0 32 200
use NOR2X1  NOR2X1_7
timestamp 1513729314
transform -1 0 2056 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_46
timestamp 1513729314
transform 1 0 2056 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_12
timestamp 1513729314
transform 1 0 2120 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_31
timestamp 1513729314
transform 1 0 2168 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_57
timestamp 1513729314
transform 1 0 2216 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_11
timestamp 1513729314
transform 1 0 2280 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_30
timestamp 1513729314
transform 1 0 2328 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_6
timestamp 1513729314
transform 1 0 2376 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_25
timestamp 1513729314
transform 1 0 2424 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_75
timestamp 1513729314
transform -1 0 2536 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_10
timestamp 1513729314
transform 1 0 2536 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_17
timestamp 1513729314
transform -1 0 2664 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_22
timestamp 1513729314
transform -1 0 2712 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_16
timestamp 1513729314
transform 1 0 2712 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_16
timestamp 1513729314
transform 1 0 2760 0 -1 210
box 0 0 64 200
use FILL  FILL_0_2_0
timestamp 1513729314
transform 1 0 2824 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1513729314
transform 1 0 2840 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_35
timestamp 1513729314
transform 1 0 2856 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_49
timestamp 1513729314
transform 1 0 2904 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_15
timestamp 1513729314
transform 1 0 2968 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_34
timestamp 1513729314
transform 1 0 3016 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_43
timestamp 1513729314
transform -1 0 3128 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_84
timestamp 1513729314
transform -1 0 3192 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_18
timestamp 1513729314
transform 1 0 3192 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_37
timestamp 1513729314
transform 1 0 3240 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_38
timestamp 1513729314
transform 1 0 3288 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_19
timestamp 1513729314
transform -1 0 3384 0 -1 210
box 0 0 48 200
use BUFX4  BUFX4_20
timestamp 1513729314
transform -1 0 3448 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_55
timestamp 1513729314
transform -1 0 3512 0 -1 210
box 0 0 64 200
use MUX2X1  MUX2X1_25
timestamp 1513729314
transform 1 0 3512 0 -1 210
box 0 0 96 200
use FILL  FILL_1_1
timestamp 1513729314
transform -1 0 3624 0 -1 210
box 0 0 16 200
use FILL  FILL_1_2
timestamp 1513729314
transform -1 0 3640 0 -1 210
box 0 0 16 200
use FILL  FILL_1_3
timestamp 1513729314
transform -1 0 3656 0 -1 210
box 0 0 16 200
<< labels >>
flabel space 996 42 1004 136 6 FreeSans 48 0 0 0 vdd
port 0 nsew
flabel space 2020 42 2028 136 6 FreeSans 48 0 0 0 gnd
port 1 nsew
flabel metal2 1232 -40 1232 -40 7 FreeSans 48 270 0 0 ULA_A<0>
port 2 nsew
flabel metal2 2224 2460 2224 2460 3 FreeSans 48 90 0 0 ULA_A<1>
port 3 nsew
flabel metal2 1568 2460 1568 2460 3 FreeSans 48 90 0 0 ULA_A<2>
port 4 nsew
flabel metal2 1280 2460 1280 2460 3 FreeSans 48 90 0 0 ULA_A<3>
port 5 nsew
flabel metal2 1696 2460 1696 2460 3 FreeSans 48 90 0 0 ULA_A<4>
port 6 nsew
flabel metal2 1504 2460 1504 2460 3 FreeSans 48 90 0 0 ULA_A<5>
port 7 nsew
flabel metal2 1632 2460 1632 2460 3 FreeSans 48 90 0 0 ULA_A<6>
port 8 nsew
flabel metal2 1808 2460 1808 2460 3 FreeSans 48 90 0 0 ULA_A<7>
port 9 nsew
flabel metal2 1728 -40 1728 -40 7 FreeSans 48 270 0 0 ULA_A<8>
port 10 nsew
flabel metal2 1536 -40 1536 -40 7 FreeSans 48 270 0 0 ULA_A<9>
port 11 nsew
flabel metal2 1920 -40 1920 -40 7 FreeSans 48 270 0 0 ULA_A<10>
port 12 nsew
flabel metal2 1376 -40 1376 -40 7 FreeSans 48 270 0 0 ULA_A<11>
port 13 nsew
flabel metal2 1792 -40 1792 -40 7 FreeSans 48 270 0 0 ULA_A<12>
port 14 nsew
flabel metal3 -48 1160 -48 1160 7 FreeSans 48 0 0 0 ULA_A<13>
port 15 nsew
flabel metal2 592 -40 592 -40 7 FreeSans 48 270 0 0 ULA_A<14>
port 16 nsew
flabel metal3 -48 980 -48 980 7 FreeSans 48 0 0 0 ULA_A<15>
port 17 nsew
flabel metal2 2144 2460 2144 2460 3 FreeSans 48 90 0 0 ULA_B<0>
port 18 nsew
flabel metal2 2592 2460 2592 2460 3 FreeSans 48 90 0 0 ULA_B<1>
port 19 nsew
flabel metal2 816 2460 816 2460 3 FreeSans 48 90 0 0 ULA_B<2>
port 20 nsew
flabel metal2 688 2460 688 2460 3 FreeSans 48 90 0 0 ULA_B<3>
port 21 nsew
flabel metal3 -48 1320 -48 1320 7 FreeSans 48 0 0 0 ULA_B<4>
port 22 nsew
flabel metal3 -48 1780 -48 1780 7 FreeSans 48 0 0 0 ULA_B<5>
port 23 nsew
flabel metal2 1136 2460 1136 2460 3 FreeSans 48 90 0 0 ULA_B<6>
port 24 nsew
flabel metal2 944 2460 944 2460 3 FreeSans 48 90 0 0 ULA_B<7>
port 25 nsew
flabel metal2 1664 -40 1664 -40 7 FreeSans 48 270 0 0 ULA_B<8>
port 26 nsew
flabel metal2 1472 -40 1472 -40 7 FreeSans 48 270 0 0 ULA_B<9>
port 27 nsew
flabel metal2 1856 -40 1856 -40 7 FreeSans 48 270 0 0 ULA_B<10>
port 28 nsew
flabel metal2 1312 -40 1312 -40 7 FreeSans 48 270 0 0 ULA_B<11>
port 29 nsew
flabel metal2 944 -40 944 -40 7 FreeSans 48 270 0 0 ULA_B<12>
port 30 nsew
flabel metal3 -48 1080 -48 1080 7 FreeSans 48 0 0 0 ULA_B<13>
port 31 nsew
flabel metal2 656 -40 656 -40 7 FreeSans 48 270 0 0 ULA_B<14>
port 32 nsew
flabel metal3 -48 920 -48 920 7 FreeSans 48 0 0 0 ULA_B<15>
port 33 nsew
flabel metal2 768 -40 768 -40 7 FreeSans 48 270 0 0 ULA_ctrl<0>
port 34 nsew
flabel metal3 -48 520 -48 520 7 FreeSans 48 0 0 0 ULA_ctrl<1>
port 35 nsew
flabel metal2 192 -40 192 -40 7 FreeSans 48 270 0 0 ULA_ctrl<2>
port 36 nsew
flabel metal3 -48 300 -48 300 7 FreeSans 48 0 0 0 ULA_ctrl<3>
port 37 nsew
flabel metal3 3712 320 3712 320 3 FreeSans 48 0 0 0 ULA_OUT<0>
port 38 nsew
flabel metal2 3280 2460 3280 2460 3 FreeSans 48 90 0 0 ULA_OUT<1>
port 39 nsew
flabel metal2 2672 -40 2672 -40 7 FreeSans 48 270 0 0 ULA_OUT<2>
port 40 nsew
flabel metal3 -48 1720 -48 1720 7 FreeSans 48 0 0 0 ULA_OUT<3>
port 41 nsew
flabel metal2 3376 2460 3376 2460 3 FreeSans 48 90 0 0 ULA_OUT<4>
port 42 nsew
flabel metal2 2464 -40 2464 -40 7 FreeSans 48 270 0 0 ULA_OUT<5>
port 43 nsew
flabel metal3 3712 920 3712 920 3 FreeSans 48 0 0 0 ULA_OUT<6>
port 44 nsew
flabel metal2 3488 2460 3488 2460 3 FreeSans 48 90 0 0 ULA_OUT<7>
port 45 nsew
flabel metal3 3712 520 3712 520 3 FreeSans 48 0 0 0 ULA_OUT<8>
port 46 nsew
flabel metal2 320 2460 320 2460 3 FreeSans 48 90 0 0 ULA_OUT<9>
port 47 nsew
flabel metal2 2368 -40 2368 -40 7 FreeSans 48 270 0 0 ULA_OUT<10>
port 48 nsew
flabel metal2 2208 -40 2208 -40 7 FreeSans 48 270 0 0 ULA_OUT<11>
port 49 nsew
flabel metal3 3712 720 3712 720 3 FreeSans 48 0 0 0 ULA_OUT<12>
port 50 nsew
flabel metal3 -48 2120 -48 2120 7 FreeSans 48 0 0 0 ULA_OUT<13>
port 51 nsew
flabel metal2 3024 -40 3024 -40 7 FreeSans 48 270 0 0 ULA_OUT<14>
port 52 nsew
flabel metal2 2864 -40 2864 -40 7 FreeSans 48 270 0 0 ULA_OUT<15>
port 53 nsew
flabel metal3 -48 2320 -48 2320 7 FreeSans 48 0 0 0 ULA_flags<0>
port 54 nsew
flabel metal2 3280 -40 3280 -40 7 FreeSans 48 270 0 0 ULA_flags<1>
port 55 nsew
flabel metal2 3344 -40 3344 -40 7 FreeSans 48 270 0 0 ULA_flags<2>
port 56 nsew
<< end >>
