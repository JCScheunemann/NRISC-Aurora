magic
tech scmos
magscale 1 4
timestamp 1515882711
<< metal1 >>
rect 2973 5577 3000 5583
rect 3213 5577 3224 5583
rect 1869 5517 1912 5523
rect 173 5497 184 5503
rect 1293 5497 1320 5503
rect 3000 5497 3027 5503
rect 3613 5503 3619 5523
rect 3581 5497 3619 5503
rect 3725 5503 3731 5523
rect 4717 5517 4771 5523
rect 4781 5517 4792 5523
rect 3656 5497 3699 5503
rect 3725 5497 3779 5503
rect 3912 5497 3939 5503
rect 4376 5497 4387 5503
rect 4541 5497 4568 5503
rect 4877 5497 4904 5503
rect 5085 5503 5091 5523
rect 5213 5517 5235 5523
rect 5085 5497 5139 5503
rect 5197 5497 5208 5503
rect 5229 5503 5235 5517
rect 5229 5497 5267 5503
rect 5608 5497 5635 5503
rect 6029 5503 6035 5523
rect 6029 5497 6115 5503
rect 6248 5497 6275 5503
rect 6456 5497 6483 5503
rect 6605 5503 6611 5523
rect 6605 5497 6659 5503
rect 6957 5503 6963 5523
rect 6925 5497 6963 5503
rect 6989 5497 7016 5503
rect 7160 5497 7187 5503
rect 7576 5497 7603 5503
rect 284 5477 324 5483
rect 781 5477 819 5483
rect 861 5477 899 5483
rect 140 5468 148 5472
rect 556 5463 564 5472
rect 556 5457 584 5463
rect 781 5457 787 5477
rect 893 5463 899 5477
rect 1704 5477 1715 5483
rect 2744 5477 2771 5483
rect 3128 5477 3139 5483
rect 3789 5477 3828 5483
rect 3820 5472 3828 5477
rect 4444 5477 4484 5483
rect 4988 5477 5016 5483
rect 4988 5472 4996 5477
rect 5976 5477 5987 5483
rect 6136 5477 6164 5483
rect 6156 5472 6164 5477
rect 7048 5477 7076 5483
rect 7068 5472 7076 5477
rect 7272 5477 7284 5483
rect 893 5457 947 5463
rect 1164 5463 1172 5472
rect 1372 5468 1380 5472
rect 1144 5457 1172 5463
rect 1468 5463 1476 5472
rect 2412 5468 2420 5472
rect 1468 5457 1496 5463
rect 3388 5466 3396 5472
rect 4300 5468 4308 5472
rect 2716 5463 2724 5466
rect 2716 5457 2755 5463
rect 5452 5466 5460 5472
rect 5756 5463 5764 5472
rect 5756 5457 5784 5463
rect 6844 5463 6852 5472
rect 6824 5457 6852 5463
rect 7964 5463 7972 5472
rect 7944 5457 7972 5463
rect 493 5437 504 5443
rect 1869 5437 1880 5443
rect 3352 5437 3363 5443
rect 5512 5437 5523 5443
rect 6360 5437 6371 5443
rect 7480 5437 7491 5443
rect 2157 5377 2168 5383
rect 2877 5377 2888 5383
rect 2941 5377 2984 5383
rect 3208 5377 3219 5383
rect 3917 5377 3928 5383
rect 4440 5377 4451 5383
rect 60 5357 88 5363
rect 60 5348 68 5357
rect 237 5357 291 5363
rect 264 5337 307 5343
rect 317 5337 376 5343
rect 413 5343 419 5363
rect 541 5357 579 5363
rect 796 5357 808 5363
rect 796 5354 804 5357
rect 413 5337 451 5343
rect 461 5337 504 5343
rect 360 5317 371 5323
rect 461 5317 467 5337
rect 877 5343 883 5363
rect 1389 5357 1400 5363
rect 1613 5357 1651 5363
rect 2397 5357 2408 5363
rect 3533 5357 3544 5363
rect 4104 5357 4116 5363
rect 4108 5354 4116 5357
rect 4540 5348 4548 5354
rect 6668 5348 6676 5354
rect 1036 5343 1044 5348
rect 877 5337 915 5343
rect 1005 5337 1044 5343
rect 1341 5337 1352 5343
rect 2349 5337 2387 5343
rect 2408 5337 2451 5343
rect 2504 5337 2515 5343
rect 3373 5337 3411 5343
rect 4312 5337 4323 5343
rect 488 5317 499 5323
rect 925 5317 968 5323
rect 1277 5317 1331 5323
rect 1277 5297 1283 5317
rect 1944 5317 2019 5323
rect 2269 5317 2307 5323
rect 2184 5297 2195 5303
rect 2301 5297 2307 5317
rect 2584 5317 2611 5323
rect 3069 5317 3096 5323
rect 3293 5317 3331 5323
rect 2381 5297 2408 5303
rect 3325 5297 3331 5317
rect 3965 5317 4035 5323
rect 4061 5317 4088 5323
rect 3805 5297 3816 5303
rect 3981 5297 4008 5303
rect 4029 5297 4035 5317
rect 4200 5317 4227 5323
rect 4333 5317 4371 5323
rect 4365 5297 4371 5317
rect 4477 5317 4488 5323
rect 4813 5323 4819 5343
rect 5768 5337 5779 5343
rect 6365 5337 6403 5343
rect 6989 5337 7000 5343
rect 7100 5343 7108 5348
rect 7048 5337 7108 5343
rect 7820 5343 7828 5348
rect 7800 5337 7828 5343
rect 4792 5317 4819 5323
rect 4941 5317 4968 5323
rect 5052 5317 5112 5323
rect 5052 5314 5060 5317
rect 5245 5317 5283 5323
rect 5277 5297 5283 5317
rect 5485 5317 5523 5323
rect 5517 5297 5523 5317
rect 5645 5317 5672 5323
rect 5805 5317 5832 5323
rect 6157 5317 6200 5323
rect 6221 5317 6259 5323
rect 5912 5297 5923 5303
rect 6253 5297 6259 5317
rect 6445 5317 6483 5323
rect 6445 5297 6451 5317
rect 6700 5317 6755 5323
rect 6700 5314 6708 5317
rect 6813 5317 6824 5323
rect 6989 5317 7027 5323
rect 6989 5297 6995 5317
rect 7192 5317 7219 5323
rect 7405 5317 7443 5323
rect 7405 5297 7411 5317
rect 7693 5317 7731 5323
rect 7693 5297 7699 5317
rect 7912 5317 7939 5323
rect 3142 5276 3144 5284
rect 2157 5237 2168 5243
rect 3181 5237 3192 5243
rect 3165 5177 3176 5183
rect 5096 5136 5098 5144
rect 7720 5136 7722 5144
rect 333 5097 344 5103
rect 429 5097 456 5103
rect 637 5097 664 5103
rect 1101 5103 1107 5123
rect 1101 5097 1155 5103
rect 1485 5103 1491 5123
rect 1485 5097 1539 5103
rect 2333 5103 2339 5123
rect 3037 5117 3064 5123
rect 2333 5097 2387 5103
rect 3261 5097 3288 5103
rect 3372 5103 3380 5106
rect 3372 5097 3384 5103
rect 3437 5103 3443 5123
rect 3405 5097 3443 5103
rect 3640 5097 3667 5103
rect 3885 5097 3896 5103
rect 4061 5103 4067 5123
rect 3997 5097 4067 5103
rect 4397 5103 4403 5123
rect 4365 5097 4403 5103
rect 4589 5103 4595 5123
rect 4536 5097 4563 5103
rect 4589 5097 4643 5103
rect 4776 5097 4803 5103
rect 4909 5097 4920 5103
rect 5144 5097 5171 5103
rect 5288 5097 5304 5103
rect 5597 5097 5608 5103
rect 5805 5097 5832 5103
rect 5981 5103 5987 5123
rect 5981 5097 6019 5103
rect 6269 5097 6296 5103
rect 6477 5097 6488 5103
rect 6653 5103 6659 5123
rect 6653 5097 6707 5103
rect 6856 5097 6867 5103
rect 7144 5097 7171 5103
rect 7293 5103 7299 5123
rect 7565 5117 7603 5123
rect 7293 5097 7347 5103
rect 7629 5097 7640 5103
rect 7768 5097 7795 5103
rect 237 5077 275 5083
rect 204 5063 212 5066
rect 204 5057 216 5063
rect 269 5063 275 5077
rect 748 5077 787 5083
rect 797 5077 808 5083
rect 748 5072 756 5077
rect 1213 5077 1252 5083
rect 1244 5072 1252 5077
rect 1597 5077 1636 5083
rect 1628 5072 1636 5077
rect 1965 5077 2008 5083
rect 2205 5077 2232 5083
rect 2333 5077 2344 5083
rect 2604 5077 2616 5083
rect 2604 5072 2612 5077
rect 3053 5077 3080 5083
rect 3372 5077 3395 5083
rect 3372 5072 3380 5077
rect 3549 5077 3560 5083
rect 3576 5077 3587 5083
rect 3901 5077 3939 5083
rect 3960 5077 3987 5083
rect 4316 5077 4328 5083
rect 4589 5077 4616 5083
rect 4664 5077 4692 5083
rect 4684 5072 4692 5077
rect 6157 5077 6168 5083
rect 6200 5077 6212 5083
rect 6717 5077 6756 5083
rect 6748 5072 6756 5077
rect 7357 5077 7368 5083
rect 7405 5077 7432 5083
rect 7645 5077 7656 5083
rect 860 5068 868 5072
rect 6348 5068 6356 5072
rect 6556 5068 6564 5072
rect 269 5057 291 5063
rect 7084 5063 7092 5072
rect 7084 5057 7112 5063
rect 1192 5037 1203 5043
rect 1576 5037 1587 5043
rect 2168 5037 2179 5043
rect 4136 5037 4147 5043
rect 5016 5037 5059 5043
rect 5528 5037 5539 5043
rect 6744 5037 6755 5043
rect 7880 5037 7891 5043
rect 477 4957 515 4963
rect 525 4957 536 4963
rect 732 4957 744 4963
rect 732 4954 740 4957
rect 813 4943 819 4963
rect 893 4957 979 4963
rect 1261 4957 1272 4963
rect 2876 4957 2915 4963
rect 2876 4954 2884 4957
rect 2572 4948 2580 4954
rect 3276 4948 3284 4954
rect 4300 4948 4308 4954
rect 7565 4957 7604 4963
rect 7596 4954 7604 4957
rect 7372 4948 7380 4952
rect 7628 4948 7636 4952
rect 813 4937 851 4943
rect 1149 4937 1176 4943
rect 1868 4943 1876 4948
rect 1868 4937 1907 4943
rect 1917 4937 1971 4943
rect 2200 4937 2211 4943
rect 2280 4937 2291 4943
rect 4077 4937 4115 4943
rect 4332 4943 4340 4948
rect 4332 4937 4371 4943
rect 4525 4937 4552 4943
rect 4605 4937 4648 4943
rect 5020 4943 5028 4948
rect 4968 4937 5028 4943
rect 5592 4937 5603 4943
rect 7772 4937 7784 4943
rect 621 4917 632 4923
rect 1133 4917 1160 4923
rect 1757 4917 1784 4923
rect 2173 4917 2228 4923
rect 2220 4916 2228 4917
rect 2333 4917 2387 4923
rect 397 4897 408 4903
rect 1416 4897 1427 4903
rect 1469 4897 1491 4903
rect 2013 4897 2024 4903
rect 2333 4897 2339 4917
rect 2653 4917 2680 4923
rect 3197 4917 3252 4923
rect 3244 4914 3252 4917
rect 3453 4917 3491 4923
rect 2904 4897 2963 4903
rect 2973 4897 3043 4903
rect 3485 4897 3491 4917
rect 3965 4917 4035 4923
rect 4061 4917 4072 4923
rect 4029 4897 4035 4917
rect 4221 4917 4248 4923
rect 4381 4917 4419 4923
rect 4413 4897 4419 4917
rect 4909 4917 4947 4923
rect 4909 4897 4915 4917
rect 5112 4917 5139 4923
rect 5357 4917 5384 4923
rect 5496 4917 5507 4923
rect 5693 4917 5731 4923
rect 5261 4897 5272 4903
rect 5725 4897 5731 4917
rect 5853 4917 5880 4923
rect 5960 4917 5971 4923
rect 6152 4917 6179 4923
rect 6301 4917 6339 4923
rect 6301 4897 6307 4917
rect 6360 4917 6387 4923
rect 6493 4917 6547 4923
rect 6493 4897 6499 4917
rect 7448 4917 7459 4923
rect 7992 4897 8019 4903
rect 109 4877 184 4883
rect 1069 4877 1108 4883
rect 1069 4857 1075 4877
rect 1432 4877 1459 4883
rect 2838 4876 2840 4884
rect 1917 4837 1944 4843
rect 3917 4837 3928 4843
rect 6056 4837 6067 4843
rect 7192 4737 7219 4743
rect 840 4717 867 4723
rect 909 4717 936 4723
rect 669 4697 696 4703
rect 1032 4697 1043 4703
rect 1069 4703 1075 4723
rect 1773 4717 1795 4723
rect 2296 4717 2307 4723
rect 3256 4717 3315 4723
rect 3389 4717 3427 4723
rect 5773 4717 5784 4723
rect 5960 4717 5971 4723
rect 7037 4717 7064 4723
rect 1069 4697 1123 4703
rect 1437 4697 1448 4703
rect 1693 4697 1704 4703
rect 1992 4697 2024 4703
rect 2648 4697 2675 4703
rect 2796 4703 2804 4708
rect 2796 4697 2824 4703
rect 2845 4697 2856 4703
rect 3740 4703 3748 4708
rect 3740 4697 3752 4703
rect 3789 4697 3827 4703
rect 3916 4703 3924 4708
rect 3916 4697 3928 4703
rect 3965 4697 3976 4703
rect 4173 4697 4184 4703
rect 4252 4703 4260 4708
rect 4252 4697 4264 4703
rect 4301 4697 4339 4703
rect 4540 4703 4548 4708
rect 4540 4697 4552 4703
rect 4648 4697 4659 4703
rect 5405 4697 5416 4703
rect 5496 4697 5507 4703
rect 5576 4697 5619 4703
rect 61 4677 72 4683
rect 1965 4677 1992 4683
rect 2424 4677 2451 4683
rect 2504 4677 2515 4683
rect 2525 4677 2564 4683
rect 2556 4672 2564 4677
rect 2989 4677 3032 4683
rect 3341 4677 3368 4683
rect 5144 4677 5155 4683
rect 5165 4677 5176 4683
rect 748 4668 756 4672
rect 77 4657 115 4663
rect 1309 4657 1347 4663
rect 1629 4657 1667 4663
rect 2236 4663 2244 4672
rect 2216 4657 2244 4663
rect 3228 4663 3236 4666
rect 3228 4657 3267 4663
rect 3644 4663 3652 4672
rect 4764 4668 4772 4672
rect 3624 4657 3652 4663
rect 5021 4657 5107 4663
rect 5165 4657 5171 4677
rect 5613 4677 5619 4697
rect 6024 4697 6067 4703
rect 6365 4697 6392 4703
rect 6456 4697 6472 4703
rect 6552 4697 6595 4703
rect 7149 4703 7155 4723
rect 7517 4717 7528 4723
rect 7128 4697 7155 4703
rect 7304 4697 7331 4703
rect 7528 4697 7555 4703
rect 7773 4703 7779 4723
rect 7773 4697 7811 4703
rect 7996 4706 8004 4712
rect 5997 4677 6040 4683
rect 6381 4677 6392 4683
rect 6413 4677 6483 4683
rect 6680 4677 6691 4683
rect 7181 4677 7220 4683
rect 7212 4672 7220 4677
rect 7693 4677 7704 4683
rect 7773 4677 7784 4683
rect 5293 4657 5304 4663
rect 5469 4657 5480 4663
rect 6456 4657 6467 4663
rect 3304 4637 3315 4643
rect 765 4577 792 4583
rect 2168 4577 2179 4583
rect 2328 4577 2339 4583
rect 3597 4577 3608 4583
rect 3661 4577 3672 4583
rect 4189 4577 4200 4583
rect 4253 4577 4264 4583
rect 5576 4577 5587 4583
rect 5720 4577 5731 4583
rect 6344 4577 6355 4583
rect 6445 4577 6472 4583
rect 7080 4577 7123 4583
rect 877 4557 920 4563
rect 1229 4557 1267 4563
rect 1741 4557 1752 4563
rect 1912 4557 1923 4563
rect 2940 4557 3011 4563
rect 2940 4554 2948 4557
rect 552 4537 568 4543
rect 861 4537 920 4543
rect 941 4523 947 4543
rect 1464 4537 1491 4543
rect 1944 4537 2035 4543
rect 2125 4537 2152 4543
rect 2189 4537 2200 4543
rect 904 4517 947 4523
rect 2253 4523 2259 4543
rect 2733 4537 2744 4543
rect 2984 4537 3027 4543
rect 3560 4537 3571 4543
rect 3624 4537 3635 4543
rect 4136 4537 4163 4543
rect 4200 4537 4227 4543
rect 4605 4537 4643 4543
rect 2072 4517 2099 4523
rect 2221 4517 2259 4523
rect 2424 4517 2451 4523
rect 2653 4517 2691 4523
rect 269 4483 275 4503
rect 269 4477 307 4483
rect 301 4457 307 4477
rect 360 4477 387 4483
rect 589 4483 595 4503
rect 1117 4497 1128 4503
rect 1352 4497 1364 4503
rect 1373 4497 1395 4503
rect 1356 4492 1364 4497
rect 2301 4497 2312 4503
rect 2685 4497 2691 4517
rect 3160 4517 3187 4523
rect 3240 4517 3251 4523
rect 4509 4517 4547 4523
rect 3021 4497 3059 4503
rect 3069 4497 3107 4503
rect 3124 4496 3128 4504
rect 3293 4497 3304 4503
rect 3357 4497 3368 4503
rect 3533 4497 3560 4503
rect 4008 4497 4035 4503
rect 4541 4497 4547 4517
rect 4605 4523 4611 4537
rect 4909 4537 4920 4543
rect 5016 4537 5075 4543
rect 5261 4543 5267 4563
rect 6013 4557 6056 4563
rect 5128 4537 5155 4543
rect 5213 4537 5267 4543
rect 5352 4537 5379 4543
rect 5677 4537 5688 4543
rect 5757 4537 5784 4543
rect 6221 4543 6227 4563
rect 6557 4557 6611 4563
rect 6717 4557 6728 4563
rect 6173 4537 6227 4543
rect 6381 4537 6408 4543
rect 6653 4537 6723 4543
rect 7053 4537 7112 4543
rect 7160 4537 7171 4543
rect 7485 4537 7496 4543
rect 7549 4537 7571 4543
rect 4584 4517 4611 4523
rect 4829 4517 4867 4523
rect 4861 4497 4867 4517
rect 5101 4517 5128 4523
rect 5421 4517 5475 4523
rect 5421 4497 5427 4517
rect 6552 4517 6595 4523
rect 7032 4517 7043 4523
rect 7565 4523 7571 4537
rect 7708 4543 7716 4548
rect 7688 4537 7716 4543
rect 7949 4537 7960 4543
rect 7565 4517 7592 4523
rect 7629 4517 7667 4523
rect 7016 4497 7027 4503
rect 7629 4497 7635 4517
rect 7800 4517 7827 4523
rect 589 4477 627 4483
rect 621 4457 627 4477
rect 696 4477 707 4483
rect 3276 4477 3315 4483
rect 3309 4457 3315 4477
rect 3368 4477 3395 4483
rect 4008 4477 4067 4483
rect 845 4377 856 4383
rect 1197 4377 1208 4383
rect 333 4337 360 4343
rect 717 4337 744 4343
rect 808 4337 835 4343
rect 3176 4337 3203 4343
rect 3533 4337 3544 4343
rect 3560 4337 3619 4343
rect 3832 4337 3875 4343
rect 6952 4337 6963 4343
rect 264 4317 291 4323
rect 909 4317 920 4323
rect 1005 4317 1016 4323
rect 1960 4317 2003 4323
rect 2045 4317 2067 4323
rect 2589 4317 2643 4323
rect 2973 4317 3000 4323
rect 4877 4317 4904 4323
rect 2157 4297 2184 4303
rect 2796 4303 2804 4304
rect 2472 4297 2499 4303
rect 2749 4297 2804 4303
rect 4168 4297 4195 4303
rect 4488 4297 4515 4303
rect 4957 4303 4963 4323
rect 5789 4317 5827 4323
rect 6013 4317 6067 4323
rect 4925 4297 4963 4303
rect 5160 4297 5187 4303
rect 5341 4297 5368 4303
rect 5480 4297 5491 4303
rect 5501 4297 5512 4303
rect 5613 4297 5640 4303
rect 5949 4297 5960 4303
rect 5997 4297 6040 4303
rect 6061 4303 6067 4317
rect 6061 4297 6099 4303
rect 6120 4297 6131 4303
rect 6429 4303 6435 4323
rect 6397 4297 6435 4303
rect 6637 4297 6664 4303
rect 6797 4303 6803 4323
rect 7421 4317 7475 4323
rect 6765 4297 6803 4303
rect 7021 4297 7032 4303
rect 7192 4297 7219 4303
rect 7304 4297 7315 4303
rect 7384 4297 7395 4303
rect 7549 4303 7555 4323
rect 7640 4317 7652 4323
rect 7644 4312 7652 4317
rect 7549 4297 7587 4303
rect 7597 4297 7624 4303
rect 7736 4297 7763 4303
rect 1224 4277 1251 4283
rect 1548 4277 1588 4283
rect 2328 4277 2339 4283
rect 2349 4277 2388 4283
rect 2669 4277 2680 4283
rect 2380 4272 2388 4277
rect 2712 4277 2723 4283
rect 2776 4277 2787 4283
rect 3293 4277 3304 4283
rect 3357 4277 3384 4283
rect 4600 4277 4627 4283
rect 4840 4277 4851 4283
rect 5032 4277 5076 4283
rect 5068 4272 5076 4277
rect 5244 4277 5284 4283
rect 6568 4277 6611 4283
rect 6680 4277 6691 4283
rect 6744 4277 6755 4283
rect 6909 4277 6936 4283
rect 7820 4277 7860 4283
rect 60 4268 68 4272
rect 1756 4263 1764 4266
rect 1756 4257 1768 4263
rect 1837 4257 1875 4263
rect 3229 4257 3276 4263
rect 3320 4257 3340 4263
rect 6157 4257 6168 4263
rect 6332 4263 6340 4272
rect 6312 4257 6340 4263
rect 1304 4237 1315 4243
rect 2200 4237 2211 4243
rect 4056 4237 4083 4243
rect 4280 4237 4291 4243
rect 4392 4237 4403 4243
rect 7064 4237 7107 4243
rect 8029 4237 8040 4243
rect 3368 4177 3379 4183
rect 3853 4177 3864 4183
rect 4920 4177 4931 4183
rect 8008 4177 8019 4183
rect 93 4157 147 4163
rect 1325 4157 1379 4163
rect 1885 4157 1923 4163
rect 2088 4157 2099 4163
rect 2616 4157 2644 4163
rect 2636 4148 2644 4157
rect 2904 4157 2915 4163
rect 1052 4143 1060 4148
rect 888 4137 915 4143
rect 1021 4137 1060 4143
rect 1869 4137 1896 4143
rect 2216 4137 2243 4143
rect 2333 4137 2360 4143
rect 3048 4137 3059 4143
rect 3661 4143 3667 4163
rect 6348 4157 6376 4163
rect 6348 4148 6356 4157
rect 7304 4157 7332 4163
rect 7324 4148 7332 4157
rect 7356 4157 7395 4163
rect 7356 4154 7364 4157
rect 3661 4137 3688 4143
rect 3864 4137 3891 4143
rect 4524 4143 4532 4148
rect 4493 4137 4532 4143
rect 4893 4137 4904 4143
rect 5100 4137 5144 4143
rect 5340 4143 5348 4148
rect 5340 4137 5352 4143
rect 5464 4137 5491 4143
rect 6157 4137 6195 4143
rect 520 4117 531 4123
rect 1720 4117 1731 4123
rect 2381 4117 2419 4123
rect 412 4103 420 4108
rect 392 4097 420 4103
rect 808 4097 819 4103
rect 1485 4097 1496 4103
rect 2413 4097 2419 4117
rect 2445 4117 2472 4123
rect 2717 4117 2744 4123
rect 2861 4117 2899 4123
rect 3085 4117 3123 4123
rect 3560 4117 3571 4123
rect 3645 4117 3688 4123
rect 3965 4117 4040 4123
rect 4125 4117 4163 4123
rect 4189 4117 4232 4123
rect 2708 4096 2712 4104
rect 3533 4097 3544 4103
rect 4008 4097 4067 4103
rect 4077 4097 4104 4103
rect 4157 4097 4163 4117
rect 4445 4117 4483 4123
rect 4269 4097 4296 4103
rect 4445 4097 4451 4117
rect 4556 4108 4564 4114
rect 4616 4117 4643 4123
rect 4813 4117 4851 4123
rect 4845 4097 4851 4117
rect 5016 4117 5043 4123
rect 5229 4117 5256 4123
rect 5437 4117 5448 4123
rect 5565 4117 5603 4123
rect 5629 4117 5656 4123
rect 5517 4097 5544 4103
rect 5597 4097 5603 4117
rect 5741 4117 5768 4123
rect 6061 4117 6072 4123
rect 6189 4123 6195 4137
rect 7469 4137 7507 4143
rect 6104 4117 6131 4123
rect 6189 4117 6200 4123
rect 6269 4117 6324 4123
rect 6316 4114 6324 4117
rect 6616 4117 6644 4123
rect 6636 4114 6644 4117
rect 6925 4117 6936 4123
rect 7053 4117 7139 4123
rect 5917 4097 5971 4103
rect 7053 4097 7059 4117
rect 7453 4117 7464 4123
rect 7608 4117 7619 4123
rect 7629 4117 7667 4123
rect 7528 4097 7571 4103
rect 7661 4097 7667 4117
rect 7736 4117 7748 4123
rect 7740 4114 7748 4117
rect 7832 4117 7859 4123
rect 765 4077 808 4083
rect 1096 4076 1098 4084
rect 1677 4077 1704 4083
rect 1677 4057 1683 4077
rect 3340 4083 3348 4088
rect 3340 4077 3352 4083
rect 3501 4077 3528 4083
rect 3852 4083 3860 4088
rect 3852 4077 3880 4083
rect 861 4037 872 4043
rect 984 4037 1011 4043
rect 3544 3937 3560 3943
rect 3784 3937 3795 3943
rect 3944 3937 3987 3943
rect 5336 3937 5347 3943
rect 6456 3937 6468 3943
rect 6460 3932 6468 3937
rect 125 3917 147 3923
rect 2605 3917 2616 3923
rect 477 3897 488 3903
rect 1757 3897 1784 3903
rect 1912 3897 1923 3903
rect 2300 3906 2308 3912
rect 2429 3897 2456 3903
rect 2568 3897 2579 3903
rect 2989 3897 3016 3903
rect 3100 3903 3108 3906
rect 3100 3897 3128 3903
rect 3245 3903 3251 3923
rect 3213 3897 3251 3903
rect 4056 3897 4067 3903
rect 4573 3903 4579 3923
rect 4541 3897 4579 3903
rect 4712 3897 4723 3903
rect 4733 3897 4760 3903
rect 5053 3903 5059 3923
rect 4872 3897 4899 3903
rect 4989 3897 5059 3903
rect 5132 3903 5140 3906
rect 5128 3897 5140 3903
rect 5224 3897 5251 3903
rect 5645 3903 5651 3923
rect 5613 3897 5651 3903
rect 5773 3897 5800 3903
rect 6109 3897 6136 3903
rect 6264 3897 6275 3903
rect 6365 3903 6371 3923
rect 6365 3897 6419 3903
rect 6653 3897 6680 3903
rect 6829 3903 6835 3923
rect 6829 3897 6867 3903
rect 7245 3903 7251 3923
rect 7608 3917 7635 3923
rect 7245 3897 7299 3903
rect 7565 3897 7592 3903
rect 7656 3897 7683 3903
rect 7773 3903 7779 3923
rect 7741 3897 7779 3903
rect 7917 3897 7944 3903
rect 861 3877 920 3883
rect 1085 3877 1123 3883
rect 440 3857 451 3863
rect 461 3857 515 3863
rect 717 3857 755 3863
rect 776 3857 792 3863
rect 877 3857 947 3863
rect 1117 3863 1123 3877
rect 1277 3877 1336 3883
rect 1544 3877 1571 3883
rect 1868 3877 1907 3883
rect 1917 3877 1971 3883
rect 1868 3872 1876 3877
rect 2125 3877 2136 3883
rect 3293 3877 3304 3883
rect 4040 3877 4051 3883
rect 4157 3877 4168 3883
rect 4237 3877 4275 3883
rect 4492 3877 4504 3883
rect 4568 3877 4579 3883
rect 6013 3877 6072 3883
rect 6120 3877 6163 3883
rect 6941 3877 6952 3883
rect 7608 3877 7619 3883
rect 1117 3857 1139 3863
rect 1272 3857 1283 3863
rect 2780 3863 2788 3872
rect 2760 3857 2788 3863
rect 4348 3866 4356 3872
rect 5420 3866 5428 3872
rect 7484 3868 7492 3872
rect 4316 3863 4324 3866
rect 5388 3863 5396 3866
rect 4285 3857 4324 3863
rect 5357 3857 5396 3863
rect 6056 3857 6083 3863
rect 6093 3857 6147 3863
rect 7996 3863 8004 3872
rect 7976 3857 8004 3863
rect 6557 3837 6568 3843
rect 1304 3777 1315 3783
rect 2845 3777 2856 3783
rect 237 3757 291 3763
rect 568 3757 579 3763
rect 776 3757 804 3763
rect 60 3748 68 3752
rect 396 3748 404 3752
rect 796 3748 804 3757
rect 568 3737 595 3743
rect 1485 3743 1491 3763
rect 1896 3757 1907 3763
rect 2184 3757 2195 3763
rect 3352 3757 3372 3763
rect 3608 3757 3619 3763
rect 3784 3757 3796 3763
rect 3788 3754 3796 3757
rect 4232 3757 4244 3763
rect 4236 3754 4244 3757
rect 4760 3757 4772 3763
rect 4764 3754 4772 3757
rect 4968 3757 4988 3763
rect 5421 3757 5460 3763
rect 5452 3754 5460 3757
rect 5100 3748 5108 3754
rect 5484 3748 5492 3754
rect 6317 3757 6328 3763
rect 6392 3757 6435 3763
rect 7005 3757 7076 3763
rect 7068 3754 7076 3757
rect 7100 3748 7108 3754
rect 1485 3737 1523 3743
rect 1661 3737 1672 3743
rect 1896 3737 1923 3743
rect 2157 3737 2211 3743
rect 2392 3737 2419 3743
rect 2520 3737 2563 3743
rect 3272 3737 3299 3743
rect 904 3717 947 3723
rect 1208 3717 1219 3723
rect 1404 3717 1416 3723
rect 1404 3712 1412 3717
rect 1725 3717 1752 3723
rect 1853 3717 1896 3723
rect 1928 3717 1939 3723
rect 2216 3717 2227 3723
rect 2429 3717 2467 3723
rect 1981 3697 1992 3703
rect 2461 3697 2467 3717
rect 2620 3717 2632 3723
rect 2620 3712 2628 3717
rect 2717 3717 2755 3723
rect 2792 3717 2808 3723
rect 2973 3717 3016 3723
rect 3117 3717 3128 3723
rect 3485 3723 3491 3743
rect 3581 3737 3592 3743
rect 3757 3737 3768 3743
rect 4412 3737 4424 3743
rect 5373 3737 5384 3743
rect 5628 3737 5640 3743
rect 5757 3737 5768 3743
rect 6253 3737 6323 3743
rect 6456 3737 6467 3743
rect 6957 3737 6995 3743
rect 7384 3737 7427 3743
rect 7501 3737 7523 3743
rect 3448 3717 3491 3723
rect 3677 3717 3715 3723
rect 2845 3697 2856 3703
rect 3496 3697 3507 3703
rect 3709 3697 3715 3717
rect 3880 3717 3907 3723
rect 4125 3717 4163 3723
rect 4157 3697 4163 3717
rect 4328 3717 4355 3723
rect 4589 3717 4627 3723
rect 4653 3717 4664 3723
rect 4541 3697 4552 3703
rect 4621 3697 4627 3717
rect 4696 3717 4707 3723
rect 4856 3717 4883 3723
rect 5016 3717 5076 3723
rect 5068 3714 5076 3717
rect 5293 3717 5331 3723
rect 4733 3697 4744 3703
rect 5325 3697 5331 3717
rect 5720 3717 5731 3723
rect 5853 3717 5880 3723
rect 6029 3717 6099 3723
rect 6029 3697 6035 3717
rect 6120 3717 6163 3723
rect 6541 3717 6547 3732
rect 7693 3717 7731 3723
rect 6056 3697 6083 3703
rect 7309 3697 7363 3703
rect 7565 3697 7619 3703
rect 7693 3697 7699 3717
rect 7932 3708 7940 3714
rect 152 3537 163 3543
rect 344 3537 355 3543
rect 1677 3537 1704 3543
rect 1736 3537 1763 3543
rect 3080 3537 3091 3543
rect 3352 3537 3363 3543
rect 6838 3536 6840 3544
rect 7576 3537 7587 3543
rect 408 3497 419 3503
rect 621 3497 648 3503
rect 1133 3503 1139 3523
rect 1720 3517 1731 3523
rect 1837 3517 1908 3523
rect 1900 3512 1908 3517
rect 4125 3517 4163 3523
rect 1133 3497 1187 3503
rect 1224 3497 1235 3503
rect 1453 3497 1480 3503
rect 1932 3506 1940 3512
rect 2140 3503 2148 3508
rect 2140 3497 2152 3503
rect 2349 3497 2360 3503
rect 2621 3497 2659 3503
rect 472 3477 515 3483
rect 765 3477 776 3483
rect 856 3477 900 3483
rect 892 3472 900 3477
rect 2200 3477 2243 3483
rect 2296 3477 2323 3483
rect 2653 3483 2659 3497
rect 3192 3497 3203 3503
rect 3928 3497 3955 3503
rect 4168 3497 4179 3503
rect 4780 3506 4788 3512
rect 4989 3503 4995 3523
rect 4957 3497 4995 3503
rect 5021 3497 5064 3503
rect 5464 3497 5475 3503
rect 5853 3497 5880 3503
rect 6029 3503 6035 3523
rect 6029 3497 6115 3503
rect 6392 3497 6403 3503
rect 6541 3497 6568 3503
rect 6621 3503 6627 3523
rect 6876 3517 6915 3523
rect 6876 3512 6884 3517
rect 6589 3497 6627 3503
rect 6765 3497 6792 3503
rect 7005 3503 7011 3523
rect 6968 3497 6979 3503
rect 7005 3497 7043 3503
rect 7053 3497 7112 3503
rect 7224 3497 7251 3503
rect 7304 3497 7315 3503
rect 7501 3503 7507 3523
rect 7469 3497 7507 3503
rect 7672 3497 7699 3503
rect 7917 3497 7944 3503
rect 2568 3477 2595 3483
rect 2653 3477 2675 3483
rect 3816 3477 3827 3483
rect 4205 3477 4216 3483
rect 4461 3477 4483 3483
rect 5688 3477 5720 3483
rect 6269 3477 6296 3483
rect 1592 3457 1603 3463
rect 2173 3457 2227 3463
rect 2541 3457 2552 3463
rect 4380 3466 4388 3472
rect 4412 3463 4420 3466
rect 4412 3457 4451 3463
rect 829 3437 856 3443
rect 2616 3377 2627 3383
rect 4264 3377 4275 3383
rect 5944 3377 5955 3383
rect 7000 3377 7011 3383
rect 669 3357 680 3363
rect 1688 3357 1700 3363
rect 1692 3354 1700 3357
rect 3448 3357 3460 3363
rect 4413 3357 4452 3363
rect 3452 3354 3460 3357
rect 4444 3354 4452 3357
rect 4476 3348 4484 3354
rect 7352 3357 7364 3363
rect 7356 3354 7364 3357
rect 40 3337 51 3343
rect 120 3337 131 3343
rect 653 3337 707 3343
rect 1037 3337 1048 3343
rect 1868 3337 1923 3343
rect 2536 3337 2563 3343
rect 2744 3337 2755 3343
rect 2861 3337 2883 3343
rect 557 3317 568 3323
rect 1176 3317 1188 3323
rect 1180 3312 1188 3317
rect 1949 3317 1992 3323
rect 2157 3317 2184 3323
rect 2333 3317 2371 3323
rect 285 3283 291 3303
rect 1480 3297 1507 3303
rect 1613 3297 1624 3303
rect 2333 3297 2339 3317
rect 2392 3317 2419 3323
rect 2440 3317 2483 3323
rect 2600 3317 2616 3323
rect 2861 3323 2867 3337
rect 4076 3343 4084 3348
rect 4076 3337 4147 3343
rect 4365 3337 4403 3343
rect 4908 3343 4916 3348
rect 4888 3337 4916 3343
rect 5224 3337 5235 3343
rect 5624 3337 5635 3343
rect 5917 3337 5944 3343
rect 6220 3337 6275 3343
rect 6365 3337 6403 3343
rect 6540 3343 6548 3348
rect 6520 3337 6548 3343
rect 7037 3337 7096 3343
rect 7597 3337 7608 3343
rect 2845 3317 2867 3323
rect 3053 3317 3091 3323
rect 2909 3297 2931 3303
rect 3085 3297 3091 3317
rect 3341 3317 3379 3323
rect 3405 3317 3432 3323
rect 3373 3297 3379 3317
rect 3560 3317 3571 3323
rect 3709 3317 3736 3323
rect 3965 3317 3992 3323
rect 4157 3317 4195 3323
rect 4189 3297 4195 3317
rect 4712 3317 4723 3323
rect 4733 3317 4744 3323
rect 4813 3317 4867 3323
rect 4669 3297 4707 3303
rect 4813 3297 4819 3317
rect 5000 3317 5027 3323
rect 5197 3317 5224 3323
rect 5324 3308 5332 3314
rect 5517 3317 5555 3323
rect 5292 3303 5300 3308
rect 5261 3297 5300 3303
rect 5549 3297 5555 3317
rect 5709 3317 5747 3323
rect 5661 3297 5688 3303
rect 5741 3297 5747 3317
rect 5784 3317 5827 3323
rect 5853 3317 5907 3323
rect 5853 3297 5859 3317
rect 6136 3317 6163 3323
rect 6301 3317 6312 3323
rect 6445 3317 6499 3323
rect 5880 3297 5891 3303
rect 6044 3303 6052 3308
rect 6008 3297 6052 3303
rect 6445 3297 6451 3317
rect 6632 3317 6659 3323
rect 6856 3317 6867 3323
rect 7181 3317 7219 3323
rect 7048 3297 7096 3303
rect 7213 3297 7219 3317
rect 7448 3317 7475 3323
rect 7597 3317 7651 3323
rect 7597 3297 7603 3317
rect 7836 3308 7844 3314
rect 7896 3317 7907 3323
rect 7933 3317 7987 3323
rect 7933 3297 7939 3317
rect 285 3277 323 3283
rect 317 3257 323 3277
rect 797 3277 836 3283
rect 797 3257 803 3277
rect 1208 3277 1219 3283
rect 2620 3283 2628 3288
rect 2616 3277 2628 3283
rect 2780 3283 2788 3288
rect 2780 3277 2792 3283
rect 6088 3276 6090 3284
rect 6968 3277 6979 3283
rect 445 3177 456 3183
rect 3144 3177 3155 3183
rect 3613 3177 3624 3183
rect 6584 3177 6595 3183
rect 7053 3177 7080 3183
rect 1517 3143 1523 3163
rect 1752 3157 1763 3163
rect 1517 3137 1555 3143
rect 61 3103 67 3123
rect 685 3117 696 3123
rect 1132 3117 1144 3123
rect 1132 3112 1140 3117
rect 1288 3117 1299 3123
rect 1405 3117 1416 3123
rect 1549 3117 1555 3137
rect 5528 3136 5530 3144
rect 6344 3137 6371 3143
rect 7896 3137 7907 3143
rect 2120 3117 2131 3123
rect 2664 3117 2675 3123
rect 2813 3117 2824 3123
rect 61 3097 72 3103
rect 269 3097 280 3103
rect 1021 3097 1032 3103
rect 1160 3097 1171 3103
rect 2440 3097 2451 3103
rect 3325 3097 3336 3103
rect 3404 3106 3412 3112
rect 3517 3103 3523 3123
rect 3677 3117 3716 3123
rect 3708 3112 3716 3117
rect 3485 3097 3523 3103
rect 3740 3106 3748 3112
rect 3965 3103 3971 3123
rect 3933 3097 3971 3103
rect 3997 3097 4040 3103
rect 4285 3103 4291 3123
rect 4696 3117 4707 3123
rect 5176 3117 5187 3123
rect 5261 3108 5267 3123
rect 5997 3117 6040 3123
rect 6253 3117 6307 3123
rect 6968 3117 6979 3123
rect 4285 3097 4339 3103
rect 4781 3097 4824 3103
rect 552 3077 563 3083
rect 920 3077 964 3083
rect 1197 3077 1208 3083
rect 2077 3077 2088 3083
rect 2157 3077 2168 3083
rect 2424 3077 2435 3083
rect 2840 3077 2867 3083
rect 3436 3077 3475 3083
rect 3436 3072 3444 3077
rect 4173 3077 4227 3083
rect 4376 3077 4388 3083
rect 4605 3077 4627 3083
rect 4813 3083 4819 3097
rect 4957 3097 4984 3103
rect 5228 3097 5256 3103
rect 5228 3092 5236 3097
rect 5592 3097 5603 3103
rect 5784 3097 5811 3103
rect 6024 3097 6067 3103
rect 6493 3097 6531 3103
rect 4813 3077 4851 3083
rect 5293 3077 5304 3083
rect 6221 3077 6259 3083
rect 6408 3077 6435 3083
rect 7453 3097 7480 3103
rect 7640 3097 7667 3103
rect 7741 3097 7779 3103
rect 7944 3097 7955 3103
rect 6712 3077 6723 3083
rect 6861 3077 6872 3083
rect 7005 3077 7016 3083
rect 7160 3077 7188 3083
rect 7180 3072 7188 3077
rect 7356 3077 7396 3083
rect 1788 3066 1796 3072
rect 1997 3057 2051 3063
rect 3592 3057 3603 3063
rect 4524 3063 4532 3072
rect 4504 3057 4532 3063
rect 4556 3063 4564 3066
rect 4556 3057 4595 3063
rect 5484 3063 5492 3066
rect 5453 3057 5492 3063
rect 6500 3057 6520 3063
rect 2184 3037 2195 3043
rect 5480 3037 5491 3043
rect 5896 3037 5907 3043
rect 6136 3037 6147 3043
rect 6296 3037 6307 3043
rect 6797 3037 6808 3043
rect 2984 2977 2995 2983
rect 4109 2977 4120 2983
rect 4744 2977 4755 2983
rect 5800 2977 5811 2983
rect 5944 2977 5955 2983
rect 93 2957 120 2963
rect 221 2957 275 2963
rect 652 2957 664 2963
rect 652 2954 660 2957
rect 733 2957 771 2963
rect 845 2957 867 2963
rect 360 2937 371 2943
rect 845 2943 851 2957
rect 1096 2957 1124 2963
rect 1116 2948 1124 2957
rect 1176 2957 1187 2963
rect 1277 2957 1315 2963
rect 1480 2957 1508 2963
rect 1500 2948 1508 2957
rect 1853 2957 1864 2963
rect 2093 2957 2115 2963
rect 813 2937 851 2943
rect 2093 2943 2099 2957
rect 2700 2957 2728 2963
rect 2700 2954 2708 2957
rect 5357 2957 5368 2963
rect 6728 2957 6740 2963
rect 6732 2954 6740 2957
rect 3164 2948 3172 2952
rect 2061 2937 2099 2943
rect 2248 2937 2259 2943
rect 2749 2937 2771 2943
rect 2941 2937 2968 2943
rect 3132 2943 3140 2948
rect 3101 2937 3140 2943
rect 3464 2937 3491 2943
rect 3581 2937 3592 2943
rect 3624 2937 3636 2943
rect 3944 2937 3960 2943
rect 3976 2937 3987 2943
rect 4056 2937 4083 2943
rect 4456 2937 4484 2943
rect 4652 2943 4660 2948
rect 4652 2937 4680 2943
rect 4845 2937 4872 2943
rect 7080 2937 7124 2943
rect 7564 2937 7576 2943
rect 45 2917 67 2923
rect 141 2917 163 2923
rect 317 2917 344 2923
rect 909 2917 920 2923
rect 1805 2917 1880 2923
rect 1980 2923 1988 2928
rect 1928 2917 1988 2923
rect 2589 2917 2616 2923
rect 2861 2917 2899 2923
rect 1880 2897 1891 2903
rect 2216 2897 2227 2903
rect 2488 2897 2499 2903
rect 2813 2897 2824 2903
rect 2893 2897 2899 2917
rect 3021 2917 3064 2923
rect 3517 2917 3528 2923
rect 3693 2917 3720 2923
rect 4013 2917 4056 2923
rect 4172 2908 4180 2914
rect 4541 2917 4568 2923
rect 4796 2923 4804 2928
rect 4796 2917 4808 2923
rect 5084 2923 5092 2928
rect 5084 2917 5123 2923
rect 3064 2897 3075 2903
rect 3085 2897 3112 2903
rect 3869 2897 3923 2903
rect 4140 2903 4148 2908
rect 4109 2897 4148 2903
rect 4381 2897 4435 2903
rect 4445 2897 4456 2903
rect 4813 2897 4819 2912
rect 5117 2908 5123 2917
rect 5224 2917 5251 2923
rect 5436 2923 5444 2928
rect 5436 2917 5464 2923
rect 5485 2917 5523 2923
rect 4909 2897 4936 2903
rect 5517 2897 5523 2917
rect 5740 2908 5748 2914
rect 5916 2923 5924 2928
rect 5916 2917 5928 2923
rect 5965 2917 6019 2923
rect 6189 2917 6200 2923
rect 6221 2917 6275 2923
rect 6269 2897 6275 2917
rect 6424 2917 6451 2923
rect 6685 2917 6712 2923
rect 6824 2917 6851 2923
rect 7016 2917 7027 2923
rect 7037 2917 7064 2923
rect 7420 2908 7428 2914
rect 7693 2917 7731 2923
rect 6285 2897 6312 2903
rect 6621 2897 6659 2903
rect 7292 2903 7300 2908
rect 7292 2897 7315 2903
rect 7725 2897 7731 2917
rect 7896 2917 7923 2923
rect 1565 2877 1576 2883
rect 2284 2883 2292 2888
rect 2284 2877 2323 2883
rect 2317 2857 2323 2877
rect 6312 2877 6339 2883
rect 7800 2877 7811 2883
rect 5384 2857 5395 2863
rect 5000 2837 5043 2843
rect 3064 2777 3075 2783
rect 4424 2777 4435 2783
rect 7832 2777 7843 2783
rect 2408 2736 2410 2744
rect 3400 2737 3411 2743
rect 6712 2736 6714 2744
rect 2205 2717 2243 2723
rect 716 2706 724 2712
rect 856 2697 867 2703
rect 2621 2703 2627 2723
rect 2589 2697 2627 2703
rect 2989 2703 2995 2723
rect 3512 2717 3539 2723
rect 2925 2697 2995 2703
rect 3469 2697 3512 2703
rect 3693 2703 3699 2723
rect 3768 2717 3780 2723
rect 3772 2712 3780 2717
rect 3661 2697 3699 2703
rect 3725 2697 3752 2703
rect 3864 2697 3891 2703
rect 3992 2697 4003 2703
rect 4232 2697 4259 2703
rect 4685 2703 4691 2723
rect 4653 2697 4691 2703
rect 4717 2697 4744 2703
rect 4813 2697 4824 2703
rect 4893 2703 4899 2723
rect 4861 2697 4899 2703
rect 4925 2697 4936 2703
rect 5004 2703 5012 2706
rect 4968 2697 5012 2703
rect 5096 2697 5123 2703
rect 5469 2703 5475 2723
rect 5437 2697 5475 2703
rect 5501 2697 5544 2703
rect 5581 2703 5587 2723
rect 5581 2697 5635 2703
rect 5725 2697 5768 2703
rect 6349 2703 6355 2723
rect 6317 2697 6355 2703
rect 6381 2697 6392 2703
rect 6461 2703 6467 2723
rect 6461 2697 6515 2703
rect 6668 2703 6676 2706
rect 6621 2697 6676 2703
rect 6989 2697 7016 2703
rect 7197 2703 7203 2723
rect 7224 2717 7235 2723
rect 7405 2717 7416 2723
rect 7444 2716 7448 2724
rect 7197 2697 7251 2703
rect 7720 2697 7747 2703
rect 7928 2697 7955 2703
rect 280 2677 307 2683
rect 568 2677 580 2683
rect 893 2677 920 2683
rect 1005 2677 1016 2683
rect 1085 2677 1112 2683
rect 3160 2677 3188 2683
rect 3180 2672 3188 2677
rect 3485 2677 3496 2683
rect 3613 2677 3624 2683
rect 4109 2677 4120 2683
rect 4344 2677 4371 2683
rect 4680 2677 4691 2683
rect 4733 2677 4760 2683
rect 4941 2677 4984 2683
rect 5464 2677 5475 2683
rect 5741 2677 5811 2683
rect 5832 2677 5843 2683
rect 5928 2677 5939 2683
rect 5960 2677 6003 2683
rect 7100 2677 7128 2683
rect 7100 2672 7108 2677
rect 7368 2677 7379 2683
rect 7533 2677 7544 2683
rect 60 2663 68 2672
rect 60 2657 88 2663
rect 716 2663 724 2672
rect 1244 2666 1252 2672
rect 2396 2668 2404 2672
rect 696 2657 724 2663
rect 1421 2657 1475 2663
rect 2732 2663 2740 2672
rect 2732 2657 2760 2663
rect 4460 2666 4468 2672
rect 5244 2668 5252 2672
rect 6700 2666 6708 2672
rect 7660 2663 7668 2672
rect 7660 2657 7688 2663
rect 360 2637 371 2643
rect 1208 2637 1219 2643
rect 6461 2637 6472 2643
rect 3656 2577 3667 2583
rect 4296 2577 4307 2583
rect 6104 2577 6115 2583
rect 301 2557 323 2563
rect 525 2557 563 2563
rect 301 2543 307 2557
rect 1293 2557 1304 2563
rect 1661 2557 1715 2563
rect 1960 2557 2028 2563
rect 2952 2557 2980 2563
rect 2972 2548 2980 2557
rect 3004 2557 3075 2563
rect 3004 2554 3012 2557
rect 5885 2557 5896 2563
rect 4540 2548 4548 2554
rect 269 2537 307 2543
rect 349 2537 360 2543
rect 1277 2537 1304 2543
rect 2461 2537 2483 2543
rect 2824 2537 2836 2543
rect 3085 2537 3107 2543
rect 3356 2543 3364 2548
rect 3356 2537 3384 2543
rect 3949 2537 3987 2543
rect 4760 2537 4771 2543
rect 6312 2537 6323 2543
rect 6440 2537 6451 2543
rect 7116 2543 7124 2548
rect 7080 2537 7124 2543
rect 7421 2537 7475 2543
rect 7741 2537 7779 2543
rect 7880 2537 7923 2543
rect 157 2517 168 2523
rect 472 2517 483 2523
rect 733 2517 744 2523
rect 1628 2517 1640 2523
rect 1628 2512 1636 2517
rect 1949 2517 2008 2523
rect 3112 2517 3123 2523
rect 3245 2517 3272 2523
rect 3469 2517 3507 2523
rect 941 2497 968 2503
rect 989 2483 995 2503
rect 1373 2497 1395 2503
rect 1501 2497 1523 2503
rect 2061 2497 2072 2503
rect 2316 2497 2328 2503
rect 2316 2492 2324 2497
rect 2525 2497 2579 2503
rect 2717 2497 2755 2503
rect 3356 2503 3364 2508
rect 3356 2497 3395 2503
rect 3501 2497 3507 2517
rect 3757 2517 3768 2523
rect 3805 2517 3843 2523
rect 3837 2497 3843 2517
rect 4008 2517 4083 2523
rect 4189 2517 4227 2523
rect 4221 2497 4227 2517
rect 4392 2517 4419 2523
rect 4733 2517 4771 2523
rect 4765 2497 4771 2517
rect 4861 2517 4899 2523
rect 4893 2497 4899 2517
rect 5144 2517 5171 2523
rect 5501 2517 5528 2523
rect 5677 2517 5715 2523
rect 5677 2497 5683 2517
rect 5736 2517 5763 2523
rect 5821 2517 5832 2523
rect 5965 2517 5992 2523
rect 6333 2517 6371 2523
rect 6365 2497 6371 2517
rect 6888 2517 6899 2523
rect 6925 2517 6936 2523
rect 6477 2497 6488 2503
rect 6893 2497 6899 2517
rect 6973 2517 7011 2523
rect 7005 2497 7011 2517
rect 7208 2517 7235 2523
rect 7405 2517 7416 2523
rect 7528 2517 7560 2523
rect 7688 2517 7715 2523
rect 7320 2497 7331 2503
rect 7341 2497 7379 2503
rect 925 2477 995 2483
rect 925 2457 931 2477
rect 2072 2477 2099 2483
rect 2205 2477 2244 2483
rect 2205 2457 2211 2477
rect 2333 2477 2372 2483
rect 2333 2457 2339 2477
rect 6152 2476 6154 2484
rect 3960 2377 4003 2383
rect 7517 2377 7528 2383
rect 1293 2343 1299 2363
rect 4264 2357 4275 2363
rect 1261 2337 1299 2343
rect 1000 2317 1027 2323
rect 1261 2317 1267 2337
rect 1660 2317 1683 2323
rect 1725 2317 1747 2323
rect 1660 2312 1668 2317
rect 1965 2317 1976 2323
rect 2317 2317 2339 2323
rect 45 2297 67 2303
rect 109 2297 120 2303
rect 61 2283 67 2297
rect 541 2297 552 2303
rect 1453 2297 1464 2303
rect 2076 2303 2084 2308
rect 2076 2297 2104 2303
rect 2301 2297 2312 2303
rect 2333 2303 2339 2317
rect 3821 2317 3875 2323
rect 4376 2317 4403 2323
rect 4888 2317 4916 2323
rect 4908 2312 4916 2317
rect 2333 2297 2371 2303
rect 2845 2297 2872 2303
rect 3080 2297 3091 2303
rect 3309 2297 3320 2303
rect 3533 2297 3544 2303
rect 4088 2297 4115 2303
rect 4344 2297 4387 2303
rect 61 2277 83 2283
rect 1096 2277 1123 2283
rect 1149 2277 1187 2283
rect 764 2268 772 2272
rect 189 2257 227 2263
rect 1149 2257 1155 2277
rect 1896 2277 1907 2283
rect 2173 2277 2200 2283
rect 3000 2277 3011 2283
rect 3160 2277 3187 2283
rect 3549 2277 3560 2283
rect 4381 2277 4387 2297
rect 4424 2297 4451 2303
rect 4813 2297 4840 2303
rect 5000 2297 5027 2303
rect 5144 2297 5155 2303
rect 5560 2297 5571 2303
rect 5677 2303 5683 2323
rect 5677 2297 5731 2303
rect 5916 2306 5924 2312
rect 6280 2297 6291 2303
rect 6328 2297 6371 2303
rect 6685 2303 6691 2323
rect 6536 2297 6547 2303
rect 6653 2297 6691 2303
rect 6936 2297 6979 2303
rect 7117 2297 7144 2303
rect 7293 2303 7299 2323
rect 7421 2303 7427 2323
rect 7293 2297 7347 2303
rect 7389 2297 7427 2303
rect 7453 2297 7464 2303
rect 7597 2303 7603 2323
rect 7565 2297 7603 2303
rect 7832 2297 7859 2303
rect 4536 2277 4564 2283
rect 4556 2272 4564 2277
rect 5084 2277 5112 2283
rect 5432 2277 5443 2283
rect 5480 2277 5491 2283
rect 5768 2277 5780 2283
rect 6461 2277 6531 2283
rect 6925 2277 6952 2283
rect 7016 2277 7060 2283
rect 7469 2277 7480 2283
rect 7736 2277 7748 2283
rect 7740 2272 7748 2277
rect 1357 2257 1411 2263
rect 1628 2263 1636 2272
rect 1608 2257 1636 2263
rect 2556 2266 2564 2272
rect 3612 2263 3620 2272
rect 6156 2268 6164 2272
rect 7196 2268 7204 2272
rect 1880 2257 1891 2263
rect 3612 2257 3640 2263
rect 3933 2257 3960 2263
rect 6317 2257 6328 2263
rect 4840 2237 4851 2243
rect 205 2177 216 2183
rect 2989 2177 3000 2183
rect 4360 2177 4371 2183
rect 412 2157 435 2163
rect 445 2157 499 2163
rect 412 2154 420 2157
rect 797 2157 851 2163
rect 1469 2157 1491 2163
rect 1164 2148 1172 2152
rect 1260 2148 1268 2152
rect 472 2137 515 2143
rect 525 2137 552 2143
rect 856 2137 867 2143
rect 1469 2143 1475 2157
rect 4205 2157 4252 2163
rect 5180 2148 5188 2154
rect 1437 2137 1475 2143
rect 1756 2143 1764 2148
rect 1624 2137 1651 2143
rect 1725 2137 1764 2143
rect 2108 2143 2116 2148
rect 2077 2137 2116 2143
rect 2392 2137 2403 2143
rect 3432 2137 3459 2143
rect 3613 2137 3651 2143
rect 4189 2137 4200 2143
rect 4877 2137 4915 2143
rect 6205 2137 6216 2143
rect 6237 2143 6243 2163
rect 6748 2157 6776 2163
rect 6412 2148 6420 2152
rect 6748 2148 6756 2157
rect 7308 2148 7316 2152
rect 6232 2137 6243 2143
rect 6621 2137 6648 2143
rect 6968 2137 6979 2143
rect 7037 2137 7107 2143
rect 301 2117 312 2123
rect 1085 2117 1112 2123
rect 2477 2117 2515 2123
rect 1196 2103 1204 2108
rect 1196 2097 1208 2103
rect 2509 2097 2515 2117
rect 2653 2117 2680 2123
rect 2829 2117 2867 2123
rect 2829 2097 2835 2117
rect 2888 2117 2915 2123
rect 3757 2117 3784 2123
rect 4589 2117 4627 2123
rect 3133 2097 3171 2103
rect 3533 2097 3571 2103
rect 3933 2097 3987 2103
rect 3997 2097 4008 2103
rect 4621 2097 4627 2117
rect 4861 2117 4872 2123
rect 5373 2117 5411 2123
rect 5405 2097 5411 2117
rect 5549 2117 5576 2123
rect 5725 2117 5779 2123
rect 5725 2097 5731 2117
rect 5960 2117 5987 2123
rect 6013 2117 6099 2123
rect 6013 2097 6019 2117
rect 6205 2117 6216 2123
rect 6296 2117 6307 2123
rect 6941 2117 6979 2123
rect 6685 2097 6696 2103
rect 6973 2097 6979 2117
rect 7037 2123 7043 2137
rect 7016 2117 7043 2123
rect 7229 2117 7284 2123
rect 7276 2114 7284 2117
rect 7533 2117 7544 2123
rect 7581 2117 7619 2123
rect 7645 2117 7656 2123
rect 7613 2097 7619 2117
rect 7688 2117 7700 2123
rect 7692 2114 7700 2117
rect 7784 2117 7811 2123
rect 3309 2077 3352 2083
rect 4092 2077 4131 2083
rect 4125 2057 4131 2077
rect 4280 2077 4323 2083
rect 205 2037 216 2043
rect 1704 2037 1715 2043
rect 2598 1936 2600 1944
rect 3384 1937 3395 1943
rect 3981 1943 3987 1963
rect 7848 1957 7859 1963
rect 3948 1937 3987 1943
rect 200 1897 227 1903
rect 365 1897 376 1903
rect 600 1897 611 1903
rect 840 1897 851 1903
rect 1160 1897 1171 1903
rect 1256 1897 1267 1903
rect 2296 1897 2323 1903
rect 2941 1903 2947 1923
rect 3544 1917 3555 1923
rect 3645 1917 3656 1923
rect 2909 1897 2947 1903
rect 3213 1897 3251 1903
rect 3581 1897 3603 1903
rect 572 1877 600 1883
rect 572 1872 580 1877
rect 1693 1877 1731 1883
rect 653 1857 691 1863
rect 876 1863 884 1872
rect 856 1857 884 1863
rect 1309 1857 1347 1863
rect 1725 1863 1731 1877
rect 2349 1877 2392 1883
rect 2824 1877 2835 1883
rect 3149 1877 3160 1883
rect 3581 1877 3587 1897
rect 3832 1897 3843 1903
rect 4040 1897 4067 1903
rect 4525 1897 4552 1903
rect 4717 1903 4723 1923
rect 4685 1897 4723 1903
rect 5245 1903 5251 1923
rect 5213 1897 5251 1903
rect 5469 1897 5491 1903
rect 5581 1897 5624 1903
rect 4429 1877 4440 1883
rect 4636 1877 4664 1883
rect 4636 1872 4644 1877
rect 4792 1877 4819 1883
rect 5293 1877 5304 1883
rect 5357 1877 5384 1883
rect 5469 1883 5475 1897
rect 6045 1903 6051 1923
rect 6045 1897 6115 1903
rect 6248 1897 6275 1903
rect 6429 1897 6440 1903
rect 6712 1897 6723 1903
rect 6973 1903 6979 1923
rect 7048 1917 7092 1923
rect 7084 1912 7092 1917
rect 6941 1897 6979 1903
rect 7176 1897 7203 1903
rect 7352 1897 7379 1903
rect 7512 1897 7523 1903
rect 7709 1903 7715 1923
rect 7677 1897 7715 1903
rect 7960 1897 7971 1903
rect 5448 1877 5475 1883
rect 5517 1877 5528 1883
rect 5565 1877 5635 1883
rect 6125 1877 6164 1883
rect 6156 1872 6164 1877
rect 6540 1877 6595 1883
rect 7325 1877 7352 1883
rect 1725 1857 1747 1863
rect 1964 1863 1972 1872
rect 5772 1868 5780 1872
rect 1944 1857 1972 1863
rect 2636 1863 2644 1866
rect 2040 1857 2067 1863
rect 2636 1857 2675 1863
rect 3277 1857 3324 1863
rect 3517 1857 3564 1863
rect 4093 1857 4140 1863
rect 6396 1863 6404 1872
rect 6396 1857 6424 1863
rect 2072 1777 2083 1783
rect 2344 1777 2355 1783
rect 4248 1777 4259 1783
rect 5805 1777 5816 1783
rect 61 1757 83 1763
rect 61 1743 67 1757
rect 29 1737 67 1743
rect 669 1757 723 1763
rect 1373 1757 1384 1763
rect 1672 1757 1683 1763
rect 1992 1757 2008 1763
rect 3101 1757 3140 1763
rect 3132 1754 3140 1757
rect 4536 1757 4548 1763
rect 4540 1754 4548 1757
rect 5624 1757 5635 1763
rect 5980 1748 5988 1754
rect 7944 1757 7972 1763
rect 6876 1748 6884 1752
rect 7964 1748 7972 1757
rect 1672 1737 1699 1743
rect 2652 1743 2660 1748
rect 2584 1737 2611 1743
rect 2621 1737 2660 1743
rect 2904 1737 2931 1743
rect 3064 1737 3091 1743
rect 4397 1737 4435 1743
rect 4765 1737 4787 1743
rect 5048 1737 5107 1743
rect 5292 1743 5300 1748
rect 5261 1737 5300 1743
rect 6216 1737 6227 1743
rect 6360 1737 6403 1743
rect 6605 1737 6616 1743
rect 7788 1737 7828 1743
rect 765 1717 776 1723
rect 1245 1717 1272 1723
rect 2184 1717 2195 1723
rect 2493 1717 2531 1723
rect 168 1677 200 1683
rect 445 1683 451 1703
rect 1453 1697 1475 1703
rect 1581 1697 1603 1703
rect 1965 1697 1976 1703
rect 2408 1697 2419 1703
rect 2525 1697 2531 1717
rect 2744 1717 2771 1723
rect 3224 1717 3251 1723
rect 3516 1717 3528 1723
rect 3516 1712 3524 1717
rect 3848 1717 3875 1723
rect 4332 1717 4344 1723
rect 4332 1712 4340 1717
rect 4632 1717 4659 1723
rect 5197 1717 5251 1723
rect 2957 1697 2984 1703
rect 4029 1697 4040 1703
rect 4157 1697 4168 1703
rect 5000 1697 5011 1703
rect 5048 1697 5123 1703
rect 5197 1697 5203 1717
rect 5384 1717 5411 1723
rect 5517 1717 5528 1723
rect 5741 1717 5752 1723
rect 5816 1717 5859 1723
rect 6189 1717 6227 1723
rect 5292 1703 5300 1708
rect 5272 1697 5300 1703
rect 5805 1697 5816 1703
rect 6221 1697 6227 1717
rect 6461 1717 6499 1723
rect 6493 1697 6499 1717
rect 7213 1717 7240 1723
rect 7352 1717 7363 1723
rect 7389 1717 7427 1723
rect 6844 1703 6852 1708
rect 6840 1697 6852 1703
rect 7389 1697 7395 1717
rect 7528 1717 7555 1723
rect 7644 1708 7652 1714
rect 7704 1717 7731 1723
rect 7928 1717 7939 1723
rect 7612 1703 7620 1708
rect 7581 1697 7620 1703
rect 445 1677 456 1683
rect 557 1677 627 1683
rect 557 1657 563 1677
rect 909 1677 995 1683
rect 1181 1677 1220 1683
rect 1181 1657 1187 1677
rect 1544 1677 1571 1683
rect 4008 1677 4067 1683
rect 4232 1677 4259 1683
rect 3016 1577 3027 1583
rect 1304 1536 1306 1544
rect 3917 1543 3923 1563
rect 3884 1537 3923 1543
rect 4012 1537 4024 1543
rect 4012 1532 4020 1537
rect 4120 1537 4132 1543
rect 4124 1532 4132 1537
rect 232 1497 243 1503
rect 797 1497 808 1503
rect 1352 1497 1379 1503
rect 1757 1503 1763 1523
rect 1832 1517 1843 1523
rect 2440 1517 2467 1523
rect 2541 1517 2552 1523
rect 1757 1497 1811 1503
rect 1821 1497 1832 1503
rect 1181 1477 1219 1483
rect 1229 1477 1268 1483
rect 1260 1472 1268 1477
rect 1485 1477 1524 1483
rect 1516 1472 1524 1477
rect 1821 1477 1827 1497
rect 1869 1497 1896 1503
rect 2461 1497 2499 1503
rect 2013 1477 2067 1483
rect 2264 1477 2291 1483
rect 2360 1477 2419 1483
rect 2429 1477 2440 1483
rect 2493 1477 2499 1497
rect 2572 1503 2580 1506
rect 2552 1497 2580 1503
rect 2664 1497 2691 1503
rect 2909 1503 2915 1523
rect 4269 1517 4280 1523
rect 2877 1497 2915 1503
rect 3160 1497 3187 1503
rect 3373 1497 3411 1503
rect 3752 1497 3779 1503
rect 4024 1497 4067 1503
rect 4604 1506 4612 1512
rect 4813 1503 4819 1523
rect 4989 1517 5060 1523
rect 5052 1512 5060 1517
rect 5293 1517 5347 1523
rect 5084 1506 5092 1512
rect 4776 1497 4787 1503
rect 4813 1497 4867 1503
rect 5533 1497 5560 1503
rect 5725 1503 5731 1523
rect 5693 1497 5731 1503
rect 5853 1503 5859 1523
rect 5821 1497 5859 1503
rect 5932 1503 5940 1506
rect 5912 1497 5940 1503
rect 5997 1497 6008 1503
rect 6221 1503 6227 1523
rect 6189 1497 6227 1503
rect 6637 1503 6643 1523
rect 6957 1517 6968 1523
rect 6637 1497 6691 1503
rect 7197 1503 7203 1523
rect 7165 1497 7203 1503
rect 7437 1503 7443 1523
rect 7656 1517 7667 1523
rect 7405 1497 7443 1503
rect 7720 1497 7731 1503
rect 7880 1497 7907 1503
rect 2856 1477 2867 1483
rect 2957 1477 3027 1483
rect 3469 1477 3496 1483
rect 3549 1477 3592 1483
rect 3976 1477 3987 1483
rect 4077 1477 4104 1483
rect 4221 1477 4275 1483
rect 4408 1477 4435 1483
rect 4888 1477 4915 1483
rect 172 1463 180 1472
rect 152 1457 180 1463
rect 3068 1463 3076 1466
rect 2008 1457 2019 1463
rect 2237 1457 2275 1463
rect 3037 1457 3076 1463
rect 3421 1457 3432 1463
rect 4093 1457 4140 1463
rect 4388 1457 4408 1463
rect 4909 1457 4915 1477
rect 5368 1477 5411 1483
rect 5644 1477 5683 1483
rect 5644 1472 5652 1477
rect 6108 1477 6152 1483
rect 6424 1477 6451 1483
rect 6701 1477 6728 1483
rect 6829 1477 6856 1483
rect 7021 1477 7048 1483
rect 7144 1477 7155 1483
rect 7309 1477 7347 1483
rect 7432 1477 7443 1483
rect 6397 1457 6408 1463
rect 7048 1457 7068 1463
rect 7357 1457 7368 1463
rect 1208 1437 1219 1443
rect 4333 1437 4344 1443
rect 4461 1437 4472 1443
rect 2584 1377 2595 1383
rect 7384 1377 7395 1383
rect 7720 1377 7731 1383
rect 7768 1377 7779 1383
rect 61 1357 83 1363
rect 61 1343 67 1357
rect 925 1357 1011 1363
rect 1272 1357 1283 1363
rect 2285 1357 2307 1363
rect 29 1337 67 1343
rect 1277 1337 1304 1343
rect 1469 1337 1496 1343
rect 1821 1337 1832 1343
rect 2285 1343 2291 1357
rect 3180 1348 3188 1354
rect 4392 1357 4412 1363
rect 2253 1337 2291 1343
rect 2333 1337 2360 1343
rect 2648 1337 2675 1343
rect 2808 1337 2819 1343
rect 3464 1337 3475 1343
rect 3992 1337 4024 1343
rect 4733 1343 4739 1363
rect 4888 1357 4900 1363
rect 5629 1357 5640 1363
rect 4892 1354 4900 1357
rect 6040 1357 6084 1363
rect 6076 1354 6084 1357
rect 4685 1337 4723 1343
rect 4733 1337 4760 1343
rect 5068 1337 5112 1343
rect 5581 1337 5619 1343
rect 5757 1337 5795 1343
rect 6285 1337 6312 1343
rect 6381 1343 6387 1363
rect 6333 1337 6387 1343
rect 6952 1337 6963 1343
rect 7960 1337 7987 1343
rect 7997 1337 8008 1343
rect 892 1317 904 1323
rect 892 1312 900 1317
rect 1165 1317 1192 1323
rect 2845 1317 2856 1323
rect 2909 1317 2963 1323
rect 317 1283 323 1303
rect 1688 1297 1715 1303
rect 1901 1297 1912 1303
rect 2584 1297 2595 1303
rect 2909 1297 2915 1317
rect 3341 1317 3363 1323
rect 3628 1317 3640 1323
rect 3628 1312 3636 1317
rect 3932 1317 3944 1323
rect 3932 1312 3940 1317
rect 3981 1317 3992 1323
rect 4024 1317 4051 1323
rect 4781 1317 4819 1323
rect 3549 1297 3560 1303
rect 4813 1297 4819 1317
rect 4984 1317 5011 1323
rect 5277 1317 5304 1323
rect 5453 1317 5507 1323
rect 5453 1297 5459 1317
rect 5544 1317 5555 1323
rect 5976 1317 5987 1323
rect 6141 1317 6152 1323
rect 6184 1317 6195 1323
rect 6824 1317 6851 1323
rect 7453 1317 7464 1323
rect 5640 1297 5667 1303
rect 5677 1297 5715 1303
rect 6541 1297 6552 1303
rect 7629 1297 7683 1303
rect 317 1277 355 1283
rect 349 1257 355 1277
rect 1564 1277 1603 1283
rect 1597 1257 1603 1277
rect 3624 1277 3652 1283
rect 3816 1277 3843 1283
rect 4456 1277 4483 1283
rect 1005 1177 1016 1183
rect 3736 1177 3747 1183
rect 157 1137 168 1143
rect 888 1137 952 1143
rect 4200 1137 4211 1143
rect 4360 1137 4372 1143
rect 4364 1132 4372 1137
rect 4408 1137 4440 1143
rect 4557 1143 4563 1163
rect 4524 1137 4563 1143
rect 4524 1132 4532 1137
rect 4680 1137 4692 1143
rect 4684 1132 4692 1137
rect 4749 1143 4755 1163
rect 4728 1137 4755 1143
rect 920 1117 963 1123
rect 1725 1117 1736 1123
rect 2301 1117 2312 1123
rect 2868 1116 2872 1124
rect 3132 1117 3160 1123
rect 3132 1112 3140 1117
rect 1757 1097 1800 1103
rect 2312 1097 2355 1103
rect 2376 1097 2419 1103
rect 2813 1097 2840 1103
rect 2877 1097 2904 1103
rect 3021 1097 3048 1103
rect 3213 1103 3219 1123
rect 3181 1097 3219 1103
rect 3389 1103 3395 1123
rect 3357 1097 3395 1103
rect 3517 1103 3523 1123
rect 3768 1117 3779 1123
rect 3992 1117 4003 1123
rect 4413 1117 4424 1123
rect 4808 1117 4819 1123
rect 3485 1097 3523 1103
rect 3896 1097 3907 1103
rect 4925 1103 4931 1123
rect 4893 1097 4931 1103
rect 4968 1097 4995 1103
rect 5085 1097 5096 1103
rect 604 1077 616 1083
rect 604 1076 612 1077
rect 701 1077 712 1083
rect 1048 1077 1059 1083
rect 1181 1077 1192 1083
rect 1437 1077 1448 1083
rect 1480 1077 1491 1083
rect 1949 1077 2020 1083
rect 2012 1072 2020 1077
rect 2237 1077 2259 1083
rect 2700 1077 2728 1083
rect 2700 1072 2708 1077
rect 3261 1077 3299 1083
rect 3672 1077 3683 1083
rect 4040 1077 4051 1083
rect 4989 1083 4995 1097
rect 5165 1103 5171 1123
rect 5133 1097 5171 1103
rect 5244 1103 5252 1106
rect 5224 1097 5252 1103
rect 5501 1103 5507 1123
rect 5336 1097 5363 1103
rect 5469 1097 5507 1103
rect 5837 1103 5843 1123
rect 5672 1097 5699 1103
rect 5805 1097 5843 1103
rect 6221 1097 6232 1103
rect 6472 1097 6483 1103
rect 6536 1097 6563 1103
rect 6589 1103 6595 1123
rect 7112 1117 7123 1123
rect 6589 1097 6643 1103
rect 7437 1103 7443 1123
rect 7405 1097 7443 1103
rect 7469 1097 7480 1103
rect 7757 1103 7763 1123
rect 7725 1097 7763 1103
rect 7901 1097 7912 1103
rect 4989 1077 5059 1083
rect 5213 1077 5224 1083
rect 5549 1077 5560 1083
rect 5756 1077 5768 1083
rect 6168 1077 6211 1083
rect 6344 1077 6387 1083
rect 7053 1077 7112 1083
rect 7485 1077 7496 1083
rect 7805 1077 7816 1083
rect 7965 1077 7987 1083
rect 717 1057 728 1063
rect 1197 1057 1208 1063
rect 1453 1057 1464 1063
rect 1613 1057 1651 1063
rect 3912 1057 3923 1063
rect 5997 1057 6083 1063
rect 6248 1057 6259 1063
rect 6828 1063 6836 1072
rect 6808 1057 6836 1063
rect 7212 1066 7220 1072
rect 7548 1066 7556 1072
rect 6888 1057 6908 1063
rect 2456 1037 2467 1043
rect 4360 1037 4371 1043
rect 4680 1037 4691 1043
rect 6952 1037 6963 1043
rect 7016 1037 7027 1043
rect 7080 1037 7123 1043
rect 248 977 259 983
rect 440 977 451 983
rect 2557 977 2568 983
rect 3944 977 3955 983
rect 7592 977 7603 983
rect 7821 977 7832 983
rect 301 957 355 963
rect 1181 957 1219 963
rect 1416 957 1427 963
rect 1672 957 1700 963
rect 60 948 68 952
rect 1692 948 1700 957
rect 2381 957 2392 963
rect 2456 957 2467 963
rect 3148 957 3160 963
rect 3148 954 3156 957
rect 4008 957 4060 963
rect 5496 957 5508 963
rect 5500 954 5508 957
rect 6445 957 6499 963
rect 6637 957 6648 963
rect 2220 948 2228 952
rect 328 937 371 943
rect 568 937 595 943
rect 1165 937 1192 943
rect 1416 937 1443 943
rect 1544 937 1556 943
rect 2008 937 2019 943
rect 2477 937 2515 943
rect 760 917 771 923
rect 1373 917 1432 923
rect 2845 937 2872 943
rect 3981 937 4024 943
rect 4557 937 4568 943
rect 4780 937 4835 943
rect 5005 937 5075 943
rect 5293 937 5331 943
rect 5368 937 5379 943
rect 6968 937 6995 943
rect 7096 937 7107 943
rect 7308 943 7316 948
rect 7288 937 7316 943
rect 7848 937 7860 943
rect 2429 917 2440 923
rect 2472 917 2483 923
rect 3037 917 3064 923
rect 3245 917 3272 923
rect 3405 917 3443 923
rect 1016 897 1027 903
rect 2808 897 2819 903
rect 3437 897 3443 917
rect 3916 917 3944 923
rect 3916 912 3924 917
rect 4492 917 4504 923
rect 4492 912 4500 917
rect 4669 917 4680 923
rect 5704 917 5715 923
rect 5848 917 5875 923
rect 6168 917 6179 923
rect 6413 917 6456 923
rect 6776 917 6787 923
rect 7112 917 7123 923
rect 7149 917 7203 923
rect 4333 897 4344 903
rect 5352 897 5395 903
rect 5405 897 5432 903
rect 7149 897 7155 917
rect 7416 917 7427 923
rect 1032 877 1059 883
rect 1686 876 1688 884
rect 3318 876 3320 884
rect 3768 877 3779 883
rect 3948 883 3956 888
rect 3928 877 3956 883
rect 4044 883 4052 888
rect 3992 877 4052 883
rect 4168 877 4195 883
rect 5096 777 5107 783
rect 1000 737 1016 743
rect 1256 737 1272 743
rect 4205 743 4211 763
rect 4205 737 4260 743
rect 4252 732 4260 737
rect 6408 737 6419 743
rect 7304 736 7306 744
rect 1277 717 1288 723
rect 1341 717 1363 723
rect 204 703 212 706
rect 204 697 216 703
rect 1400 697 1416 703
rect 2333 697 2360 703
rect 2749 697 2776 703
rect 2860 703 2868 706
rect 2860 697 2888 703
rect 2957 697 3016 703
rect 3133 703 3139 723
rect 3388 717 3427 723
rect 3437 717 3475 723
rect 3388 712 3396 717
rect 4216 717 4227 723
rect 4408 717 4451 723
rect 4552 717 4564 723
rect 4556 712 4564 717
rect 3101 697 3139 703
rect 3356 706 3364 712
rect 3576 697 3619 703
rect 3656 697 3667 703
rect 3741 697 3768 703
rect 4488 697 4499 703
rect 4973 703 4979 723
rect 4973 697 5027 703
rect 5192 697 5219 703
rect 5501 703 5507 723
rect 7128 717 7139 723
rect 7149 717 7187 723
rect 7256 717 7268 723
rect 7260 712 7268 717
rect 5469 697 5507 703
rect 5672 697 5699 703
rect 6253 697 6280 703
rect 6504 697 6531 703
rect 7352 697 7379 703
rect 7644 703 7652 706
rect 7644 697 7656 703
rect 7901 697 7928 703
rect 7980 706 7988 712
rect 264 677 307 683
rect 328 677 387 683
rect 824 677 851 683
rect 1528 677 1539 683
rect 1613 677 1652 683
rect 1644 672 1652 677
rect 1933 677 2004 683
rect 1996 672 2004 677
rect 2493 677 2520 683
rect 3016 677 3027 683
rect 3821 677 3832 683
rect 4024 677 4083 683
rect 4349 677 4387 683
rect 4861 677 4899 683
rect 5037 677 5108 683
rect 5100 672 5108 677
rect 5341 677 5352 683
rect 5549 677 5560 683
rect 5933 677 5944 683
rect 6013 677 6024 683
rect 6845 677 6899 683
rect 204 663 212 666
rect 492 663 500 666
rect 204 657 227 663
rect 237 657 291 663
rect 413 657 451 663
rect 461 657 500 663
rect 524 663 532 672
rect 524 657 552 663
rect 749 657 787 663
rect 877 657 915 663
rect 925 657 952 663
rect 2444 663 2452 666
rect 2444 657 2483 663
rect 3848 657 3859 663
rect 4248 657 4268 663
rect 5304 657 5324 663
rect 6893 657 6899 677
rect 4525 637 4536 643
rect 5976 637 5987 643
rect 1960 577 2003 583
rect 2984 577 3011 583
rect 4168 577 4179 583
rect 4856 577 4867 583
rect 6040 577 6083 583
rect 349 543 355 563
rect 1112 557 1140 563
rect 1132 548 1140 557
rect 1256 557 1267 563
rect 1661 557 1699 563
rect 2892 557 2931 563
rect 2892 554 2900 557
rect 3384 557 3412 563
rect 3404 548 3412 557
rect 3800 557 3812 563
rect 3804 554 3812 557
rect 5896 557 5924 563
rect 5916 548 5924 557
rect 6824 557 6852 563
rect 6844 548 6852 557
rect 349 537 387 543
rect 552 537 568 543
rect 1261 537 1315 543
rect 1464 537 1475 543
rect 1645 537 1672 543
rect 2120 537 2147 543
rect 2344 537 2355 543
rect 2445 537 2467 543
rect 856 517 867 523
rect 2077 517 2136 523
rect 2445 523 2451 537
rect 2520 537 2531 543
rect 3176 537 3187 543
rect 3565 537 3576 543
rect 4744 537 4755 543
rect 5036 537 5064 543
rect 5197 537 5208 543
rect 5576 537 5587 543
rect 5688 537 5699 543
rect 6941 537 6952 543
rect 7132 543 7140 548
rect 7080 537 7140 543
rect 7725 537 7763 543
rect 2429 517 2451 523
rect 2541 517 2579 523
rect 204 503 212 508
rect 204 497 227 503
rect 461 483 467 503
rect 461 477 499 483
rect 493 457 499 477
rect 589 483 595 503
rect 1805 497 1827 503
rect 2573 497 2579 517
rect 3549 517 3560 523
rect 3896 517 3923 523
rect 4140 517 4152 523
rect 4140 512 4148 517
rect 4252 517 4264 523
rect 4252 512 4260 517
rect 4301 517 4339 523
rect 2648 497 2659 503
rect 2920 497 2947 503
rect 3048 497 3059 503
rect 3485 497 3523 503
rect 3540 496 3544 504
rect 3672 497 3683 503
rect 3693 497 3731 503
rect 4333 497 4339 517
rect 4504 517 4531 523
rect 4653 517 4707 523
rect 4653 497 4659 517
rect 5117 517 5155 523
rect 5149 497 5155 517
rect 5245 517 5283 523
rect 5277 497 5283 517
rect 5688 517 5715 523
rect 6184 517 6195 523
rect 7021 517 7059 523
rect 7021 497 7027 517
rect 7224 517 7251 523
rect 7672 517 7699 523
rect 589 477 627 483
rect 621 457 627 477
rect 1126 476 1128 484
rect 1133 377 1144 383
rect 2152 377 2163 383
rect 3016 377 3043 383
rect 93 337 104 343
rect 1080 337 1123 343
rect 1336 337 1379 343
rect 392 317 403 323
rect 573 317 595 323
rect 1080 317 1091 323
rect 1336 317 1347 323
rect 1837 297 1848 303
rect 1901 303 1907 323
rect 2077 303 2083 323
rect 1901 297 1955 303
rect 2045 297 2083 303
rect 2508 303 2516 304
rect 2296 297 2323 303
rect 2461 297 2516 303
rect 2717 303 2723 323
rect 2685 297 2723 303
rect 3116 306 3124 312
rect 3357 303 3363 312
rect 3320 297 3363 303
rect 3677 297 3688 303
rect 3869 297 3880 303
rect 3912 297 3923 303
rect 4072 297 4083 303
rect 4136 297 4147 303
rect 4301 303 4307 323
rect 4493 317 4520 323
rect 4301 297 4355 303
rect 4413 297 4424 303
rect 4557 303 4563 323
rect 4440 297 4467 303
rect 4557 297 4584 303
rect 88 277 104 283
rect 701 277 712 283
rect 1837 277 1859 283
rect 1965 277 2024 283
rect 2125 277 2163 283
rect 2173 277 2212 283
rect 2204 272 2212 277
rect 2488 277 2499 283
rect 2568 277 2611 283
rect 3352 277 3379 283
rect 3416 277 3443 283
rect 3693 277 3704 283
rect 4429 277 4440 283
rect 4461 277 4467 297
rect 4684 306 4692 312
rect 4909 303 4915 323
rect 4877 297 4915 303
rect 5085 297 5112 303
rect 5261 303 5267 323
rect 5421 317 5459 323
rect 6669 317 6723 323
rect 5261 297 5315 303
rect 5736 297 5763 303
rect 6173 297 6200 303
rect 6284 303 6292 306
rect 6284 297 6328 303
rect 6493 297 6520 303
rect 6856 297 6883 303
rect 7085 303 7091 323
rect 7085 297 7155 303
rect 7288 297 7315 303
rect 7565 303 7571 323
rect 7533 297 7571 303
rect 7677 303 7683 323
rect 7645 297 7683 303
rect 4541 277 4552 283
rect 4957 277 5000 283
rect 5336 277 5363 283
rect 717 257 755 263
rect 828 263 836 272
rect 828 257 856 263
rect 1213 257 1251 263
rect 1485 257 1539 263
rect 1644 266 1652 272
rect 2972 263 2980 266
rect 2972 257 3016 263
rect 5357 257 5363 277
rect 5565 277 5603 283
rect 5624 277 5652 283
rect 5820 277 5832 283
rect 5644 272 5652 277
rect 5885 277 5939 283
rect 6776 277 6787 283
rect 7085 277 7128 283
rect 7176 277 7204 283
rect 7196 272 7204 277
rect 7372 277 7400 283
rect 7736 277 7747 283
rect 5613 257 5624 263
rect 4109 237 4120 243
rect 4173 237 4184 243
rect 1352 177 1363 183
rect 1944 177 1987 183
rect 3864 177 3875 183
rect 4456 177 4467 183
rect 4760 177 4771 183
rect 7560 177 7571 183
rect 7768 177 7779 183
rect 269 157 291 163
rect 60 148 68 152
rect 269 143 275 157
rect 397 157 419 163
rect 237 137 275 143
rect 397 143 403 157
rect 616 157 644 163
rect 636 148 644 157
rect 328 137 355 143
rect 365 137 403 143
rect 264 117 291 123
rect 349 117 355 137
rect 989 143 995 163
rect 1272 157 1300 163
rect 1292 148 1300 157
rect 3276 157 3315 163
rect 3276 154 3284 157
rect 4632 157 4660 163
rect 4652 148 4660 157
rect 5752 157 5764 163
rect 5756 154 5764 157
rect 6088 157 6132 163
rect 6124 154 6132 157
rect 6776 157 6804 163
rect 6796 148 6804 157
rect 6984 157 7028 163
rect 7020 154 7028 157
rect 7480 157 7508 163
rect 7500 148 7508 157
rect 989 137 1027 143
rect 1144 137 1156 143
rect 1404 143 1412 148
rect 1373 137 1412 143
rect 2028 143 2036 148
rect 1997 137 2036 143
rect 2412 143 2420 148
rect 2381 137 2420 143
rect 2744 137 2755 143
rect 3389 137 3411 143
rect 461 117 472 123
rect 904 117 947 123
rect 1645 117 1699 123
rect 1645 97 1651 117
rect 2269 117 2323 123
rect 2269 97 2275 117
rect 2653 117 2707 123
rect 2957 117 3027 123
rect 2296 97 2307 103
rect 2653 97 2659 117
rect 3021 97 3027 117
rect 3389 123 3395 137
rect 5260 137 5300 143
rect 6061 137 6104 143
rect 6557 137 6568 143
rect 3373 117 3395 123
rect 3528 117 3539 123
rect 3976 117 3987 123
rect 4296 117 4307 123
rect 4856 117 4883 123
rect 5357 117 5384 123
rect 5645 117 5683 123
rect 5533 97 5587 103
rect 5677 97 5683 117
rect 5848 117 5875 123
rect 6216 117 6243 123
rect 6365 117 6403 123
rect 5981 97 6019 103
rect 6365 97 6371 117
rect 6557 117 6611 123
rect 6557 97 6563 117
rect 7112 117 7139 123
rect 7245 117 7283 123
rect 6877 97 6915 103
rect 7277 97 7283 117
rect 7656 117 7683 123
rect 7880 117 7891 123
<< m2contact >>
rect 925 5602 961 5618
rect 2957 5602 2993 5618
rect 5021 5602 5057 5618
rect 7053 5602 7089 5618
rect 2872 5572 2888 5588
rect 2920 5572 2936 5588
rect 3000 5572 3016 5588
rect 3048 5572 3064 5588
rect 3096 5572 3112 5588
rect 3224 5572 3240 5588
rect 3320 5572 3336 5588
rect 4136 5572 4152 5588
rect 4184 5572 4200 5588
rect 4232 5572 4248 5588
rect 1640 5512 1656 5528
rect 1912 5512 1928 5528
rect 2120 5512 2136 5528
rect 2216 5512 2248 5528
rect 2456 5512 2472 5528
rect 3592 5512 3608 5528
rect 72 5492 88 5508
rect 184 5492 200 5508
rect 232 5490 248 5506
rect 376 5492 392 5508
rect 648 5490 664 5506
rect 728 5492 744 5508
rect 824 5492 856 5508
rect 952 5492 968 5508
rect 984 5492 1000 5508
rect 1064 5490 1080 5506
rect 1320 5492 1336 5508
rect 1560 5490 1576 5506
rect 1800 5492 1816 5508
rect 2056 5490 2072 5506
rect 2136 5492 2168 5508
rect 2328 5492 2344 5508
rect 2472 5492 2504 5508
rect 2584 5490 2600 5506
rect 2792 5492 2808 5508
rect 2840 5492 2856 5508
rect 2888 5492 2904 5508
rect 2936 5492 2952 5508
rect 2984 5492 3000 5508
rect 3064 5492 3080 5508
rect 3160 5492 3192 5508
rect 3240 5492 3256 5508
rect 3288 5492 3304 5508
rect 3480 5490 3496 5506
rect 3628 5512 3644 5528
rect 3640 5492 3656 5508
rect 3752 5512 3768 5528
rect 4792 5512 4808 5528
rect 3896 5492 3912 5508
rect 4056 5492 4072 5508
rect 4104 5492 4120 5508
rect 4152 5492 4168 5508
rect 4200 5492 4216 5508
rect 4360 5492 4376 5508
rect 4568 5492 4584 5508
rect 4680 5492 4712 5508
rect 4904 5492 4920 5508
rect 5048 5492 5080 5508
rect 5112 5512 5128 5528
rect 5176 5492 5192 5508
rect 5208 5492 5224 5508
rect 5240 5512 5256 5528
rect 5912 5512 5928 5528
rect 5368 5492 5384 5508
rect 5592 5492 5608 5508
rect 5848 5490 5864 5506
rect 5928 5492 5960 5508
rect 5992 5492 6024 5508
rect 6088 5512 6104 5528
rect 6232 5492 6248 5508
rect 6440 5492 6456 5508
rect 6568 5492 6600 5508
rect 6632 5512 6648 5528
rect 6936 5512 6952 5528
rect 6744 5490 6760 5506
rect 7720 5512 7752 5528
rect 6968 5492 6984 5508
rect 7016 5492 7032 5508
rect 7144 5492 7160 5508
rect 7336 5492 7352 5508
rect 7560 5492 7576 5508
rect 7688 5492 7704 5508
rect 7752 5492 7784 5508
rect 7864 5490 7880 5506
rect 632 5472 648 5488
rect 744 5472 776 5488
rect 136 5452 152 5468
rect 584 5452 600 5468
rect 792 5452 808 5468
rect 872 5452 888 5468
rect 968 5472 984 5488
rect 1096 5472 1112 5488
rect 1304 5472 1320 5488
rect 1592 5472 1608 5488
rect 1672 5472 1704 5488
rect 1832 5472 1848 5488
rect 2088 5472 2104 5488
rect 2168 5472 2184 5488
rect 2200 5472 2216 5488
rect 2280 5472 2296 5488
rect 2504 5472 2520 5488
rect 2728 5472 2744 5488
rect 2824 5472 2840 5488
rect 3112 5472 3128 5488
rect 3272 5472 3288 5488
rect 3384 5472 3400 5488
rect 3448 5472 3464 5488
rect 3560 5472 3576 5488
rect 3656 5472 3688 5488
rect 3720 5472 3736 5488
rect 3976 5472 3992 5488
rect 4088 5472 4104 5488
rect 4328 5472 4344 5488
rect 4552 5472 4568 5488
rect 4648 5472 4680 5488
rect 4744 5472 4760 5488
rect 4888 5472 4904 5488
rect 5016 5472 5048 5488
rect 5144 5472 5176 5488
rect 5272 5472 5288 5488
rect 5384 5472 5400 5488
rect 5448 5472 5464 5488
rect 5608 5472 5624 5488
rect 5880 5472 5896 5488
rect 5960 5472 5976 5488
rect 6120 5472 6136 5488
rect 6248 5472 6264 5488
rect 6456 5472 6472 5488
rect 6552 5472 6568 5488
rect 6664 5472 6680 5488
rect 6712 5472 6728 5488
rect 6904 5472 6920 5488
rect 7000 5472 7016 5488
rect 7032 5472 7048 5488
rect 7224 5472 7240 5488
rect 7256 5472 7272 5488
rect 7432 5472 7448 5488
rect 7672 5472 7688 5488
rect 7784 5472 7800 5488
rect 7832 5472 7848 5488
rect 1128 5452 1144 5468
rect 1368 5452 1384 5468
rect 1496 5452 1512 5468
rect 2408 5452 2424 5468
rect 2584 5452 2600 5468
rect 4296 5452 4312 5468
rect 5784 5452 5800 5468
rect 6808 5452 6824 5468
rect 7608 5452 7624 5468
rect 7928 5452 7944 5468
rect 40 5432 56 5448
rect 504 5432 520 5448
rect 1640 5432 1656 5448
rect 1720 5432 1736 5448
rect 1768 5432 1784 5448
rect 1880 5432 1896 5448
rect 1928 5432 1944 5448
rect 3336 5432 3352 5448
rect 3816 5432 3832 5448
rect 5496 5432 5512 5448
rect 6344 5432 6360 5448
rect 7464 5432 7480 5448
rect 7720 5432 7736 5448
rect 1949 5402 1985 5418
rect 3997 5402 4033 5418
rect 6045 5402 6081 5418
rect 392 5372 408 5388
rect 520 5372 536 5388
rect 1432 5372 1448 5388
rect 1528 5372 1544 5388
rect 1592 5372 1608 5388
rect 1688 5372 1704 5388
rect 2088 5372 2104 5388
rect 2168 5372 2184 5388
rect 2200 5372 2216 5388
rect 2296 5372 2312 5388
rect 2632 5372 2648 5388
rect 2888 5372 2904 5388
rect 2984 5372 3000 5388
rect 3192 5372 3208 5388
rect 3928 5372 3944 5388
rect 4360 5372 4376 5388
rect 4424 5372 4440 5388
rect 5512 5372 5528 5388
rect 5608 5372 5624 5388
rect 5848 5372 5864 5388
rect 5912 5372 5928 5388
rect 5992 5372 6008 5388
rect 6248 5372 6264 5388
rect 6360 5372 6376 5388
rect 7336 5372 7352 5388
rect 7400 5372 7416 5388
rect 7624 5372 7640 5388
rect 88 5352 104 5368
rect 216 5352 232 5368
rect 184 5332 200 5348
rect 248 5332 264 5348
rect 376 5332 392 5348
rect 424 5352 440 5368
rect 584 5352 600 5368
rect 808 5352 824 5368
rect 88 5312 104 5328
rect 152 5314 168 5330
rect 248 5312 264 5328
rect 328 5312 360 5328
rect 504 5332 520 5348
rect 632 5332 648 5348
rect 840 5332 856 5348
rect 888 5352 904 5368
rect 984 5352 1000 5368
rect 1400 5352 1416 5368
rect 1656 5352 1672 5368
rect 2136 5352 2152 5368
rect 2408 5352 2424 5368
rect 3416 5352 3432 5368
rect 3544 5352 3560 5368
rect 4088 5352 4104 5368
rect 4632 5352 4648 5368
rect 6568 5352 6584 5368
rect 7688 5352 7704 5368
rect 1224 5332 1240 5348
rect 1352 5332 1384 5348
rect 1480 5332 1496 5348
rect 1576 5332 1592 5348
rect 1784 5332 1800 5348
rect 1928 5332 1944 5348
rect 2024 5332 2040 5348
rect 2216 5332 2232 5348
rect 2248 5332 2264 5348
rect 2392 5332 2408 5348
rect 2488 5332 2504 5348
rect 2680 5332 2696 5348
rect 2808 5332 2824 5348
rect 3016 5332 3032 5348
rect 3272 5332 3288 5348
rect 3432 5332 3448 5348
rect 3480 5332 3496 5348
rect 3720 5332 3736 5348
rect 3768 5332 3784 5348
rect 3864 5332 3880 5348
rect 3944 5332 3960 5348
rect 4072 5332 4088 5348
rect 4168 5332 4184 5348
rect 4264 5332 4280 5348
rect 4296 5332 4312 5348
rect 4408 5332 4424 5348
rect 4536 5332 4552 5348
rect 472 5312 488 5328
rect 552 5312 568 5328
rect 680 5312 696 5328
rect 728 5312 744 5328
rect 824 5312 840 5328
rect 856 5312 872 5328
rect 968 5312 984 5328
rect 1096 5312 1112 5328
rect 1160 5314 1176 5330
rect 1240 5312 1256 5328
rect 1252 5292 1268 5308
rect 1464 5312 1480 5328
rect 1496 5312 1512 5328
rect 1560 5312 1576 5328
rect 1624 5312 1640 5328
rect 1816 5314 1832 5330
rect 1896 5312 1944 5328
rect 2056 5312 2072 5328
rect 1304 5292 1320 5308
rect 1528 5292 1544 5308
rect 1880 5292 1896 5308
rect 1992 5292 2008 5308
rect 2168 5292 2184 5308
rect 2280 5292 2296 5308
rect 2328 5312 2344 5328
rect 2472 5312 2488 5328
rect 2552 5312 2584 5328
rect 2840 5312 2856 5328
rect 2904 5312 2920 5328
rect 3096 5312 3112 5328
rect 3240 5312 3256 5328
rect 2408 5292 2424 5308
rect 2776 5292 2792 5308
rect 3304 5292 3320 5308
rect 3336 5312 3368 5328
rect 3464 5312 3480 5328
rect 3688 5314 3704 5330
rect 3832 5312 3848 5328
rect 3880 5312 3896 5328
rect 3432 5292 3448 5308
rect 3816 5292 3832 5308
rect 4008 5292 4024 5308
rect 4088 5312 4104 5328
rect 4184 5312 4200 5328
rect 4044 5292 4060 5308
rect 4344 5292 4360 5308
rect 4392 5312 4408 5328
rect 4488 5312 4504 5328
rect 4632 5314 4648 5330
rect 4712 5312 4744 5328
rect 4776 5312 4792 5328
rect 4888 5332 4904 5348
rect 5224 5332 5240 5348
rect 5272 5332 5288 5348
rect 5320 5332 5336 5348
rect 5464 5332 5480 5348
rect 5560 5332 5576 5348
rect 5752 5332 5768 5348
rect 5944 5332 5960 5348
rect 6200 5332 6216 5348
rect 6296 5332 6312 5348
rect 6488 5332 6504 5348
rect 6664 5332 6680 5348
rect 6936 5332 6952 5348
rect 7000 5332 7016 5348
rect 7032 5332 7048 5348
rect 7256 5332 7272 5348
rect 7288 5332 7304 5348
rect 7352 5332 7368 5348
rect 7448 5332 7480 5348
rect 7592 5332 7608 5348
rect 7640 5332 7656 5348
rect 7736 5332 7768 5348
rect 7784 5332 7800 5348
rect 7976 5332 7992 5348
rect 4968 5312 5000 5328
rect 5112 5312 5144 5328
rect 5176 5312 5208 5328
rect 4840 5292 4856 5308
rect 5256 5292 5272 5308
rect 5304 5312 5320 5328
rect 5368 5312 5384 5328
rect 5416 5312 5448 5328
rect 5496 5292 5512 5308
rect 5544 5312 5560 5328
rect 5672 5312 5688 5328
rect 5832 5312 5848 5328
rect 5880 5312 5896 5328
rect 6024 5312 6040 5328
rect 6088 5312 6120 5328
rect 6200 5312 6216 5328
rect 5896 5292 5912 5308
rect 6232 5292 6248 5308
rect 6280 5312 6296 5328
rect 6328 5312 6344 5328
rect 6408 5312 6424 5328
rect 6420 5292 6436 5308
rect 6568 5314 6584 5330
rect 6792 5312 6808 5328
rect 6824 5312 6840 5328
rect 6856 5312 6872 5328
rect 6904 5312 6936 5328
rect 6952 5312 6968 5328
rect 6456 5292 6472 5308
rect 7176 5312 7192 5328
rect 7304 5312 7320 5328
rect 7368 5312 7384 5328
rect 7000 5292 7016 5308
rect 7336 5292 7352 5308
rect 7480 5312 7512 5328
rect 7544 5312 7560 5328
rect 7656 5312 7672 5328
rect 7416 5292 7432 5308
rect 7624 5292 7640 5308
rect 7896 5312 7912 5328
rect 7704 5292 7720 5308
rect 7784 5292 7800 5308
rect 3144 5272 3160 5288
rect 2168 5232 2184 5248
rect 2728 5232 2744 5248
rect 2792 5232 2808 5248
rect 3192 5232 3208 5248
rect 3512 5232 3528 5248
rect 3560 5232 3576 5248
rect 3784 5232 3800 5248
rect 4760 5232 4776 5248
rect 4824 5232 4840 5248
rect 5160 5232 5176 5248
rect 5400 5232 5416 5248
rect 5608 5232 5624 5248
rect 5704 5232 5720 5248
rect 5848 5232 5864 5248
rect 6136 5232 6152 5248
rect 6776 5232 6792 5248
rect 6872 5232 6888 5248
rect 7528 5232 7544 5248
rect 7768 5232 7784 5248
rect 925 5202 961 5218
rect 2957 5202 2993 5218
rect 5021 5202 5057 5218
rect 7053 5202 7089 5218
rect 2952 5172 2968 5188
rect 3176 5172 3192 5188
rect 3784 5172 3800 5188
rect 3832 5172 3848 5188
rect 7384 5172 7400 5188
rect 7976 5172 7992 5188
rect 1944 5152 1960 5168
rect 5080 5132 5096 5148
rect 7704 5132 7720 5148
rect 280 5112 296 5128
rect 88 5092 104 5108
rect 136 5092 152 5108
rect 216 5092 232 5108
rect 344 5092 360 5108
rect 456 5092 472 5108
rect 664 5092 680 5108
rect 952 5090 968 5106
rect 1064 5092 1096 5108
rect 1128 5112 1144 5128
rect 1368 5090 1384 5106
rect 1448 5092 1480 5108
rect 1512 5112 1528 5128
rect 1844 5112 1860 5128
rect 1864 5112 1880 5128
rect 2056 5112 2072 5128
rect 2168 5112 2184 5128
rect 2264 5112 2280 5128
rect 1752 5090 1768 5106
rect 1832 5092 1848 5108
rect 2088 5092 2104 5108
rect 2296 5092 2312 5108
rect 2360 5112 2376 5128
rect 2664 5112 2680 5128
rect 2760 5112 2776 5128
rect 3016 5112 3032 5128
rect 3064 5112 3096 5128
rect 3416 5112 3432 5128
rect 2488 5092 2504 5108
rect 2744 5092 2760 5108
rect 2792 5092 2808 5108
rect 2840 5092 2856 5108
rect 2920 5092 2936 5108
rect 3128 5092 3144 5108
rect 3288 5092 3304 5108
rect 3384 5092 3400 5108
rect 3496 5112 3512 5128
rect 3608 5112 3624 5128
rect 3640 5112 3656 5128
rect 3848 5112 3864 5128
rect 4008 5112 4024 5128
rect 3464 5092 3480 5108
rect 3528 5092 3544 5108
rect 3624 5092 3640 5108
rect 3704 5092 3720 5108
rect 3752 5092 3768 5108
rect 3800 5092 3816 5108
rect 3896 5092 3912 5108
rect 4376 5112 4392 5128
rect 4088 5092 4104 5108
rect 4264 5090 4280 5106
rect 4408 5092 4440 5108
rect 4472 5092 4488 5108
rect 4520 5092 4536 5108
rect 4616 5112 4632 5128
rect 4872 5112 4888 5128
rect 4936 5112 4952 5128
rect 5240 5112 5256 5128
rect 4744 5092 4776 5108
rect 4888 5092 4904 5108
rect 4920 5092 4936 5108
rect 4952 5092 4984 5108
rect 5128 5092 5144 5108
rect 5256 5092 5288 5108
rect 5304 5092 5320 5108
rect 5368 5090 5384 5106
rect 5432 5092 5448 5108
rect 5608 5092 5624 5108
rect 5640 5092 5656 5108
rect 5832 5092 5848 5108
rect 5912 5092 5928 5108
rect 5944 5092 5960 5108
rect 5992 5112 6008 5128
rect 6088 5092 6120 5108
rect 6152 5092 6168 5108
rect 6296 5092 6328 5108
rect 6488 5092 6504 5108
rect 6616 5092 6632 5108
rect 6680 5112 6696 5128
rect 6936 5112 6952 5128
rect 6808 5092 6824 5108
rect 6840 5092 6856 5108
rect 6952 5092 6984 5108
rect 7128 5092 7144 5108
rect 7256 5092 7272 5108
rect 7320 5112 7336 5128
rect 7368 5112 7384 5128
rect 7544 5112 7560 5128
rect 7880 5112 7896 5128
rect 7448 5092 7464 5108
rect 7496 5092 7528 5108
rect 7608 5092 7624 5108
rect 7640 5092 7656 5108
rect 7752 5092 7768 5108
rect 7944 5092 7960 5108
rect 40 5072 56 5088
rect 216 5052 232 5068
rect 248 5052 264 5068
rect 312 5072 328 5088
rect 376 5072 392 5088
rect 584 5072 600 5088
rect 808 5072 824 5088
rect 984 5072 1000 5088
rect 1048 5072 1064 5088
rect 1160 5072 1176 5088
rect 1336 5072 1352 5088
rect 1432 5072 1448 5088
rect 1544 5072 1560 5088
rect 1736 5072 1752 5088
rect 1784 5072 1800 5088
rect 1816 5072 1832 5088
rect 2008 5072 2040 5088
rect 2232 5072 2248 5088
rect 2280 5072 2296 5088
rect 2344 5072 2360 5088
rect 2392 5072 2408 5088
rect 2440 5072 2456 5088
rect 2536 5072 2552 5088
rect 2616 5072 2648 5088
rect 2808 5072 2824 5088
rect 2872 5072 2888 5088
rect 3080 5072 3096 5088
rect 3112 5072 3128 5088
rect 3208 5072 3224 5088
rect 3304 5072 3320 5088
rect 3432 5072 3448 5088
rect 3480 5072 3496 5088
rect 3560 5072 3576 5088
rect 3672 5072 3688 5088
rect 3736 5072 3752 5088
rect 3944 5072 3960 5088
rect 4056 5072 4072 5088
rect 4104 5072 4120 5088
rect 4328 5072 4360 5088
rect 4440 5072 4456 5088
rect 4504 5072 4520 5088
rect 4536 5072 4552 5088
rect 4616 5072 4632 5088
rect 4648 5072 4664 5088
rect 4840 5072 4856 5088
rect 4920 5072 4936 5088
rect 4984 5072 5000 5088
rect 5208 5072 5224 5088
rect 5288 5072 5304 5088
rect 5336 5072 5352 5088
rect 5752 5072 5768 5088
rect 5928 5072 5944 5088
rect 5960 5072 5976 5088
rect 6024 5072 6040 5088
rect 6168 5072 6200 5088
rect 6600 5072 6616 5088
rect 6648 5072 6664 5088
rect 6984 5072 7000 5088
rect 7208 5072 7224 5088
rect 7240 5072 7256 5088
rect 7368 5072 7384 5088
rect 7432 5072 7464 5088
rect 7576 5072 7592 5088
rect 7656 5072 7688 5088
rect 7832 5072 7848 5088
rect 7912 5072 7928 5088
rect 7976 5072 7992 5088
rect 616 5052 632 5068
rect 856 5052 872 5068
rect 3944 5052 3960 5068
rect 6344 5052 6360 5068
rect 6456 5052 6472 5068
rect 6552 5052 6568 5068
rect 7112 5052 7128 5068
rect 536 5032 552 5048
rect 1176 5032 1192 5048
rect 1560 5032 1576 5048
rect 2056 5032 2072 5048
rect 2120 5032 2136 5048
rect 2152 5032 2168 5048
rect 2248 5032 2264 5048
rect 2648 5032 2664 5048
rect 2712 5032 2728 5048
rect 2760 5032 2776 5048
rect 3096 5032 3112 5048
rect 3496 5032 3512 5048
rect 3592 5032 3608 5048
rect 3848 5032 3864 5048
rect 4120 5032 4136 5048
rect 5000 5032 5016 5048
rect 5496 5032 5528 5048
rect 6728 5032 6744 5048
rect 7288 5032 7304 5048
rect 7864 5032 7880 5048
rect 1949 5002 1985 5018
rect 3997 5002 4033 5018
rect 6045 5002 6081 5018
rect 40 4972 56 4988
rect 456 4972 472 4988
rect 984 4972 1000 4988
rect 1240 4972 1256 4988
rect 2136 4972 2152 4988
rect 3144 4972 3160 4988
rect 3784 4972 3800 4988
rect 4712 4972 4728 4988
rect 5240 4972 5256 4988
rect 5720 4972 5736 4988
rect 5816 4972 5832 4988
rect 5896 4972 5912 4988
rect 6296 4972 6312 4988
rect 6408 4972 6424 4988
rect 6488 4972 6504 4988
rect 6616 4972 6632 4988
rect 6808 4972 6824 4988
rect 6888 4972 6904 4988
rect 6936 4972 6952 4988
rect 7800 4972 7816 4988
rect 536 4952 552 4968
rect 744 4952 760 4968
rect 440 4932 456 4948
rect 616 4932 632 4948
rect 776 4932 808 4948
rect 824 4952 840 4968
rect 856 4952 888 4968
rect 1272 4952 1288 4968
rect 1480 4952 1496 4968
rect 1736 4952 1752 4968
rect 2072 4952 2088 4968
rect 3480 4952 3496 4968
rect 4120 4952 4136 4968
rect 4648 4952 4664 4968
rect 5144 4952 5160 4968
rect 5336 4952 5352 4968
rect 6184 4952 6200 4968
rect 7272 4952 7288 4968
rect 7368 4952 7384 4968
rect 7624 4952 7640 4968
rect 1000 4932 1016 4948
rect 1112 4932 1128 4948
rect 1176 4932 1192 4948
rect 1224 4932 1240 4948
rect 1528 4932 1544 4948
rect 2184 4932 2200 4948
rect 2264 4932 2280 4948
rect 2392 4932 2408 4948
rect 2440 4932 2456 4948
rect 2568 4932 2584 4948
rect 2664 4932 2680 4948
rect 2712 4932 2728 4948
rect 2984 4932 3000 4948
rect 3080 4932 3096 4948
rect 3208 4932 3224 4948
rect 3272 4932 3288 4948
rect 3400 4932 3416 4948
rect 3432 4932 3448 4948
rect 3528 4932 3560 4948
rect 3944 4932 3960 4948
rect 4024 4932 4040 4948
rect 4168 4932 4184 4948
rect 4296 4932 4312 4948
rect 4408 4932 4424 4948
rect 4456 4932 4472 4948
rect 4552 4932 4568 4948
rect 4648 4932 4664 4948
rect 4728 4932 4744 4948
rect 4856 4932 4872 4948
rect 4904 4932 4920 4948
rect 4952 4932 4968 4948
rect 5224 4932 5240 4948
rect 5576 4932 5592 4948
rect 5672 4932 5688 4948
rect 5768 4932 5784 4948
rect 5944 4932 5960 4948
rect 5992 4932 6008 4948
rect 6248 4932 6264 4948
rect 6344 4932 6360 4948
rect 6440 4932 6456 4948
rect 6552 4932 6568 4948
rect 6968 4932 6984 4948
rect 7688 4932 7704 4948
rect 7784 4932 7800 4948
rect 7832 4932 7864 4948
rect 7880 4932 7896 4948
rect 7912 4932 7928 4948
rect 7992 4932 8008 4948
rect 72 4912 88 4928
rect 120 4912 136 4928
rect 168 4912 184 4928
rect 248 4912 264 4928
rect 312 4912 328 4928
rect 376 4912 392 4928
rect 424 4912 440 4928
rect 488 4912 504 4928
rect 632 4912 648 4928
rect 760 4912 776 4928
rect 856 4912 872 4928
rect 904 4912 920 4928
rect 1016 4912 1032 4928
rect 1064 4912 1080 4928
rect 1160 4912 1176 4928
rect 1224 4912 1240 4928
rect 1304 4912 1320 4928
rect 1384 4912 1400 4928
rect 1432 4912 1448 4928
rect 1512 4912 1528 4928
rect 1576 4912 1592 4928
rect 1640 4912 1656 4928
rect 1784 4912 1816 4928
rect 1976 4912 2008 4928
rect 2040 4912 2056 4928
rect 2296 4912 2328 4928
rect 136 4892 168 4908
rect 264 4892 280 4908
rect 328 4892 344 4908
rect 408 4892 424 4908
rect 1080 4892 1096 4908
rect 1288 4892 1304 4908
rect 1400 4892 1416 4908
rect 1592 4892 1608 4908
rect 1656 4892 1672 4908
rect 2024 4892 2040 4908
rect 2472 4914 2488 4930
rect 2632 4912 2648 4928
rect 2680 4912 2696 4928
rect 2744 4914 2760 4930
rect 3064 4912 3080 4928
rect 3112 4912 3128 4928
rect 3304 4912 3320 4928
rect 3352 4912 3368 4928
rect 2360 4892 2376 4908
rect 2616 4892 2632 4908
rect 2888 4892 2904 4908
rect 3160 4892 3176 4908
rect 3464 4892 3480 4908
rect 3512 4912 3528 4928
rect 3560 4912 3592 4928
rect 3640 4912 3656 4928
rect 3688 4912 3704 4928
rect 3752 4912 3768 4928
rect 3832 4912 3848 4928
rect 3880 4912 3896 4928
rect 3592 4892 3608 4908
rect 3656 4892 3672 4908
rect 3720 4892 3736 4908
rect 3848 4892 3880 4908
rect 3976 4892 3992 4908
rect 4072 4912 4088 4928
rect 4248 4912 4264 4928
rect 4392 4892 4408 4908
rect 4440 4912 4456 4928
rect 4488 4912 4504 4928
rect 4568 4912 4584 4928
rect 4760 4912 4792 4928
rect 4824 4912 4840 4928
rect 4856 4912 4888 4928
rect 4696 4892 4712 4908
rect 5096 4912 5112 4928
rect 5384 4912 5400 4928
rect 5480 4912 5496 4928
rect 5512 4912 5528 4928
rect 5560 4912 5576 4928
rect 5592 4912 5640 4928
rect 4920 4892 4936 4908
rect 5272 4892 5288 4908
rect 5640 4892 5656 4908
rect 5704 4892 5720 4908
rect 5752 4912 5768 4928
rect 5880 4912 5896 4928
rect 5928 4912 5960 4928
rect 6136 4912 6152 4928
rect 6264 4912 6280 4928
rect 5992 4892 6008 4908
rect 6344 4912 6360 4928
rect 6456 4912 6472 4928
rect 6312 4892 6328 4908
rect 6584 4912 6600 4928
rect 6664 4912 6696 4928
rect 6728 4912 6744 4928
rect 6776 4912 6792 4928
rect 6856 4912 6872 4928
rect 7000 4912 7016 4928
rect 7112 4912 7144 4928
rect 7176 4912 7192 4928
rect 7288 4912 7304 4928
rect 7336 4912 7352 4928
rect 7432 4912 7448 4928
rect 7496 4912 7528 4928
rect 7720 4914 7736 4930
rect 7864 4912 7880 4928
rect 7928 4912 7944 4928
rect 6520 4892 6536 4908
rect 6936 4892 6952 4908
rect 7800 4892 7816 4908
rect 7896 4892 7912 4908
rect 7940 4892 7956 4908
rect 7960 4892 7992 4908
rect 8024 4892 8040 4908
rect 184 4872 200 4888
rect 232 4872 248 4888
rect 296 4872 312 4888
rect 360 4872 376 4888
rect 1048 4872 1064 4888
rect 312 4852 328 4868
rect 1320 4872 1336 4888
rect 1368 4872 1384 4888
rect 1416 4872 1432 4888
rect 1560 4872 1576 4888
rect 1624 4872 1640 4888
rect 2840 4872 2856 4888
rect 3624 4872 3640 4888
rect 3688 4872 3704 4888
rect 3816 4872 3832 4888
rect 3896 4872 3912 4888
rect 6408 4852 6424 4868
rect 40 4832 56 4848
rect 120 4832 136 4848
rect 200 4832 216 4848
rect 248 4832 264 4848
rect 376 4832 392 4848
rect 1336 4832 1352 4848
rect 1384 4832 1400 4848
rect 1576 4832 1592 4848
rect 1608 4832 1624 4848
rect 1944 4832 1960 4848
rect 2216 4832 2232 4848
rect 3064 4832 3080 4848
rect 3192 4832 3208 4848
rect 3640 4832 3656 4848
rect 3704 4832 3720 4848
rect 3832 4832 3848 4848
rect 3928 4832 3944 4848
rect 4664 4832 4680 4848
rect 4808 4832 4824 4848
rect 5464 4832 5480 4848
rect 5528 4832 5544 4848
rect 6040 4832 6056 4848
rect 6696 4832 6712 4848
rect 7032 4832 7048 4848
rect 7144 4832 7160 4848
rect 7464 4832 7480 4848
rect 7544 4832 7560 4848
rect 925 4802 961 4818
rect 2957 4802 2993 4818
rect 5021 4802 5057 4818
rect 7053 4802 7089 4818
rect 360 4772 376 4788
rect 408 4772 424 4788
rect 2776 4772 2792 4788
rect 2904 4772 2920 4788
rect 3688 4772 3704 4788
rect 4072 4772 4088 4788
rect 4200 4772 4216 4788
rect 4376 4772 4392 4788
rect 4488 4772 4504 4788
rect 4600 4772 4616 4788
rect 5624 4772 5640 4788
rect 5976 4772 5992 4788
rect 7688 4772 7704 4788
rect 536 4752 552 4768
rect 792 4752 808 4768
rect 984 4752 1000 4768
rect 3864 4752 3880 4768
rect 168 4732 184 4748
rect 232 4732 248 4748
rect 280 4732 296 4748
rect 344 4732 360 4748
rect 424 4732 440 4748
rect 488 4732 504 4748
rect 552 4732 568 4748
rect 808 4732 824 4748
rect 888 4732 904 4748
rect 968 4732 984 4748
rect 1752 4732 1768 4748
rect 2760 4732 2776 4748
rect 2888 4732 2904 4748
rect 3704 4732 3720 4748
rect 3880 4732 3896 4748
rect 4056 4732 4072 4748
rect 4504 4732 4520 4748
rect 5256 4732 5272 4748
rect 5384 4732 5400 4748
rect 6232 4732 6248 4748
rect 6936 4732 6952 4748
rect 7176 4732 7192 4748
rect 136 4712 152 4728
rect 200 4712 216 4728
rect 312 4712 328 4728
rect 376 4712 408 4728
rect 456 4712 472 4728
rect 520 4712 536 4728
rect 824 4712 840 4728
rect 936 4712 952 4728
rect 1000 4712 1016 4728
rect 24 4692 40 4708
rect 88 4692 104 4708
rect 152 4692 168 4708
rect 216 4692 232 4708
rect 248 4692 264 4708
rect 280 4692 296 4708
rect 360 4692 376 4708
rect 408 4692 424 4708
rect 472 4692 488 4708
rect 536 4692 552 4708
rect 696 4692 712 4708
rect 824 4692 840 4708
rect 872 4692 888 4708
rect 984 4692 1000 4708
rect 1016 4692 1032 4708
rect 1048 4692 1064 4708
rect 1096 4712 1112 4728
rect 1144 4712 1160 4728
rect 1336 4712 1352 4728
rect 1400 4712 1416 4728
rect 1464 4712 1480 4728
rect 1656 4712 1672 4728
rect 1720 4712 1736 4728
rect 1848 4712 1864 4728
rect 1912 4712 1928 4728
rect 2056 4712 2072 4728
rect 2280 4712 2296 4728
rect 2344 4712 2360 4728
rect 2364 4712 2380 4728
rect 2856 4712 2872 4728
rect 2936 4712 2952 4728
rect 3240 4712 3256 4728
rect 3368 4712 3384 4728
rect 3800 4712 3816 4728
rect 3928 4712 3944 4728
rect 3948 4712 3964 4728
rect 4088 4712 4104 4728
rect 4184 4712 4200 4728
rect 4216 4712 4232 4728
rect 4312 4712 4328 4728
rect 4392 4712 4408 4728
rect 4936 4712 4952 4728
rect 5448 4712 5464 4728
rect 5640 4712 5656 4728
rect 5704 4712 5720 4728
rect 5784 4712 5800 4728
rect 5816 4712 5832 4728
rect 5944 4712 5960 4728
rect 6328 4712 6344 4728
rect 6348 4712 6364 4728
rect 6568 4712 6584 4728
rect 7064 4712 7096 4728
rect 1176 4692 1192 4708
rect 1272 4692 1288 4708
rect 1368 4692 1384 4708
rect 1448 4692 1464 4708
rect 1496 4692 1512 4708
rect 1592 4692 1608 4708
rect 1704 4692 1720 4708
rect 1736 4692 1752 4708
rect 1816 4692 1832 4708
rect 1880 4692 1896 4708
rect 1944 4692 1960 4708
rect 1976 4692 1992 4708
rect 2024 4692 2056 4708
rect 2136 4690 2152 4706
rect 2376 4692 2392 4708
rect 2472 4692 2488 4708
rect 2616 4692 2648 4708
rect 2760 4692 2776 4708
rect 2824 4692 2840 4708
rect 2856 4692 2872 4708
rect 2888 4692 2904 4708
rect 2920 4692 2936 4708
rect 2952 4692 2984 4708
rect 3096 4690 3112 4706
rect 3160 4692 3176 4708
rect 3432 4692 3464 4708
rect 3544 4690 3560 4706
rect 3720 4692 3736 4708
rect 3752 4692 3768 4708
rect 3832 4692 3848 4708
rect 3896 4692 3912 4708
rect 3928 4692 3944 4708
rect 3976 4692 3992 4708
rect 4056 4692 4072 4708
rect 4088 4692 4104 4708
rect 4120 4692 4136 4708
rect 4152 4692 4168 4708
rect 4184 4692 4200 4708
rect 4232 4692 4248 4708
rect 4264 4692 4296 4708
rect 4392 4692 4408 4708
rect 4424 4692 4472 4708
rect 4504 4692 4520 4708
rect 4552 4692 4584 4708
rect 4632 4692 4648 4708
rect 4840 4692 4856 4708
rect 4984 4692 5000 4708
rect 5080 4692 5096 4708
rect 5128 4692 5144 4708
rect 5192 4692 5208 4708
rect 5224 4692 5240 4708
rect 5256 4692 5272 4708
rect 5304 4692 5320 4708
rect 5368 4692 5384 4708
rect 5416 4692 5448 4708
rect 5480 4692 5496 4708
rect 5512 4692 5528 4708
rect 5560 4692 5576 4708
rect 40 4672 56 4688
rect 72 4672 88 4688
rect 616 4672 632 4688
rect 1016 4672 1032 4688
rect 1128 4672 1144 4688
rect 1160 4672 1176 4688
rect 1192 4672 1208 4688
rect 1256 4672 1288 4688
rect 1384 4672 1400 4688
rect 1448 4672 1464 4688
rect 1512 4672 1528 4688
rect 1608 4672 1624 4688
rect 1704 4672 1720 4688
rect 1832 4672 1848 4688
rect 1896 4672 1912 4688
rect 1992 4672 2024 4688
rect 2104 4672 2120 4688
rect 2328 4672 2344 4688
rect 2392 4672 2424 4688
rect 2488 4672 2504 4688
rect 2824 4672 2840 4688
rect 3032 4672 3048 4688
rect 3368 4672 3384 4688
rect 3400 4672 3416 4688
rect 3464 4672 3480 4688
rect 3512 4672 3528 4688
rect 3768 4672 3784 4688
rect 3848 4672 3864 4688
rect 3976 4672 3992 4688
rect 4136 4672 4152 4688
rect 4264 4672 4280 4688
rect 4344 4672 4360 4688
rect 5000 4672 5016 4688
rect 5128 4672 5144 4688
rect 120 4652 136 4668
rect 280 4652 296 4668
rect 504 4652 520 4668
rect 744 4652 760 4668
rect 1848 4652 1864 4668
rect 2200 4652 2216 4668
rect 3096 4652 3112 4668
rect 3608 4652 3624 4668
rect 3752 4652 3768 4668
rect 4024 4652 4040 4668
rect 4360 4652 4376 4668
rect 4472 4652 4488 4668
rect 4760 4652 4776 4668
rect 4856 4652 4872 4668
rect 5112 4652 5128 4668
rect 5176 4672 5192 4688
rect 5240 4672 5256 4688
rect 5352 4672 5368 4688
rect 5416 4672 5432 4688
rect 5672 4692 5704 4708
rect 5736 4692 5752 4708
rect 5848 4692 5864 4708
rect 5880 4692 5896 4708
rect 6008 4692 6024 4708
rect 6072 4692 6088 4708
rect 6120 4692 6136 4708
rect 6168 4692 6184 4708
rect 6200 4692 6216 4708
rect 6232 4692 6248 4708
rect 6312 4692 6328 4708
rect 6392 4692 6408 4708
rect 6424 4692 6456 4708
rect 6472 4692 6504 4708
rect 6536 4692 6552 4708
rect 6600 4692 6616 4708
rect 6632 4692 6648 4708
rect 6696 4692 6744 4708
rect 6760 4692 6776 4708
rect 6808 4692 6824 4708
rect 6872 4692 6888 4708
rect 6904 4692 6920 4708
rect 6936 4692 6952 4708
rect 7000 4692 7032 4708
rect 7096 4692 7128 4708
rect 7160 4712 7176 4728
rect 7400 4712 7416 4728
rect 7528 4712 7544 4728
rect 7288 4692 7304 4708
rect 7432 4692 7448 4708
rect 7512 4692 7528 4708
rect 7560 4692 7576 4708
rect 7608 4692 7624 4708
rect 7656 4692 7672 4708
rect 7736 4692 7752 4708
rect 7784 4712 7800 4728
rect 7992 4712 8008 4728
rect 7912 4692 7928 4708
rect 5656 4672 5672 4688
rect 5720 4672 5736 4688
rect 6040 4672 6056 4688
rect 6152 4672 6168 4688
rect 6216 4672 6232 4688
rect 6392 4672 6408 4688
rect 6616 4672 6632 4688
rect 6664 4672 6680 4688
rect 6744 4672 6760 4688
rect 6856 4672 6872 4688
rect 6888 4672 6904 4688
rect 6920 4672 6936 4688
rect 6984 4672 7000 4688
rect 7128 4672 7144 4688
rect 7336 4672 7352 4688
rect 7448 4672 7464 4688
rect 7480 4672 7496 4688
rect 7704 4672 7736 4688
rect 7784 4672 7800 4688
rect 7816 4672 7832 4688
rect 7864 4672 7880 4688
rect 5224 4652 5240 4668
rect 5304 4652 5320 4668
rect 5336 4652 5352 4668
rect 5480 4652 5496 4668
rect 5528 4652 5544 4668
rect 6264 4652 6296 4668
rect 6392 4652 6408 4668
rect 6440 4652 6456 4668
rect 6664 4652 6680 4668
rect 6792 4652 6808 4668
rect 6840 4652 6856 4668
rect 6968 4652 6984 4668
rect 7576 4652 7592 4668
rect 184 4632 200 4648
rect 1400 4632 1416 4648
rect 1464 4632 1480 4648
rect 1608 4632 1624 4648
rect 1784 4632 1800 4648
rect 1912 4632 1928 4648
rect 2296 4632 2312 4648
rect 3288 4632 3304 4648
rect 4680 4632 4696 4648
rect 5320 4632 5336 4648
rect 5768 4632 5784 4648
rect 5912 4632 5928 4648
rect 6088 4632 6104 4648
rect 6200 4632 6216 4648
rect 6296 4632 6312 4648
rect 6472 4632 6488 4648
rect 6648 4632 6664 4648
rect 6776 4632 6792 4648
rect 6824 4632 6840 4648
rect 7400 4632 7416 4648
rect 7496 4632 7512 4648
rect 1949 4602 1985 4618
rect 3997 4602 4033 4618
rect 6045 4602 6081 4618
rect 376 4572 392 4588
rect 456 4572 472 4588
rect 792 4572 808 4588
rect 856 4572 872 4588
rect 1048 4572 1064 4588
rect 1208 4572 1224 4588
rect 1384 4572 1400 4588
rect 1720 4572 1736 4588
rect 1768 4572 1784 4588
rect 1880 4572 1896 4588
rect 2152 4572 2168 4588
rect 2312 4572 2328 4588
rect 3608 4572 3624 4588
rect 3672 4572 3688 4588
rect 3704 4572 3720 4588
rect 3896 4572 3912 4588
rect 4104 4572 4120 4588
rect 4200 4572 4216 4588
rect 4264 4572 4280 4588
rect 4856 4572 4872 4588
rect 4968 4572 4984 4588
rect 5064 4572 5080 4588
rect 5272 4572 5288 4588
rect 5496 4572 5512 4588
rect 5560 4572 5576 4588
rect 5704 4572 5720 4588
rect 5784 4572 5800 4588
rect 5864 4572 5880 4588
rect 5960 4572 5976 4588
rect 6232 4572 6248 4588
rect 6328 4572 6344 4588
rect 6472 4572 6488 4588
rect 6712 4572 6728 4588
rect 6936 4572 6952 4588
rect 7064 4572 7080 4588
rect 7416 4572 7432 4588
rect 920 4552 936 4568
rect 1112 4552 1128 4568
rect 1464 4552 1480 4568
rect 1752 4552 1768 4568
rect 1896 4552 1912 4568
rect 3208 4552 3224 4568
rect 3912 4552 3928 4568
rect 4120 4552 4136 4568
rect 4408 4552 4424 4568
rect 4728 4552 4744 4568
rect 5224 4552 5240 4568
rect 40 4532 56 4548
rect 568 4532 584 4548
rect 744 4532 760 4548
rect 920 4532 936 4548
rect 72 4514 88 4530
rect 136 4512 152 4528
rect 248 4512 264 4528
rect 296 4512 312 4528
rect 360 4512 376 4528
rect 424 4512 440 4528
rect 504 4512 520 4528
rect 568 4512 584 4528
rect 616 4512 632 4528
rect 680 4512 696 4528
rect 840 4512 856 4528
rect 888 4512 904 4528
rect 968 4532 984 4548
rect 1000 4532 1016 4548
rect 1064 4532 1080 4548
rect 1192 4532 1208 4548
rect 1304 4532 1320 4548
rect 1432 4532 1464 4548
rect 1704 4532 1720 4548
rect 1816 4532 1832 4548
rect 1912 4532 1944 4548
rect 2152 4532 2168 4548
rect 2200 4532 2216 4548
rect 2232 4532 2248 4548
rect 952 4512 968 4528
rect 1016 4512 1032 4528
rect 1080 4512 1096 4528
rect 1192 4512 1208 4528
rect 1288 4512 1304 4528
rect 1352 4512 1368 4528
rect 1416 4512 1432 4528
rect 1496 4512 1512 4528
rect 1608 4512 1624 4528
rect 1704 4512 1720 4528
rect 1800 4512 1816 4528
rect 1896 4512 1912 4528
rect 2056 4512 2072 4528
rect 2296 4532 2312 4548
rect 2440 4532 2456 4548
rect 2536 4532 2552 4548
rect 2632 4532 2648 4548
rect 2744 4532 2760 4548
rect 2776 4532 2792 4548
rect 2968 4532 2984 4548
rect 3080 4532 3096 4548
rect 3144 4532 3176 4548
rect 3224 4532 3240 4548
rect 3544 4532 3560 4548
rect 3608 4532 3624 4548
rect 3752 4532 3768 4548
rect 3800 4532 3832 4548
rect 3864 4532 3880 4548
rect 4120 4532 4136 4548
rect 4184 4532 4200 4548
rect 4296 4532 4312 4548
rect 4488 4532 4504 4548
rect 4536 4532 4552 4548
rect 4584 4532 4600 4548
rect 2264 4512 2280 4528
rect 2408 4512 2424 4528
rect 200 4492 216 4508
rect 232 4472 248 4488
rect 280 4492 296 4508
rect 344 4492 360 4508
rect 408 4492 424 4508
rect 520 4492 536 4508
rect 248 4452 264 4468
rect 312 4472 328 4488
rect 344 4472 360 4488
rect 440 4472 456 4488
rect 488 4472 504 4488
rect 552 4472 568 4488
rect 600 4492 616 4508
rect 664 4492 680 4508
rect 984 4492 1000 4508
rect 1048 4492 1064 4508
rect 1128 4492 1144 4508
rect 1256 4492 1272 4508
rect 1320 4492 1352 4508
rect 1544 4492 1560 4508
rect 1624 4492 1640 4508
rect 1768 4492 1784 4508
rect 2312 4492 2328 4508
rect 2664 4492 2680 4508
rect 2696 4512 2728 4528
rect 2808 4514 2824 4530
rect 3128 4512 3160 4528
rect 3224 4512 3240 4528
rect 3256 4512 3272 4528
rect 3320 4512 3336 4528
rect 3368 4512 3384 4528
rect 3432 4512 3448 4528
rect 3496 4512 3512 4528
rect 3736 4512 3752 4528
rect 3768 4512 3784 4528
rect 3832 4512 3848 4528
rect 3880 4512 3896 4528
rect 3944 4512 3960 4528
rect 3976 4512 3992 4528
rect 4040 4512 4056 4528
rect 4072 4512 4104 4528
rect 4408 4514 4424 4530
rect 3128 4492 3144 4508
rect 3208 4492 3224 4508
rect 3304 4492 3320 4508
rect 3368 4492 3384 4508
rect 3416 4492 3432 4508
rect 3560 4492 3576 4508
rect 3800 4492 3816 4508
rect 3864 4492 3880 4508
rect 3928 4492 3944 4508
rect 3992 4492 4008 4508
rect 4520 4492 4536 4508
rect 4568 4512 4584 4528
rect 4680 4532 4696 4548
rect 4792 4532 4824 4548
rect 4920 4532 4936 4548
rect 5000 4532 5016 4548
rect 5112 4532 5128 4548
rect 5416 4552 5432 4568
rect 5992 4552 6008 4568
rect 6056 4552 6072 4568
rect 6184 4552 6200 4568
rect 5272 4532 5288 4548
rect 5336 4532 5352 4548
rect 5480 4532 5496 4548
rect 5544 4532 5560 4548
rect 5608 4532 5624 4548
rect 5688 4532 5704 4548
rect 5784 4532 5800 4548
rect 5816 4532 5832 4548
rect 6072 4532 6088 4548
rect 6136 4532 6152 4548
rect 6616 4552 6632 4568
rect 6664 4552 6680 4568
rect 6728 4552 6744 4568
rect 7832 4552 7848 4568
rect 6232 4532 6248 4548
rect 6408 4532 6424 4548
rect 6536 4532 6552 4548
rect 6808 4532 6824 4548
rect 6872 4532 6888 4548
rect 6984 4532 7000 4548
rect 7112 4532 7128 4548
rect 7144 4532 7160 4548
rect 7208 4532 7224 4548
rect 7304 4532 7320 4548
rect 7432 4532 7448 4548
rect 7496 4532 7512 4548
rect 4664 4512 4680 4528
rect 4696 4512 4712 4528
rect 4728 4492 4744 4508
rect 4760 4492 4776 4508
rect 4840 4492 4856 4508
rect 4888 4512 4904 4528
rect 4936 4512 4952 4528
rect 5128 4512 5144 4528
rect 5176 4512 5208 4528
rect 5288 4512 5304 4528
rect 5384 4512 5400 4528
rect 5528 4512 5544 4528
rect 5640 4512 5656 4528
rect 5896 4512 5912 4528
rect 5928 4512 5944 4528
rect 6024 4512 6040 4528
rect 6088 4512 6104 4528
rect 6120 4512 6136 4528
rect 6152 4512 6168 4528
rect 6248 4512 6264 4528
rect 6520 4512 6552 4528
rect 6632 4512 6648 4528
rect 6728 4512 6744 4528
rect 6824 4512 6856 4528
rect 6888 4512 6920 4528
rect 6968 4512 6984 4528
rect 7016 4512 7032 4528
rect 7192 4512 7208 4528
rect 7304 4512 7320 4528
rect 7464 4512 7480 4528
rect 7512 4512 7528 4528
rect 7576 4532 7592 4548
rect 7624 4532 7640 4548
rect 7672 4532 7688 4548
rect 7960 4532 7976 4548
rect 7592 4512 7608 4528
rect 5448 4492 5464 4508
rect 5496 4492 5512 4508
rect 5576 4492 5592 4508
rect 5720 4492 5736 4508
rect 5784 4492 5800 4508
rect 6344 4492 6360 4508
rect 6440 4492 6456 4508
rect 6856 4492 6872 4508
rect 6920 4492 6952 4508
rect 7000 4492 7016 4508
rect 7112 4492 7128 4508
rect 7160 4492 7176 4508
rect 7432 4492 7448 4508
rect 7784 4512 7800 4528
rect 7976 4512 7992 4528
rect 7640 4492 7656 4508
rect 7912 4492 7928 4508
rect 632 4472 648 4488
rect 680 4472 696 4488
rect 1352 4472 1368 4488
rect 1592 4472 1608 4488
rect 1608 4452 1624 4468
rect 3320 4472 3336 4488
rect 3352 4472 3368 4488
rect 3448 4472 3464 4488
rect 3496 4472 3512 4488
rect 3592 4472 3608 4488
rect 3656 4472 3672 4488
rect 3960 4472 3976 4488
rect 3992 4472 4008 4488
rect 4184 4472 4200 4488
rect 4248 4472 4264 4488
rect 3400 4452 3416 4468
rect 504 4432 520 4448
rect 712 4432 728 4448
rect 2216 4432 2232 4448
rect 2584 4432 2600 4448
rect 3432 4432 3448 4448
rect 3512 4432 3528 4448
rect 4776 4432 4792 4448
rect 5864 4432 5880 4448
rect 5960 4432 5976 4448
rect 6104 4432 6120 4448
rect 6472 4432 6488 4448
rect 7928 4432 7944 4448
rect 8008 4432 8024 4448
rect 925 4402 961 4418
rect 2957 4402 2993 4418
rect 5021 4402 5057 4418
rect 7053 4402 7089 4418
rect 392 4372 408 4388
rect 504 4372 520 4388
rect 584 4372 600 4388
rect 856 4372 872 4388
rect 888 4372 904 4388
rect 984 4372 1000 4388
rect 1032 4372 1048 4388
rect 1128 4372 1144 4388
rect 1208 4372 1224 4388
rect 2824 4372 2840 4388
rect 2856 4372 2872 4388
rect 2920 4372 2936 4388
rect 3096 4372 3112 4388
rect 3160 4372 3176 4388
rect 3400 4372 3416 4388
rect 3480 4372 3496 4388
rect 3544 4372 3560 4388
rect 3592 4372 3608 4388
rect 3656 4372 3672 4388
rect 3800 4372 3816 4388
rect 3848 4372 3864 4388
rect 3928 4372 3944 4388
rect 4008 4372 4024 4388
rect 4856 4372 4872 4388
rect 6680 4372 6696 4388
rect 6888 4372 6904 4388
rect 7336 4372 7352 4388
rect 424 4352 440 4368
rect 616 4352 632 4368
rect 1928 4352 1944 4368
rect 232 4332 248 4348
rect 312 4332 328 4348
rect 360 4332 392 4348
rect 440 4332 456 4348
rect 488 4332 504 4348
rect 568 4332 584 4348
rect 632 4332 648 4348
rect 696 4332 712 4348
rect 744 4332 776 4348
rect 792 4332 808 4348
rect 904 4332 920 4348
rect 968 4332 984 4348
rect 1048 4332 1064 4348
rect 1112 4332 1128 4348
rect 1176 4332 1192 4348
rect 1912 4332 1928 4348
rect 2024 4332 2040 4348
rect 3144 4332 3176 4348
rect 3464 4332 3480 4348
rect 3544 4332 3560 4348
rect 3672 4332 3688 4348
rect 3784 4332 3800 4348
rect 3816 4332 3832 4348
rect 3912 4332 3928 4348
rect 3976 4332 4008 4348
rect 6536 4332 6552 4348
rect 6936 4332 6952 4348
rect 248 4312 264 4328
rect 344 4312 360 4328
rect 408 4312 424 4328
rect 520 4312 552 4328
rect 600 4312 616 4328
rect 664 4312 680 4328
rect 728 4312 744 4328
rect 776 4312 808 4328
rect 920 4312 936 4328
rect 1016 4312 1032 4328
rect 1080 4312 1096 4328
rect 1144 4312 1160 4328
rect 1304 4312 1320 4328
rect 1944 4312 1960 4328
rect 2120 4312 2136 4328
rect 2200 4312 2216 4328
rect 2296 4312 2312 4328
rect 2872 4312 2888 4328
rect 2904 4312 2920 4328
rect 2936 4312 2952 4328
rect 3000 4312 3016 4328
rect 3080 4312 3096 4328
rect 3112 4312 3128 4328
rect 3176 4312 3192 4328
rect 3256 4312 3272 4328
rect 3320 4312 3336 4328
rect 3496 4312 3512 4328
rect 3560 4312 3592 4328
rect 3640 4312 3656 4328
rect 3704 4312 3720 4328
rect 3816 4312 3848 4328
rect 3944 4312 3976 4328
rect 4312 4312 4328 4328
rect 4904 4312 4920 4328
rect 4936 4312 4952 4328
rect 152 4290 168 4306
rect 248 4292 264 4308
rect 296 4292 312 4308
rect 360 4292 376 4308
rect 424 4292 440 4308
rect 504 4292 520 4308
rect 552 4292 568 4308
rect 616 4292 632 4308
rect 680 4292 696 4308
rect 744 4292 760 4308
rect 808 4292 824 4308
rect 984 4292 1000 4308
rect 1032 4292 1048 4308
rect 1096 4292 1112 4308
rect 1160 4292 1176 4308
rect 1272 4292 1288 4308
rect 1432 4292 1448 4308
rect 1480 4292 1496 4308
rect 1640 4292 1656 4308
rect 1784 4292 1800 4308
rect 1848 4292 1864 4308
rect 1928 4292 1944 4308
rect 2008 4292 2024 4308
rect 2088 4292 2104 4308
rect 2184 4292 2200 4308
rect 2264 4292 2296 4308
rect 2440 4292 2472 4308
rect 2888 4292 2904 4308
rect 2952 4292 2968 4308
rect 3016 4292 3048 4308
rect 3096 4292 3112 4308
rect 3144 4292 3160 4308
rect 3192 4292 3208 4308
rect 3432 4292 3448 4308
rect 3480 4292 3496 4308
rect 3528 4292 3544 4308
rect 3608 4292 3624 4308
rect 3656 4292 3672 4308
rect 3736 4292 3752 4308
rect 3800 4292 3816 4308
rect 3848 4292 3864 4308
rect 3928 4292 3944 4308
rect 3976 4292 3992 4308
rect 4152 4292 4168 4308
rect 4344 4292 4360 4308
rect 4472 4292 4488 4308
rect 4648 4292 4664 4308
rect 4680 4292 4696 4308
rect 4808 4292 4824 4308
rect 5464 4312 5480 4328
rect 5720 4312 5736 4328
rect 5832 4312 5848 4328
rect 4968 4292 5000 4308
rect 5144 4292 5160 4308
rect 5368 4292 5384 4308
rect 5464 4292 5480 4308
rect 5512 4292 5528 4308
rect 5640 4292 5672 4308
rect 5752 4292 5784 4308
rect 5880 4292 5896 4308
rect 5928 4292 5944 4308
rect 5960 4292 5992 4308
rect 6040 4292 6056 4308
rect 6072 4312 6088 4328
rect 6136 4312 6152 4328
rect 6408 4312 6424 4328
rect 6104 4292 6120 4308
rect 6232 4290 6248 4306
rect 6776 4312 6792 4328
rect 6456 4292 6472 4308
rect 6504 4292 6520 4308
rect 6664 4292 6680 4308
rect 6712 4292 6728 4308
rect 6872 4312 6888 4328
rect 6968 4312 7000 4328
rect 7480 4312 7496 4328
rect 6824 4292 6840 4308
rect 7000 4292 7016 4308
rect 7032 4292 7048 4308
rect 7176 4292 7192 4308
rect 7288 4292 7304 4308
rect 7368 4292 7384 4308
rect 7400 4292 7416 4308
rect 7496 4292 7528 4308
rect 7560 4312 7576 4328
rect 7624 4312 7640 4328
rect 7624 4292 7640 4308
rect 7720 4292 7736 4308
rect 7896 4290 7912 4306
rect 7960 4292 7976 4308
rect 136 4272 152 4288
rect 232 4272 248 4288
rect 872 4272 888 4288
rect 1208 4272 1224 4288
rect 1336 4272 1352 4288
rect 1800 4272 1832 4288
rect 2104 4272 2120 4288
rect 2168 4272 2184 4288
rect 2232 4272 2264 4288
rect 2312 4272 2328 4288
rect 2680 4272 2712 4288
rect 2760 4272 2776 4288
rect 3304 4272 3320 4288
rect 3384 4272 3400 4288
rect 3720 4272 3736 4288
rect 3752 4272 3768 4288
rect 4232 4272 4248 4288
rect 4360 4272 4376 4288
rect 4504 4272 4520 4288
rect 4584 4272 4600 4288
rect 4824 4272 4840 4288
rect 4904 4272 4920 4288
rect 5000 4272 5032 4288
rect 5176 4272 5192 4288
rect 5512 4272 5528 4288
rect 5736 4272 5752 4288
rect 5800 4272 5816 4288
rect 5960 4272 5976 4288
rect 6104 4272 6120 4288
rect 6376 4272 6392 4288
rect 6472 4272 6488 4288
rect 6552 4272 6568 4288
rect 6664 4272 6680 4288
rect 6728 4272 6744 4288
rect 6840 4272 6856 4288
rect 6936 4272 6952 4288
rect 7032 4272 7048 4288
rect 7368 4272 7384 4288
rect 7448 4272 7464 4288
rect 7496 4272 7512 4288
rect 7544 4272 7560 4288
rect 7608 4272 7624 4288
rect 56 4252 72 4268
rect 1768 4252 1784 4268
rect 1880 4252 1896 4268
rect 2600 4252 2616 4268
rect 3048 4252 3064 4268
rect 3304 4252 3320 4268
rect 4296 4252 4328 4268
rect 6168 4252 6184 4268
rect 6232 4252 6248 4268
rect 6296 4252 6312 4268
rect 7224 4252 7240 4268
rect 7896 4252 7912 4268
rect 904 4232 920 4248
rect 1288 4232 1304 4248
rect 1368 4232 1384 4248
rect 2056 4232 2072 4248
rect 2120 4232 2136 4248
rect 2184 4232 2200 4248
rect 2584 4232 2600 4248
rect 2648 4232 2664 4248
rect 3400 4232 3416 4248
rect 4040 4232 4056 4248
rect 4264 4232 4280 4248
rect 4376 4232 4392 4248
rect 4712 4232 4728 4248
rect 4776 4232 4792 4248
rect 5448 4232 5464 4248
rect 5912 4232 5928 4248
rect 6424 4232 6440 4248
rect 6792 4232 6808 4248
rect 7048 4232 7064 4248
rect 8040 4232 8056 4248
rect 1949 4202 1985 4218
rect 3997 4202 4033 4218
rect 6045 4202 6081 4218
rect 152 4172 168 4188
rect 344 4172 360 4188
rect 728 4172 744 4188
rect 1384 4172 1400 4188
rect 1608 4172 1624 4188
rect 1864 4172 1880 4188
rect 2136 4172 2152 4188
rect 2296 4172 2312 4188
rect 3128 4172 3144 4188
rect 3320 4172 3336 4188
rect 3352 4172 3368 4188
rect 3704 4172 3720 4188
rect 3784 4172 3800 4188
rect 3864 4172 3880 4188
rect 3896 4172 3912 4188
rect 4360 4172 4376 4188
rect 4904 4172 4920 4188
rect 5496 4172 5512 4188
rect 5912 4172 5928 4188
rect 6024 4172 6040 4188
rect 6856 4172 6872 4188
rect 6984 4172 7000 4188
rect 7400 4172 7432 4188
rect 7992 4172 8008 4188
rect 72 4152 88 4168
rect 1304 4152 1320 4168
rect 2008 4152 2024 4168
rect 2072 4152 2088 4168
rect 2536 4152 2552 4168
rect 2600 4152 2616 4168
rect 2888 4152 2904 4168
rect 2920 4152 2936 4168
rect 3144 4152 3160 4168
rect 168 4132 184 4148
rect 696 4132 712 4148
rect 872 4132 888 4148
rect 1208 4132 1224 4148
rect 1240 4132 1256 4148
rect 1272 4132 1288 4148
rect 1400 4132 1416 4148
rect 1752 4132 1768 4148
rect 1896 4132 1912 4148
rect 1960 4132 1976 4148
rect 2056 4132 2072 4148
rect 2120 4132 2136 4148
rect 2200 4132 2216 4148
rect 2360 4132 2376 4148
rect 2456 4132 2472 4148
rect 2568 4132 2584 4148
rect 2728 4132 2744 4148
rect 2824 4132 2840 4148
rect 3032 4132 3048 4148
rect 3304 4132 3320 4148
rect 3400 4132 3416 4148
rect 4376 4152 4392 4168
rect 5720 4152 5736 4168
rect 5848 4152 5864 4168
rect 6376 4152 6392 4168
rect 7224 4152 7240 4168
rect 7288 4152 7304 4168
rect 7512 4152 7528 4168
rect 3688 4132 3704 4148
rect 3736 4132 3752 4148
rect 3816 4132 3832 4148
rect 3848 4132 3864 4148
rect 3928 4132 3944 4148
rect 3976 4132 3992 4148
rect 4040 4132 4056 4148
rect 4104 4132 4120 4148
rect 4168 4132 4184 4148
rect 4200 4132 4216 4148
rect 4232 4132 4264 4148
rect 4296 4132 4312 4148
rect 4392 4132 4408 4148
rect 4440 4132 4456 4148
rect 4680 4132 4696 4148
rect 4760 4132 4776 4148
rect 4792 4132 4808 4148
rect 4904 4132 4920 4148
rect 5144 4132 5160 4148
rect 5176 4132 5192 4148
rect 5352 4132 5368 4148
rect 5448 4132 5464 4148
rect 5544 4132 5560 4148
rect 5592 4132 5608 4148
rect 5640 4132 5656 4148
rect 5864 4132 5880 4148
rect 5944 4132 5960 4148
rect 40 4112 56 4128
rect 104 4112 136 4128
rect 184 4112 232 4128
rect 248 4112 264 4128
rect 296 4112 312 4128
rect 360 4112 376 4128
rect 472 4112 488 4128
rect 504 4112 520 4128
rect 664 4112 680 4128
rect 776 4112 792 4128
rect 824 4112 840 4128
rect 936 4112 952 4128
rect 1160 4112 1176 4128
rect 1256 4112 1272 4128
rect 1336 4112 1352 4128
rect 1416 4112 1432 4128
rect 1464 4112 1480 4128
rect 1512 4112 1528 4128
rect 1576 4112 1592 4128
rect 1672 4112 1688 4128
rect 1704 4112 1720 4128
rect 1848 4112 1864 4128
rect 1944 4112 1960 4128
rect 2040 4112 2056 4128
rect 2120 4112 2136 4128
rect 2264 4112 2280 4128
rect 56 4092 72 4108
rect 312 4092 328 4108
rect 376 4092 392 4108
rect 632 4092 648 4108
rect 728 4092 744 4108
rect 792 4092 808 4108
rect 1288 4092 1304 4108
rect 1496 4092 1512 4108
rect 1656 4092 1672 4108
rect 1688 4092 1704 4108
rect 1912 4092 1928 4108
rect 2008 4092 2024 4108
rect 2296 4092 2312 4108
rect 2392 4092 2408 4108
rect 2424 4112 2440 4128
rect 2472 4112 2488 4128
rect 2536 4114 2552 4130
rect 2744 4112 2760 4128
rect 2808 4112 2824 4128
rect 2840 4112 2856 4128
rect 2984 4112 3000 4128
rect 3064 4112 3080 4128
rect 3176 4112 3192 4128
rect 3240 4112 3256 4128
rect 3432 4112 3448 4128
rect 3480 4112 3512 4128
rect 3544 4112 3560 4128
rect 3688 4112 3704 4128
rect 3752 4112 3768 4128
rect 4040 4112 4056 4128
rect 2680 4092 2696 4108
rect 2712 4092 2728 4108
rect 2872 4092 2888 4108
rect 3096 4092 3112 4108
rect 3160 4092 3176 4108
rect 3224 4092 3240 4108
rect 3416 4092 3432 4108
rect 3544 4092 3560 4108
rect 3720 4092 3736 4108
rect 3784 4092 3800 4108
rect 3928 4092 3944 4108
rect 3992 4092 4008 4108
rect 4104 4092 4120 4108
rect 4136 4092 4152 4108
rect 4232 4112 4248 4128
rect 4408 4112 4424 4128
rect 4296 4092 4312 4108
rect 4328 4092 4344 4108
rect 4600 4112 4616 4128
rect 4456 4092 4472 4108
rect 4552 4092 4568 4108
rect 4728 4092 4744 4108
rect 4824 4092 4840 4108
rect 4856 4112 4888 4128
rect 5000 4112 5016 4128
rect 5256 4112 5288 4128
rect 5368 4112 5400 4128
rect 5448 4112 5464 4128
rect 5544 4092 5560 4108
rect 5576 4092 5592 4108
rect 5656 4112 5672 4128
rect 5768 4112 5784 4128
rect 5880 4112 5896 4128
rect 6072 4112 6104 4128
rect 6472 4132 6488 4148
rect 6744 4132 6760 4148
rect 6840 4132 6856 4148
rect 6936 4132 6968 4148
rect 7000 4132 7016 4148
rect 7048 4132 7064 4148
rect 7144 4132 7160 4148
rect 7544 4132 7560 4148
rect 7592 4132 7608 4148
rect 7672 4132 7688 4148
rect 7704 4132 7720 4148
rect 7896 4132 7912 4148
rect 7928 4132 7944 4148
rect 8040 4132 8056 4148
rect 6200 4112 6232 4128
rect 6424 4112 6440 4128
rect 6520 4112 6552 4128
rect 6584 4112 6616 4128
rect 6760 4114 6776 4130
rect 6936 4112 6952 4128
rect 7016 4112 7032 4128
rect 5976 4092 5992 4108
rect 6872 4092 6904 4108
rect 6908 4092 6924 4108
rect 6984 4092 7000 4108
rect 7224 4114 7240 4130
rect 7288 4112 7304 4128
rect 7464 4112 7480 4128
rect 7592 4112 7608 4128
rect 7112 4092 7128 4108
rect 7416 4092 7432 4108
rect 7512 4092 7528 4108
rect 7576 4092 7592 4108
rect 7640 4092 7656 4108
rect 7688 4112 7704 4128
rect 7720 4112 7736 4128
rect 7816 4112 7832 4128
rect 7944 4112 7960 4128
rect 7976 4092 7992 4108
rect 8008 4092 8024 4108
rect 24 4072 40 4088
rect 232 4072 248 4088
rect 280 4072 296 4088
rect 344 4072 360 4088
rect 808 4072 824 4088
rect 840 4072 856 4088
rect 1080 4072 1096 4088
rect 1448 4072 1464 4088
rect 1528 4072 1544 4088
rect 1704 4072 1720 4088
rect 3192 4072 3208 4088
rect 3256 4072 3272 4088
rect 3352 4072 3384 4088
rect 3448 4072 3464 4088
rect 3528 4072 3544 4088
rect 3880 4072 3896 4088
rect 3912 4072 3928 4088
rect 3176 4052 3192 4068
rect 3240 4052 3256 4068
rect 3432 4052 3448 4068
rect 8 4032 24 4048
rect 264 4032 280 4048
rect 712 4032 728 4048
rect 776 4032 792 4048
rect 872 4032 888 4048
rect 968 4032 984 4048
rect 1464 4032 1480 4048
rect 1512 4032 1528 4048
rect 2776 4032 2792 4048
rect 3016 4032 3032 4048
rect 3592 4032 3608 4048
rect 4312 4032 4328 4048
rect 4744 4032 4760 4048
rect 5416 4032 5432 4048
rect 6248 4032 6264 4048
rect 6552 4032 6568 4048
rect 7944 4032 7960 4048
rect 925 4002 961 4018
rect 2957 4002 2993 4018
rect 5021 4002 5057 4018
rect 7053 4002 7089 4018
rect 248 3972 264 3988
rect 312 3972 328 3988
rect 360 3972 376 3988
rect 504 3972 520 3988
rect 1560 3972 1576 3988
rect 1640 3972 1656 3988
rect 2856 3972 2872 3988
rect 3336 3972 3352 3988
rect 3416 3972 3432 3988
rect 3480 3972 3496 3988
rect 3544 3972 3560 3988
rect 3640 3972 3656 3988
rect 3800 3972 3816 3988
rect 3848 3972 3864 3988
rect 3912 3972 3928 3988
rect 3960 3972 3976 3988
rect 4776 3972 4792 3988
rect 5736 3972 5752 3988
rect 5832 3972 5848 3988
rect 6920 3972 6936 3988
rect 8024 3972 8040 3988
rect 1352 3952 1368 3968
rect 24 3932 40 3948
rect 88 3932 104 3948
rect 152 3932 168 3948
rect 232 3932 248 3948
rect 296 3932 312 3948
rect 344 3932 360 3948
rect 600 3932 616 3948
rect 1624 3932 1640 3948
rect 3496 3932 3512 3948
rect 3528 3932 3544 3948
rect 3560 3932 3576 3948
rect 3720 3932 3736 3948
rect 3768 3932 3784 3948
rect 3832 3932 3848 3948
rect 3896 3932 3912 3948
rect 3928 3932 3944 3948
rect 5320 3932 5336 3948
rect 6440 3932 6456 3948
rect 8 3912 24 3928
rect 56 3912 72 3928
rect 184 3912 216 3928
rect 264 3912 280 3928
rect 376 3912 392 3928
rect 936 3912 952 3928
rect 1000 3912 1016 3928
rect 1448 3912 1464 3928
rect 1512 3912 1528 3928
rect 1656 3912 1672 3928
rect 1988 3912 2004 3928
rect 2008 3912 2024 3928
rect 2072 3912 2088 3928
rect 2104 3912 2120 3928
rect 2296 3912 2312 3928
rect 2616 3912 2632 3928
rect 3160 3912 3176 3928
rect 3224 3912 3240 3928
rect 40 3892 56 3908
rect 104 3892 120 3908
rect 168 3892 184 3908
rect 216 3892 232 3908
rect 280 3892 296 3908
rect 360 3892 376 3908
rect 424 3892 440 3908
rect 488 3892 504 3908
rect 552 3892 568 3908
rect 632 3892 648 3908
rect 664 3892 680 3908
rect 728 3892 744 3908
rect 840 3892 856 3908
rect 968 3892 984 3908
rect 1032 3892 1048 3908
rect 1064 3892 1080 3908
rect 1176 3892 1192 3908
rect 1256 3892 1272 3908
rect 1384 3892 1400 3908
rect 1416 3892 1432 3908
rect 1480 3892 1496 3908
rect 1592 3892 1608 3908
rect 1640 3892 1656 3908
rect 1784 3892 1816 3908
rect 1896 3892 1912 3908
rect 1976 3892 1992 3908
rect 2040 3892 2056 3908
rect 2200 3890 2216 3906
rect 2456 3892 2472 3908
rect 2552 3892 2568 3908
rect 2584 3892 2600 3908
rect 2680 3890 2696 3906
rect 2856 3892 2872 3908
rect 3016 3892 3032 3908
rect 3128 3892 3144 3908
rect 3464 3912 3480 3928
rect 3528 3912 3544 3928
rect 3752 3912 3768 3928
rect 3864 3912 3880 3928
rect 3928 3912 3960 3928
rect 4088 3912 4104 3928
rect 4184 3912 4200 3928
rect 4552 3912 4568 3928
rect 3256 3892 3288 3908
rect 3368 3892 3384 3908
rect 3448 3892 3464 3908
rect 3480 3892 3496 3908
rect 3544 3892 3560 3908
rect 3608 3892 3624 3908
rect 3688 3892 3704 3908
rect 3768 3892 3784 3908
rect 3832 3892 3848 3908
rect 3912 3892 3928 3908
rect 3960 3892 3976 3908
rect 4040 3892 4056 3908
rect 4072 3892 4088 3908
rect 4120 3892 4136 3908
rect 4216 3892 4232 3908
rect 4440 3890 4456 3906
rect 4632 3912 4648 3928
rect 4696 3912 4712 3928
rect 5000 3912 5016 3928
rect 4600 3892 4616 3908
rect 4648 3892 4680 3908
rect 4696 3892 4712 3908
rect 4760 3892 4776 3908
rect 4856 3892 4872 3908
rect 5068 3912 5084 3928
rect 5624 3912 5640 3928
rect 5080 3892 5096 3908
rect 5112 3892 5128 3908
rect 5208 3892 5224 3908
rect 5512 3890 5528 3906
rect 5896 3912 5912 3928
rect 6296 3912 6312 3928
rect 5672 3892 5688 3908
rect 5800 3892 5816 3908
rect 5880 3892 5896 3908
rect 5912 3892 5928 3908
rect 5944 3892 5960 3908
rect 6024 3892 6040 3908
rect 6136 3892 6152 3908
rect 6168 3892 6184 3908
rect 6248 3892 6264 3908
rect 6280 3892 6296 3908
rect 6328 3892 6344 3908
rect 6392 3912 6408 3928
rect 6456 3912 6488 3928
rect 6552 3912 6568 3928
rect 6760 3912 6776 3928
rect 6520 3892 6536 3908
rect 6680 3892 6696 3908
rect 6792 3892 6824 3908
rect 6840 3912 6856 3928
rect 6904 3912 6920 3928
rect 7220 3912 7236 3928
rect 6872 3892 6888 3908
rect 7016 3890 7032 3906
rect 7208 3892 7224 3908
rect 7272 3912 7288 3928
rect 7528 3912 7544 3928
rect 7592 3912 7608 3928
rect 7640 3912 7656 3928
rect 7752 3912 7768 3928
rect 7400 3892 7416 3908
rect 7448 3892 7464 3908
rect 7592 3892 7608 3908
rect 7640 3892 7656 3908
rect 7720 3892 7736 3908
rect 7800 3892 7816 3908
rect 7944 3892 7960 3908
rect 88 3872 104 3888
rect 536 3872 552 3888
rect 680 3872 696 3888
rect 920 3872 936 3888
rect 984 3872 1000 3888
rect 1016 3872 1032 3888
rect 1048 3872 1064 3888
rect 392 3852 408 3868
rect 424 3852 440 3868
rect 760 3852 776 3868
rect 792 3852 808 3868
rect 1096 3852 1112 3868
rect 1144 3872 1176 3888
rect 1336 3872 1352 3888
rect 1400 3872 1416 3888
rect 1432 3872 1448 3888
rect 1464 3872 1480 3888
rect 1512 3872 1544 3888
rect 2024 3872 2040 3888
rect 2072 3872 2088 3888
rect 2136 3872 2152 3888
rect 2168 3872 2184 3888
rect 2440 3872 2456 3888
rect 2552 3872 2568 3888
rect 2648 3872 2664 3888
rect 2936 3872 2952 3888
rect 3112 3872 3128 3888
rect 3144 3872 3160 3888
rect 3192 3872 3208 3888
rect 3304 3872 3320 3888
rect 4024 3872 4040 3888
rect 4168 3872 4200 3888
rect 4344 3872 4360 3888
rect 4424 3872 4440 3888
rect 4504 3872 4536 3888
rect 4552 3872 4568 3888
rect 4616 3872 4632 3888
rect 4680 3872 4696 3888
rect 4744 3872 4760 3888
rect 4856 3872 4872 3888
rect 4936 3872 4952 3888
rect 4968 3872 4984 3888
rect 5096 3872 5112 3888
rect 5192 3872 5208 3888
rect 5288 3872 5304 3888
rect 5416 3872 5432 3888
rect 5592 3872 5608 3888
rect 5640 3872 5656 3888
rect 5688 3872 5704 3888
rect 5864 3872 5880 3888
rect 5928 3872 5944 3888
rect 6072 3872 6088 3888
rect 6104 3872 6120 3888
rect 6248 3872 6264 3888
rect 6312 3872 6328 3888
rect 6344 3872 6360 3888
rect 6424 3872 6440 3888
rect 6488 3872 6520 3888
rect 6776 3872 6792 3888
rect 6888 3872 6904 3888
rect 6952 3872 6968 3888
rect 6984 3872 7000 3888
rect 7192 3872 7208 3888
rect 7304 3872 7320 3888
rect 7528 3872 7544 3888
rect 7576 3872 7608 3888
rect 7704 3872 7720 3888
rect 7816 3872 7832 3888
rect 7896 3872 7912 3888
rect 1256 3852 1272 3868
rect 2744 3852 2760 3868
rect 2824 3852 2840 3868
rect 5512 3852 5528 3868
rect 5976 3852 6008 3868
rect 6040 3852 6056 3868
rect 6632 3852 6648 3868
rect 7480 3852 7496 3868
rect 7688 3852 7704 3868
rect 7960 3852 7976 3868
rect 408 3832 424 3848
rect 696 3832 712 3848
rect 856 3832 872 3848
rect 1272 3832 1288 3848
rect 2536 3832 2552 3848
rect 5960 3832 5976 3848
rect 6152 3832 6168 3848
rect 6568 3832 6584 3848
rect 7144 3832 7160 3848
rect 7768 3832 7784 3848
rect 1949 3802 1985 3818
rect 3997 3802 4033 3818
rect 6045 3802 6081 3818
rect 840 3772 856 3788
rect 968 3772 984 3788
rect 1096 3772 1112 3788
rect 1288 3772 1304 3788
rect 1688 3772 1704 3788
rect 2056 3772 2072 3788
rect 2232 3772 2248 3788
rect 2456 3772 2472 3788
rect 2632 3772 2648 3788
rect 2760 3772 2776 3788
rect 2856 3772 2872 3788
rect 3160 3772 3176 3788
rect 3400 3772 3416 3788
rect 3544 3772 3560 3788
rect 4040 3772 4056 3788
rect 4456 3772 4472 3788
rect 4520 3772 4536 3788
rect 4728 3772 4744 3788
rect 6024 3772 6040 3788
rect 6184 3772 6200 3788
rect 6312 3772 6328 3788
rect 6504 3772 6520 3788
rect 6664 3772 6680 3788
rect 6824 3772 6840 3788
rect 6888 3772 6920 3788
rect 8008 3772 8024 3788
rect 56 3752 72 3768
rect 216 3752 232 3768
rect 296 3752 312 3768
rect 392 3752 408 3768
rect 552 3752 568 3768
rect 760 3752 776 3768
rect 136 3732 152 3748
rect 312 3732 328 3748
rect 472 3732 488 3748
rect 552 3732 568 3748
rect 600 3732 616 3748
rect 1256 3732 1272 3748
rect 1448 3732 1464 3748
rect 1496 3752 1512 3768
rect 1880 3752 1896 3768
rect 2168 3752 2184 3768
rect 2536 3752 2552 3768
rect 2776 3752 2792 3768
rect 2936 3752 2952 3768
rect 3240 3752 3256 3768
rect 3336 3752 3352 3768
rect 3592 3752 3608 3768
rect 3624 3752 3640 3768
rect 3768 3752 3784 3768
rect 3912 3752 3928 3768
rect 4216 3752 4232 3768
rect 4744 3752 4760 3768
rect 4888 3752 4904 3768
rect 4952 3752 4968 3768
rect 5832 3752 5848 3768
rect 6264 3752 6280 3768
rect 6328 3752 6344 3768
rect 6376 3752 6392 3768
rect 6440 3752 6456 3768
rect 6568 3752 6584 3768
rect 7480 3752 7496 3768
rect 1672 3732 1688 3748
rect 1736 3732 1768 3748
rect 1800 3732 1816 3748
rect 1832 3732 1848 3748
rect 1864 3732 1896 3748
rect 2088 3732 2120 3748
rect 2376 3732 2392 3748
rect 2504 3732 2520 3748
rect 2664 3732 2696 3748
rect 2792 3732 2808 3748
rect 3016 3732 3032 3748
rect 3128 3732 3144 3748
rect 3256 3732 3272 3748
rect 3384 3732 3400 3748
rect 3448 3732 3464 3748
rect 152 3714 168 3730
rect 248 3712 264 3728
rect 328 3712 344 3728
rect 424 3712 440 3728
rect 488 3714 504 3730
rect 616 3712 632 3728
rect 696 3714 712 3730
rect 760 3712 776 3728
rect 872 3712 904 3728
rect 1064 3712 1080 3728
rect 1192 3712 1208 3728
rect 1336 3712 1352 3728
rect 1384 3712 1400 3728
rect 1416 3712 1448 3728
rect 1528 3712 1544 3728
rect 1576 3712 1608 3728
rect 1624 3712 1640 3728
rect 1752 3712 1768 3728
rect 1784 3712 1800 3728
rect 1896 3712 1928 3728
rect 2120 3712 2136 3728
rect 2200 3712 2216 3728
rect 1368 3692 1384 3708
rect 1560 3692 1576 3708
rect 1688 3692 1704 3708
rect 1752 3692 1768 3708
rect 1816 3692 1832 3708
rect 1992 3692 2008 3708
rect 2040 3692 2072 3708
rect 2152 3692 2168 3708
rect 2440 3692 2456 3708
rect 2488 3712 2504 3728
rect 2600 3712 2616 3728
rect 2632 3712 2648 3728
rect 2696 3712 2712 3728
rect 2776 3712 2792 3728
rect 2808 3712 2824 3728
rect 2872 3712 2888 3728
rect 2952 3712 2968 3728
rect 3016 3712 3048 3728
rect 3096 3712 3112 3728
rect 3128 3712 3144 3728
rect 3176 3712 3240 3728
rect 3320 3712 3336 3728
rect 3432 3712 3448 3728
rect 3592 3732 3608 3748
rect 3656 3732 3672 3748
rect 3768 3732 3784 3748
rect 4104 3732 4120 3748
rect 4152 3732 4168 3748
rect 4200 3732 4216 3748
rect 4424 3732 4456 3748
rect 4504 3732 4520 3748
rect 4568 3732 4584 3748
rect 4616 3732 4632 3748
rect 4664 3732 4696 3748
rect 5000 3732 5016 3748
rect 5096 3732 5112 3748
rect 5144 3732 5160 3748
rect 5224 3732 5240 3748
rect 5272 3732 5288 3748
rect 5320 3732 5336 3748
rect 5384 3732 5400 3748
rect 5480 3732 5496 3748
rect 5640 3732 5672 3748
rect 5768 3732 5784 3748
rect 5960 3732 5992 3748
rect 6104 3732 6120 3748
rect 6440 3732 6456 3748
rect 6520 3732 6552 3748
rect 6584 3732 6600 3748
rect 6696 3732 6712 3748
rect 6760 3732 6792 3748
rect 6840 3732 6856 3748
rect 7096 3732 7112 3748
rect 7256 3732 7272 3748
rect 7336 3732 7352 3748
rect 7368 3732 7384 3748
rect 7544 3732 7560 3748
rect 7592 3732 7608 3748
rect 7640 3732 7656 3748
rect 7688 3732 7704 3748
rect 7752 3732 7768 3748
rect 7800 3732 7816 3748
rect 2632 3692 2648 3708
rect 2728 3692 2744 3708
rect 2856 3692 2872 3708
rect 3044 3692 3060 3708
rect 3064 3692 3096 3708
rect 3400 3692 3416 3708
rect 3480 3692 3496 3708
rect 3512 3692 3528 3708
rect 3688 3692 3704 3708
rect 3720 3712 3752 3728
rect 3864 3712 3880 3728
rect 4072 3712 4088 3728
rect 4136 3692 4152 3708
rect 4184 3712 4200 3728
rect 4296 3712 4328 3728
rect 4472 3692 4488 3708
rect 4552 3692 4568 3708
rect 4600 3692 4616 3708
rect 4664 3712 4696 3728
rect 4840 3712 4856 3728
rect 5000 3712 5016 3728
rect 5176 3712 5192 3728
rect 4744 3692 4760 3708
rect 4968 3692 4984 3708
rect 5304 3692 5320 3708
rect 5352 3712 5368 3728
rect 5512 3712 5528 3728
rect 5576 3714 5592 3730
rect 5704 3712 5720 3728
rect 5736 3712 5752 3728
rect 5880 3712 5896 3728
rect 5992 3712 6008 3728
rect 5672 3692 5720 3708
rect 6104 3712 6120 3728
rect 6200 3712 6248 3728
rect 6328 3712 6344 3728
rect 6408 3712 6424 3728
rect 6472 3712 6488 3728
rect 6504 3712 6520 3728
rect 6552 3712 6568 3728
rect 6600 3712 6616 3728
rect 6792 3712 6808 3728
rect 6856 3712 6872 3728
rect 6936 3712 6952 3728
rect 7128 3712 7144 3728
rect 7176 3712 7192 3728
rect 7272 3712 7304 3728
rect 7448 3712 7464 3728
rect 7528 3712 7544 3728
rect 7656 3712 7672 3728
rect 6040 3692 6056 3708
rect 6612 3692 6628 3708
rect 6632 3692 6648 3708
rect 6664 3692 6680 3708
rect 6728 3692 6760 3708
rect 6824 3692 6840 3708
rect 6888 3692 6920 3708
rect 7368 3692 7384 3708
rect 7624 3692 7640 3708
rect 7736 3712 7752 3728
rect 7848 3712 7864 3728
rect 8040 3712 8056 3728
rect 7704 3692 7720 3708
rect 7928 3692 7944 3708
rect 2568 3672 2600 3688
rect 3160 3672 3176 3688
rect 3352 3672 3368 3688
rect 3544 3672 3560 3688
rect 1352 3652 1368 3668
rect 1544 3652 1560 3668
rect 1032 3632 1048 3648
rect 1480 3632 1496 3648
rect 2360 3632 2376 3648
rect 2904 3632 2920 3648
rect 5400 3632 5416 3648
rect 925 3602 961 3618
rect 2957 3602 2993 3618
rect 5021 3602 5057 3618
rect 7053 3602 7089 3618
rect 88 3572 104 3588
rect 296 3572 312 3588
rect 440 3572 456 3588
rect 584 3572 600 3588
rect 1560 3572 1576 3588
rect 1688 3572 1704 3588
rect 1736 3572 1752 3588
rect 1816 3572 1832 3588
rect 2120 3572 2136 3588
rect 2312 3572 2328 3588
rect 2808 3572 2824 3588
rect 2872 3572 2888 3588
rect 3096 3572 3112 3588
rect 3128 3572 3144 3588
rect 3272 3572 3288 3588
rect 3336 3572 3352 3588
rect 3400 3572 3416 3588
rect 3448 3572 3464 3588
rect 3560 3572 3576 3588
rect 3592 3572 3608 3588
rect 3832 3572 3848 3588
rect 3896 3572 3912 3588
rect 3976 3572 3992 3588
rect 4056 3572 4072 3588
rect 4696 3572 4712 3588
rect 5496 3572 5512 3588
rect 6504 3572 6520 3588
rect 6920 3572 6936 3588
rect 7160 3572 7176 3588
rect 7816 3572 7832 3588
rect 7880 3572 7896 3588
rect 200 3552 216 3568
rect 5128 3552 5144 3568
rect 8 3532 24 3548
rect 136 3532 152 3548
rect 328 3532 344 3548
rect 1704 3532 1736 3548
rect 1800 3532 1816 3548
rect 2104 3532 2120 3548
rect 2824 3532 2840 3548
rect 2888 3532 2904 3548
rect 3064 3532 3080 3548
rect 3144 3532 3160 3548
rect 3288 3532 3304 3548
rect 3336 3532 3352 3548
rect 3416 3532 3432 3548
rect 3464 3532 3480 3548
rect 3544 3532 3560 3548
rect 3608 3532 3624 3548
rect 6840 3532 6856 3548
rect 6904 3532 6920 3548
rect 7560 3532 7576 3548
rect 1108 3512 1124 3528
rect 40 3492 56 3508
rect 120 3492 136 3508
rect 184 3492 200 3508
rect 232 3492 248 3508
rect 264 3492 280 3508
rect 376 3492 408 3508
rect 536 3492 552 3508
rect 648 3492 664 3508
rect 696 3492 712 3508
rect 728 3492 744 3508
rect 1016 3490 1032 3506
rect 1096 3492 1112 3508
rect 1160 3512 1176 3528
rect 1704 3512 1720 3528
rect 1928 3512 1944 3528
rect 2136 3512 2152 3528
rect 2488 3512 2504 3528
rect 2520 3512 2536 3528
rect 2856 3512 2872 3528
rect 2920 3512 2936 3528
rect 3016 3512 3032 3528
rect 3048 3512 3064 3528
rect 3112 3512 3128 3528
rect 3224 3512 3240 3528
rect 3256 3512 3272 3528
rect 3320 3512 3336 3528
rect 3384 3512 3400 3528
rect 3496 3512 3528 3528
rect 3576 3512 3592 3528
rect 3688 3512 3704 3528
rect 3848 3512 3864 3528
rect 3912 3512 3928 3528
rect 4104 3512 4120 3528
rect 4500 3512 4516 3528
rect 4520 3512 4536 3528
rect 4664 3512 4680 3528
rect 4776 3512 4792 3528
rect 4968 3512 4984 3528
rect 1208 3492 1224 3508
rect 1304 3492 1320 3508
rect 1480 3492 1512 3508
rect 1640 3492 1656 3508
rect 1688 3492 1704 3508
rect 1736 3492 1768 3508
rect 1816 3492 1832 3508
rect 1960 3492 1976 3508
rect 2024 3490 2040 3506
rect 2120 3492 2136 3508
rect 2152 3492 2168 3508
rect 2184 3492 2200 3508
rect 2264 3492 2280 3508
rect 2360 3492 2376 3508
rect 2424 3492 2440 3508
rect 2504 3492 2520 3508
rect 456 3472 472 3488
rect 776 3472 792 3488
rect 808 3472 824 3488
rect 840 3472 856 3488
rect 968 3472 984 3488
rect 1000 3472 1016 3488
rect 1080 3472 1096 3488
rect 1192 3472 1208 3488
rect 1624 3472 1640 3488
rect 2184 3472 2200 3488
rect 2248 3472 2264 3488
rect 2280 3472 2296 3488
rect 2456 3472 2472 3488
rect 2552 3472 2568 3488
rect 2696 3492 2712 3508
rect 2840 3492 2856 3508
rect 2904 3492 2920 3508
rect 2984 3492 3000 3508
rect 3080 3492 3096 3508
rect 3128 3492 3144 3508
rect 3176 3492 3192 3508
rect 3272 3492 3288 3508
rect 3352 3492 3368 3508
rect 3416 3492 3432 3508
rect 3480 3492 3496 3508
rect 3528 3492 3544 3508
rect 3592 3492 3608 3508
rect 3656 3492 3672 3508
rect 3736 3492 3752 3508
rect 3912 3492 3928 3508
rect 4152 3492 4168 3508
rect 4184 3492 4200 3508
rect 4280 3490 4296 3506
rect 4488 3492 4504 3508
rect 4600 3492 4616 3508
rect 4872 3490 4888 3506
rect 5004 3512 5020 3528
rect 5320 3512 5336 3528
rect 5384 3512 5400 3528
rect 5960 3512 5976 3528
rect 5064 3492 5080 3508
rect 5096 3492 5112 3508
rect 5224 3492 5240 3508
rect 5256 3492 5272 3508
rect 5336 3492 5368 3508
rect 5416 3492 5432 3508
rect 5448 3492 5464 3508
rect 5544 3492 5560 3508
rect 5624 3492 5640 3508
rect 5752 3492 5768 3508
rect 5880 3492 5896 3508
rect 5992 3492 6008 3508
rect 6088 3512 6104 3528
rect 6424 3512 6440 3528
rect 6600 3512 6616 3528
rect 6200 3492 6216 3508
rect 6232 3492 6248 3508
rect 6312 3492 6328 3508
rect 6376 3492 6392 3508
rect 6472 3492 6504 3508
rect 6568 3492 6584 3508
rect 6648 3492 6664 3508
rect 6792 3492 6808 3508
rect 6952 3492 6968 3508
rect 7016 3512 7032 3528
rect 7252 3512 7268 3528
rect 7272 3512 7288 3528
rect 7336 3512 7352 3528
rect 7416 3512 7432 3528
rect 7480 3512 7496 3528
rect 7112 3492 7128 3508
rect 7144 3492 7160 3508
rect 7192 3492 7224 3508
rect 7288 3492 7304 3508
rect 7448 3492 7464 3508
rect 7516 3512 7532 3528
rect 7976 3512 7992 3528
rect 7528 3492 7544 3508
rect 7656 3492 7672 3508
rect 7784 3492 7800 3508
rect 7944 3492 7960 3508
rect 2792 3472 2808 3488
rect 3800 3472 3816 3488
rect 3880 3472 3896 3488
rect 4136 3472 4152 3488
rect 4216 3472 4232 3488
rect 4296 3472 4328 3488
rect 4376 3472 4392 3488
rect 4568 3472 4584 3488
rect 4632 3472 4648 3488
rect 4856 3472 4872 3488
rect 4936 3472 4952 3488
rect 5032 3472 5048 3488
rect 5368 3472 5384 3488
rect 5432 3472 5448 3488
rect 5656 3472 5688 3488
rect 5720 3472 5736 3488
rect 5800 3472 5816 3488
rect 5976 3472 5992 3488
rect 6024 3472 6040 3488
rect 6120 3472 6136 3488
rect 6296 3472 6312 3488
rect 6568 3472 6584 3488
rect 6632 3472 6648 3488
rect 6664 3472 6680 3488
rect 6712 3472 6728 3488
rect 6936 3472 6968 3488
rect 6984 3472 7000 3488
rect 7064 3472 7080 3488
rect 7224 3472 7240 3488
rect 7384 3472 7400 3488
rect 7432 3472 7448 3488
rect 7544 3472 7560 3488
rect 7672 3472 7688 3488
rect 1576 3452 1592 3468
rect 2152 3452 2168 3468
rect 2552 3452 2568 3468
rect 4072 3452 4088 3468
rect 4712 3452 4728 3468
rect 5384 3452 5400 3468
rect 6168 3452 6184 3468
rect 7400 3452 7416 3468
rect 88 3432 104 3448
rect 584 3432 600 3448
rect 664 3432 680 3448
rect 856 3432 872 3448
rect 1256 3432 1272 3448
rect 1336 3432 1352 3448
rect 1608 3432 1624 3448
rect 2392 3432 2408 3448
rect 2472 3432 2488 3448
rect 2664 3432 2680 3448
rect 2776 3432 2792 3448
rect 3768 3432 3784 3448
rect 4664 3432 4680 3448
rect 5192 3432 5208 3448
rect 5288 3432 5304 3448
rect 5496 3432 5512 3448
rect 5576 3432 5592 3448
rect 6344 3432 6360 3448
rect 1949 3402 1985 3418
rect 3997 3402 4033 3418
rect 6045 3402 6081 3418
rect 648 3372 664 3388
rect 1352 3372 1368 3388
rect 1400 3372 1416 3388
rect 1576 3372 1592 3388
rect 1656 3372 1672 3388
rect 1912 3372 1928 3388
rect 2024 3372 2040 3388
rect 2504 3372 2520 3388
rect 2600 3372 2616 3388
rect 2760 3372 2776 3388
rect 3080 3372 3096 3388
rect 3192 3372 3208 3388
rect 3256 3372 3272 3388
rect 3672 3372 3688 3388
rect 3848 3372 3864 3388
rect 4072 3372 4088 3388
rect 4248 3372 4264 3388
rect 5240 3372 5256 3388
rect 5640 3372 5656 3388
rect 5928 3372 5944 3388
rect 6360 3372 6376 3388
rect 6744 3372 6760 3388
rect 6984 3372 7000 3388
rect 7096 3372 7112 3388
rect 680 3352 696 3368
rect 824 3352 840 3368
rect 1064 3352 1080 3368
rect 1592 3352 1608 3368
rect 1672 3352 1688 3368
rect 2136 3352 2152 3368
rect 2680 3352 2696 3368
rect 2888 3352 2904 3368
rect 3432 3352 3448 3368
rect 5544 3352 5560 3368
rect 6952 3352 6968 3368
rect 7336 3352 7352 3368
rect 7480 3352 7496 3368
rect 7736 3352 7752 3368
rect 24 3332 40 3348
rect 104 3332 120 3348
rect 184 3332 200 3348
rect 744 3332 760 3348
rect 872 3332 888 3348
rect 936 3332 952 3348
rect 1000 3332 1016 3348
rect 1048 3332 1064 3348
rect 1080 3332 1096 3348
rect 1112 3332 1128 3348
rect 1288 3332 1304 3348
rect 2264 3332 2296 3348
rect 2376 3332 2408 3348
rect 2456 3332 2472 3348
rect 2520 3332 2536 3348
rect 2648 3332 2664 3348
rect 2728 3332 2744 3348
rect 72 3312 88 3328
rect 152 3312 168 3328
rect 200 3312 232 3328
rect 264 3312 280 3328
rect 312 3312 328 3328
rect 376 3312 392 3328
rect 456 3312 472 3328
rect 568 3312 584 3328
rect 632 3312 648 3328
rect 728 3312 744 3328
rect 792 3312 808 3328
rect 856 3312 872 3328
rect 904 3312 936 3328
rect 1016 3312 1032 3328
rect 1096 3312 1112 3328
rect 1160 3312 1176 3328
rect 1192 3312 1208 3328
rect 1256 3312 1272 3328
rect 1320 3312 1336 3328
rect 1384 3312 1400 3328
rect 1464 3312 1480 3328
rect 1512 3312 1528 3328
rect 1560 3312 1576 3328
rect 1624 3312 1640 3328
rect 1800 3312 1816 3328
rect 1992 3312 2008 3328
rect 2056 3312 2072 3328
rect 2184 3312 2200 3328
rect 2296 3312 2328 3328
rect 184 3272 200 3288
rect 248 3272 264 3288
rect 296 3292 312 3308
rect 360 3292 376 3308
rect 424 3292 440 3308
rect 696 3292 712 3308
rect 808 3292 824 3308
rect 888 3292 904 3308
rect 984 3292 1000 3308
rect 1240 3292 1256 3308
rect 1304 3292 1320 3308
rect 1368 3292 1384 3308
rect 1464 3292 1480 3308
rect 1624 3292 1640 3308
rect 2376 3312 2392 3328
rect 2424 3312 2440 3328
rect 2584 3312 2600 3328
rect 2616 3312 2632 3328
rect 2696 3312 2712 3328
rect 2808 3312 2824 3328
rect 3032 3332 3048 3348
rect 3128 3332 3144 3348
rect 3320 3332 3336 3348
rect 3416 3332 3432 3348
rect 3608 3332 3624 3348
rect 3960 3332 3976 3348
rect 4184 3332 4200 3348
rect 4232 3332 4248 3348
rect 4312 3332 4328 3348
rect 4472 3332 4488 3348
rect 4600 3332 4616 3348
rect 4680 3332 4696 3348
rect 4744 3332 4776 3348
rect 4808 3332 4824 3348
rect 4872 3332 4888 3348
rect 5064 3332 5080 3348
rect 5208 3332 5224 3348
rect 5352 3332 5368 3348
rect 5448 3332 5464 3348
rect 5496 3332 5512 3348
rect 5592 3332 5624 3348
rect 5688 3332 5704 3348
rect 5784 3332 5816 3348
rect 5848 3332 5864 3348
rect 5944 3332 5960 3348
rect 5976 3332 5992 3348
rect 6440 3332 6456 3348
rect 6504 3332 6520 3348
rect 7096 3332 7112 3348
rect 7128 3332 7144 3348
rect 7160 3332 7176 3348
rect 7256 3332 7272 3348
rect 7320 3332 7336 3348
rect 7544 3332 7560 3348
rect 7608 3332 7624 3348
rect 7656 3332 7672 3348
rect 7880 3332 7896 3348
rect 7912 3332 7928 3348
rect 7992 3332 8008 3348
rect 2936 3312 2952 3328
rect 2344 3292 2360 3308
rect 2440 3292 2456 3308
rect 2504 3292 2520 3308
rect 2712 3292 2728 3308
rect 2792 3292 2808 3308
rect 2968 3292 2984 3308
rect 3064 3292 3080 3308
rect 3112 3312 3128 3328
rect 3160 3312 3176 3328
rect 3288 3312 3304 3328
rect 3352 3292 3368 3308
rect 3432 3312 3448 3328
rect 3544 3312 3560 3328
rect 3736 3312 3752 3328
rect 3784 3312 3800 3328
rect 3816 3312 3832 3328
rect 3992 3312 4008 3328
rect 3388 3292 3404 3308
rect 4168 3292 4184 3308
rect 4216 3312 4232 3328
rect 4296 3312 4312 3328
rect 4344 3312 4360 3328
rect 4568 3314 4584 3330
rect 4696 3312 4712 3328
rect 4744 3312 4760 3328
rect 4776 3312 4792 3328
rect 4312 3292 4328 3308
rect 4648 3292 4664 3308
rect 4984 3312 5000 3328
rect 5224 3312 5240 3328
rect 5400 3312 5416 3328
rect 4840 3292 4856 3308
rect 5320 3292 5336 3308
rect 5528 3292 5544 3308
rect 5576 3312 5592 3328
rect 5688 3292 5704 3308
rect 5720 3292 5736 3308
rect 5768 3312 5784 3328
rect 5756 3292 5772 3308
rect 6120 3312 6136 3328
rect 6312 3312 6344 3328
rect 6408 3312 6424 3328
rect 5864 3292 5880 3308
rect 5944 3292 5960 3308
rect 5992 3292 6008 3308
rect 6600 3312 6632 3328
rect 6808 3312 6824 3328
rect 6840 3312 6856 3328
rect 6472 3292 6488 3308
rect 7000 3292 7016 3308
rect 7032 3292 7048 3308
rect 7096 3292 7112 3308
rect 7192 3292 7208 3308
rect 7240 3312 7256 3328
rect 7304 3312 7320 3328
rect 7432 3312 7448 3328
rect 7560 3312 7576 3328
rect 7228 3292 7244 3308
rect 7272 3292 7288 3308
rect 7752 3312 7768 3328
rect 7880 3312 7896 3328
rect 7624 3292 7640 3308
rect 7832 3292 7848 3308
rect 7960 3292 7976 3308
rect 328 3272 344 3288
rect 392 3272 408 3288
rect 456 3272 472 3288
rect 776 3272 792 3288
rect 520 3252 536 3268
rect 1192 3272 1208 3288
rect 1272 3272 1288 3288
rect 1336 3272 1352 3288
rect 1400 3272 1416 3288
rect 1448 3272 1464 3288
rect 1528 3272 1544 3288
rect 1640 3272 1656 3288
rect 2600 3272 2616 3288
rect 2680 3272 2696 3288
rect 2792 3272 2808 3288
rect 2824 3272 2840 3288
rect 2936 3272 2952 3288
rect 3848 3272 3864 3288
rect 6072 3272 6088 3288
rect 6952 3272 6968 3288
rect 1224 3252 1240 3268
rect 1464 3252 1480 3268
rect 40 3232 56 3248
rect 264 3232 280 3248
rect 376 3232 392 3248
rect 440 3232 456 3248
rect 1544 3232 1560 3248
rect 1912 3232 1928 3248
rect 3672 3232 3688 3248
rect 3752 3232 3768 3248
rect 5160 3232 5176 3248
rect 7304 3232 7320 3248
rect 925 3202 961 3218
rect 2957 3202 2993 3218
rect 5021 3202 5057 3218
rect 7053 3202 7089 3218
rect 152 3172 168 3188
rect 456 3172 472 3188
rect 488 3172 504 3188
rect 568 3172 584 3188
rect 664 3172 680 3188
rect 728 3172 744 3188
rect 808 3172 824 3188
rect 888 3172 904 3188
rect 1256 3172 1272 3188
rect 1304 3172 1320 3188
rect 1352 3172 1368 3188
rect 1432 3172 1448 3188
rect 1592 3172 1608 3188
rect 1624 3172 1640 3188
rect 1688 3172 1704 3188
rect 2136 3172 2152 3188
rect 2504 3172 2520 3188
rect 2584 3172 2600 3188
rect 2648 3172 2664 3188
rect 2792 3172 2808 3188
rect 3048 3172 3064 3188
rect 3112 3172 3144 3188
rect 3624 3172 3640 3188
rect 4712 3172 4728 3188
rect 4920 3172 4936 3188
rect 5000 3172 5016 3188
rect 5128 3172 5144 3188
rect 5336 3172 5352 3188
rect 5432 3172 5448 3188
rect 5688 3172 5704 3188
rect 6088 3172 6104 3188
rect 6424 3172 6440 3188
rect 6568 3172 6584 3188
rect 6664 3172 6680 3188
rect 6728 3172 6744 3188
rect 6920 3172 6936 3188
rect 6984 3172 7000 3188
rect 7080 3172 7096 3188
rect 7128 3172 7144 3188
rect 7912 3172 7928 3188
rect 7976 3172 7992 3188
rect 136 3132 152 3148
rect 424 3132 440 3148
rect 648 3132 664 3148
rect 792 3132 808 3148
rect 872 3132 888 3148
rect 1240 3132 1256 3148
rect 1320 3132 1336 3148
rect 1368 3132 1384 3148
rect 1448 3132 1464 3148
rect 1496 3132 1512 3148
rect 1736 3152 1752 3168
rect 168 3112 184 3128
rect 392 3112 408 3128
rect 696 3112 712 3128
rect 824 3112 856 3128
rect 1144 3112 1160 3128
rect 1272 3112 1288 3128
rect 1416 3112 1432 3128
rect 1528 3112 1544 3128
rect 1576 3132 1592 3148
rect 1640 3132 1656 3148
rect 1704 3132 1720 3148
rect 2520 3132 2536 3148
rect 2568 3132 2584 3148
rect 2632 3132 2648 3148
rect 2776 3132 2792 3148
rect 5512 3132 5528 3148
rect 6328 3132 6344 3148
rect 7560 3132 7576 3148
rect 7752 3132 7768 3148
rect 7880 3132 7896 3148
rect 1608 3112 1624 3128
rect 1672 3112 1688 3128
rect 2104 3112 2120 3128
rect 2392 3112 2408 3128
rect 2472 3112 2504 3128
rect 2600 3112 2616 3128
rect 2648 3112 2664 3128
rect 2824 3112 2840 3128
rect 3064 3112 3080 3128
rect 3224 3112 3240 3128
rect 3400 3112 3416 3128
rect 3496 3112 3512 3128
rect 72 3092 88 3108
rect 152 3092 168 3108
rect 280 3092 296 3108
rect 312 3092 328 3108
rect 408 3092 424 3108
rect 520 3092 536 3108
rect 664 3092 680 3108
rect 760 3092 776 3108
rect 808 3092 824 3108
rect 856 3092 872 3108
rect 1032 3092 1048 3108
rect 1144 3092 1160 3108
rect 1208 3092 1224 3108
rect 1256 3092 1272 3108
rect 1304 3092 1320 3108
rect 1384 3092 1400 3108
rect 1432 3092 1448 3108
rect 1512 3092 1528 3108
rect 1560 3092 1576 3108
rect 1624 3092 1640 3108
rect 1688 3092 1704 3108
rect 1864 3092 1880 3108
rect 2008 3092 2024 3108
rect 2040 3092 2056 3108
rect 2088 3092 2104 3108
rect 2296 3092 2312 3108
rect 2408 3092 2440 3108
rect 2456 3092 2472 3108
rect 2504 3092 2520 3108
rect 2584 3092 2600 3108
rect 2648 3092 2664 3108
rect 2744 3092 2760 3108
rect 2792 3092 2808 3108
rect 2888 3092 2904 3108
rect 2920 3092 2936 3108
rect 3112 3092 3128 3108
rect 3336 3092 3352 3108
rect 3736 3112 3752 3128
rect 3944 3112 3960 3128
rect 3544 3092 3560 3108
rect 3832 3090 3848 3106
rect 4104 3112 4136 3128
rect 4260 3112 4276 3128
rect 3976 3092 3992 3108
rect 4040 3092 4056 3108
rect 4136 3092 4168 3108
rect 4248 3092 4264 3108
rect 4312 3112 4328 3128
rect 4664 3112 4696 3128
rect 4744 3112 4760 3128
rect 5160 3112 5176 3128
rect 5320 3112 5336 3128
rect 6040 3112 6056 3128
rect 6136 3112 6152 3128
rect 6184 3112 6200 3128
rect 6504 3112 6520 3128
rect 6648 3112 6664 3128
rect 6744 3112 6760 3128
rect 6792 3112 6808 3128
rect 6952 3112 6968 3128
rect 7144 3112 7160 3128
rect 7624 3112 7640 3128
rect 7688 3112 7704 3128
rect 7800 3112 7816 3128
rect 7864 3112 7880 3128
rect 4424 3090 4440 3106
rect 4488 3092 4504 3108
rect 4632 3092 4648 3108
rect 24 3072 40 3088
rect 88 3072 104 3088
rect 360 3072 376 3088
rect 536 3072 552 3088
rect 584 3072 600 3088
rect 904 3072 920 3088
rect 968 3072 984 3088
rect 1208 3072 1224 3088
rect 1784 3072 1800 3088
rect 1912 3072 1928 3088
rect 2088 3072 2104 3088
rect 2168 3072 2184 3088
rect 2344 3072 2360 3088
rect 2408 3072 2424 3088
rect 2824 3072 2840 3088
rect 3032 3072 3048 3088
rect 3192 3072 3208 3088
rect 3272 3072 3288 3088
rect 3512 3072 3528 3088
rect 3560 3072 3576 3088
rect 3640 3072 3656 3088
rect 3864 3072 3880 3088
rect 3912 3072 3928 3088
rect 4008 3072 4024 3088
rect 4072 3072 4088 3088
rect 4232 3072 4248 3088
rect 4344 3072 4376 3088
rect 4728 3072 4744 3088
rect 4792 3072 4808 3088
rect 4824 3092 4840 3108
rect 4872 3092 4888 3108
rect 4984 3092 5000 3108
rect 5032 3092 5048 3108
rect 5096 3092 5112 3108
rect 5208 3092 5224 3108
rect 5256 3092 5272 3108
rect 5384 3092 5416 3108
rect 5576 3092 5592 3108
rect 5768 3092 5784 3108
rect 5928 3092 5944 3108
rect 6008 3092 6024 3108
rect 6456 3092 6472 3108
rect 6536 3092 6552 3108
rect 6632 3092 6648 3108
rect 6888 3092 6904 3108
rect 5304 3072 5320 3088
rect 5352 3072 5368 3088
rect 5640 3072 5656 3088
rect 5848 3072 5864 3088
rect 5944 3072 5960 3088
rect 5976 3072 5992 3088
rect 6168 3072 6184 3088
rect 6328 3072 6344 3088
rect 6392 3072 6408 3088
rect 6472 3072 6488 3088
rect 6616 3076 6632 3092
rect 7304 3090 7320 3106
rect 7480 3092 7496 3108
rect 7592 3092 7640 3108
rect 7672 3092 7688 3108
rect 7832 3092 7848 3108
rect 7896 3092 7912 3108
rect 7928 3092 7944 3108
rect 6680 3072 6712 3088
rect 6760 3072 6776 3088
rect 6840 3072 6856 3088
rect 6872 3072 6888 3088
rect 7016 3072 7032 3088
rect 7112 3072 7128 3088
rect 7144 3072 7160 3088
rect 7240 3072 7256 3088
rect 7448 3072 7464 3088
rect 7576 3072 7592 3088
rect 7640 3072 7656 3088
rect 7784 3072 7800 3088
rect 7848 3072 7864 3088
rect 40 3052 56 3068
rect 104 3052 120 3068
rect 1160 3052 1176 3068
rect 1976 3052 1992 3068
rect 2376 3052 2392 3068
rect 3080 3052 3096 3068
rect 3160 3052 3176 3068
rect 3576 3052 3592 3068
rect 4200 3052 4216 3068
rect 4488 3052 4504 3068
rect 5272 3052 5288 3068
rect 5368 3052 5384 3068
rect 6264 3052 6280 3068
rect 6376 3052 6392 3068
rect 6520 3052 6536 3068
rect 6552 3052 6568 3068
rect 7032 3052 7048 3068
rect 7704 3052 7720 3068
rect 728 3032 744 3048
rect 2168 3032 2184 3048
rect 2712 3032 2728 3048
rect 2952 3032 2968 3048
rect 3208 3032 3224 3048
rect 3656 3032 3672 3048
rect 4104 3032 4120 3048
rect 4664 3032 4680 3048
rect 4744 3032 4760 3048
rect 5128 3032 5144 3048
rect 5464 3032 5480 3048
rect 5880 3032 5896 3048
rect 6088 3032 6104 3048
rect 6120 3032 6136 3048
rect 6184 3032 6200 3048
rect 6280 3032 6296 3048
rect 6664 3032 6680 3048
rect 6808 3032 6824 3048
rect 6920 3032 6936 3048
rect 7720 3032 7736 3048
rect 7800 3032 7816 3048
rect 7896 3032 7912 3048
rect 1949 3002 1985 3018
rect 3997 3002 4033 3018
rect 6045 3002 6081 3018
rect 72 2972 88 2988
rect 280 2972 296 2988
rect 424 2972 440 2988
rect 712 2972 728 2988
rect 1144 2972 1160 2988
rect 1560 2972 1576 2988
rect 1656 2972 1672 2988
rect 1720 2972 1736 2988
rect 2024 2972 2040 2988
rect 2120 2972 2136 2988
rect 2280 2972 2296 2988
rect 2392 2972 2408 2988
rect 2456 2972 2472 2988
rect 2808 2972 2824 2988
rect 2968 2972 2984 2988
rect 3800 2972 3816 2988
rect 4120 2972 4136 2988
rect 4712 2972 4744 2988
rect 4968 2972 4984 2988
rect 5112 2972 5128 2988
rect 5512 2972 5528 2988
rect 5784 2972 5800 2988
rect 5864 2972 5880 2988
rect 5928 2972 5944 2988
rect 6040 2972 6056 2988
rect 6136 2972 6152 2988
rect 6648 2972 6664 2988
rect 6968 2972 6984 2988
rect 8024 2972 8040 2988
rect 24 2952 40 2968
rect 120 2952 136 2968
rect 168 2952 216 2968
rect 440 2952 456 2968
rect 664 2952 680 2968
rect 776 2952 792 2968
rect 824 2952 840 2968
rect 296 2932 312 2948
rect 344 2932 360 2948
rect 552 2932 568 2948
rect 696 2932 712 2948
rect 1080 2952 1096 2968
rect 1160 2952 1176 2968
rect 1192 2952 1208 2968
rect 1320 2952 1336 2968
rect 1400 2952 1416 2968
rect 1464 2952 1480 2968
rect 1768 2952 1784 2968
rect 1864 2952 1880 2968
rect 1896 2952 1912 2968
rect 2072 2952 2088 2968
rect 888 2932 904 2948
rect 1016 2932 1032 2948
rect 1240 2932 1256 2948
rect 1912 2932 1928 2948
rect 2184 2952 2200 2968
rect 2728 2952 2744 2968
rect 3160 2952 3176 2968
rect 3256 2952 3272 2968
rect 5192 2952 5208 2968
rect 5224 2952 5240 2968
rect 5272 2952 5288 2968
rect 5368 2952 5384 2968
rect 6152 2952 6168 2968
rect 6232 2952 6248 2968
rect 6520 2952 6536 2968
rect 6712 2952 6728 2968
rect 8008 2952 8024 2968
rect 2136 2932 2152 2948
rect 2232 2932 2248 2948
rect 2536 2932 2552 2948
rect 2840 2932 2856 2948
rect 2888 2932 2904 2948
rect 2968 2932 2984 2948
rect 3032 2932 3048 2948
rect 3368 2932 3384 2948
rect 3432 2932 3464 2948
rect 3592 2932 3624 2948
rect 3816 2932 3832 2948
rect 3896 2932 3912 2948
rect 3928 2932 3944 2948
rect 3960 2932 3976 2948
rect 4040 2932 4056 2948
rect 4296 2932 4312 2948
rect 4328 2932 4344 2948
rect 4408 2932 4424 2948
rect 4440 2932 4456 2948
rect 4552 2932 4568 2948
rect 4680 2932 4696 2948
rect 4872 2932 4888 2948
rect 4936 2932 4952 2948
rect 5144 2932 5160 2948
rect 5176 2932 5192 2948
rect 5464 2932 5480 2948
rect 5560 2932 5576 2948
rect 5608 2932 5624 2948
rect 5832 2932 5848 2948
rect 5976 2932 5992 2948
rect 6104 2932 6120 2948
rect 6296 2932 6312 2948
rect 6456 2932 6472 2948
rect 6536 2932 6552 2948
rect 6632 2932 6648 2948
rect 6696 2932 6712 2948
rect 6888 2932 6904 2948
rect 7000 2932 7016 2948
rect 7064 2932 7080 2948
rect 7304 2932 7320 2948
rect 7352 2932 7368 2948
rect 7448 2932 7464 2948
rect 7576 2932 7592 2948
rect 7608 2932 7624 2948
rect 7656 2932 7672 2948
rect 7768 2932 7784 2948
rect 232 2912 248 2928
rect 344 2912 360 2928
rect 392 2912 424 2928
rect 536 2912 552 2928
rect 680 2912 696 2928
rect 744 2912 760 2928
rect 792 2912 808 2928
rect 872 2912 888 2928
rect 920 2912 936 2928
rect 1032 2912 1048 2928
rect 1160 2912 1176 2928
rect 1224 2912 1240 2928
rect 1272 2912 1304 2928
rect 1400 2914 1416 2930
rect 1576 2912 1592 2928
rect 1624 2912 1640 2928
rect 1752 2912 1768 2928
rect 1784 2912 1800 2928
rect 1880 2912 1896 2928
rect 1912 2912 1928 2928
rect 1992 2912 2008 2928
rect 2040 2912 2056 2928
rect 2152 2912 2168 2928
rect 2200 2912 2216 2928
rect 2328 2912 2344 2928
rect 2424 2912 2440 2928
rect 2472 2912 2488 2928
rect 2616 2912 2648 2928
rect 2776 2912 2792 2928
rect 1592 2892 1608 2908
rect 1864 2892 1880 2908
rect 2200 2892 2216 2908
rect 2296 2892 2312 2908
rect 2472 2892 2488 2908
rect 2824 2892 2840 2908
rect 2872 2892 2888 2908
rect 2920 2912 2936 2928
rect 3064 2912 3080 2928
rect 3192 2912 3208 2928
rect 3256 2914 3272 2930
rect 3336 2912 3368 2928
rect 3400 2912 3432 2928
rect 3528 2912 3560 2928
rect 3720 2912 3752 2928
rect 3832 2912 3864 2928
rect 4056 2912 4072 2928
rect 4264 2914 4280 2930
rect 4344 2912 4376 2928
rect 4568 2912 4584 2928
rect 4776 2912 4792 2928
rect 4808 2912 4824 2928
rect 5064 2912 5080 2928
rect 2984 2892 3000 2908
rect 3048 2892 3064 2908
rect 3112 2892 3128 2908
rect 3320 2892 3336 2908
rect 3384 2892 3400 2908
rect 3928 2892 3944 2908
rect 4168 2892 4184 2908
rect 4456 2892 4472 2908
rect 4712 2892 4728 2908
rect 5208 2912 5224 2928
rect 5256 2912 5272 2928
rect 5304 2912 5336 2928
rect 5416 2912 5432 2928
rect 5464 2912 5480 2928
rect 4936 2892 4952 2908
rect 4968 2892 4984 2908
rect 5112 2892 5128 2908
rect 5208 2892 5224 2908
rect 5288 2892 5304 2908
rect 5336 2892 5352 2908
rect 5496 2892 5512 2908
rect 5544 2912 5560 2928
rect 5640 2914 5656 2930
rect 5896 2912 5912 2928
rect 5928 2912 5944 2928
rect 6200 2912 6216 2928
rect 5736 2892 5752 2908
rect 5800 2892 5816 2908
rect 5944 2892 5960 2908
rect 6136 2892 6152 2908
rect 6168 2892 6184 2908
rect 6216 2892 6232 2908
rect 6408 2912 6424 2928
rect 6712 2912 6728 2928
rect 6808 2912 6824 2928
rect 6936 2912 6952 2928
rect 7000 2912 7016 2928
rect 7064 2912 7080 2928
rect 7160 2914 7176 2930
rect 7224 2912 7240 2928
rect 7336 2912 7352 2928
rect 7496 2912 7512 2928
rect 7640 2912 7656 2928
rect 7672 2912 7688 2928
rect 6312 2892 6328 2908
rect 6600 2892 6616 2908
rect 7048 2892 7064 2908
rect 7416 2892 7432 2908
rect 7704 2892 7720 2908
rect 7736 2912 7768 2928
rect 7864 2912 7896 2928
rect 1576 2872 1592 2888
rect 2184 2872 2200 2888
rect 2328 2872 2344 2888
rect 2456 2872 2472 2888
rect 6296 2872 6312 2888
rect 7304 2872 7320 2888
rect 7784 2872 7800 2888
rect 5368 2852 5384 2868
rect 56 2832 72 2848
rect 360 2832 376 2848
rect 1656 2832 1672 2848
rect 1720 2832 1736 2848
rect 2024 2832 2040 2848
rect 4824 2832 4840 2848
rect 4888 2832 4904 2848
rect 4984 2832 5000 2848
rect 5192 2832 5208 2848
rect 5816 2832 5832 2848
rect 5960 2832 5976 2848
rect 6040 2832 6056 2848
rect 6568 2832 6584 2848
rect 6728 2832 6744 2848
rect 6968 2832 6984 2848
rect 925 2802 961 2818
rect 2957 2802 2993 2818
rect 5021 2802 5057 2818
rect 7053 2802 7089 2818
rect 296 2772 312 2788
rect 792 2772 808 2788
rect 1768 2772 1784 2788
rect 3048 2772 3064 2788
rect 4408 2772 4424 2788
rect 7320 2772 7336 2788
rect 7816 2772 7832 2788
rect 2056 2732 2072 2748
rect 2120 2732 2136 2748
rect 2184 2732 2200 2748
rect 2312 2732 2328 2748
rect 2392 2732 2408 2748
rect 3384 2732 3400 2748
rect 6696 2732 6712 2748
rect 712 2712 728 2728
rect 2088 2712 2104 2728
rect 2152 2712 2168 2728
rect 2280 2712 2296 2728
rect 2600 2712 2616 2728
rect 152 2690 168 2706
rect 248 2692 264 2708
rect 328 2692 344 2708
rect 472 2692 488 2708
rect 616 2690 632 2706
rect 680 2692 696 2708
rect 824 2692 856 2708
rect 968 2692 984 2708
rect 1048 2692 1064 2708
rect 1128 2692 1144 2708
rect 1320 2692 1336 2708
rect 1432 2692 1448 2708
rect 1512 2692 1528 2708
rect 1672 2690 1688 2706
rect 1800 2692 1816 2708
rect 1832 2692 1848 2708
rect 1960 2692 1976 2708
rect 2024 2692 2040 2708
rect 2104 2692 2120 2708
rect 2168 2692 2184 2708
rect 2296 2692 2312 2708
rect 2488 2690 2504 2706
rect 2936 2712 2952 2728
rect 2632 2692 2664 2708
rect 2824 2690 2840 2706
rect 3004 2712 3020 2728
rect 3144 2712 3160 2728
rect 3416 2712 3448 2728
rect 3496 2712 3512 2728
rect 3544 2712 3576 2728
rect 3672 2712 3688 2728
rect 3016 2692 3032 2708
rect 3304 2690 3320 2706
rect 3448 2692 3464 2708
rect 3512 2692 3528 2708
rect 3576 2692 3608 2708
rect 3752 2712 3768 2728
rect 4008 2712 4024 2728
rect 4104 2712 4120 2728
rect 4664 2712 4680 2728
rect 3752 2692 3768 2708
rect 3848 2692 3864 2708
rect 3976 2692 3992 2708
rect 4072 2692 4088 2708
rect 4216 2692 4232 2708
rect 4392 2692 4408 2708
rect 4552 2690 4568 2706
rect 4776 2712 4792 2728
rect 4872 2712 4888 2728
rect 4744 2692 4760 2708
rect 4824 2692 4840 2708
rect 5448 2712 5464 2728
rect 4904 2692 4920 2708
rect 4936 2692 4968 2708
rect 5080 2692 5096 2708
rect 5336 2690 5352 2706
rect 5544 2692 5576 2708
rect 5608 2712 5624 2728
rect 6152 2712 6168 2728
rect 6216 2712 6232 2728
rect 6248 2712 6280 2728
rect 6328 2712 6344 2728
rect 5768 2692 5800 2708
rect 5848 2692 5864 2708
rect 5880 2692 5896 2708
rect 5944 2692 5960 2708
rect 5992 2692 6008 2708
rect 6040 2692 6072 2708
rect 6120 2692 6136 2708
rect 6184 2692 6216 2708
rect 6360 2692 6376 2708
rect 6392 2692 6408 2708
rect 6424 2692 6440 2708
rect 6488 2712 6504 2728
rect 6888 2712 6904 2728
rect 7172 2712 7188 2728
rect 6552 2692 6584 2708
rect 6792 2690 6808 2706
rect 7016 2692 7048 2708
rect 7160 2692 7176 2708
rect 7208 2712 7224 2728
rect 7416 2712 7432 2728
rect 7448 2712 7464 2728
rect 7480 2712 7496 2728
rect 7592 2712 7608 2728
rect 7288 2692 7304 2708
rect 7448 2692 7464 2708
rect 7496 2692 7528 2708
rect 7704 2692 7720 2708
rect 7912 2692 7928 2708
rect 184 2672 200 2688
rect 264 2672 280 2688
rect 520 2672 536 2688
rect 552 2672 568 2688
rect 920 2672 936 2688
rect 1016 2672 1032 2688
rect 1112 2672 1128 2688
rect 1240 2672 1256 2688
rect 1368 2672 1384 2688
rect 1496 2672 1512 2688
rect 1560 2672 1576 2688
rect 1640 2672 1656 2688
rect 2264 2672 2280 2688
rect 2520 2672 2536 2688
rect 2568 2672 2584 2688
rect 2664 2672 2680 2688
rect 2808 2672 2824 2688
rect 2904 2672 2920 2688
rect 3032 2672 3048 2688
rect 3112 2672 3128 2688
rect 3144 2672 3160 2688
rect 3272 2672 3288 2688
rect 3384 2672 3400 2688
rect 3496 2672 3528 2688
rect 3624 2672 3656 2688
rect 3704 2672 3720 2688
rect 3736 2672 3752 2688
rect 3832 2672 3848 2688
rect 3864 2672 3880 2688
rect 3976 2672 3992 2688
rect 4056 2672 4072 2688
rect 4120 2672 4136 2688
rect 4296 2672 4312 2688
rect 4328 2672 4344 2688
rect 4456 2672 4472 2688
rect 4584 2672 4600 2688
rect 4632 2672 4648 2688
rect 4664 2672 4680 2688
rect 4760 2672 4776 2688
rect 4840 2672 4856 2688
rect 4984 2672 5000 2688
rect 5064 2672 5080 2688
rect 5160 2672 5176 2688
rect 5272 2672 5288 2688
rect 5416 2672 5432 2688
rect 5448 2672 5464 2688
rect 5512 2672 5544 2688
rect 5640 2672 5656 2688
rect 5816 2672 5832 2688
rect 5896 2672 5928 2688
rect 5944 2672 5960 2688
rect 6104 2672 6120 2688
rect 6136 2672 6152 2688
rect 6168 2672 6184 2688
rect 6280 2672 6312 2688
rect 6392 2672 6424 2688
rect 6520 2672 6536 2688
rect 6696 2672 6712 2688
rect 6824 2672 6840 2688
rect 6856 2672 6872 2688
rect 7128 2672 7160 2688
rect 7256 2672 7272 2688
rect 7352 2672 7368 2688
rect 7464 2672 7480 2688
rect 7544 2672 7576 2688
rect 7784 2672 7800 2688
rect 7992 2672 8008 2688
rect 88 2652 104 2668
rect 216 2652 232 2668
rect 680 2652 696 2668
rect 1400 2652 1416 2668
rect 1480 2652 1496 2668
rect 1864 2652 1880 2668
rect 2312 2652 2328 2668
rect 2392 2652 2408 2668
rect 2760 2652 2776 2668
rect 3080 2652 3096 2668
rect 5240 2652 5256 2668
rect 5336 2652 5352 2668
rect 5752 2652 5768 2668
rect 5816 2652 5832 2668
rect 5912 2652 5928 2668
rect 6584 2652 6600 2668
rect 7688 2652 7704 2668
rect 232 2632 248 2648
rect 344 2632 360 2648
rect 1160 2632 1176 2648
rect 1192 2632 1208 2648
rect 1928 2632 1944 2648
rect 2056 2632 2072 2648
rect 2120 2632 2136 2648
rect 2232 2632 2248 2648
rect 3144 2632 3160 2648
rect 4136 2632 4152 2648
rect 5704 2632 5720 2648
rect 5880 2632 5896 2648
rect 6472 2632 6488 2648
rect 6872 2632 6888 2648
rect 7400 2632 7416 2648
rect 7592 2632 7608 2648
rect 1949 2602 1985 2618
rect 3997 2602 4033 2618
rect 6045 2602 6081 2618
rect 40 2572 56 2588
rect 120 2572 136 2588
rect 216 2572 232 2588
rect 328 2572 344 2588
rect 504 2572 520 2588
rect 632 2572 648 2588
rect 696 2572 712 2588
rect 1272 2572 1288 2588
rect 1720 2572 1736 2588
rect 2632 2572 2648 2588
rect 3640 2572 3656 2588
rect 3896 2572 3912 2588
rect 4104 2572 4120 2588
rect 4280 2572 4296 2588
rect 5000 2572 5016 2588
rect 5384 2572 5400 2588
rect 6088 2572 6104 2588
rect 6456 2572 6472 2588
rect 6680 2572 6696 2588
rect 6888 2572 6904 2588
rect 7480 2572 7496 2588
rect 7576 2572 7592 2588
rect 7672 2572 7688 2588
rect 232 2552 248 2568
rect 280 2552 296 2568
rect 200 2532 216 2548
rect 568 2552 584 2568
rect 1304 2552 1320 2568
rect 1368 2552 1384 2568
rect 1640 2552 1656 2568
rect 1912 2552 1928 2568
rect 1944 2552 1960 2568
rect 2152 2552 2168 2568
rect 2360 2552 2376 2568
rect 2440 2552 2456 2568
rect 2936 2552 2952 2568
rect 3672 2552 3688 2568
rect 3720 2552 3736 2568
rect 3992 2552 4008 2568
rect 5896 2552 5912 2568
rect 6360 2552 6376 2568
rect 7448 2552 7464 2568
rect 7784 2552 7800 2568
rect 360 2532 376 2548
rect 488 2532 504 2548
rect 1304 2532 1336 2548
rect 1448 2532 1464 2548
rect 1480 2532 1496 2548
rect 1736 2532 1752 2548
rect 2040 2532 2056 2548
rect 2232 2532 2248 2548
rect 2280 2532 2296 2548
rect 2408 2532 2440 2548
rect 2504 2532 2520 2548
rect 2552 2532 2568 2548
rect 2728 2532 2744 2548
rect 2792 2532 2824 2548
rect 3256 2532 3288 2548
rect 3384 2532 3400 2548
rect 3416 2532 3432 2548
rect 3448 2532 3464 2548
rect 3496 2532 3512 2548
rect 3544 2532 3560 2548
rect 3784 2532 3800 2548
rect 3880 2532 3896 2548
rect 4056 2532 4072 2548
rect 4136 2532 4152 2548
rect 4168 2532 4184 2548
rect 4232 2532 4248 2548
rect 4264 2532 4280 2548
rect 4424 2532 4440 2548
rect 4536 2532 4552 2548
rect 4584 2532 4600 2548
rect 4616 2532 4632 2548
rect 4712 2532 4728 2548
rect 4744 2532 4760 2548
rect 4808 2532 4824 2548
rect 4840 2532 4856 2548
rect 4936 2532 4952 2548
rect 5112 2532 5128 2548
rect 5496 2532 5512 2548
rect 5608 2532 5640 2548
rect 5720 2532 5736 2548
rect 5816 2532 5832 2548
rect 6264 2532 6280 2548
rect 6296 2532 6312 2548
rect 6408 2532 6440 2548
rect 6520 2532 6536 2548
rect 6744 2532 6760 2548
rect 6936 2532 6968 2548
rect 7048 2532 7080 2548
rect 7224 2532 7240 2548
rect 7352 2532 7368 2548
rect 7528 2532 7544 2548
rect 7624 2532 7640 2548
rect 7864 2532 7880 2548
rect 72 2512 88 2528
rect 168 2512 200 2528
rect 248 2512 264 2528
rect 360 2512 376 2528
rect 440 2512 472 2528
rect 536 2512 552 2528
rect 600 2512 616 2528
rect 744 2512 776 2528
rect 856 2512 872 2528
rect 920 2512 936 2528
rect 1000 2512 1016 2528
rect 1064 2512 1080 2528
rect 1176 2512 1192 2528
rect 1256 2512 1272 2528
rect 1336 2512 1352 2528
rect 1416 2512 1432 2528
rect 1464 2512 1480 2528
rect 1544 2512 1560 2528
rect 1608 2512 1624 2528
rect 1640 2512 1656 2528
rect 1672 2512 1688 2528
rect 1752 2512 1768 2528
rect 1832 2512 1848 2528
rect 1880 2512 1896 2528
rect 1928 2512 1944 2528
rect 2008 2512 2024 2528
rect 2088 2512 2104 2528
rect 2120 2512 2136 2528
rect 2200 2512 2216 2528
rect 2264 2512 2280 2528
rect 2312 2512 2328 2528
rect 2392 2512 2408 2528
rect 2488 2512 2504 2528
rect 2664 2512 2680 2528
rect 2760 2512 2792 2528
rect 2872 2514 2888 2530
rect 2936 2512 2952 2528
rect 3096 2512 3112 2528
rect 3272 2512 3288 2528
rect 792 2492 808 2508
rect 872 2492 888 2508
rect 968 2492 984 2508
rect 840 2472 856 2488
rect 904 2472 920 2488
rect 1032 2492 1064 2508
rect 1432 2492 1448 2508
rect 1560 2492 1576 2508
rect 1624 2492 1640 2508
rect 1864 2492 1880 2508
rect 1896 2492 1912 2508
rect 2072 2492 2088 2508
rect 2216 2492 2232 2508
rect 2328 2492 2360 2508
rect 2584 2492 2600 2508
rect 2696 2492 2712 2508
rect 3124 2492 3140 2508
rect 3144 2492 3160 2508
rect 3480 2492 3496 2508
rect 3528 2512 3544 2528
rect 3624 2512 3640 2528
rect 3768 2512 3784 2528
rect 3816 2492 3832 2508
rect 3848 2512 3896 2528
rect 3928 2512 3944 2528
rect 3992 2512 4008 2528
rect 3896 2492 3912 2508
rect 4088 2492 4120 2508
rect 4200 2492 4216 2508
rect 4248 2512 4264 2528
rect 4376 2512 4392 2528
rect 4568 2512 4584 2528
rect 4632 2514 4648 2530
rect 4744 2492 4760 2508
rect 4792 2512 4808 2528
rect 4872 2492 4888 2508
rect 4920 2512 4936 2528
rect 4968 2512 4984 2528
rect 5080 2512 5096 2528
rect 5128 2512 5144 2528
rect 5240 2512 5272 2528
rect 5304 2512 5320 2528
rect 5352 2512 5368 2528
rect 5528 2512 5544 2528
rect 5640 2512 5672 2528
rect 4908 2492 4924 2508
rect 5720 2512 5736 2528
rect 5768 2512 5784 2528
rect 5832 2512 5864 2528
rect 5992 2512 6008 2528
rect 6040 2512 6056 2528
rect 6216 2512 6232 2528
rect 5688 2492 5704 2508
rect 6344 2492 6360 2508
rect 6392 2512 6408 2528
rect 6568 2512 6584 2528
rect 6712 2512 6728 2528
rect 6792 2512 6824 2528
rect 6856 2512 6888 2528
rect 6488 2492 6504 2508
rect 6936 2512 6952 2528
rect 6984 2492 7000 2508
rect 7016 2512 7048 2528
rect 7192 2512 7208 2528
rect 7416 2512 7432 2528
rect 7512 2512 7528 2528
rect 7560 2512 7576 2528
rect 7608 2512 7624 2528
rect 7640 2512 7656 2528
rect 7672 2512 7688 2528
rect 7720 2512 7752 2528
rect 7816 2512 7832 2528
rect 7944 2512 7960 2528
rect 8024 2512 8040 2528
rect 7304 2492 7320 2508
rect 7388 2492 7404 2508
rect 7480 2492 7496 2508
rect 7672 2492 7704 2508
rect 1016 2472 1032 2488
rect 1080 2472 1096 2488
rect 1400 2472 1416 2488
rect 1528 2472 1544 2488
rect 1592 2472 1608 2488
rect 2008 2472 2024 2488
rect 2056 2472 2072 2488
rect 2184 2472 2200 2488
rect 2312 2472 2328 2488
rect 6008 2472 6024 2488
rect 6136 2472 6152 2488
rect 40 2432 56 2448
rect 408 2432 424 2448
rect 632 2432 648 2448
rect 856 2432 872 2448
rect 1064 2432 1080 2448
rect 1144 2432 1160 2448
rect 1608 2432 1624 2448
rect 1800 2432 1816 2448
rect 1880 2432 1896 2448
rect 2072 2432 2088 2448
rect 2120 2432 2136 2448
rect 3400 2432 3416 2448
rect 3592 2432 3608 2448
rect 5000 2432 5016 2448
rect 5192 2432 5208 2448
rect 5288 2432 5304 2448
rect 5848 2432 5864 2448
rect 5928 2432 5944 2448
rect 6824 2432 6840 2448
rect 7848 2432 7864 2448
rect 7992 2432 8008 2448
rect 925 2402 961 2418
rect 2957 2402 2993 2418
rect 5021 2402 5057 2418
rect 7053 2402 7089 2418
rect 424 2372 440 2388
rect 1032 2372 1048 2388
rect 2632 2372 2648 2388
rect 3912 2372 3928 2388
rect 3944 2372 3960 2388
rect 4216 2372 4232 2388
rect 4776 2372 4792 2388
rect 5224 2372 5240 2388
rect 5592 2372 5608 2388
rect 6584 2372 6600 2388
rect 7528 2372 7544 2388
rect 7688 2372 7704 2388
rect 7976 2372 7992 2388
rect 984 2352 1000 2368
rect 1240 2352 1256 2368
rect 8 2332 24 2348
rect 440 2332 456 2348
rect 968 2332 984 2348
rect 1048 2332 1064 2348
rect 1224 2332 1240 2348
rect 2712 2352 2728 2368
rect 4248 2352 4264 2368
rect 408 2312 424 2328
rect 984 2312 1000 2328
rect 1304 2332 1320 2348
rect 1704 2332 1720 2348
rect 2024 2332 2040 2348
rect 2152 2332 2168 2348
rect 5448 2332 5464 2348
rect 1272 2312 1288 2328
rect 1800 2312 1816 2328
rect 1976 2312 1992 2328
rect 2040 2312 2056 2328
rect 120 2292 152 2308
rect 200 2292 216 2308
rect 312 2292 328 2308
rect 392 2292 408 2308
rect 424 2292 440 2308
rect 552 2292 584 2308
rect 696 2292 712 2308
rect 840 2292 856 2308
rect 984 2292 1000 2308
rect 1032 2292 1048 2308
rect 1096 2292 1112 2308
rect 1192 2292 1208 2308
rect 1240 2292 1256 2308
rect 1288 2292 1304 2308
rect 1368 2292 1384 2308
rect 1464 2292 1480 2308
rect 1544 2292 1560 2308
rect 1688 2292 1704 2308
rect 1768 2292 1784 2308
rect 1816 2292 1848 2308
rect 1912 2292 1928 2308
rect 2056 2292 2072 2308
rect 2104 2292 2120 2308
rect 2248 2292 2264 2308
rect 2280 2292 2296 2308
rect 2312 2292 2328 2308
rect 2344 2312 2360 2328
rect 3000 2312 3016 2328
rect 3432 2312 3448 2328
rect 3496 2312 3512 2328
rect 3880 2312 3896 2328
rect 4200 2312 4216 2328
rect 4232 2312 4248 2328
rect 4296 2312 4312 2328
rect 4360 2312 4376 2328
rect 4408 2312 4424 2328
rect 4488 2312 4504 2328
rect 4840 2312 4856 2328
rect 4872 2312 4888 2328
rect 5464 2312 5496 2328
rect 2472 2292 2488 2308
rect 2520 2292 2536 2308
rect 2664 2292 2696 2308
rect 2744 2292 2760 2308
rect 2872 2292 2888 2308
rect 3032 2292 3048 2308
rect 3064 2292 3080 2308
rect 3208 2292 3224 2308
rect 3320 2292 3336 2308
rect 3352 2292 3368 2308
rect 3464 2292 3480 2308
rect 3544 2292 3560 2308
rect 3640 2292 3656 2308
rect 3704 2290 3720 2306
rect 3784 2292 3816 2308
rect 4056 2292 4088 2308
rect 4200 2292 4216 2308
rect 4328 2292 4344 2308
rect 152 2272 168 2288
rect 360 2272 376 2288
rect 824 2272 840 2288
rect 1080 2272 1096 2288
rect 232 2252 248 2268
rect 760 2252 776 2268
rect 1432 2272 1448 2288
rect 1496 2272 1512 2288
rect 1752 2272 1768 2288
rect 1784 2272 1800 2288
rect 1848 2272 1864 2288
rect 1880 2272 1896 2288
rect 2200 2272 2216 2288
rect 2264 2272 2280 2288
rect 2376 2272 2392 2288
rect 2552 2272 2568 2288
rect 2792 2272 2808 2288
rect 2984 2272 3000 2288
rect 3048 2272 3064 2288
rect 3112 2272 3128 2288
rect 3144 2272 3160 2288
rect 3256 2272 3272 2288
rect 3432 2272 3448 2288
rect 3480 2272 3496 2288
rect 3560 2272 3576 2288
rect 3736 2272 3752 2288
rect 3768 2272 3784 2288
rect 3848 2272 3864 2288
rect 4344 2272 4360 2288
rect 4408 2292 4424 2308
rect 4616 2292 4632 2308
rect 4680 2290 4696 2306
rect 4840 2292 4856 2308
rect 4984 2292 5000 2308
rect 5128 2292 5144 2308
rect 5352 2290 5368 2306
rect 5512 2292 5528 2308
rect 5544 2292 5560 2308
rect 5640 2292 5672 2308
rect 5704 2312 5720 2328
rect 5912 2312 5928 2328
rect 6232 2312 6248 2328
rect 6664 2312 6680 2328
rect 5816 2290 5832 2306
rect 5880 2292 5896 2308
rect 6072 2292 6088 2308
rect 6216 2292 6232 2308
rect 6248 2292 6280 2308
rect 6296 2292 6328 2308
rect 6408 2292 6456 2308
rect 6520 2292 6536 2308
rect 6772 2312 6788 2328
rect 6792 2312 6808 2328
rect 6856 2312 6872 2328
rect 6888 2312 6920 2328
rect 6984 2312 7000 2328
rect 6712 2292 6728 2308
rect 6760 2292 6776 2308
rect 6824 2292 6856 2308
rect 6920 2292 6936 2308
rect 7144 2292 7176 2308
rect 7256 2292 7288 2308
rect 7320 2312 7336 2328
rect 7400 2312 7416 2328
rect 7576 2312 7592 2328
rect 7464 2292 7480 2308
rect 7672 2312 7688 2328
rect 7608 2292 7640 2308
rect 7816 2292 7832 2308
rect 7944 2292 7960 2308
rect 4520 2272 4536 2288
rect 4872 2272 4888 2288
rect 5064 2272 5080 2288
rect 5112 2272 5128 2288
rect 5336 2272 5352 2288
rect 5384 2272 5400 2288
rect 5416 2272 5432 2288
rect 5464 2272 5480 2288
rect 5528 2272 5544 2288
rect 5624 2272 5640 2288
rect 5736 2272 5768 2288
rect 6024 2272 6040 2288
rect 6200 2272 6216 2288
rect 6264 2272 6280 2288
rect 6632 2272 6648 2288
rect 6728 2272 6760 2288
rect 6808 2272 6824 2288
rect 6952 2272 6968 2288
rect 7000 2272 7016 2288
rect 7240 2272 7256 2288
rect 7352 2272 7384 2288
rect 7432 2272 7448 2288
rect 7480 2272 7496 2288
rect 7544 2272 7560 2288
rect 7640 2272 7656 2288
rect 7704 2272 7736 2288
rect 7848 2272 7864 2288
rect 1160 2252 1176 2268
rect 1336 2252 1352 2268
rect 1592 2252 1608 2268
rect 1864 2252 1880 2268
rect 3640 2252 3656 2268
rect 3960 2252 3976 2268
rect 4280 2252 4296 2268
rect 4456 2252 4472 2268
rect 6152 2252 6168 2268
rect 6328 2252 6344 2268
rect 6392 2252 6408 2268
rect 6472 2252 6488 2268
rect 6504 2252 6520 2268
rect 7192 2252 7208 2268
rect 7496 2252 7512 2268
rect 168 2232 184 2248
rect 280 2232 296 2248
rect 504 2232 520 2248
rect 600 2232 616 2248
rect 664 2232 680 2248
rect 1128 2232 1144 2248
rect 1416 2232 1432 2248
rect 2216 2232 2232 2248
rect 2632 2232 2648 2248
rect 2712 2232 2728 2248
rect 2952 2232 2968 2248
rect 3416 2232 3432 2248
rect 3496 2232 3512 2248
rect 4296 2232 4312 2248
rect 4504 2232 4520 2248
rect 4776 2232 4792 2248
rect 4824 2232 4840 2248
rect 5176 2232 5192 2248
rect 5592 2232 5608 2248
rect 6680 2232 6696 2248
rect 7976 2232 7992 2248
rect 1949 2202 1985 2218
rect 3997 2202 4033 2218
rect 6045 2202 6081 2218
rect 216 2172 232 2188
rect 744 2172 760 2188
rect 1496 2172 1512 2188
rect 2056 2172 2072 2188
rect 2936 2172 2952 2188
rect 3000 2172 3016 2188
rect 3464 2172 3480 2188
rect 4344 2172 4360 2188
rect 4680 2172 4696 2188
rect 5832 2172 5848 2188
rect 6008 2172 6024 2188
rect 6248 2172 6264 2188
rect 7096 2172 7112 2188
rect 776 2152 792 2168
rect 1160 2152 1176 2168
rect 1256 2152 1272 2168
rect 1448 2152 1464 2168
rect 296 2132 312 2148
rect 456 2132 472 2148
rect 552 2132 568 2148
rect 840 2132 856 2148
rect 872 2132 888 2148
rect 1032 2132 1048 2148
rect 1384 2132 1400 2148
rect 3656 2152 3672 2168
rect 3736 2152 3752 2168
rect 4312 2152 4328 2168
rect 4920 2152 4936 2168
rect 1512 2132 1528 2148
rect 1608 2132 1624 2148
rect 1912 2132 1928 2148
rect 1976 2132 1992 2148
rect 2296 2132 2312 2148
rect 2376 2132 2392 2148
rect 2456 2132 2472 2148
rect 2552 2132 2568 2148
rect 2600 2132 2616 2148
rect 2760 2132 2792 2148
rect 2872 2132 2904 2148
rect 2952 2132 2968 2148
rect 3144 2132 3160 2148
rect 3208 2132 3224 2148
rect 3416 2132 3432 2148
rect 3544 2132 3560 2148
rect 3864 2132 3896 2148
rect 3960 2132 3976 2148
rect 4040 2132 4056 2148
rect 4088 2132 4104 2148
rect 4200 2132 4216 2148
rect 4264 2132 4280 2148
rect 4424 2132 4440 2148
rect 4472 2132 4488 2148
rect 4568 2132 4584 2148
rect 4616 2132 4632 2148
rect 4664 2132 4680 2148
rect 4728 2132 4744 2148
rect 4792 2132 4808 2148
rect 5096 2132 5112 2148
rect 5176 2132 5192 2148
rect 5304 2132 5320 2148
rect 5352 2132 5368 2148
rect 5400 2132 5416 2148
rect 5448 2132 5464 2148
rect 5496 2132 5512 2148
rect 5528 2132 5544 2148
rect 5656 2132 5688 2148
rect 5784 2132 5800 2148
rect 5960 2132 5976 2148
rect 6104 2132 6120 2148
rect 6216 2132 6232 2148
rect 6408 2152 6424 2168
rect 6776 2152 6792 2168
rect 6840 2152 6856 2168
rect 7304 2152 7320 2168
rect 7400 2152 7416 2168
rect 6536 2132 6552 2148
rect 6648 2132 6664 2148
rect 6920 2132 6936 2148
rect 6952 2132 6968 2148
rect 7016 2132 7032 2148
rect 88 2112 104 2128
rect 136 2112 152 2128
rect 312 2112 328 2128
rect 456 2112 472 2128
rect 536 2112 552 2128
rect 568 2112 584 2128
rect 664 2112 680 2128
rect 712 2112 728 2128
rect 808 2112 824 2128
rect 888 2112 904 2128
rect 952 2112 968 2128
rect 1112 2112 1128 2128
rect 1288 2112 1304 2128
rect 1352 2114 1368 2130
rect 1416 2112 1432 2128
rect 1528 2112 1544 2128
rect 1560 2112 1576 2128
rect 1672 2112 1688 2128
rect 1880 2114 1896 2130
rect 1992 2112 2024 2128
rect 2168 2112 2184 2128
rect 2216 2112 2232 2128
rect 2312 2112 2344 2128
rect 2424 2112 2440 2128
rect 680 2092 696 2108
rect 936 2092 952 2108
rect 1208 2092 1224 2108
rect 1544 2092 1560 2108
rect 2024 2092 2040 2108
rect 2344 2092 2360 2108
rect 2488 2092 2504 2108
rect 2536 2112 2552 2128
rect 2680 2112 2696 2128
rect 2792 2112 2808 2128
rect 2524 2092 2540 2108
rect 2804 2092 2820 2108
rect 2872 2112 2888 2128
rect 3048 2112 3064 2128
rect 3192 2112 3208 2128
rect 3256 2112 3272 2128
rect 3320 2112 3336 2128
rect 3368 2112 3384 2128
rect 3576 2112 3608 2128
rect 3784 2112 3800 2128
rect 3896 2112 3928 2128
rect 4056 2112 4072 2128
rect 4136 2112 4152 2128
rect 4168 2112 4184 2128
rect 4296 2112 4312 2128
rect 4488 2114 4504 2130
rect 2840 2092 2856 2108
rect 2936 2092 2952 2108
rect 2984 2092 3000 2108
rect 3032 2092 3048 2108
rect 3112 2092 3128 2108
rect 3272 2092 3288 2108
rect 3336 2092 3352 2108
rect 3480 2092 3496 2108
rect 3512 2092 3528 2108
rect 4008 2092 4024 2108
rect 4104 2092 4120 2108
rect 4280 2092 4296 2108
rect 4600 2092 4616 2108
rect 4648 2112 4664 2128
rect 4712 2112 4728 2128
rect 4760 2112 4776 2128
rect 4872 2112 4888 2128
rect 4936 2112 4968 2128
rect 5064 2112 5080 2128
rect 5272 2114 5288 2130
rect 4680 2092 4696 2108
rect 4824 2092 4840 2108
rect 4844 2092 4860 2108
rect 5384 2092 5400 2108
rect 5432 2112 5448 2128
rect 5576 2112 5592 2128
rect 5688 2112 5720 2128
rect 5864 2112 5880 2128
rect 5896 2112 5912 2128
rect 5944 2112 5960 2128
rect 5752 2092 5768 2108
rect 6136 2112 6168 2128
rect 6216 2112 6232 2128
rect 6264 2112 6296 2128
rect 6440 2112 6456 2128
rect 6504 2114 6520 2130
rect 6840 2114 6856 2130
rect 6072 2092 6088 2108
rect 6696 2092 6712 2108
rect 6952 2092 6968 2108
rect 7000 2112 7016 2128
rect 7496 2132 7512 2148
rect 7544 2132 7560 2148
rect 7656 2132 7672 2148
rect 7848 2132 7864 2148
rect 7880 2132 7896 2148
rect 7128 2112 7144 2128
rect 7160 2112 7192 2128
rect 7400 2114 7416 2130
rect 7544 2112 7576 2128
rect 7592 2092 7608 2108
rect 7656 2112 7688 2128
rect 7768 2112 7784 2128
rect 7896 2112 7928 2128
rect 7944 2112 7976 2128
rect 7628 2092 7644 2108
rect 7928 2092 7944 2108
rect 600 2072 616 2088
rect 648 2072 664 2088
rect 968 2072 984 2088
rect 1576 2072 1592 2088
rect 3064 2072 3080 2088
rect 3240 2072 3256 2088
rect 3352 2072 3368 2088
rect 4136 2072 4152 2088
rect 4232 2072 4248 2088
rect 4264 2072 4280 2088
rect 6584 2072 6600 2088
rect 216 2032 232 2048
rect 408 2032 424 2048
rect 632 2032 648 2048
rect 744 2032 760 2048
rect 984 2032 1000 2048
rect 1560 2032 1576 2048
rect 1688 2032 1704 2048
rect 3048 2032 3064 2048
rect 3192 2032 3208 2048
rect 3224 2032 3240 2048
rect 3320 2032 3336 2048
rect 3400 2032 3416 2048
rect 4984 2032 5000 2048
rect 5656 2032 5672 2048
rect 5832 2032 5848 2048
rect 5928 2032 5944 2048
rect 6328 2032 6344 2048
rect 6600 2032 6616 2048
rect 6664 2032 6680 2048
rect 6712 2032 6728 2048
rect 7096 2032 7112 2048
rect 7192 2032 7208 2048
rect 7992 2032 8008 2048
rect 925 2002 961 2018
rect 2957 2002 2993 2018
rect 5021 2002 5057 2018
rect 7053 2002 7089 2018
rect 984 1972 1000 1988
rect 2184 1972 2200 1988
rect 2344 1972 2360 1988
rect 2408 1972 2424 1988
rect 2680 1972 2696 1988
rect 2760 1972 2776 1988
rect 2824 1972 2840 1988
rect 3704 1972 3720 1988
rect 4248 1972 4264 1988
rect 6152 1972 6168 1988
rect 7400 1972 7416 1988
rect 7784 1972 7800 1988
rect 3368 1952 3384 1968
rect 328 1932 344 1948
rect 2600 1932 2616 1948
rect 3304 1932 3320 1948
rect 3352 1932 3384 1948
rect 3448 1932 3464 1948
rect 3608 1932 3624 1948
rect 3864 1932 3880 1948
rect 7832 1952 7848 1968
rect 3992 1932 4008 1948
rect 4200 1932 4216 1948
rect 4264 1932 4280 1948
rect 1528 1912 1544 1928
rect 2392 1912 2408 1928
rect 2920 1912 2936 1928
rect 72 1892 88 1908
rect 184 1892 200 1908
rect 376 1892 392 1908
rect 456 1892 472 1908
rect 504 1892 520 1908
rect 584 1892 600 1908
rect 664 1892 680 1908
rect 792 1892 808 1908
rect 824 1892 840 1908
rect 1016 1892 1032 1908
rect 1112 1892 1128 1908
rect 1144 1892 1160 1908
rect 1240 1892 1256 1908
rect 1320 1892 1336 1908
rect 1384 1892 1400 1908
rect 1512 1892 1528 1908
rect 1560 1892 1576 1908
rect 1656 1892 1688 1908
rect 1752 1892 1768 1908
rect 1784 1892 1800 1908
rect 1864 1890 1880 1906
rect 2104 1892 2120 1908
rect 2280 1892 2296 1908
rect 2520 1892 2536 1908
rect 2856 1892 2872 1908
rect 3032 1912 3048 1928
rect 3224 1912 3240 1928
rect 3352 1912 3368 1928
rect 3416 1912 3432 1928
rect 3464 1912 3480 1928
rect 3528 1912 3544 1928
rect 3656 1912 3672 1928
rect 3960 1912 3976 1928
rect 4120 1912 4136 1928
rect 4168 1912 4184 1928
rect 4232 1912 4248 1928
rect 4328 1912 4344 1928
rect 4392 1912 4408 1928
rect 4696 1912 4712 1928
rect 2968 1892 2984 1908
rect 3048 1892 3080 1908
rect 3112 1892 3128 1908
rect 3192 1892 3208 1908
rect 3384 1892 3400 1908
rect 3432 1892 3448 1908
rect 3480 1892 3496 1908
rect 264 1872 280 1888
rect 600 1872 632 1888
rect 1272 1872 1288 1888
rect 1576 1872 1592 1888
rect 696 1852 712 1868
rect 840 1852 856 1868
rect 1352 1852 1368 1868
rect 1480 1852 1496 1868
rect 1704 1852 1720 1868
rect 1768 1872 1784 1888
rect 1832 1872 1848 1888
rect 2088 1872 2104 1888
rect 2136 1872 2152 1888
rect 2392 1872 2408 1888
rect 2424 1872 2440 1888
rect 2520 1872 2536 1888
rect 2776 1872 2792 1888
rect 2808 1872 2824 1888
rect 2888 1872 2904 1888
rect 2952 1872 2968 1888
rect 2984 1872 3000 1888
rect 3080 1872 3096 1888
rect 3160 1872 3192 1888
rect 3336 1872 3352 1888
rect 3624 1892 3640 1908
rect 3672 1892 3688 1908
rect 3752 1892 3768 1908
rect 3816 1892 3832 1908
rect 3912 1892 3928 1908
rect 3976 1892 3992 1908
rect 4024 1892 4040 1908
rect 4184 1892 4200 1908
rect 4216 1892 4232 1908
rect 4248 1892 4264 1908
rect 4360 1892 4376 1908
rect 4552 1892 4584 1908
rect 5224 1912 5240 1928
rect 4728 1892 4760 1908
rect 4840 1892 4856 1908
rect 4872 1892 4888 1908
rect 5096 1892 5112 1908
rect 5928 1912 5944 1928
rect 5948 1912 5964 1928
rect 5256 1892 5304 1908
rect 5320 1892 5336 1908
rect 5400 1892 5416 1908
rect 3896 1872 3912 1888
rect 3944 1872 3960 1888
rect 4152 1872 4168 1888
rect 4440 1872 4456 1888
rect 4472 1872 4488 1888
rect 4664 1872 4680 1888
rect 4760 1872 4792 1888
rect 4904 1872 4920 1888
rect 5112 1872 5128 1888
rect 5192 1872 5208 1888
rect 5304 1872 5320 1888
rect 5384 1872 5400 1888
rect 5432 1872 5448 1888
rect 5624 1892 5656 1908
rect 5864 1890 5880 1906
rect 5960 1892 5976 1908
rect 6008 1892 6024 1908
rect 6088 1912 6104 1928
rect 6632 1912 6648 1928
rect 6696 1912 6712 1928
rect 6904 1912 6920 1928
rect 6952 1912 6968 1928
rect 6232 1892 6248 1908
rect 6440 1892 6456 1908
rect 6488 1890 6504 1906
rect 6616 1892 6632 1908
rect 6664 1892 6680 1908
rect 6696 1892 6712 1908
rect 6728 1892 6744 1908
rect 6776 1892 6808 1908
rect 6840 1892 6856 1908
rect 7032 1912 7048 1928
rect 7480 1912 7496 1928
rect 7624 1912 7640 1928
rect 7688 1912 7704 1928
rect 7000 1892 7016 1908
rect 7160 1892 7176 1908
rect 7288 1892 7304 1908
rect 7336 1892 7352 1908
rect 7496 1892 7512 1908
rect 7656 1892 7672 1908
rect 7816 1912 7832 1928
rect 7720 1892 7752 1908
rect 7784 1892 7800 1908
rect 7944 1892 7960 1908
rect 5528 1872 5544 1888
rect 5896 1872 5912 1888
rect 5976 1872 6008 1888
rect 6040 1872 6056 1888
rect 6312 1872 6328 1888
rect 6680 1872 6696 1888
rect 6744 1872 6760 1888
rect 6840 1872 6856 1888
rect 6872 1872 6888 1888
rect 6920 1872 6936 1888
rect 6984 1872 7000 1888
rect 7016 1872 7032 1888
rect 7352 1872 7368 1888
rect 7448 1872 7464 1888
rect 7592 1872 7608 1888
rect 7640 1872 7656 1888
rect 7752 1872 7784 1888
rect 7912 1872 7928 1888
rect 7976 1872 7992 1888
rect 1928 1852 1944 1868
rect 2024 1852 2040 1868
rect 5544 1852 5560 1868
rect 5608 1852 5624 1868
rect 5768 1852 5784 1868
rect 6424 1852 6440 1868
rect 6632 1852 6648 1868
rect 7208 1852 7224 1868
rect 40 1832 56 1848
rect 104 1832 120 1848
rect 632 1832 648 1848
rect 1224 1832 1240 1848
rect 1288 1832 1304 1848
rect 1416 1832 1432 1848
rect 1528 1832 1544 1848
rect 1624 1832 1640 1848
rect 2072 1832 2088 1848
rect 2248 1832 2264 1848
rect 3256 1832 3272 1848
rect 3496 1832 3512 1848
rect 3784 1832 3800 1848
rect 4072 1832 4088 1848
rect 4408 1832 4424 1848
rect 4984 1832 5000 1848
rect 5624 1832 5640 1848
rect 6904 1832 6920 1848
rect 7464 1832 7480 1848
rect 7544 1832 7560 1848
rect 7608 1832 7624 1848
rect 1949 1802 1985 1818
rect 3997 1802 4033 1818
rect 6045 1802 6081 1818
rect 88 1772 104 1788
rect 728 1772 744 1788
rect 1720 1772 1736 1788
rect 2024 1772 2040 1788
rect 2056 1772 2072 1788
rect 2328 1772 2344 1788
rect 2936 1772 2952 1788
rect 3368 1772 3384 1788
rect 3656 1772 3672 1788
rect 4232 1772 4248 1788
rect 4968 1772 4984 1788
rect 5816 1772 5832 1788
rect 6328 1772 6344 1788
rect 6488 1772 6504 1788
rect 6664 1772 6680 1788
rect 40 1752 56 1768
rect 104 1732 120 1748
rect 376 1738 392 1754
rect 648 1752 664 1768
rect 1384 1752 1400 1768
rect 1592 1752 1608 1768
rect 1656 1752 1672 1768
rect 1976 1752 1992 1768
rect 2008 1752 2024 1768
rect 4440 1752 4456 1768
rect 4520 1752 4536 1768
rect 4744 1752 4760 1768
rect 5480 1752 5496 1768
rect 5608 1752 5624 1768
rect 5640 1752 5656 1768
rect 5704 1752 5720 1768
rect 6872 1752 6888 1768
rect 7032 1752 7048 1768
rect 7928 1752 7944 1768
rect 744 1732 760 1748
rect 1096 1732 1112 1748
rect 1224 1732 1240 1748
rect 1256 1732 1272 1748
rect 1320 1732 1352 1748
rect 1512 1732 1528 1748
rect 1640 1732 1672 1748
rect 2168 1732 2184 1748
rect 2376 1732 2392 1748
rect 2440 1732 2456 1748
rect 2472 1732 2488 1748
rect 2568 1732 2584 1748
rect 2760 1732 2776 1748
rect 2856 1732 2872 1748
rect 2888 1732 2904 1748
rect 3016 1732 3032 1748
rect 3048 1732 3064 1748
rect 3256 1732 3272 1748
rect 4504 1732 4520 1748
rect 4632 1732 4648 1748
rect 4808 1732 4824 1748
rect 4920 1732 4936 1748
rect 5032 1732 5048 1748
rect 5144 1732 5160 1748
rect 5192 1732 5208 1748
rect 5528 1732 5544 1748
rect 5592 1732 5608 1748
rect 5768 1732 5784 1748
rect 5976 1732 5992 1748
rect 6104 1732 6120 1748
rect 6168 1732 6184 1748
rect 6200 1732 6216 1748
rect 6264 1732 6280 1748
rect 6344 1732 6360 1748
rect 6440 1732 6456 1748
rect 6536 1732 6552 1748
rect 6616 1732 6632 1748
rect 7000 1732 7016 1748
rect 7080 1732 7096 1748
rect 7160 1732 7176 1748
rect 7208 1732 7224 1748
rect 7336 1732 7352 1748
rect 7368 1732 7384 1748
rect 7448 1732 7480 1748
rect 7528 1732 7544 1748
rect 8 1712 24 1728
rect 120 1712 136 1728
rect 168 1712 184 1728
rect 216 1712 232 1728
rect 248 1712 264 1728
rect 296 1712 312 1728
rect 344 1712 360 1728
rect 424 1712 440 1728
rect 472 1712 488 1728
rect 552 1712 568 1728
rect 600 1712 616 1728
rect 680 1712 696 1728
rect 776 1712 808 1728
rect 872 1712 888 1728
rect 968 1712 984 1728
rect 1032 1712 1048 1728
rect 1176 1712 1192 1728
rect 1272 1712 1288 1728
rect 1336 1712 1352 1728
rect 1416 1712 1432 1728
rect 1496 1712 1512 1728
rect 1544 1712 1560 1728
rect 1624 1712 1640 1728
rect 1704 1712 1720 1728
rect 1816 1712 1832 1728
rect 1880 1712 1896 1728
rect 1944 1712 1960 1728
rect 2040 1712 2056 1728
rect 2136 1712 2152 1728
rect 2168 1712 2184 1728
rect 2280 1712 2296 1728
rect 184 1692 216 1708
rect 312 1692 344 1708
rect 152 1672 168 1688
rect 200 1672 216 1688
rect 232 1672 248 1688
rect 280 1672 296 1688
rect 360 1672 376 1688
rect 408 1672 424 1688
rect 456 1692 472 1708
rect 568 1692 600 1708
rect 856 1692 872 1708
rect 952 1692 968 1708
rect 1016 1692 1032 1708
rect 1128 1692 1144 1708
rect 1192 1692 1208 1708
rect 1400 1692 1416 1708
rect 1484 1692 1500 1708
rect 1528 1692 1544 1708
rect 1832 1692 1848 1708
rect 1896 1692 1912 1708
rect 1976 1692 1992 1708
rect 2264 1692 2280 1708
rect 2344 1692 2360 1708
rect 2392 1692 2408 1708
rect 2504 1692 2520 1708
rect 2536 1712 2568 1728
rect 2728 1712 2744 1728
rect 3032 1712 3048 1728
rect 3208 1712 3224 1728
rect 3336 1712 3352 1728
rect 3416 1712 3432 1728
rect 3448 1712 3464 1728
rect 3496 1712 3512 1728
rect 3528 1712 3560 1728
rect 3624 1712 3640 1728
rect 3704 1712 3720 1728
rect 3832 1712 3848 1728
rect 3960 1712 3976 1728
rect 4056 1712 4072 1728
rect 4104 1712 4120 1728
rect 4152 1712 4184 1728
rect 4248 1712 4264 1728
rect 4296 1712 4312 1728
rect 4344 1712 4392 1728
rect 4472 1712 4504 1728
rect 4616 1712 4632 1728
rect 4792 1712 4808 1728
rect 4904 1712 4920 1728
rect 4936 1712 4952 1728
rect 5160 1712 5176 1728
rect 2872 1692 2904 1708
rect 2984 1692 3016 1708
rect 3976 1692 3992 1708
rect 4040 1692 4056 1708
rect 4088 1692 4104 1708
rect 4168 1692 4184 1708
rect 4216 1692 4232 1708
rect 4296 1692 4312 1708
rect 4344 1692 4360 1708
rect 4456 1692 4472 1708
rect 4824 1692 4840 1708
rect 4968 1692 5000 1708
rect 5016 1692 5048 1708
rect 5128 1692 5144 1708
rect 5352 1712 5384 1728
rect 5528 1712 5592 1728
rect 5608 1712 5624 1728
rect 5672 1712 5704 1728
rect 5752 1712 5768 1728
rect 5800 1712 5816 1728
rect 5896 1712 5928 1728
rect 6008 1712 6024 1728
rect 6072 1714 6088 1730
rect 5224 1692 5240 1708
rect 5256 1692 5272 1708
rect 5496 1692 5512 1708
rect 5816 1692 5832 1708
rect 6200 1692 6216 1708
rect 6248 1712 6264 1728
rect 6296 1712 6312 1728
rect 6424 1712 6440 1728
rect 6472 1692 6488 1708
rect 6520 1712 6536 1728
rect 6568 1712 6584 1728
rect 6696 1712 6712 1728
rect 6744 1712 6760 1728
rect 6792 1712 6824 1728
rect 6952 1712 6968 1728
rect 7064 1712 7080 1728
rect 7240 1712 7256 1728
rect 7336 1712 7352 1728
rect 6824 1692 6840 1708
rect 7032 1692 7048 1708
rect 7320 1692 7336 1708
rect 7432 1712 7448 1728
rect 7480 1712 7496 1728
rect 7512 1712 7528 1728
rect 7688 1712 7704 1728
rect 7880 1712 7896 1728
rect 7912 1712 7928 1728
rect 7400 1692 7416 1708
rect 7492 1692 7508 1708
rect 7512 1692 7528 1708
rect 7640 1692 7656 1708
rect 456 1672 472 1688
rect 488 1672 504 1688
rect 536 1672 552 1688
rect 168 1652 184 1668
rect 296 1652 312 1668
rect 424 1652 440 1668
rect 472 1652 488 1668
rect 888 1672 904 1688
rect 1048 1672 1064 1688
rect 1160 1672 1176 1688
rect 1032 1652 1048 1668
rect 1432 1672 1448 1688
rect 1528 1672 1544 1688
rect 1800 1672 1816 1688
rect 1864 1672 1880 1688
rect 1928 1672 1944 1688
rect 2296 1672 2312 1688
rect 3416 1672 3432 1688
rect 3480 1672 3496 1688
rect 3800 1672 3816 1688
rect 3944 1672 3960 1688
rect 3992 1672 4008 1688
rect 4120 1672 4136 1688
rect 4184 1672 4200 1688
rect 4216 1672 4232 1688
rect 7544 1672 7560 1688
rect 3736 1652 3752 1668
rect 632 1632 648 1648
rect 824 1632 840 1648
rect 1000 1632 1016 1648
rect 1112 1632 1128 1648
rect 1816 1632 1832 1648
rect 1880 1632 1896 1648
rect 1944 1632 1960 1648
rect 2312 1632 2328 1648
rect 2424 1632 2440 1648
rect 3432 1632 3448 1648
rect 3496 1632 3512 1648
rect 3576 1632 3592 1648
rect 3656 1632 3672 1648
rect 3896 1632 3912 1648
rect 3960 1632 3976 1648
rect 4072 1632 4088 1648
rect 4104 1632 4120 1648
rect 4200 1632 4216 1648
rect 4312 1632 4328 1648
rect 4872 1632 4888 1648
rect 5880 1632 5896 1648
rect 6392 1632 6408 1648
rect 6664 1632 6680 1648
rect 6776 1632 6792 1648
rect 7992 1632 8008 1648
rect 925 1602 961 1618
rect 2957 1602 2993 1618
rect 5021 1602 5057 1618
rect 7053 1602 7089 1618
rect 344 1572 360 1588
rect 392 1572 408 1588
rect 456 1572 472 1588
rect 600 1572 616 1588
rect 1464 1572 1480 1588
rect 3000 1572 3016 1588
rect 3368 1572 3384 1588
rect 3464 1572 3480 1588
rect 3704 1572 3720 1588
rect 4200 1572 4216 1588
rect 4920 1572 4936 1588
rect 4968 1572 4984 1588
rect 408 1532 424 1548
rect 472 1532 488 1548
rect 616 1532 632 1548
rect 1288 1532 1304 1548
rect 3608 1532 3624 1548
rect 3928 1532 3944 1548
rect 4024 1532 4040 1548
rect 4104 1532 4120 1548
rect 376 1512 392 1528
rect 440 1512 456 1528
rect 584 1512 600 1528
rect 1128 1512 1144 1528
rect 88 1492 104 1508
rect 136 1492 152 1508
rect 216 1492 232 1508
rect 312 1492 328 1508
rect 392 1492 408 1508
rect 456 1492 472 1508
rect 568 1492 584 1508
rect 600 1492 616 1508
rect 712 1492 728 1508
rect 808 1492 824 1508
rect 952 1490 968 1506
rect 1064 1492 1080 1508
rect 1144 1492 1176 1508
rect 1336 1492 1352 1508
rect 1640 1490 1656 1506
rect 1720 1492 1752 1508
rect 1784 1512 1800 1528
rect 1816 1512 1832 1528
rect 2056 1512 2072 1528
rect 2120 1512 2136 1528
rect 2232 1512 2248 1528
rect 2392 1512 2408 1528
rect 2424 1512 2440 1528
rect 2552 1512 2568 1528
rect 2808 1512 2824 1528
rect 2888 1512 2904 1528
rect 984 1472 1000 1488
rect 1416 1472 1432 1488
rect 1624 1472 1640 1488
rect 1672 1472 1688 1488
rect 1704 1472 1720 1488
rect 1832 1492 1848 1508
rect 1896 1492 1912 1508
rect 1992 1492 2008 1508
rect 2088 1492 2104 1508
rect 2152 1492 2168 1508
rect 2200 1492 2216 1508
rect 2296 1492 2312 1508
rect 1880 1472 1896 1488
rect 2104 1472 2120 1488
rect 2168 1472 2200 1488
rect 2248 1472 2264 1488
rect 2344 1472 2360 1488
rect 2440 1472 2456 1488
rect 2472 1472 2488 1488
rect 2504 1492 2520 1508
rect 2536 1492 2552 1508
rect 2648 1492 2664 1508
rect 2776 1492 2792 1508
rect 3480 1512 3496 1528
rect 3896 1512 3912 1528
rect 4184 1512 4200 1528
rect 4280 1512 4296 1528
rect 4392 1512 4408 1528
rect 4456 1512 4472 1528
rect 4600 1512 4616 1528
rect 2920 1492 2952 1508
rect 3128 1492 3160 1508
rect 3320 1492 3336 1508
rect 3512 1492 3528 1508
rect 3736 1492 3752 1508
rect 3848 1492 3864 1508
rect 3912 1492 3928 1508
rect 4008 1492 4024 1508
rect 4296 1492 4312 1508
rect 4488 1492 4504 1508
rect 4632 1492 4648 1508
rect 4696 1490 4712 1506
rect 4760 1492 4776 1508
rect 4840 1512 4856 1528
rect 5080 1512 5096 1528
rect 5268 1512 5284 1528
rect 5352 1512 5368 1528
rect 5704 1512 5720 1528
rect 5112 1492 5128 1508
rect 5176 1490 5192 1506
rect 5256 1492 5272 1508
rect 5432 1492 5448 1508
rect 5560 1492 5592 1508
rect 5832 1512 5848 1528
rect 5736 1492 5768 1508
rect 6200 1512 6216 1528
rect 5880 1492 5912 1508
rect 6008 1492 6024 1508
rect 6056 1490 6072 1506
rect 6312 1512 6328 1528
rect 6536 1512 6552 1528
rect 6232 1492 6264 1508
rect 6296 1492 6312 1508
rect 6328 1492 6344 1508
rect 6360 1492 6376 1508
rect 6440 1492 6456 1508
rect 6488 1492 6520 1508
rect 6600 1492 6616 1508
rect 6664 1512 6680 1528
rect 6760 1512 6776 1528
rect 6792 1512 6808 1528
rect 6888 1512 6904 1528
rect 6968 1512 7000 1528
rect 7048 1512 7064 1528
rect 7176 1512 7192 1528
rect 6920 1492 6936 1508
rect 7256 1512 7272 1528
rect 7416 1512 7432 1528
rect 7224 1492 7240 1508
rect 7288 1492 7304 1508
rect 7576 1512 7592 1528
rect 7640 1512 7656 1528
rect 7732 1512 7748 1528
rect 7752 1512 7768 1528
rect 7992 1512 8008 1528
rect 7464 1492 7480 1508
rect 7512 1492 7528 1508
rect 7608 1492 7624 1508
rect 7704 1492 7720 1508
rect 7848 1492 7880 1508
rect 2536 1472 2552 1488
rect 2728 1472 2744 1488
rect 2840 1472 2856 1488
rect 3448 1472 3464 1488
rect 3496 1472 3512 1488
rect 3592 1472 3608 1488
rect 3656 1472 3672 1488
rect 3832 1472 3848 1488
rect 3880 1472 3896 1488
rect 3960 1472 3976 1488
rect 4104 1472 4120 1488
rect 4152 1472 4168 1488
rect 4360 1472 4376 1488
rect 4392 1472 4408 1488
rect 4680 1472 4696 1488
rect 4760 1472 4776 1488
rect 4792 1472 4808 1488
rect 4872 1472 4888 1488
rect 72 1452 88 1468
rect 136 1452 152 1468
rect 1992 1452 2008 1468
rect 3336 1452 3352 1468
rect 3432 1452 3448 1468
rect 4248 1452 4264 1468
rect 4408 1452 4424 1468
rect 4952 1472 4968 1488
rect 5240 1472 5256 1488
rect 5320 1472 5336 1488
rect 5352 1472 5368 1488
rect 5768 1472 5784 1488
rect 5800 1472 5816 1488
rect 5864 1472 5880 1488
rect 5896 1472 5912 1488
rect 6152 1472 6184 1488
rect 6264 1472 6296 1488
rect 6344 1472 6360 1488
rect 6408 1472 6424 1488
rect 6568 1472 6600 1488
rect 6632 1472 6648 1488
rect 6728 1472 6744 1488
rect 6856 1472 6872 1488
rect 6904 1472 6920 1488
rect 6936 1472 6952 1488
rect 7048 1472 7064 1488
rect 7080 1472 7096 1488
rect 7128 1472 7144 1488
rect 7240 1472 7272 1488
rect 7384 1472 7400 1488
rect 7416 1472 7432 1488
rect 7480 1472 7496 1488
rect 7624 1472 7640 1488
rect 7688 1472 7720 1488
rect 7800 1472 7816 1488
rect 8024 1472 8040 1488
rect 6376 1452 6392 1468
rect 6408 1452 6424 1468
rect 7032 1452 7048 1468
rect 7368 1452 7384 1468
rect 264 1432 280 1448
rect 536 1432 552 1448
rect 680 1432 696 1448
rect 760 1432 776 1448
rect 824 1432 840 1448
rect 1096 1432 1112 1448
rect 1192 1432 1208 1448
rect 1832 1432 1848 1448
rect 2008 1432 2024 1448
rect 2120 1432 2136 1448
rect 2312 1432 2328 1448
rect 3288 1432 3304 1448
rect 3704 1432 3720 1448
rect 3800 1432 3816 1448
rect 3992 1432 4008 1448
rect 4344 1432 4360 1448
rect 4472 1432 4488 1448
rect 4520 1432 4536 1448
rect 5640 1432 5656 1448
rect 6552 1432 6568 1448
rect 6760 1432 6776 1448
rect 6808 1432 6824 1448
rect 6888 1432 6904 1448
rect 7000 1432 7016 1448
rect 7192 1432 7208 1448
rect 7544 1432 7560 1448
rect 7576 1432 7592 1448
rect 7672 1432 7688 1448
rect 8008 1432 8024 1448
rect 1949 1402 1985 1418
rect 3997 1402 4033 1418
rect 6045 1402 6081 1418
rect 88 1372 104 1388
rect 1016 1372 1032 1388
rect 1064 1372 1080 1388
rect 1272 1372 1288 1388
rect 1464 1372 1480 1388
rect 1560 1372 1576 1388
rect 2568 1372 2584 1388
rect 3256 1372 3272 1388
rect 3368 1372 3384 1388
rect 3416 1372 3432 1388
rect 3496 1372 3512 1388
rect 4232 1372 4248 1388
rect 5848 1372 5864 1388
rect 5944 1372 5960 1388
rect 6392 1372 6408 1388
rect 6744 1372 6760 1388
rect 7064 1372 7080 1388
rect 7368 1372 7384 1388
rect 7704 1372 7720 1388
rect 7752 1372 7768 1388
rect 40 1352 56 1368
rect 904 1352 920 1368
rect 1256 1352 1272 1368
rect 1464 1352 1480 1368
rect 2264 1352 2280 1368
rect 104 1332 120 1348
rect 1032 1332 1048 1348
rect 1112 1332 1128 1348
rect 1144 1332 1160 1348
rect 1176 1332 1192 1348
rect 1304 1332 1320 1348
rect 1496 1332 1528 1348
rect 1832 1332 1848 1348
rect 2088 1332 2104 1348
rect 2200 1332 2216 1348
rect 2376 1352 2392 1368
rect 3320 1352 3336 1368
rect 3384 1352 3416 1368
rect 3864 1352 3880 1368
rect 3944 1352 3960 1368
rect 4216 1352 4232 1368
rect 4376 1352 4392 1368
rect 2360 1332 2376 1348
rect 2536 1332 2552 1348
rect 2616 1332 2648 1348
rect 2712 1332 2728 1348
rect 2744 1332 2760 1348
rect 2792 1332 2808 1348
rect 2856 1332 2872 1348
rect 2968 1332 2984 1348
rect 3048 1332 3064 1348
rect 3176 1332 3192 1348
rect 3448 1332 3464 1348
rect 3560 1332 3576 1348
rect 3640 1332 3656 1348
rect 3688 1332 3704 1348
rect 3976 1332 3992 1348
rect 4024 1332 4040 1348
rect 4424 1332 4440 1348
rect 4632 1332 4648 1348
rect 4872 1352 4888 1368
rect 5640 1352 5656 1368
rect 5800 1352 5816 1368
rect 6008 1352 6040 1368
rect 6264 1352 6280 1368
rect 6344 1352 6360 1368
rect 4760 1332 4776 1348
rect 4856 1332 4872 1348
rect 5112 1332 5128 1348
rect 5224 1332 5240 1348
rect 5384 1332 5416 1348
rect 5512 1332 5528 1348
rect 5688 1332 5720 1348
rect 6312 1332 6328 1348
rect 6616 1352 6632 1368
rect 7304 1352 7320 1368
rect 7736 1352 7752 1368
rect 6392 1332 6408 1348
rect 6488 1332 6504 1348
rect 6536 1332 6552 1348
rect 6808 1332 6824 1348
rect 6872 1332 6888 1348
rect 6936 1332 6952 1348
rect 7160 1332 7176 1348
rect 7224 1332 7240 1348
rect 7544 1332 7560 1348
rect 7576 1332 7592 1348
rect 7656 1332 7672 1348
rect 7800 1332 7832 1348
rect 7880 1332 7896 1348
rect 7944 1332 7960 1348
rect 8008 1332 8024 1348
rect 8 1312 24 1328
rect 120 1312 136 1328
rect 168 1312 200 1328
rect 232 1312 248 1328
rect 296 1312 312 1328
rect 344 1312 360 1328
rect 408 1312 424 1328
rect 472 1312 488 1328
rect 536 1312 552 1328
rect 600 1312 616 1328
rect 664 1312 680 1328
rect 728 1312 744 1328
rect 808 1312 824 1328
rect 872 1312 888 1328
rect 904 1312 920 1328
rect 936 1312 952 1328
rect 1048 1312 1064 1328
rect 1096 1312 1112 1328
rect 1192 1312 1208 1328
rect 1256 1312 1272 1328
rect 1336 1312 1352 1328
rect 1448 1312 1464 1328
rect 1528 1312 1544 1328
rect 1592 1312 1608 1328
rect 1672 1312 1688 1328
rect 1720 1312 1736 1328
rect 1784 1312 1800 1328
rect 1880 1312 1896 1328
rect 1928 1312 1944 1328
rect 2072 1312 2088 1328
rect 2104 1312 2120 1328
rect 2168 1312 2184 1328
rect 2232 1312 2248 1328
rect 2312 1312 2328 1328
rect 2344 1312 2360 1328
rect 2488 1312 2504 1328
rect 2696 1312 2712 1328
rect 2728 1312 2744 1328
rect 2856 1312 2888 1328
rect 248 1292 264 1308
rect 152 1272 168 1288
rect 216 1272 232 1288
rect 280 1272 296 1288
rect 328 1292 344 1308
rect 392 1292 408 1308
rect 456 1292 472 1308
rect 520 1292 536 1308
rect 584 1292 600 1308
rect 648 1292 664 1308
rect 712 1292 728 1308
rect 824 1292 840 1308
rect 888 1292 904 1308
rect 1064 1292 1080 1308
rect 1128 1292 1144 1308
rect 1320 1292 1336 1308
rect 1576 1292 1592 1308
rect 1672 1292 1688 1308
rect 1912 1292 1928 1308
rect 2116 1292 2132 1308
rect 2136 1292 2152 1308
rect 2568 1292 2584 1308
rect 2760 1292 2776 1308
rect 2884 1292 2900 1308
rect 3080 1314 3096 1330
rect 3288 1312 3304 1328
rect 3432 1312 3448 1328
rect 3608 1312 3624 1328
rect 3640 1312 3656 1328
rect 3672 1312 3688 1328
rect 3736 1312 3752 1328
rect 3800 1312 3816 1328
rect 3832 1312 3848 1328
rect 3912 1312 3928 1328
rect 3944 1312 3960 1328
rect 3992 1312 4024 1328
rect 4056 1312 4072 1328
rect 4104 1312 4120 1328
rect 4136 1312 4152 1328
rect 4168 1312 4184 1328
rect 4248 1312 4264 1328
rect 4296 1312 4312 1328
rect 4360 1312 4376 1328
rect 4472 1312 4488 1328
rect 4520 1312 4536 1328
rect 4600 1312 4616 1328
rect 4664 1312 4680 1328
rect 2936 1292 2952 1308
rect 3496 1292 3512 1308
rect 3528 1292 3544 1308
rect 3560 1292 3576 1308
rect 3624 1292 3640 1308
rect 3752 1292 3768 1308
rect 3784 1292 3800 1308
rect 3816 1292 3832 1308
rect 3960 1292 3976 1308
rect 4072 1292 4088 1308
rect 4152 1292 4168 1308
rect 4312 1292 4328 1308
rect 4424 1292 4456 1308
rect 4504 1292 4520 1308
rect 4616 1292 4648 1308
rect 4792 1292 4808 1308
rect 4840 1312 4856 1328
rect 4952 1312 4984 1328
rect 5176 1312 5192 1328
rect 5304 1312 5320 1328
rect 5416 1312 5448 1328
rect 4828 1292 4844 1308
rect 5528 1312 5544 1328
rect 5560 1312 5576 1328
rect 5736 1312 5752 1328
rect 5880 1312 5896 1328
rect 5912 1312 5928 1328
rect 5960 1312 5976 1328
rect 6152 1312 6184 1328
rect 6296 1312 6328 1328
rect 6408 1312 6424 1328
rect 6504 1312 6520 1328
rect 6616 1314 6632 1330
rect 6776 1312 6824 1328
rect 6856 1312 6872 1328
rect 6920 1312 6936 1328
rect 6968 1312 7000 1328
rect 7176 1312 7192 1328
rect 7272 1312 7304 1328
rect 7336 1312 7352 1328
rect 7464 1312 7480 1328
rect 7512 1314 7528 1330
rect 7592 1312 7624 1328
rect 7832 1312 7848 1328
rect 7896 1312 7928 1328
rect 5480 1292 5496 1308
rect 5528 1292 5544 1308
rect 5624 1292 5640 1308
rect 5992 1292 6008 1308
rect 6552 1292 6568 1308
rect 6760 1292 6776 1308
rect 6824 1292 6840 1308
rect 6888 1292 6904 1308
rect 6908 1292 6924 1308
rect 7000 1292 7016 1308
rect 7688 1292 7704 1308
rect 7768 1292 7784 1308
rect 7864 1292 7880 1308
rect 7928 1292 7944 1308
rect 7960 1292 7976 1308
rect 168 1252 184 1268
rect 232 1252 248 1268
rect 360 1272 376 1288
rect 424 1272 440 1288
rect 488 1272 504 1288
rect 552 1272 568 1288
rect 616 1272 632 1288
rect 680 1272 696 1288
rect 744 1272 760 1288
rect 792 1272 808 1288
rect 856 1272 872 1288
rect 1352 1272 1368 1288
rect 840 1252 856 1268
rect 1608 1272 1624 1288
rect 1640 1272 1672 1288
rect 1736 1272 1752 1288
rect 1864 1272 1880 1288
rect 1944 1272 1960 1288
rect 2040 1272 2056 1288
rect 3592 1272 3624 1288
rect 3720 1272 3736 1288
rect 3800 1272 3816 1288
rect 3896 1272 3912 1288
rect 4104 1272 4120 1288
rect 4184 1272 4200 1288
rect 4280 1272 4296 1288
rect 4392 1272 4408 1288
rect 4440 1272 4456 1288
rect 4536 1272 4552 1288
rect 4584 1272 4600 1288
rect 1928 1252 1944 1268
rect 4168 1252 4184 1268
rect 4520 1252 4536 1268
rect 296 1232 312 1248
rect 408 1232 424 1248
rect 504 1232 520 1248
rect 536 1232 552 1248
rect 600 1232 616 1248
rect 664 1232 680 1248
rect 728 1232 744 1248
rect 776 1232 792 1248
rect 1336 1232 1352 1248
rect 1720 1232 1736 1248
rect 1848 1232 1864 1248
rect 2664 1232 2680 1248
rect 3256 1232 3272 1248
rect 3608 1232 3624 1248
rect 3736 1232 3752 1248
rect 3800 1232 3816 1248
rect 3880 1232 3896 1248
rect 4120 1232 4136 1248
rect 4296 1232 4312 1248
rect 4328 1232 4344 1248
rect 4488 1232 4504 1248
rect 4600 1232 4616 1248
rect 5144 1232 5160 1248
rect 7832 1232 7848 1248
rect 925 1202 961 1218
rect 2957 1202 2993 1218
rect 5021 1202 5057 1218
rect 7053 1202 7089 1218
rect 168 1172 184 1188
rect 360 1172 376 1188
rect 888 1172 904 1188
rect 1016 1172 1032 1188
rect 1928 1172 1944 1188
rect 2744 1172 2760 1188
rect 3720 1172 3736 1188
rect 4616 1172 4632 1188
rect 4824 1172 4840 1188
rect 5944 1172 5960 1188
rect 7512 1172 7528 1188
rect 7848 1172 7864 1188
rect 40 1152 56 1168
rect 488 1152 504 1168
rect 24 1132 40 1148
rect 88 1132 104 1148
rect 168 1132 184 1148
rect 232 1132 248 1148
rect 296 1132 328 1148
rect 344 1132 360 1148
rect 408 1132 424 1148
rect 472 1132 488 1148
rect 536 1132 552 1148
rect 600 1132 616 1148
rect 872 1132 888 1148
rect 952 1132 1000 1148
rect 2232 1132 2248 1148
rect 3960 1132 3976 1148
rect 4184 1132 4200 1148
rect 4248 1132 4264 1148
rect 4344 1132 4360 1148
rect 4392 1132 4408 1148
rect 4440 1132 4456 1148
rect 4568 1132 4584 1148
rect 4632 1132 4648 1148
rect 4664 1132 4680 1148
rect 4712 1132 4728 1148
rect 4760 1132 4776 1148
rect 56 1112 72 1128
rect 120 1112 136 1128
rect 184 1112 216 1128
rect 248 1112 280 1128
rect 376 1112 392 1128
rect 440 1112 456 1128
rect 504 1112 520 1128
rect 568 1112 584 1128
rect 632 1112 648 1128
rect 904 1112 920 1128
rect 1272 1112 1288 1128
rect 1316 1112 1332 1128
rect 1336 1112 1352 1128
rect 1528 1112 1544 1128
rect 1736 1112 1752 1128
rect 1832 1112 1848 1128
rect 1896 1112 1912 1128
rect 2312 1112 2344 1128
rect 2392 1112 2408 1128
rect 2456 1112 2472 1128
rect 2760 1112 2776 1128
rect 2824 1112 2856 1128
rect 2872 1112 2888 1128
rect 3160 1112 3176 1128
rect 3192 1112 3208 1128
rect 40 1092 56 1108
rect 104 1092 120 1108
rect 168 1092 184 1108
rect 216 1092 232 1108
rect 280 1092 296 1108
rect 360 1092 376 1108
rect 424 1092 440 1108
rect 488 1092 504 1108
rect 552 1092 568 1108
rect 616 1092 632 1108
rect 664 1092 680 1108
rect 792 1092 808 1108
rect 840 1092 856 1108
rect 872 1092 888 1108
rect 968 1092 984 1108
rect 1080 1092 1096 1108
rect 1160 1092 1176 1108
rect 1240 1092 1256 1108
rect 1304 1092 1320 1108
rect 1416 1092 1432 1108
rect 1496 1092 1512 1108
rect 1560 1092 1576 1108
rect 1624 1092 1640 1108
rect 1688 1092 1704 1108
rect 1800 1092 1832 1108
rect 1864 1092 1880 1108
rect 2120 1092 2136 1108
rect 2264 1092 2280 1108
rect 2296 1092 2312 1108
rect 2360 1092 2376 1108
rect 2584 1092 2600 1108
rect 2792 1092 2808 1108
rect 2840 1092 2856 1108
rect 2904 1092 2920 1108
rect 3048 1092 3080 1108
rect 3228 1112 3244 1128
rect 3368 1112 3384 1128
rect 3240 1092 3256 1108
rect 3404 1112 3420 1128
rect 3496 1112 3512 1128
rect 3416 1092 3432 1108
rect 3624 1112 3640 1128
rect 3752 1112 3768 1128
rect 3860 1112 3876 1128
rect 3880 1112 3896 1128
rect 3944 1112 3960 1128
rect 3976 1112 3992 1128
rect 4088 1112 4104 1128
rect 4168 1112 4184 1128
rect 4216 1112 4232 1128
rect 4424 1112 4440 1128
rect 4536 1112 4552 1128
rect 4600 1112 4616 1128
rect 4728 1112 4744 1128
rect 4792 1112 4808 1128
rect 4904 1112 4920 1128
rect 3544 1092 3560 1108
rect 3592 1092 3608 1108
rect 3704 1092 3720 1108
rect 3800 1092 3816 1108
rect 3848 1092 3864 1108
rect 3880 1092 3896 1108
rect 3976 1092 3992 1108
rect 4056 1092 4072 1108
rect 4120 1092 4136 1108
rect 4184 1092 4200 1108
rect 4264 1092 4328 1108
rect 4408 1092 4440 1108
rect 4568 1092 4584 1108
rect 4616 1092 4632 1108
rect 4760 1092 4776 1108
rect 5144 1112 5160 1128
rect 4952 1092 4968 1108
rect 536 1072 552 1088
rect 616 1072 632 1088
rect 680 1072 696 1088
rect 712 1072 728 1088
rect 760 1072 776 1088
rect 1032 1072 1048 1088
rect 1192 1072 1208 1088
rect 1224 1072 1240 1088
rect 1256 1072 1272 1088
rect 1288 1072 1304 1088
rect 1448 1072 1480 1088
rect 1512 1072 1528 1088
rect 1576 1072 1592 1088
rect 1672 1072 1688 1088
rect 1768 1072 1800 1088
rect 1848 1072 1864 1088
rect 2120 1072 2136 1088
rect 2216 1072 2232 1088
rect 2360 1072 2376 1088
rect 2424 1072 2440 1088
rect 2488 1072 2504 1088
rect 2536 1072 2552 1088
rect 2728 1072 2744 1088
rect 2776 1072 2792 1088
rect 2888 1072 2904 1088
rect 2968 1072 2984 1088
rect 3160 1072 3176 1088
rect 3336 1072 3352 1088
rect 3432 1072 3448 1088
rect 3464 1072 3480 1088
rect 3560 1072 3592 1088
rect 3656 1072 3672 1088
rect 3784 1072 3800 1088
rect 3816 1072 3848 1088
rect 4024 1072 4040 1088
rect 4088 1072 4104 1088
rect 4392 1072 4408 1088
rect 4488 1072 4504 1088
rect 4712 1072 4728 1088
rect 4840 1072 4856 1088
rect 4872 1072 4888 1088
rect 4968 1072 4984 1088
rect 5096 1092 5112 1108
rect 5480 1112 5496 1128
rect 5192 1092 5224 1108
rect 5304 1092 5336 1108
rect 5816 1112 5832 1128
rect 5512 1092 5544 1108
rect 5640 1092 5672 1108
rect 5864 1092 5880 1108
rect 5912 1092 5928 1108
rect 6008 1092 6024 1108
rect 6104 1092 6120 1108
rect 6232 1092 6248 1108
rect 6280 1092 6296 1108
rect 6360 1092 6376 1108
rect 6408 1092 6424 1108
rect 6456 1092 6472 1108
rect 6520 1092 6536 1108
rect 6568 1092 6584 1108
rect 6616 1112 6632 1128
rect 6888 1112 6904 1128
rect 6952 1112 6968 1128
rect 7016 1112 7032 1128
rect 7096 1112 7112 1128
rect 7416 1112 7432 1128
rect 6728 1090 6744 1106
rect 7304 1090 7320 1106
rect 7736 1112 7752 1128
rect 7448 1092 7464 1108
rect 7480 1092 7496 1108
rect 7640 1090 7656 1106
rect 7864 1112 7880 1128
rect 8024 1112 8040 1128
rect 7768 1092 7816 1108
rect 7848 1092 7864 1108
rect 7880 1092 7896 1108
rect 7912 1092 7928 1108
rect 7992 1092 8008 1108
rect 5112 1072 5128 1088
rect 5176 1072 5192 1088
rect 5224 1072 5240 1088
rect 5368 1072 5384 1088
rect 5448 1072 5464 1088
rect 5560 1072 5592 1088
rect 5768 1072 5800 1088
rect 5880 1072 5896 1088
rect 6088 1072 6104 1088
rect 6152 1072 6168 1088
rect 6264 1072 6280 1088
rect 6328 1072 6344 1088
rect 6536 1072 6552 1088
rect 6648 1072 6664 1088
rect 6696 1072 6712 1088
rect 6920 1072 6936 1088
rect 6984 1072 7000 1088
rect 7112 1072 7128 1088
rect 7144 1072 7160 1088
rect 7208 1072 7224 1088
rect 7336 1072 7352 1088
rect 7384 1072 7400 1088
rect 7496 1072 7512 1088
rect 7544 1072 7560 1088
rect 7608 1072 7624 1088
rect 7704 1072 7720 1088
rect 7816 1072 7832 1088
rect 7912 1072 7928 1088
rect 8024 1072 8040 1088
rect 88 1052 104 1068
rect 728 1052 744 1068
rect 808 1052 840 1068
rect 1208 1052 1224 1068
rect 1464 1052 1480 1068
rect 1656 1052 1672 1068
rect 1720 1052 1736 1068
rect 2296 1052 2312 1068
rect 3304 1052 3320 1068
rect 3752 1052 3768 1068
rect 3896 1052 3912 1068
rect 3928 1052 3944 1068
rect 4328 1052 4344 1068
rect 4440 1052 4456 1068
rect 5976 1052 5992 1068
rect 6184 1052 6200 1068
rect 6232 1052 6248 1068
rect 6392 1052 6408 1068
rect 6440 1052 6456 1068
rect 6792 1052 6808 1068
rect 6872 1052 6888 1068
rect 7816 1052 7832 1068
rect 7944 1052 7960 1068
rect 408 1032 424 1048
rect 1176 1032 1192 1048
rect 1432 1032 1448 1048
rect 1592 1032 1608 1048
rect 1896 1032 1912 1048
rect 2440 1032 2456 1048
rect 3512 1032 3528 1048
rect 3624 1032 3640 1048
rect 4152 1032 4168 1048
rect 4248 1032 4264 1048
rect 4344 1032 4360 1048
rect 4504 1032 4520 1048
rect 4664 1032 4680 1048
rect 4920 1032 4936 1048
rect 5832 1032 5848 1048
rect 6088 1032 6104 1048
rect 6264 1032 6280 1048
rect 6424 1032 6440 1048
rect 6504 1032 6520 1048
rect 6936 1032 6952 1048
rect 7000 1032 7016 1048
rect 7064 1032 7080 1048
rect 1949 1002 1985 1018
rect 3997 1002 4033 1018
rect 6045 1002 6081 1018
rect 232 972 248 988
rect 424 972 440 988
rect 872 972 888 988
rect 1160 972 1176 988
rect 2296 972 2312 988
rect 2360 972 2376 988
rect 2568 972 2584 988
rect 2600 972 2616 988
rect 2696 972 2712 988
rect 2744 972 2760 988
rect 2808 972 2824 988
rect 2888 972 2904 988
rect 3352 972 3368 988
rect 3928 972 3944 988
rect 4552 972 4568 988
rect 4600 972 4616 988
rect 4952 972 4968 988
rect 5208 972 5224 988
rect 5464 972 5480 988
rect 5736 972 5752 988
rect 6024 972 6040 988
rect 6872 972 6888 988
rect 7256 972 7272 988
rect 7544 972 7560 988
rect 7576 972 7592 988
rect 7832 972 7848 988
rect 56 952 72 968
rect 280 952 296 968
rect 1336 952 1352 968
rect 1400 952 1416 968
rect 1656 952 1672 968
rect 2120 952 2136 968
rect 2216 952 2232 968
rect 2392 952 2424 968
rect 2440 952 2456 968
rect 3160 952 3176 968
rect 3656 952 3672 968
rect 3992 952 4008 968
rect 4120 952 4136 968
rect 4248 952 4264 968
rect 4424 952 4440 968
rect 5080 952 5096 968
rect 5240 952 5256 968
rect 5336 952 5352 968
rect 5480 952 5496 968
rect 5624 952 5640 968
rect 6040 952 6056 968
rect 6200 952 6248 968
rect 6504 952 6520 968
rect 6648 952 6664 968
rect 6680 952 6696 968
rect 7608 952 7624 968
rect 136 932 152 948
rect 312 932 328 948
rect 376 932 392 948
rect 552 932 568 948
rect 808 932 824 948
rect 1192 932 1208 948
rect 1256 932 1288 948
rect 1320 932 1336 948
rect 1384 932 1416 948
rect 1528 932 1544 948
rect 1640 932 1656 948
rect 1768 932 1784 948
rect 1992 932 2008 948
rect 88 912 104 928
rect 152 914 168 930
rect 232 912 248 928
rect 312 912 328 928
rect 392 912 408 928
rect 424 912 440 928
rect 536 912 552 928
rect 616 912 632 928
rect 712 912 728 928
rect 744 912 760 928
rect 904 912 920 928
rect 984 912 1000 928
rect 1032 912 1048 928
rect 1144 912 1160 928
rect 1240 912 1256 928
rect 1304 912 1320 928
rect 1432 912 1464 928
rect 1592 914 1608 930
rect 1816 912 1832 928
rect 1880 914 1896 930
rect 2520 928 2536 944
rect 2664 932 2680 948
rect 2872 932 2888 948
rect 2984 932 3000 948
rect 3240 932 3256 948
rect 3384 932 3400 948
rect 3432 932 3448 948
rect 3480 932 3496 948
rect 4024 932 4040 948
rect 4072 932 4088 948
rect 4568 932 4584 948
rect 5144 932 5160 948
rect 5352 932 5368 948
rect 5432 932 5448 948
rect 5928 932 5944 948
rect 5960 932 5976 948
rect 5992 932 6008 948
rect 6088 932 6104 948
rect 6152 932 6168 948
rect 6264 932 6280 948
rect 6328 932 6344 948
rect 6392 932 6408 948
rect 6424 932 6440 948
rect 6520 932 6536 948
rect 6584 932 6600 948
rect 6696 932 6712 948
rect 6728 932 6744 948
rect 6760 932 6776 948
rect 6824 932 6840 948
rect 6888 932 6904 948
rect 6952 932 6968 948
rect 7080 932 7096 948
rect 7144 932 7160 948
rect 7208 932 7224 948
rect 7272 932 7288 948
rect 7464 932 7480 948
rect 7720 932 7736 948
rect 7832 932 7848 948
rect 8008 932 8024 948
rect 2040 912 2056 928
rect 2136 912 2152 928
rect 2184 912 2200 928
rect 2328 912 2360 928
rect 2440 912 2472 928
rect 2632 912 2648 928
rect 2776 912 2792 928
rect 3064 912 3080 928
rect 3272 912 3288 928
rect 216 892 232 908
rect 408 892 424 908
rect 1000 892 1016 908
rect 1208 892 1224 908
rect 1272 892 1288 908
rect 1336 892 1352 908
rect 1496 892 1512 908
rect 2696 892 2712 908
rect 2792 892 2808 908
rect 2904 892 2920 908
rect 3416 892 3432 908
rect 3464 912 3480 928
rect 3528 912 3544 928
rect 3592 912 3608 928
rect 3624 912 3656 928
rect 3688 912 3704 928
rect 3768 912 3784 928
rect 3816 912 3832 928
rect 3896 912 3912 928
rect 3944 912 3960 928
rect 4120 912 4136 928
rect 4168 912 4184 928
rect 4216 912 4232 928
rect 4296 912 4312 928
rect 4344 912 4360 928
rect 4392 912 4424 928
rect 4456 912 4472 928
rect 4504 912 4536 928
rect 4680 912 4696 928
rect 4728 914 4744 930
rect 4856 912 4872 928
rect 4888 912 4904 928
rect 4984 912 5000 928
rect 5176 912 5192 928
rect 5272 912 5288 928
rect 5608 912 5624 928
rect 5688 912 5704 928
rect 5784 912 5800 928
rect 5832 912 5848 928
rect 5944 912 5960 928
rect 5976 912 5992 928
rect 6008 912 6024 928
rect 6104 912 6120 928
rect 6136 912 6168 928
rect 6248 912 6264 928
rect 6280 912 6296 928
rect 6312 912 6328 928
rect 6456 912 6488 928
rect 6536 912 6584 928
rect 6600 912 6616 928
rect 6648 912 6664 928
rect 6712 912 6728 928
rect 6760 912 6776 928
rect 6792 912 6808 928
rect 6840 912 6856 928
rect 6904 912 6936 928
rect 6984 912 7000 928
rect 7032 912 7064 928
rect 7096 912 7112 928
rect 3544 892 3560 908
rect 3576 892 3592 908
rect 3608 892 3624 908
rect 3672 892 3688 908
rect 3736 892 3752 908
rect 3800 892 3816 908
rect 3880 892 3896 908
rect 4088 892 4104 908
rect 4152 892 4168 908
rect 4232 892 4248 908
rect 4264 892 4280 908
rect 4344 892 4360 908
rect 4952 892 4968 908
rect 5112 892 5144 908
rect 5240 892 5256 908
rect 5336 892 5352 908
rect 5432 892 5448 908
rect 5464 892 5480 908
rect 6296 892 6312 908
rect 6616 892 6632 908
rect 6744 892 6760 908
rect 6808 892 6824 908
rect 6872 892 6888 908
rect 6936 892 6952 908
rect 7400 912 7416 928
rect 7512 912 7528 928
rect 7704 912 7720 928
rect 7896 914 7912 930
rect 7960 912 7976 928
rect 7176 892 7192 908
rect 7240 892 7256 908
rect 248 872 264 888
rect 440 872 456 888
rect 968 872 984 888
rect 1016 872 1032 888
rect 1064 872 1080 888
rect 1688 872 1704 888
rect 3320 872 3336 888
rect 3512 872 3528 888
rect 3704 872 3720 888
rect 3752 872 3768 888
rect 3832 872 3848 888
rect 3912 872 3928 888
rect 3976 872 3992 888
rect 4120 872 4136 888
rect 4152 872 4168 888
rect 4296 872 4312 888
rect 4360 872 4376 888
rect 4456 872 4472 888
rect 984 852 1000 868
rect 6120 852 6136 868
rect 504 832 520 848
rect 584 832 600 848
rect 2744 832 2760 848
rect 3528 832 3544 848
rect 3592 832 3608 848
rect 3688 832 3704 848
rect 3752 832 3768 848
rect 3816 832 3832 848
rect 3896 832 3912 848
rect 4168 832 4184 848
rect 4280 832 4296 848
rect 4344 832 4360 848
rect 4472 832 4488 848
rect 4920 832 4936 848
rect 5208 832 5224 848
rect 5816 832 5832 848
rect 5896 832 5912 848
rect 6168 832 6184 848
rect 6664 832 6680 848
rect 7544 832 7560 848
rect 925 802 961 818
rect 2957 802 2993 818
rect 5021 802 5057 818
rect 7053 802 7089 818
rect 1256 772 1272 788
rect 1528 772 1544 788
rect 1912 772 1928 788
rect 2568 772 2584 788
rect 2904 772 2920 788
rect 3912 772 3928 788
rect 3976 772 3992 788
rect 5080 772 5096 788
rect 6104 772 6120 788
rect 6648 772 6664 788
rect 6760 772 6776 788
rect 7048 772 7064 788
rect 7640 772 7656 788
rect 7704 772 7720 788
rect 1064 752 1080 768
rect 4120 752 4136 768
rect 984 732 1000 748
rect 1016 732 1032 748
rect 1048 732 1064 748
rect 1240 732 1256 748
rect 1272 732 1288 748
rect 1320 732 1336 748
rect 3896 732 3912 748
rect 3960 732 3976 748
rect 4056 732 4072 748
rect 4136 732 4152 748
rect 4184 732 4200 748
rect 6392 732 6408 748
rect 7288 732 7304 748
rect 408 712 424 728
rect 1016 712 1032 728
rect 1080 712 1112 728
rect 1160 712 1176 728
rect 1288 712 1304 728
rect 1372 712 1388 728
rect 1880 712 1896 728
rect 2232 712 2248 728
rect 2648 712 2664 728
rect 2968 712 2984 728
rect 3048 712 3064 728
rect 3112 712 3128 728
rect 88 692 104 708
rect 136 692 152 708
rect 216 692 232 708
rect 248 692 264 708
rect 328 692 344 708
rect 360 692 376 708
rect 424 692 440 708
rect 600 692 616 708
rect 696 692 712 708
rect 760 692 776 708
rect 824 692 840 708
rect 888 692 904 708
rect 1000 692 1016 708
rect 1064 692 1080 708
rect 1128 692 1144 708
rect 1192 692 1208 708
rect 1256 692 1272 708
rect 1304 692 1320 708
rect 1384 692 1400 708
rect 1416 692 1432 708
rect 1480 692 1496 708
rect 1560 692 1576 708
rect 1768 690 1784 706
rect 1848 692 1880 708
rect 2120 690 2136 706
rect 2200 692 2232 708
rect 2360 692 2376 708
rect 2616 692 2648 708
rect 2776 692 2792 708
rect 2888 692 2904 708
rect 2936 692 2952 708
rect 3016 692 3032 708
rect 3352 712 3368 728
rect 3484 712 3500 728
rect 3528 712 3544 728
rect 3548 712 3564 728
rect 3620 712 3636 728
rect 3640 712 3656 728
rect 3752 712 3768 728
rect 3816 712 3832 728
rect 3928 712 3944 728
rect 3992 712 4008 728
rect 4104 712 4120 728
rect 4200 712 4216 728
rect 4296 712 4312 728
rect 4392 712 4408 728
rect 4456 712 4472 728
rect 4536 712 4552 728
rect 4792 712 4824 728
rect 3144 692 3176 708
rect 3256 690 3272 706
rect 3320 692 3336 708
rect 3496 692 3512 708
rect 3560 692 3576 708
rect 3640 692 3656 708
rect 3720 692 3736 708
rect 3768 692 3800 708
rect 3832 692 3848 708
rect 3912 692 3928 708
rect 3960 692 3976 708
rect 4136 692 4152 708
rect 4200 692 4232 708
rect 4312 692 4344 708
rect 4472 692 4488 708
rect 4664 692 4680 708
rect 4840 692 4856 708
rect 4936 692 4952 708
rect 5000 712 5016 728
rect 5304 712 5320 728
rect 5480 712 5496 728
rect 5176 692 5192 708
rect 5416 692 5432 708
rect 5576 712 5592 728
rect 5976 712 5992 728
rect 6216 712 6232 728
rect 6264 712 6280 728
rect 6312 712 6344 728
rect 7112 712 7128 728
rect 7196 712 7212 728
rect 7240 712 7256 728
rect 7800 712 7816 728
rect 7976 712 7992 728
rect 5528 692 5544 708
rect 5656 692 5672 708
rect 5784 692 5800 708
rect 5864 692 5896 708
rect 5928 692 5944 708
rect 6072 692 6104 708
rect 6136 692 6152 708
rect 6280 692 6296 708
rect 6360 692 6376 708
rect 6488 692 6504 708
rect 6616 692 6648 708
rect 6680 692 6696 708
rect 6728 692 6760 708
rect 6792 692 6808 708
rect 6824 692 6840 708
rect 6920 692 6936 708
rect 7016 692 7032 708
rect 7208 692 7224 708
rect 7320 692 7352 708
rect 7512 690 7528 706
rect 7656 692 7704 708
rect 7736 692 7752 708
rect 7928 692 7944 708
rect 248 672 264 688
rect 312 672 328 688
rect 648 672 664 688
rect 712 672 728 688
rect 808 672 824 688
rect 984 672 1000 688
rect 1144 672 1160 688
rect 1208 672 1224 688
rect 1400 672 1416 688
rect 1512 672 1528 688
rect 1592 672 1608 688
rect 1800 672 1816 688
rect 1832 672 1848 688
rect 1912 672 1928 688
rect 2152 672 2168 688
rect 2184 672 2200 688
rect 2280 672 2296 688
rect 2520 672 2536 688
rect 2584 672 2616 688
rect 2744 672 2760 688
rect 2920 672 2936 688
rect 3000 672 3016 688
rect 3080 672 3096 688
rect 3176 672 3192 688
rect 3448 672 3464 688
rect 3512 672 3528 688
rect 3576 672 3608 688
rect 3704 672 3720 688
rect 3768 672 3784 688
rect 3832 672 3848 688
rect 4008 672 4024 688
rect 4088 672 4104 688
rect 4280 672 4296 688
rect 4424 672 4440 688
rect 4680 672 4696 688
rect 4760 672 4776 688
rect 4808 672 4824 688
rect 4920 672 4936 688
rect 4968 672 4984 688
rect 5208 672 5224 688
rect 5352 672 5368 688
rect 5448 672 5464 688
rect 5512 672 5528 688
rect 5560 672 5576 688
rect 5736 672 5752 688
rect 5816 672 5832 688
rect 5944 672 5960 688
rect 6024 672 6040 688
rect 6184 672 6200 688
rect 6232 672 6248 688
rect 6280 672 6296 688
rect 6344 672 6360 688
rect 6376 672 6392 688
rect 6504 672 6520 688
rect 552 652 568 668
rect 792 652 808 668
rect 952 652 968 668
rect 2888 652 2904 668
rect 3256 652 3272 668
rect 3688 652 3704 668
rect 3832 652 3848 668
rect 3864 652 3880 668
rect 4232 652 4248 668
rect 4392 652 4408 668
rect 4904 652 4920 668
rect 5288 652 5304 668
rect 5704 652 5720 668
rect 6856 652 6872 668
rect 6904 672 6920 688
rect 7160 672 7176 688
rect 7224 672 7240 688
rect 7416 672 7432 688
rect 7544 672 7560 688
rect 7768 672 7784 688
rect 7848 672 7864 688
rect 728 632 744 648
rect 856 632 872 648
rect 1096 632 1112 648
rect 1160 632 1176 648
rect 1448 632 1464 648
rect 2904 632 2920 648
rect 3032 632 3048 648
rect 3672 632 3688 648
rect 4536 632 4552 648
rect 4792 632 4808 648
rect 5384 632 5400 648
rect 5960 632 5976 648
rect 6200 632 6216 648
rect 6312 632 6328 648
rect 6904 632 6920 648
rect 7784 632 7800 648
rect 1949 602 1985 618
rect 3997 602 4033 618
rect 6045 602 6081 618
rect 200 572 216 588
rect 920 572 936 588
rect 1256 572 1272 588
rect 1640 572 1656 588
rect 1944 572 1960 588
rect 2264 572 2280 588
rect 2648 572 2664 588
rect 2968 572 2984 588
rect 4152 572 4168 588
rect 4648 572 4664 588
rect 4776 572 4792 588
rect 4840 572 4856 588
rect 6024 572 6040 588
rect 6584 572 6600 588
rect 6648 572 6664 588
rect 7624 572 7640 588
rect 8008 572 8024 588
rect 312 532 344 548
rect 360 552 376 568
rect 1096 552 1112 568
rect 1240 552 1256 568
rect 1368 552 1384 568
rect 1448 552 1464 568
rect 2120 552 2136 568
rect 3048 552 3064 568
rect 3368 552 3384 568
rect 3784 552 3800 568
rect 4184 552 4200 568
rect 4408 552 4424 568
rect 4760 552 4776 568
rect 5432 552 5448 568
rect 5880 552 5896 568
rect 6808 552 6824 568
rect 568 532 584 548
rect 1064 532 1080 548
rect 1352 532 1368 548
rect 1416 532 1432 548
rect 1448 532 1464 548
rect 1672 532 1688 548
rect 1736 532 1752 548
rect 1816 532 1832 548
rect 1864 532 1880 548
rect 1928 532 1944 548
rect 2024 532 2040 548
rect 2056 532 2072 548
rect 2088 532 2120 548
rect 2328 532 2344 548
rect 88 512 104 528
rect 136 512 152 528
rect 232 512 248 528
rect 296 512 312 528
rect 392 512 408 528
rect 440 512 456 528
rect 488 512 504 528
rect 568 512 584 528
rect 616 512 632 528
rect 680 512 696 528
rect 792 514 808 530
rect 840 512 856 528
rect 1032 514 1048 530
rect 1240 512 1256 528
rect 1336 512 1352 528
rect 1400 512 1416 528
rect 1480 512 1496 528
rect 1624 512 1640 528
rect 1720 512 1736 528
rect 1768 512 1784 528
rect 1848 512 1864 528
rect 1896 512 1928 528
rect 2136 512 2168 528
rect 2296 512 2312 528
rect 2376 512 2392 528
rect 2504 532 2520 548
rect 2616 532 2632 548
rect 2680 532 2696 548
rect 2728 532 2744 548
rect 3032 532 3048 548
rect 3096 532 3112 548
rect 3128 532 3144 548
rect 3160 532 3176 548
rect 3224 532 3240 548
rect 3272 532 3288 548
rect 3496 532 3512 548
rect 3576 532 3592 548
rect 3704 532 3720 548
rect 3768 532 3784 548
rect 4280 532 4296 548
rect 4344 532 4360 548
rect 4376 532 4392 548
rect 4504 532 4520 548
rect 4600 532 4616 548
rect 4712 532 4744 548
rect 4824 532 4840 548
rect 5016 532 5032 548
rect 5064 532 5080 548
rect 5096 532 5112 548
rect 5144 532 5160 548
rect 5208 532 5240 548
rect 5272 532 5288 548
rect 5320 532 5352 548
rect 5368 532 5384 548
rect 5528 532 5544 548
rect 5560 532 5576 548
rect 5640 532 5656 548
rect 5672 532 5688 548
rect 5736 532 5752 548
rect 5784 532 5800 548
rect 6008 532 6024 548
rect 6088 532 6104 548
rect 6184 532 6200 548
rect 6312 532 6328 548
rect 6376 532 6392 548
rect 6472 532 6488 548
rect 6712 532 6728 548
rect 6952 532 6984 548
rect 7016 532 7032 548
rect 7064 532 7080 548
rect 7288 532 7304 548
rect 7320 532 7336 548
rect 7368 532 7384 548
rect 7416 532 7432 548
rect 7800 532 7816 548
rect 7848 532 7864 548
rect 7896 532 7912 548
rect 2488 512 2504 528
rect 248 472 264 488
rect 424 472 440 488
rect 472 492 488 508
rect 440 452 456 468
rect 504 472 520 488
rect 552 472 568 488
rect 600 492 616 508
rect 664 492 680 508
rect 1304 492 1320 508
rect 1368 492 1384 508
rect 1688 492 1704 508
rect 1752 492 1768 508
rect 1880 492 1896 508
rect 1992 492 2008 508
rect 2040 492 2056 508
rect 2552 492 2568 508
rect 2600 512 2616 528
rect 2760 514 2776 530
rect 3080 512 3096 528
rect 3192 512 3208 528
rect 3304 514 3320 530
rect 3560 512 3576 528
rect 3640 512 3656 528
rect 3736 512 3768 528
rect 3864 512 3896 528
rect 4040 512 4056 528
rect 4072 512 4088 528
rect 4104 512 4120 528
rect 4152 512 4168 528
rect 4216 512 4232 528
rect 4264 512 4280 528
rect 2588 492 2604 508
rect 2632 492 2648 508
rect 2904 492 2920 508
rect 3000 492 3016 508
rect 3032 492 3048 508
rect 3160 492 3176 508
rect 3224 492 3240 508
rect 3464 492 3480 508
rect 3544 492 3560 508
rect 3656 492 3672 508
rect 4040 492 4056 508
rect 4312 492 4328 508
rect 4360 512 4376 528
rect 4488 512 4504 528
rect 4616 512 4632 528
rect 4808 512 4824 528
rect 4920 512 4936 528
rect 4968 512 4984 528
rect 4680 492 4696 508
rect 4776 492 4792 508
rect 5128 492 5144 508
rect 5176 512 5192 528
rect 5256 492 5272 508
rect 5304 512 5320 528
rect 5352 512 5368 528
rect 5464 512 5480 528
rect 5608 512 5624 528
rect 5672 512 5688 528
rect 5816 514 5832 530
rect 5976 512 6008 528
rect 6168 512 6184 528
rect 6280 512 6312 528
rect 6360 512 6376 528
rect 6456 514 6472 530
rect 6616 512 6632 528
rect 6744 514 6760 530
rect 6904 512 6920 528
rect 6984 512 7000 528
rect 5384 492 5400 508
rect 5496 492 5528 508
rect 5656 492 5688 508
rect 5736 492 5752 508
rect 5960 492 5976 508
rect 6264 492 6280 508
rect 6328 492 6344 508
rect 6348 492 6364 508
rect 7208 512 7224 528
rect 7336 512 7352 528
rect 7448 514 7464 530
rect 7656 512 7672 528
rect 7768 512 7784 528
rect 7880 514 7896 530
rect 7032 492 7048 508
rect 7368 492 7384 508
rect 7800 492 7816 508
rect 632 472 648 488
rect 696 472 712 488
rect 1128 472 1144 488
rect 1784 472 1800 488
rect 2200 472 2216 488
rect 3144 472 3160 488
rect 4104 472 4120 488
rect 4216 472 4232 488
rect 1528 452 1544 468
rect 232 432 248 448
rect 680 432 696 448
rect 2392 432 2408 448
rect 3608 432 3624 448
rect 4056 432 4072 448
rect 4120 432 4136 448
rect 4232 432 4248 448
rect 7576 432 7592 448
rect 7720 432 7736 448
rect 925 402 961 418
rect 2957 402 2993 418
rect 5021 402 5057 418
rect 7053 402 7089 418
rect 168 372 184 388
rect 248 372 264 388
rect 312 372 328 388
rect 360 372 376 388
rect 456 372 472 388
rect 552 372 568 388
rect 600 372 616 388
rect 1144 372 1160 388
rect 1304 372 1320 388
rect 1352 372 1368 388
rect 1432 372 1448 388
rect 2136 372 2152 388
rect 2536 372 2552 388
rect 3000 372 3016 388
rect 3544 372 3560 388
rect 3672 372 3688 388
rect 5368 372 5384 388
rect 5880 372 5896 388
rect 6344 372 6360 388
rect 6600 372 6616 388
rect 6904 372 6920 388
rect 7000 372 7016 388
rect 7432 372 7448 388
rect 7992 372 8008 388
rect 40 352 56 368
rect 1048 352 1064 368
rect 2424 352 2440 368
rect 3432 352 3448 368
rect 24 332 40 348
rect 104 332 120 348
rect 152 332 168 348
rect 232 332 248 348
rect 296 332 312 348
rect 344 332 360 348
rect 424 332 456 348
rect 472 332 488 348
rect 536 332 552 348
rect 616 332 632 348
rect 1032 332 1048 348
rect 1064 332 1080 348
rect 1288 332 1304 348
rect 1320 332 1336 348
rect 1416 332 1432 348
rect 56 312 72 328
rect 184 312 216 328
rect 264 312 280 328
rect 376 312 392 328
rect 504 312 520 328
rect 1064 312 1080 328
rect 1320 312 1336 328
rect 1448 312 1464 328
rect 40 292 56 308
rect 104 292 136 308
rect 168 292 184 308
rect 216 292 232 308
rect 280 292 296 308
rect 360 292 376 308
rect 408 292 424 308
rect 488 292 504 308
rect 552 292 568 308
rect 584 292 616 308
rect 664 292 680 308
rect 728 292 744 308
rect 920 290 936 306
rect 1048 292 1064 308
rect 1096 292 1112 308
rect 1160 292 1176 308
rect 1224 292 1240 308
rect 1304 292 1320 308
rect 1352 292 1368 308
rect 1432 292 1448 308
rect 1496 292 1512 308
rect 1576 292 1592 308
rect 1720 292 1736 308
rect 1848 292 1896 308
rect 1928 312 1944 328
rect 2056 312 2072 328
rect 2696 312 2712 328
rect 2088 292 2120 308
rect 2280 292 2296 308
rect 2632 292 2648 308
rect 3112 312 3128 328
rect 3272 312 3288 328
rect 3352 312 3368 328
rect 3640 312 3656 328
rect 3880 312 3896 328
rect 3960 312 3976 328
rect 2728 292 2760 308
rect 2840 290 2856 306
rect 3192 292 3208 308
rect 3304 292 3320 308
rect 3464 292 3480 308
rect 3592 292 3608 308
rect 3688 292 3704 308
rect 3720 292 3736 308
rect 3816 292 3832 308
rect 3880 292 3912 308
rect 3992 292 4008 308
rect 4056 292 4072 308
rect 4120 292 4136 308
rect 4232 292 4248 308
rect 4264 292 4280 308
rect 4328 312 4344 328
rect 4376 312 4392 328
rect 4520 312 4536 328
rect 4392 292 4408 308
rect 4424 292 4440 308
rect 4616 312 4632 328
rect 4680 312 4696 328
rect 4888 312 4904 328
rect 104 272 120 288
rect 680 272 696 288
rect 712 272 728 288
rect 952 272 968 288
rect 1176 272 1192 288
rect 1560 272 1576 288
rect 1640 272 1656 288
rect 1768 272 1784 288
rect 1816 272 1832 288
rect 2024 272 2040 288
rect 2328 272 2344 288
rect 2472 272 2488 288
rect 2552 272 2568 288
rect 2664 272 2680 288
rect 2760 272 2776 288
rect 2808 272 2824 288
rect 2904 272 2920 288
rect 3240 272 3256 288
rect 3272 272 3288 288
rect 3320 272 3352 288
rect 3384 272 3416 288
rect 3496 272 3512 288
rect 3704 272 3720 288
rect 3848 272 3864 288
rect 4008 272 4024 288
rect 4248 272 4264 288
rect 4360 272 4376 288
rect 4440 272 4456 288
rect 4584 292 4600 308
rect 4760 292 4776 308
rect 4936 292 4952 308
rect 5112 292 5128 308
rect 5192 292 5208 308
rect 5224 292 5256 308
rect 5288 312 5304 328
rect 5400 312 5416 328
rect 5468 312 5484 328
rect 5512 312 5528 328
rect 5960 312 5976 328
rect 6728 312 6744 328
rect 7016 312 7032 328
rect 5480 292 5496 308
rect 5528 292 5560 308
rect 5704 292 5736 308
rect 5848 292 5864 308
rect 5992 292 6008 308
rect 6200 292 6216 308
rect 6328 292 6344 308
rect 6376 292 6408 308
rect 6520 292 6536 308
rect 6632 292 6664 308
rect 6776 292 6792 308
rect 6824 292 6856 308
rect 6888 292 6904 308
rect 6936 292 6952 308
rect 7048 292 7064 308
rect 7128 312 7144 328
rect 7544 312 7560 328
rect 7272 292 7288 308
rect 7416 292 7432 308
rect 7464 292 7496 308
rect 7656 312 7672 328
rect 7592 292 7608 308
rect 7784 312 7800 328
rect 7704 292 7720 308
rect 7752 292 7784 308
rect 7864 290 7880 306
rect 4472 272 4488 288
rect 4520 272 4536 288
rect 4552 272 4584 288
rect 4808 272 4824 288
rect 4856 272 4872 288
rect 4904 272 4920 288
rect 5000 272 5016 288
rect 5064 272 5080 288
rect 5208 272 5224 288
rect 5320 272 5336 288
rect 760 252 776 268
rect 856 252 872 268
rect 1256 252 1272 268
rect 1464 252 1480 268
rect 1544 252 1560 268
rect 3016 252 3032 268
rect 3048 252 3064 268
rect 5432 272 5448 288
rect 5496 272 5512 288
rect 5608 272 5624 288
rect 5832 272 5848 288
rect 6152 272 6168 288
rect 6440 272 6456 288
rect 6472 272 6488 288
rect 6600 272 6632 288
rect 6696 272 6712 288
rect 6760 272 6776 288
rect 6984 272 7000 288
rect 7032 272 7048 288
rect 7128 272 7144 288
rect 7160 272 7176 288
rect 7288 272 7304 288
rect 7400 272 7416 288
rect 7512 272 7528 288
rect 7608 272 7640 288
rect 7720 272 7736 288
rect 7896 272 7912 288
rect 5624 252 5640 268
rect 5944 252 5960 268
rect 6024 252 6040 268
rect 1192 232 1208 248
rect 3624 232 3640 248
rect 3752 232 3768 248
rect 3784 232 3800 248
rect 3944 232 3976 248
rect 4120 232 4136 248
rect 4184 232 4216 248
rect 4296 232 4312 248
rect 4616 232 4632 248
rect 7560 232 7576 248
rect 7672 232 7688 248
rect 7992 232 8008 248
rect 1949 202 1985 218
rect 3997 202 4033 218
rect 6045 202 6081 218
rect 872 172 888 188
rect 968 172 984 188
rect 1336 172 1352 188
rect 1736 172 1752 188
rect 1928 172 1944 188
rect 2792 172 2808 188
rect 2856 172 2872 188
rect 3480 172 3496 188
rect 3720 172 3736 188
rect 3848 172 3864 188
rect 4440 172 4456 188
rect 4744 172 4760 188
rect 5000 172 5016 188
rect 5080 172 5096 188
rect 6360 172 6376 188
rect 6456 172 6472 188
rect 7544 172 7560 188
rect 7752 172 7768 188
rect 7976 172 7992 188
rect 56 152 72 168
rect 248 152 264 168
rect 136 132 152 148
rect 376 152 392 168
rect 312 132 328 148
rect 600 152 616 168
rect 152 114 168 130
rect 216 112 232 128
rect 248 112 264 128
rect 328 112 344 128
rect 440 132 456 148
rect 504 132 520 148
rect 776 132 792 148
rect 952 132 968 148
rect 1000 152 1016 168
rect 1256 152 1272 168
rect 2360 152 2376 168
rect 4472 152 4488 168
rect 4616 152 4632 168
rect 5528 152 5544 168
rect 5736 152 5752 168
rect 6072 152 6088 168
rect 6696 152 6712 168
rect 6760 152 6776 168
rect 6968 152 6984 168
rect 7400 152 7416 168
rect 7464 152 7480 168
rect 7896 152 7912 168
rect 7992 152 8008 168
rect 1080 132 1096 148
rect 1128 132 1144 148
rect 1256 132 1272 148
rect 1496 132 1512 148
rect 1592 132 1608 148
rect 1704 132 1720 148
rect 1896 132 1912 148
rect 2184 132 2200 148
rect 2216 132 2232 148
rect 2328 132 2344 148
rect 2504 132 2520 148
rect 2600 132 2616 148
rect 2632 132 2648 148
rect 2712 132 2744 148
rect 2840 132 2856 148
rect 2936 132 2952 148
rect 3064 132 3080 148
rect 3112 132 3128 148
rect 3208 132 3224 148
rect 424 112 440 128
rect 472 112 488 128
rect 536 114 552 130
rect 744 114 760 130
rect 888 112 904 128
rect 1032 112 1048 128
rect 1112 112 1128 128
rect 1192 114 1208 130
rect 1512 112 1528 128
rect 1608 112 1640 128
rect 1848 112 1864 128
rect 2152 114 2168 130
rect 2232 112 2248 128
rect 1672 92 1688 108
rect 2244 92 2260 108
rect 2536 114 2552 130
rect 2616 112 2632 128
rect 2280 92 2296 108
rect 2680 92 2696 108
rect 2968 92 2984 108
rect 3032 112 3064 128
rect 3144 114 3160 130
rect 3496 132 3512 148
rect 3560 132 3576 148
rect 3976 132 3992 148
rect 4328 132 4344 148
rect 4520 132 4536 148
rect 4920 132 4936 148
rect 5176 132 5192 148
rect 5464 132 5496 148
rect 5560 132 5576 148
rect 5624 132 5640 148
rect 5720 132 5736 148
rect 5848 132 5864 148
rect 5992 132 6008 148
rect 6104 132 6120 148
rect 6216 132 6232 148
rect 6312 132 6328 148
rect 6408 132 6424 148
rect 6504 132 6520 148
rect 6568 132 6584 148
rect 6616 132 6632 148
rect 6888 132 6904 148
rect 6920 132 6936 148
rect 6952 132 6968 148
rect 7176 132 7192 148
rect 7224 132 7240 148
rect 7320 132 7336 148
rect 7720 132 7736 148
rect 7832 132 7848 148
rect 3432 112 3448 128
rect 3512 112 3528 128
rect 3608 112 3640 128
rect 3688 112 3704 128
rect 3752 112 3768 128
rect 3800 112 3816 128
rect 3960 112 3976 128
rect 4120 112 4136 128
rect 4168 112 4184 128
rect 4216 112 4232 128
rect 4264 112 4296 128
rect 4344 112 4360 128
rect 4392 112 4408 128
rect 4552 114 4568 130
rect 4728 112 4744 128
rect 4840 112 4856 128
rect 4968 112 4984 128
rect 5208 114 5224 130
rect 5384 112 5400 128
rect 5496 112 5512 128
rect 3320 92 3336 108
rect 3464 92 3480 108
rect 5592 92 5608 108
rect 5656 92 5672 108
rect 5688 112 5720 128
rect 5832 112 5848 128
rect 6040 112 6056 128
rect 6200 112 6216 128
rect 6328 112 6344 128
rect 5960 92 5976 108
rect 6028 92 6044 108
rect 6488 112 6504 128
rect 6520 112 6536 128
rect 6376 92 6392 108
rect 6712 112 6728 128
rect 6936 112 6952 128
rect 7096 112 7112 128
rect 6584 92 6600 108
rect 6856 92 6872 108
rect 7256 92 7272 108
rect 7288 112 7320 128
rect 7416 112 7432 128
rect 7640 112 7656 128
rect 7864 112 7880 128
rect 3336 32 3352 48
rect 3576 32 3592 48
rect 3656 32 3672 48
rect 3784 32 3800 48
rect 3832 32 3848 48
rect 4088 32 4104 48
rect 4136 32 4152 48
rect 4184 32 4200 48
rect 4232 32 4248 48
rect 4376 32 4392 48
rect 4424 32 4440 48
rect 4696 32 4712 48
rect 925 2 961 18
rect 2957 2 2993 18
rect 5021 2 5057 18
rect 7053 2 7089 18
<< metal2 >>
rect 77 5488 83 5492
rect 45 5328 51 5432
rect 141 5388 147 5452
rect 189 5348 195 5492
rect 237 5488 243 5490
rect 157 5330 163 5332
rect 45 5088 51 5312
rect 29 4708 35 5012
rect 45 4988 51 5032
rect 77 4928 83 5232
rect 93 5108 99 5112
rect 45 4708 51 4832
rect 93 4708 99 5072
rect 93 4688 99 4692
rect 45 4548 51 4552
rect 77 4530 83 4672
rect 29 4088 35 4372
rect 45 4128 51 4272
rect 61 4163 67 4252
rect 61 4157 72 4163
rect 109 4128 115 5312
rect 221 5088 227 5092
rect 157 4908 163 4952
rect 253 4948 259 5052
rect 173 4883 179 4912
rect 157 4877 179 4883
rect 125 4708 131 4832
rect 141 4748 147 4752
rect 141 4728 147 4732
rect 157 4708 163 4877
rect 189 4828 195 4872
rect 205 4808 211 4832
rect 173 4748 179 4752
rect 125 4508 131 4652
rect 157 4628 163 4692
rect 141 4288 147 4512
rect 173 4388 179 4732
rect 205 4728 211 4732
rect 221 4708 227 4912
rect 269 4908 275 5352
rect 349 5328 355 5392
rect 397 5388 403 5472
rect 429 5368 435 5372
rect 509 5368 515 5432
rect 525 5388 531 5492
rect 653 5488 659 5490
rect 637 5348 643 5472
rect 733 5408 739 5492
rect 749 5488 755 5492
rect 381 5328 387 5332
rect 509 5328 515 5332
rect 333 5028 339 5312
rect 349 5108 355 5312
rect 381 5048 387 5072
rect 445 4948 451 5072
rect 461 4988 467 5092
rect 477 4988 483 5312
rect 733 5148 739 5312
rect 589 5088 595 5092
rect 477 4948 483 4972
rect 541 4968 547 5032
rect 253 4788 259 4832
rect 285 4748 291 4772
rect 221 4688 227 4692
rect 189 4528 195 4632
rect 237 4488 243 4692
rect 301 4608 307 4872
rect 317 4868 323 4872
rect 381 4863 387 4912
rect 365 4857 387 4863
rect 365 4788 371 4857
rect 317 4708 323 4712
rect 349 4648 355 4732
rect 397 4728 403 4932
rect 429 4928 435 4932
rect 445 4928 451 4932
rect 413 4788 419 4892
rect 493 4748 499 4792
rect 541 4788 547 4952
rect 621 4948 627 5052
rect 541 4748 547 4752
rect 557 4748 563 4752
rect 365 4688 371 4692
rect 365 4528 371 4672
rect 381 4588 387 4692
rect 397 4503 403 4712
rect 429 4708 435 4732
rect 413 4688 419 4692
rect 429 4548 435 4612
rect 461 4588 467 4712
rect 477 4708 483 4732
rect 541 4628 547 4692
rect 621 4688 627 4932
rect 637 4928 643 4932
rect 765 4928 771 5012
rect 781 4948 787 5492
rect 797 5008 803 5452
rect 845 5348 851 5492
rect 829 5068 835 5312
rect 829 5028 835 5052
rect 861 4968 867 5052
rect 781 4928 787 4932
rect 429 4528 435 4532
rect 397 4497 408 4503
rect 349 4468 355 4472
rect 333 4457 344 4463
rect 237 4348 243 4372
rect 253 4328 259 4352
rect 317 4328 323 4332
rect 13 3948 19 4032
rect 13 3528 19 3532
rect 29 3348 35 3932
rect 45 3908 51 4112
rect 61 4108 67 4112
rect 93 3928 99 3932
rect 45 3888 51 3892
rect 45 3768 51 3872
rect 61 3788 67 3912
rect 109 3908 115 3932
rect 93 3888 99 3892
rect 61 3768 67 3772
rect 93 3588 99 3752
rect 125 3543 131 4112
rect 141 3748 147 4272
rect 157 4188 163 4290
rect 237 4288 243 4292
rect 253 4288 259 4292
rect 173 3968 179 4132
rect 221 4128 227 4232
rect 253 4228 259 4272
rect 301 4248 307 4292
rect 189 4008 195 4112
rect 157 3928 163 3932
rect 173 3888 179 3892
rect 189 3868 195 3912
rect 205 3788 211 3912
rect 221 3908 227 4112
rect 237 4088 243 4092
rect 253 3988 259 4072
rect 221 3768 227 3772
rect 157 3730 163 3752
rect 253 3728 259 3952
rect 301 3948 307 4072
rect 317 3988 323 4092
rect 333 4088 339 4457
rect 397 4388 403 4432
rect 429 4348 435 4352
rect 445 4348 451 4372
rect 349 4188 355 4312
rect 365 4308 371 4332
rect 365 4128 371 4272
rect 413 4268 419 4312
rect 429 4248 435 4292
rect 365 3988 371 4072
rect 269 3868 275 3912
rect 109 3537 131 3543
rect 93 3368 99 3432
rect 109 3348 115 3537
rect 125 3508 131 3512
rect 141 3508 147 3532
rect 189 3508 195 3632
rect 237 3508 243 3532
rect 253 3448 259 3712
rect 285 3708 291 3892
rect 301 3848 307 3932
rect 349 3928 355 3932
rect 365 3908 371 3952
rect 381 3928 387 4092
rect 445 3948 451 4332
rect 477 4248 483 4512
rect 493 4488 499 4592
rect 493 4388 499 4472
rect 509 4388 515 4412
rect 541 4408 547 4492
rect 557 4448 563 4472
rect 573 4428 579 4512
rect 669 4508 675 4772
rect 685 4528 691 4612
rect 749 4548 755 4652
rect 797 4588 803 4612
rect 637 4468 643 4472
rect 493 4368 499 4372
rect 493 4328 499 4332
rect 525 4328 531 4392
rect 621 4348 627 4352
rect 669 4328 675 4392
rect 685 4323 691 4472
rect 685 4317 707 4323
rect 317 3728 323 3732
rect 301 3588 307 3672
rect 269 3488 275 3492
rect 189 3328 195 3332
rect 221 3328 227 3332
rect 317 3328 323 3352
rect 77 3263 83 3312
rect 61 3257 83 3263
rect 45 3148 51 3232
rect 29 3088 35 3112
rect 61 3083 67 3257
rect 157 3188 163 3252
rect 77 3108 83 3152
rect 93 3088 99 3092
rect 61 3077 83 3083
rect 29 2968 35 3072
rect 77 2988 83 3077
rect 109 3068 115 3112
rect 125 2968 131 3152
rect 141 3148 147 3152
rect 205 3148 211 3312
rect 253 3268 259 3272
rect 157 3108 163 3132
rect 173 3108 179 3112
rect 157 2948 163 3092
rect 173 3008 179 3092
rect 173 2968 179 2972
rect 189 2968 195 3112
rect 205 2968 211 2992
rect 45 2588 51 2932
rect 61 2483 67 2832
rect 157 2648 163 2690
rect 189 2688 195 2732
rect 221 2668 227 3032
rect 285 2988 291 3092
rect 301 3048 307 3292
rect 333 3268 339 3272
rect 317 3108 323 3252
rect 301 2928 307 2932
rect 301 2788 307 2912
rect 253 2708 259 2712
rect 173 2528 179 2592
rect 221 2588 227 2632
rect 237 2568 243 2632
rect 77 2508 83 2512
rect 61 2477 83 2483
rect 13 2328 19 2332
rect 45 1908 51 2432
rect 77 1968 83 2477
rect 125 2308 131 2312
rect 141 2308 147 2472
rect 157 2288 163 2292
rect 173 2288 179 2512
rect 205 2448 211 2532
rect 253 2528 259 2692
rect 269 2308 275 2672
rect 221 2257 232 2263
rect 173 2128 179 2232
rect 221 2188 227 2257
rect 141 2088 147 2112
rect 77 1908 83 1952
rect 45 1808 51 1832
rect 93 1788 99 1872
rect 109 1788 115 1832
rect 45 1768 51 1772
rect 109 1728 115 1732
rect 125 1728 131 1852
rect 109 1588 115 1712
rect 61 968 67 1112
rect 77 1003 83 1452
rect 93 1388 99 1492
rect 109 1348 115 1572
rect 141 1508 147 2072
rect 157 1688 163 1792
rect 173 1728 179 1892
rect 189 1888 195 1892
rect 189 1708 195 1772
rect 221 1743 227 2032
rect 285 1948 291 2232
rect 301 2148 307 2732
rect 317 2508 323 2972
rect 349 2948 355 3892
rect 365 3628 371 3892
rect 381 3888 387 3912
rect 429 3868 435 3872
rect 397 3768 403 3852
rect 413 3828 419 3832
rect 477 3748 483 4112
rect 493 4108 499 4312
rect 509 4288 515 4292
rect 509 3988 515 4112
rect 541 4088 547 4312
rect 605 4268 611 4312
rect 621 4228 627 4292
rect 685 4228 691 4292
rect 701 4148 707 4317
rect 717 4308 723 4432
rect 749 4357 787 4363
rect 749 4348 755 4357
rect 781 4343 787 4357
rect 813 4348 819 4732
rect 829 4728 835 4952
rect 877 4788 883 4952
rect 893 4868 899 5352
rect 973 5348 979 5472
rect 989 5408 995 5492
rect 973 5328 979 5332
rect 1101 5328 1107 5472
rect 1325 5388 1331 5492
rect 1229 5348 1235 5352
rect 957 5048 963 5090
rect 989 5088 995 5132
rect 989 4988 995 5032
rect 1021 4988 1027 5212
rect 1101 5148 1107 5312
rect 1165 5308 1171 5314
rect 1309 5308 1315 5312
rect 1309 5288 1315 5292
rect 1133 5108 1139 5112
rect 1069 5088 1075 5092
rect 1133 5088 1139 5092
rect 1165 5088 1171 5232
rect 1341 5088 1347 5472
rect 1373 5348 1379 5452
rect 1437 5388 1443 5472
rect 1565 5468 1571 5490
rect 1677 5488 1683 5663
rect 1805 5508 1811 5663
rect 1501 5368 1507 5452
rect 1597 5388 1603 5452
rect 1677 5448 1683 5472
rect 1485 5348 1491 5352
rect 1357 5248 1363 5332
rect 1469 5268 1475 5312
rect 1373 5106 1379 5112
rect 1469 5108 1475 5112
rect 1005 4928 1011 4932
rect 1021 4928 1027 4972
rect 1069 4928 1075 4932
rect 1085 4908 1091 4912
rect 1005 4748 1011 4852
rect 973 4728 979 4732
rect 1005 4728 1011 4732
rect 1101 4728 1107 5072
rect 1181 5048 1187 5072
rect 1181 4963 1187 5032
rect 1165 4957 1187 4963
rect 1165 4928 1171 4957
rect 1192 4937 1203 4943
rect 1149 4728 1155 4752
rect 1021 4708 1027 4712
rect 781 4337 792 4343
rect 733 4188 739 4252
rect 749 4228 755 4292
rect 669 4088 675 4112
rect 557 3968 563 3992
rect 557 3908 563 3952
rect 541 3888 547 3892
rect 557 3768 563 3812
rect 429 3728 435 3732
rect 493 3730 499 3732
rect 381 3508 387 3652
rect 445 3588 451 3612
rect 397 3508 403 3512
rect 461 3488 467 3692
rect 589 3588 595 3992
rect 701 3928 707 4132
rect 733 4108 739 4112
rect 605 3748 611 3892
rect 621 3788 627 3892
rect 621 3728 627 3772
rect 637 3768 643 3892
rect 701 3730 707 3832
rect 541 3488 547 3492
rect 381 3308 387 3312
rect 397 3288 403 3312
rect 429 3308 435 3332
rect 461 3328 467 3472
rect 472 3277 483 3283
rect 381 3123 387 3232
rect 445 3128 451 3232
rect 461 3188 467 3212
rect 477 3148 483 3277
rect 493 3188 499 3392
rect 573 3188 579 3312
rect 589 3288 595 3432
rect 653 3388 659 3392
rect 669 3328 675 3432
rect 701 3323 707 3492
rect 717 3348 723 4032
rect 765 4008 771 4332
rect 797 4308 803 4312
rect 813 4308 819 4312
rect 797 4128 803 4212
rect 781 3948 787 4032
rect 749 3828 755 3892
rect 797 3868 803 4092
rect 813 4088 819 4232
rect 829 4228 835 4692
rect 893 4528 899 4632
rect 845 4448 851 4512
rect 861 4388 867 4432
rect 877 4288 883 4452
rect 893 4388 899 4512
rect 909 4348 915 4692
rect 1021 4628 1027 4672
rect 957 4528 963 4572
rect 1069 4548 1075 4592
rect 1133 4568 1139 4672
rect 1181 4568 1187 4692
rect 1197 4688 1203 4937
rect 1229 4848 1235 4912
rect 1309 4908 1315 4912
rect 1389 4908 1395 4912
rect 1405 4908 1411 4992
rect 1325 4868 1331 4872
rect 1197 4648 1203 4672
rect 1245 4663 1251 4672
rect 1277 4663 1283 4672
rect 1245 4657 1283 4663
rect 1197 4548 1203 4572
rect 1309 4563 1315 4732
rect 1325 4683 1331 4852
rect 1341 4748 1347 4832
rect 1341 4708 1347 4712
rect 1325 4677 1347 4683
rect 1309 4557 1331 4563
rect 1005 4528 1011 4532
rect 1021 4528 1027 4532
rect 1085 4528 1091 4532
rect 1293 4528 1299 4532
rect 989 4388 995 4492
rect 973 4348 979 4352
rect 925 4308 931 4312
rect 877 4128 883 4132
rect 845 4088 851 4092
rect 765 3768 771 3852
rect 765 3528 771 3712
rect 781 3488 787 3532
rect 701 3317 723 3323
rect 637 3248 643 3312
rect 669 3188 675 3292
rect 717 3268 723 3317
rect 733 3188 739 3192
rect 653 3148 659 3152
rect 381 3117 392 3123
rect 413 3108 419 3112
rect 669 3108 675 3152
rect 365 3088 371 3092
rect 397 2928 403 3092
rect 541 3068 547 3072
rect 333 2708 339 2752
rect 365 2728 371 2832
rect 333 2588 339 2672
rect 349 2568 355 2632
rect 365 2548 371 2712
rect 397 2548 403 2912
rect 413 2908 419 2912
rect 317 2328 323 2492
rect 365 2488 371 2512
rect 317 2308 323 2312
rect 317 2128 323 2132
rect 333 1948 339 2432
rect 365 2288 371 2292
rect 381 1908 387 2532
rect 413 2388 419 2432
rect 429 2388 435 2932
rect 541 2928 547 2972
rect 445 2528 451 2592
rect 461 2528 467 2912
rect 557 2748 563 2932
rect 589 2848 595 3072
rect 701 2963 707 3112
rect 765 3108 771 3452
rect 781 3288 787 3472
rect 797 3328 803 3572
rect 813 3548 819 4072
rect 877 3928 883 4032
rect 909 3848 915 4232
rect 925 4128 931 4292
rect 1005 4268 1011 4512
rect 1037 4497 1048 4503
rect 1037 4388 1043 4497
rect 1133 4388 1139 4492
rect 1197 4388 1203 4512
rect 1325 4508 1331 4557
rect 1341 4508 1347 4677
rect 1357 4528 1363 4892
rect 1373 4848 1379 4872
rect 1389 4828 1395 4832
rect 1405 4728 1411 4732
rect 1389 4688 1395 4712
rect 1389 4608 1395 4672
rect 1421 4608 1427 4872
rect 1453 4708 1459 5072
rect 1485 4983 1491 5332
rect 1629 5328 1635 5332
rect 1501 5288 1507 5312
rect 1565 5228 1571 5312
rect 1645 5308 1651 5432
rect 1693 5388 1699 5472
rect 1517 5108 1523 5112
rect 1517 4988 1523 5092
rect 1549 5088 1555 5172
rect 1565 5088 1571 5212
rect 1485 4977 1507 4983
rect 1469 4728 1475 4792
rect 1501 4708 1507 4977
rect 1565 4948 1571 5032
rect 1517 4928 1523 4932
rect 1533 4728 1539 4932
rect 1581 4908 1587 4912
rect 1565 4868 1571 4872
rect 1581 4868 1587 4892
rect 1437 4677 1448 4683
rect 1437 4628 1443 4677
rect 1421 4528 1427 4552
rect 1437 4548 1443 4612
rect 1453 4548 1459 4572
rect 1469 4568 1475 4632
rect 1517 4548 1523 4672
rect 1533 4548 1539 4712
rect 1437 4528 1443 4532
rect 1357 4508 1363 4512
rect 1549 4508 1555 4792
rect 1581 4728 1587 4832
rect 1613 4768 1619 4832
rect 1597 4668 1603 4692
rect 1613 4688 1619 4692
rect 1213 4388 1219 4492
rect 1117 4348 1123 4352
rect 1021 4168 1027 4312
rect 1037 4228 1043 4292
rect 941 4108 947 4112
rect 973 3948 979 4032
rect 941 3928 947 3932
rect 973 3908 979 3932
rect 1037 3908 1043 3932
rect 1053 3888 1059 3912
rect 1069 3888 1075 3892
rect 925 3868 931 3872
rect 845 3788 851 3792
rect 861 3748 867 3832
rect 877 3728 883 3792
rect 893 3468 899 3712
rect 861 3368 867 3432
rect 861 3328 867 3352
rect 877 3348 883 3392
rect 909 3348 915 3832
rect 989 3828 995 3872
rect 1021 3868 1027 3872
rect 973 3788 979 3812
rect 797 3168 803 3312
rect 909 3308 915 3312
rect 824 3297 835 3303
rect 813 3188 819 3272
rect 701 2957 723 2963
rect 477 2688 483 2692
rect 557 2688 563 2732
rect 509 2588 515 2612
rect 493 2528 499 2532
rect 413 2328 419 2332
rect 397 2288 403 2292
rect 269 1888 275 1892
rect 381 1848 387 1892
rect 221 1737 243 1743
rect 237 1703 243 1737
rect 237 1697 259 1703
rect 173 1668 179 1672
rect 141 1368 147 1452
rect 109 1328 115 1332
rect 125 1188 131 1312
rect 157 1288 163 1392
rect 189 1328 195 1332
rect 157 1168 163 1272
rect 173 1268 179 1292
rect 205 1283 211 1672
rect 237 1448 243 1672
rect 253 1468 259 1697
rect 301 1668 307 1672
rect 317 1668 323 1692
rect 365 1688 371 1812
rect 413 1708 419 2032
rect 445 1988 451 2332
rect 461 1848 467 1892
rect 493 1888 499 2512
rect 557 2308 563 2592
rect 573 2288 579 2292
rect 509 2088 515 2232
rect 541 2128 547 2152
rect 557 2128 563 2132
rect 589 2123 595 2832
rect 637 2588 643 2812
rect 685 2788 691 2912
rect 701 2868 707 2932
rect 717 2728 723 2957
rect 733 2948 739 3032
rect 765 3028 771 3092
rect 797 3083 803 3132
rect 829 3128 835 3297
rect 893 3188 899 3292
rect 877 3148 883 3152
rect 829 3088 835 3112
rect 973 3088 979 3472
rect 989 3408 995 3812
rect 1037 3588 1043 3632
rect 1005 3488 1011 3512
rect 1021 3506 1027 3532
rect 1021 3328 1027 3352
rect 1053 3348 1059 3872
rect 1069 3708 1075 3712
rect 1085 3528 1091 4072
rect 1149 3988 1155 4312
rect 1165 4228 1171 4292
rect 1181 4248 1187 4332
rect 1309 4328 1315 4392
rect 1357 4388 1363 4472
rect 1357 4348 1363 4372
rect 1277 4308 1283 4312
rect 1213 4288 1219 4292
rect 1213 4148 1219 4272
rect 1341 4243 1347 4272
rect 1341 4237 1363 4243
rect 1165 4128 1171 4132
rect 1101 3868 1107 3972
rect 1181 3908 1187 3952
rect 1165 3888 1171 3892
rect 1101 3788 1107 3852
rect 1197 3728 1203 3872
rect 1213 3688 1219 4072
rect 1245 3948 1251 4132
rect 1293 4108 1299 4232
rect 1341 4128 1347 4192
rect 1357 4188 1363 4237
rect 1261 3908 1267 4032
rect 1357 3988 1363 4172
rect 1373 4168 1379 4232
rect 1389 4188 1395 4272
rect 1405 4028 1411 4132
rect 1421 3968 1427 4112
rect 1453 4088 1459 4372
rect 1469 4128 1475 4492
rect 1597 4488 1603 4592
rect 1613 4488 1619 4512
rect 1629 4508 1635 4592
rect 1645 4488 1651 4912
rect 1661 4908 1667 5352
rect 1725 5348 1731 5432
rect 1773 5268 1779 5432
rect 1789 5348 1795 5472
rect 1757 5106 1763 5112
rect 1789 5088 1795 5332
rect 1805 5228 1811 5492
rect 1837 5488 1843 5663
rect 1885 5308 1891 5432
rect 1917 5328 1923 5512
rect 1933 5368 1939 5432
rect 1869 5128 1875 5132
rect 1917 5128 1923 5312
rect 1933 5148 1939 5312
rect 1997 5288 2003 5292
rect 1997 5108 2003 5272
rect 2013 5248 2019 5452
rect 2093 5388 2099 5472
rect 2125 5428 2131 5512
rect 2205 5488 2211 5663
rect 2269 5628 2275 5663
rect 2237 5508 2243 5512
rect 2173 5388 2179 5472
rect 2205 5468 2211 5472
rect 1709 4948 1715 5012
rect 1741 4968 1747 5072
rect 1821 5028 1827 5072
rect 1661 4728 1667 4812
rect 1709 4708 1715 4932
rect 1805 4888 1811 4912
rect 1725 4728 1731 4772
rect 1709 4548 1715 4652
rect 1725 4608 1731 4712
rect 1741 4708 1747 4852
rect 1757 4748 1763 4832
rect 1821 4708 1827 4772
rect 1837 4708 1843 5092
rect 2013 5088 2019 5232
rect 2029 5188 2035 5332
rect 2189 5328 2195 5432
rect 2205 5388 2211 5412
rect 2061 5268 2067 5312
rect 2029 5048 2035 5072
rect 1981 4928 1987 4932
rect 2045 4928 2051 5252
rect 2061 5108 2067 5112
rect 2093 5108 2099 5252
rect 2173 5108 2179 5112
rect 1917 4728 1923 4752
rect 1949 4728 1955 4832
rect 1885 4708 1891 4712
rect 1949 4708 1955 4712
rect 1981 4708 1987 4912
rect 2061 4728 2067 5032
rect 2125 4888 2131 5032
rect 2141 4988 2147 5052
rect 2157 4908 2163 5032
rect 2173 4948 2179 5092
rect 2189 5048 2195 5312
rect 2237 5308 2243 5492
rect 2301 5388 2307 5392
rect 2253 5328 2259 5332
rect 2285 5308 2291 5312
rect 2317 5303 2323 5663
rect 2333 5408 2339 5492
rect 2397 5348 2403 5392
rect 2413 5368 2419 5452
rect 2397 5328 2403 5332
rect 2317 5297 2339 5303
rect 2237 5088 2243 5132
rect 2269 5048 2275 5072
rect 2285 5068 2291 5072
rect 2189 4948 2195 5032
rect 2125 4783 2131 4872
rect 2221 4828 2227 4832
rect 2109 4777 2131 4783
rect 1757 4568 1763 4632
rect 1821 4563 1827 4692
rect 1805 4557 1827 4563
rect 1805 4528 1811 4557
rect 1821 4528 1827 4532
rect 1597 4368 1603 4472
rect 1485 4288 1491 4292
rect 1597 4168 1603 4352
rect 1645 4288 1651 4292
rect 1613 4188 1619 4192
rect 1517 4128 1523 4132
rect 1469 4108 1475 4112
rect 1453 4008 1459 4072
rect 1389 3908 1395 3912
rect 1341 3888 1347 3892
rect 1405 3888 1411 3932
rect 1469 3923 1475 4032
rect 1464 3917 1475 3923
rect 1485 3908 1491 3912
rect 1437 3868 1443 3872
rect 1293 3788 1299 3792
rect 1117 3528 1123 3532
rect 1101 3488 1107 3492
rect 1165 3488 1171 3512
rect 1197 3488 1203 3552
rect 1213 3508 1219 3672
rect 1085 3368 1091 3472
rect 1069 3348 1075 3352
rect 1085 3308 1091 3332
rect 1165 3328 1171 3372
rect 1181 3317 1192 3323
rect 989 3288 995 3292
rect 797 3077 819 3083
rect 749 2868 755 2912
rect 685 2708 691 2712
rect 685 2568 691 2652
rect 749 2628 755 2852
rect 701 2588 707 2612
rect 605 2528 611 2532
rect 637 2208 643 2432
rect 701 2328 707 2552
rect 765 2543 771 3012
rect 781 2968 787 3072
rect 797 2908 803 2912
rect 797 2828 803 2892
rect 749 2537 771 2543
rect 749 2528 755 2537
rect 749 2408 755 2512
rect 765 2488 771 2512
rect 717 2328 723 2352
rect 701 2308 707 2312
rect 669 2248 675 2272
rect 669 2128 675 2232
rect 717 2128 723 2292
rect 749 2188 755 2332
rect 765 2163 771 2252
rect 781 2168 787 2172
rect 765 2157 776 2163
rect 584 2117 595 2123
rect 509 1908 515 2072
rect 541 1868 547 2112
rect 557 1948 563 2112
rect 429 1728 435 1732
rect 461 1708 467 1772
rect 477 1728 483 1732
rect 253 1308 259 1452
rect 269 1428 275 1432
rect 301 1308 307 1312
rect 333 1308 339 1472
rect 365 1388 371 1672
rect 381 1528 387 1692
rect 413 1668 419 1672
rect 429 1668 435 1692
rect 541 1688 547 1792
rect 557 1728 563 1912
rect 589 1868 595 1892
rect 605 1868 611 1872
rect 637 1863 643 2032
rect 669 1928 675 2112
rect 765 2108 771 2157
rect 669 1888 675 1892
rect 621 1857 643 1863
rect 397 1588 403 1652
rect 413 1548 419 1632
rect 461 1588 467 1672
rect 413 1508 419 1532
rect 477 1528 483 1532
rect 461 1508 467 1512
rect 205 1277 216 1283
rect 173 1188 179 1192
rect 93 1148 99 1152
rect 173 1148 179 1152
rect 205 1148 211 1277
rect 381 1283 387 1492
rect 397 1488 403 1492
rect 397 1308 403 1452
rect 413 1328 419 1332
rect 493 1303 499 1672
rect 557 1548 563 1712
rect 573 1708 579 1752
rect 557 1488 563 1532
rect 573 1508 579 1592
rect 589 1568 595 1652
rect 605 1588 611 1712
rect 621 1708 627 1857
rect 733 1788 739 1832
rect 749 1828 755 2032
rect 781 1808 787 2112
rect 797 1928 803 2492
rect 813 2348 819 3077
rect 893 2808 899 2932
rect 845 2568 851 2692
rect 909 2688 915 3072
rect 925 2928 931 2992
rect 973 2708 979 2872
rect 1021 2728 1027 2932
rect 861 2528 867 2572
rect 877 2508 883 2532
rect 925 2528 931 2672
rect 973 2608 979 2692
rect 1021 2688 1027 2712
rect 1053 2708 1059 3252
rect 1101 3248 1107 3312
rect 1021 2648 1027 2672
rect 1053 2628 1059 2692
rect 845 2488 851 2492
rect 909 2488 915 2492
rect 845 2388 851 2472
rect 829 2288 835 2372
rect 861 2368 867 2432
rect 973 2428 979 2492
rect 1005 2468 1011 2512
rect 1053 2508 1059 2532
rect 1069 2528 1075 2972
rect 1117 2688 1123 3132
rect 1133 2708 1139 3292
rect 1149 2988 1155 3052
rect 1165 2968 1171 3052
rect 1181 3048 1187 3317
rect 1213 3308 1219 3492
rect 1261 3468 1267 3732
rect 1341 3688 1347 3712
rect 1373 3708 1379 3732
rect 1341 3448 1347 3512
rect 1261 3428 1267 3432
rect 1229 3283 1235 3392
rect 1261 3368 1267 3412
rect 1341 3368 1347 3432
rect 1357 3388 1363 3612
rect 1389 3548 1395 3712
rect 1405 3388 1411 3792
rect 1421 3728 1427 3832
rect 1437 3728 1443 3772
rect 1469 3768 1475 3872
rect 1501 3768 1507 4092
rect 1533 4068 1539 4072
rect 1517 3928 1523 4032
rect 1565 3988 1571 4012
rect 1581 3908 1587 4112
rect 1597 4048 1603 4152
rect 1629 3948 1635 4232
rect 1661 4108 1667 4152
rect 1677 4148 1683 4472
rect 1709 4448 1715 4512
rect 1773 4468 1779 4492
rect 1805 4288 1811 4292
rect 1677 4128 1683 4132
rect 1645 3988 1651 4052
rect 1517 3888 1523 3892
rect 1437 3588 1443 3712
rect 1501 3648 1507 3752
rect 1533 3748 1539 3872
rect 1629 3748 1635 3932
rect 1661 3928 1667 4072
rect 1533 3728 1539 3732
rect 1597 3728 1603 3732
rect 1565 3708 1571 3712
rect 1485 3508 1491 3632
rect 1565 3588 1571 3632
rect 1581 3608 1587 3712
rect 1629 3708 1635 3712
rect 1645 3668 1651 3892
rect 1661 3723 1667 3912
rect 1677 3748 1683 4092
rect 1693 4088 1699 4092
rect 1709 3728 1715 4032
rect 1805 4028 1811 4272
rect 1789 3908 1795 3932
rect 1837 3888 1843 4672
rect 1901 4628 1907 4672
rect 1901 4548 1907 4552
rect 1917 4548 1923 4632
rect 1933 4548 1939 4692
rect 1933 4408 1939 4532
rect 1901 4148 1907 4232
rect 1933 4148 1939 4292
rect 1949 4268 1955 4312
rect 1949 4128 1955 4132
rect 1853 3808 1859 4112
rect 1869 3768 1875 4052
rect 1901 3788 1907 3892
rect 1965 3888 1971 4132
rect 1997 4068 2003 4672
rect 2013 4568 2019 4672
rect 2029 4488 2035 4692
rect 2109 4688 2115 4777
rect 2253 4728 2259 5032
rect 2269 4948 2275 5032
rect 2301 4928 2307 5092
rect 2285 4708 2291 4712
rect 2061 4508 2067 4512
rect 2109 4408 2115 4672
rect 2157 4588 2163 4672
rect 2205 4548 2211 4652
rect 2237 4548 2243 4572
rect 2157 4528 2163 4532
rect 2285 4528 2291 4692
rect 2333 4688 2339 5297
rect 2365 5108 2371 5112
rect 2365 4908 2371 5092
rect 2397 5088 2403 5092
rect 2445 5088 2451 5472
rect 2493 5408 2499 5492
rect 2589 5348 2595 5452
rect 2685 5348 2691 5663
rect 2813 5508 2819 5663
rect 2877 5588 2883 5663
rect 2925 5588 2931 5663
rect 2973 5657 3011 5663
rect 3005 5588 3011 5657
rect 3021 5628 3027 5663
rect 3053 5588 3059 5612
rect 3101 5588 3107 5663
rect 3181 5628 3187 5663
rect 3229 5588 3235 5663
rect 3325 5588 3331 5663
rect 3789 5657 3811 5663
rect 2829 5497 2840 5503
rect 2477 5068 2483 5312
rect 2573 5188 2579 5312
rect 2493 5088 2499 5092
rect 2397 4688 2403 4772
rect 2413 4688 2419 4972
rect 2541 4968 2547 5072
rect 2445 4948 2451 4952
rect 2301 4563 2307 4632
rect 2301 4557 2323 4563
rect 2317 4508 2323 4557
rect 2029 4328 2035 4332
rect 2013 4288 2019 4292
rect 2093 4288 2099 4292
rect 2109 4288 2115 4372
rect 2125 4328 2131 4352
rect 2045 4128 2051 4132
rect 2061 4128 2067 4132
rect 2013 4088 2019 4092
rect 1997 3928 2003 3932
rect 2013 3928 2019 4032
rect 2061 3917 2072 3923
rect 1981 3888 1987 3892
rect 2029 3888 2035 3912
rect 2045 3888 2051 3892
rect 1885 3768 1891 3772
rect 1661 3717 1683 3723
rect 1501 3468 1507 3492
rect 1533 3428 1539 3472
rect 1304 3337 1347 3343
rect 1341 3323 1347 3337
rect 1341 3317 1384 3323
rect 1245 3308 1251 3312
rect 1261 3308 1267 3312
rect 1213 3277 1235 3283
rect 1197 2968 1203 3112
rect 1213 3108 1219 3277
rect 1261 3188 1267 3232
rect 1309 3188 1315 3292
rect 1325 3268 1331 3312
rect 1352 3277 1363 3283
rect 1357 3188 1363 3277
rect 1373 3248 1379 3292
rect 1405 3268 1411 3272
rect 1437 3188 1443 3252
rect 1357 3148 1363 3152
rect 1245 3088 1251 3132
rect 1325 3128 1331 3132
rect 1421 3128 1427 3152
rect 1165 2908 1171 2912
rect 1213 2908 1219 3072
rect 1229 2928 1235 2992
rect 1261 2988 1267 3092
rect 1309 3048 1315 3092
rect 1389 3048 1395 3092
rect 1405 2968 1411 2972
rect 1293 2868 1299 2912
rect 1021 2448 1027 2472
rect 1037 2388 1043 2452
rect 989 2348 995 2352
rect 1053 2348 1059 2452
rect 1117 2408 1123 2672
rect 813 2128 819 2192
rect 829 2148 835 2272
rect 845 2148 851 2292
rect 989 2248 995 2292
rect 1037 2288 1043 2292
rect 877 2148 883 2192
rect 829 1908 835 2132
rect 941 2108 947 2172
rect 957 2128 963 2232
rect 957 2048 963 2112
rect 973 2088 979 2172
rect 797 1848 803 1892
rect 749 1728 755 1732
rect 781 1728 787 1792
rect 845 1768 851 1852
rect 845 1723 851 1752
rect 877 1748 883 2032
rect 989 2003 995 2032
rect 973 1997 995 2003
rect 877 1728 883 1732
rect 845 1717 867 1723
rect 685 1588 691 1712
rect 861 1708 867 1717
rect 893 1688 899 1912
rect 973 1743 979 1997
rect 957 1737 979 1743
rect 957 1708 963 1737
rect 1037 1728 1043 1732
rect 973 1688 979 1712
rect 1021 1668 1027 1692
rect 1037 1668 1043 1672
rect 829 1628 835 1632
rect 589 1528 595 1552
rect 1005 1548 1011 1632
rect 605 1508 611 1532
rect 541 1408 547 1432
rect 477 1297 499 1303
rect 376 1277 387 1283
rect 221 1268 227 1272
rect 237 1268 243 1272
rect 301 1168 307 1232
rect 365 1188 371 1232
rect 413 1148 419 1232
rect 429 1148 435 1272
rect 328 1137 344 1143
rect 93 1083 99 1132
rect 445 1128 451 1212
rect 93 1077 115 1083
rect 77 997 99 1003
rect 93 928 99 997
rect 93 688 99 692
rect 93 528 99 532
rect 109 428 115 1077
rect 173 1068 179 1092
rect 189 1088 195 1112
rect 237 988 243 1072
rect 269 968 275 1112
rect 365 1108 371 1112
rect 285 1088 291 1092
rect 381 1048 387 1112
rect 141 708 147 932
rect 157 930 163 932
rect 381 928 387 932
rect 397 928 403 1052
rect 413 968 419 1032
rect 429 988 435 1032
rect 221 708 227 892
rect 141 528 147 692
rect 237 528 243 912
rect 397 728 403 912
rect 461 883 467 1272
rect 477 1248 483 1297
rect 557 1288 563 1372
rect 605 1348 611 1492
rect 621 1448 627 1532
rect 1069 1508 1075 2292
rect 1085 2108 1091 2272
rect 1101 2168 1107 2292
rect 1117 2188 1123 2392
rect 1133 2308 1139 2692
rect 1245 2688 1251 2692
rect 1149 2268 1155 2432
rect 1165 2368 1171 2632
rect 1197 2548 1203 2632
rect 1133 2123 1139 2232
rect 1165 2168 1171 2252
rect 1181 2228 1187 2512
rect 1261 2508 1267 2512
rect 1293 2448 1299 2852
rect 1453 2808 1459 3132
rect 1469 2968 1475 3232
rect 1501 3128 1507 3132
rect 1501 2868 1507 3112
rect 1517 3108 1523 3312
rect 1533 3288 1539 3412
rect 1581 3388 1587 3452
rect 1629 3448 1635 3472
rect 1613 3348 1619 3432
rect 1645 3408 1651 3492
rect 1661 3388 1667 3692
rect 1677 3368 1683 3717
rect 1693 3588 1699 3692
rect 1709 3548 1715 3712
rect 1725 3548 1731 3732
rect 1741 3728 1747 3732
rect 1789 3728 1795 3732
rect 1741 3697 1752 3703
rect 1741 3588 1747 3697
rect 1693 3368 1699 3492
rect 1613 3317 1624 3323
rect 1517 3048 1523 3092
rect 1533 3068 1539 3112
rect 1549 3103 1555 3232
rect 1597 3188 1603 3312
rect 1613 3268 1619 3317
rect 1629 3188 1635 3292
rect 1693 3188 1699 3272
rect 1709 3248 1715 3512
rect 1757 3508 1763 3652
rect 1821 3588 1827 3692
rect 1805 3528 1811 3532
rect 1725 3497 1736 3503
rect 1549 3097 1560 3103
rect 1581 3083 1587 3132
rect 1565 3077 1587 3083
rect 1565 2988 1571 3077
rect 1613 3068 1619 3112
rect 1645 3088 1651 3132
rect 1581 2928 1587 3032
rect 1661 2988 1667 3112
rect 1677 3068 1683 3112
rect 1677 2908 1683 3052
rect 1437 2708 1443 2772
rect 1325 2668 1331 2692
rect 1405 2668 1411 2692
rect 1501 2688 1507 2772
rect 1325 2548 1331 2592
rect 1197 2308 1203 2432
rect 1245 2348 1251 2352
rect 1261 2323 1267 2412
rect 1309 2348 1315 2392
rect 1325 2328 1331 2532
rect 1341 2448 1347 2512
rect 1261 2317 1272 2323
rect 1245 2308 1251 2312
rect 1197 2128 1203 2292
rect 1261 2288 1267 2317
rect 1261 2168 1267 2272
rect 1293 2248 1299 2292
rect 1373 2288 1379 2292
rect 1341 2268 1347 2272
rect 1293 2128 1299 2132
rect 1128 2117 1139 2123
rect 1117 1848 1123 1892
rect 1133 1708 1139 1952
rect 1117 1523 1123 1632
rect 1133 1568 1139 1692
rect 1149 1628 1155 1892
rect 1245 1868 1251 1892
rect 1197 1788 1203 1852
rect 1229 1828 1235 1832
rect 1165 1668 1171 1672
rect 1117 1517 1128 1523
rect 1165 1508 1171 1552
rect 589 1308 595 1332
rect 605 1328 611 1332
rect 669 1328 675 1332
rect 477 1148 483 1232
rect 509 1228 515 1232
rect 541 1163 547 1232
rect 525 1157 547 1163
rect 493 1148 499 1152
rect 525 1108 531 1157
rect 557 1108 563 1192
rect 573 1128 579 1152
rect 589 1128 595 1292
rect 685 1288 691 1432
rect 765 1288 771 1432
rect 829 1308 835 1432
rect 1021 1388 1027 1492
rect 1181 1468 1187 1712
rect 1197 1708 1203 1772
rect 1229 1748 1235 1752
rect 1245 1708 1251 1852
rect 1261 1748 1267 2072
rect 1325 1908 1331 2252
rect 1373 2208 1379 2272
rect 1389 2148 1395 2592
rect 1405 2488 1411 2612
rect 1485 2548 1491 2552
rect 1469 2508 1475 2512
rect 1448 2497 1459 2503
rect 1405 2468 1411 2472
rect 1421 2148 1427 2232
rect 1453 2188 1459 2497
rect 1469 2308 1475 2452
rect 1453 2168 1459 2172
rect 1469 2148 1475 2292
rect 1501 2288 1507 2632
rect 1517 2468 1523 2692
rect 1533 2488 1539 2792
rect 1581 2728 1587 2872
rect 1549 2528 1555 2692
rect 1565 2508 1571 2672
rect 1581 2623 1587 2712
rect 1661 2708 1667 2832
rect 1709 2808 1715 3132
rect 1725 3128 1731 3497
rect 1805 3328 1811 3332
rect 1725 2988 1731 3072
rect 1757 2928 1763 3192
rect 1837 3148 1843 3212
rect 1773 2948 1779 2952
rect 1757 2848 1763 2912
rect 1725 2768 1731 2832
rect 1837 2708 1843 3132
rect 1581 2617 1603 2623
rect 1597 2488 1603 2617
rect 1645 2608 1651 2672
rect 1677 2648 1683 2690
rect 1645 2528 1651 2552
rect 1613 2488 1619 2512
rect 1597 2388 1603 2472
rect 1613 2388 1619 2432
rect 1661 2428 1667 2592
rect 1725 2588 1731 2632
rect 1549 2248 1555 2292
rect 1501 2188 1507 2232
rect 1357 2130 1363 2132
rect 1517 2128 1523 2132
rect 1533 2128 1539 2132
rect 1517 1908 1523 1972
rect 1533 1928 1539 1932
rect 1277 1888 1283 1892
rect 1357 1828 1363 1852
rect 1533 1828 1539 1832
rect 1341 1748 1347 1752
rect 1101 1428 1107 1432
rect 861 1288 867 1352
rect 877 1328 883 1332
rect 909 1328 915 1352
rect 1101 1348 1107 1412
rect 1117 1348 1123 1352
rect 621 1268 627 1272
rect 605 1148 611 1232
rect 637 1128 643 1252
rect 669 1128 675 1232
rect 685 1148 691 1272
rect 733 1208 739 1232
rect 749 1228 755 1272
rect 781 1168 787 1232
rect 877 1148 883 1212
rect 893 1188 899 1272
rect 973 1148 979 1332
rect 1037 1328 1043 1332
rect 1021 1188 1027 1292
rect 1053 1188 1059 1312
rect 1069 1288 1075 1292
rect 1181 1188 1187 1332
rect 1197 1328 1203 1432
rect 1261 1408 1267 1732
rect 1277 1708 1283 1712
rect 1277 1388 1283 1572
rect 1293 1548 1299 1612
rect 1357 1528 1363 1812
rect 1389 1768 1395 1812
rect 1405 1708 1411 1772
rect 1437 1688 1443 1772
rect 1517 1748 1523 1752
rect 1549 1743 1555 2092
rect 1581 2088 1587 2352
rect 1597 2188 1603 2252
rect 1613 2148 1619 2212
rect 1613 2128 1619 2132
rect 1565 1948 1571 2032
rect 1565 1908 1571 1912
rect 1533 1737 1555 1743
rect 1469 1708 1475 1732
rect 1501 1728 1507 1732
rect 1469 1588 1475 1692
rect 1469 1528 1475 1572
rect 1261 1368 1267 1372
rect 1053 1168 1059 1172
rect 621 1108 627 1112
rect 797 1108 803 1112
rect 845 1108 851 1112
rect 909 1108 915 1112
rect 493 1088 499 1092
rect 541 1088 547 1092
rect 493 928 499 1072
rect 669 1068 675 1092
rect 541 928 547 932
rect 557 928 563 932
rect 717 928 723 1072
rect 456 877 467 883
rect 333 708 339 712
rect 317 688 323 692
rect 317 548 323 672
rect 365 668 371 692
rect 365 568 371 572
rect 397 528 403 692
rect 461 548 467 877
rect 509 708 515 832
rect 445 528 451 532
rect 29 348 35 352
rect 45 348 51 352
rect 109 348 115 412
rect 45 308 51 312
rect 61 168 67 312
rect 109 308 115 312
rect 141 208 147 512
rect 173 388 179 392
rect 237 368 243 432
rect 189 328 195 352
rect 205 308 211 312
rect 173 288 179 292
rect 141 148 147 192
rect 269 168 275 312
rect 285 308 291 512
rect 301 368 307 512
rect 477 508 483 572
rect 557 568 563 652
rect 317 388 323 452
rect 333 288 339 352
rect 349 348 355 432
rect 365 388 371 492
rect 509 488 515 532
rect 589 528 595 832
rect 605 708 611 712
rect 701 708 707 812
rect 653 628 659 672
rect 557 488 563 492
rect 429 468 435 472
rect 509 468 515 472
rect 573 463 579 512
rect 557 457 579 463
rect 461 388 467 432
rect 429 348 435 352
rect 365 308 371 312
rect 221 128 227 132
rect 333 128 339 272
rect 381 168 387 312
rect 493 308 499 372
rect 509 328 515 352
rect 541 348 547 412
rect 557 388 563 457
rect 589 323 595 512
rect 605 508 611 552
rect 621 428 627 512
rect 669 508 675 552
rect 701 508 707 692
rect 701 468 707 472
rect 621 348 627 372
rect 685 368 691 432
rect 589 317 611 323
rect 557 308 563 312
rect 605 308 611 317
rect 717 308 723 672
rect 733 528 739 632
rect 749 628 755 912
rect 765 708 771 1072
rect 813 1068 819 1092
rect 813 948 819 1052
rect 877 988 883 1092
rect 877 928 883 972
rect 909 928 915 992
rect 957 883 963 1132
rect 1085 1108 1091 1132
rect 973 1088 979 1092
rect 1197 1088 1203 1092
rect 1229 1088 1235 1352
rect 1245 1108 1251 1132
rect 1277 1128 1283 1272
rect 1293 1088 1299 1192
rect 1309 1143 1315 1332
rect 1325 1308 1331 1512
rect 1341 1328 1347 1452
rect 1485 1423 1491 1652
rect 1517 1508 1523 1732
rect 1533 1708 1539 1737
rect 1565 1728 1571 1892
rect 1581 1888 1587 1992
rect 1549 1688 1555 1712
rect 1469 1417 1491 1423
rect 1469 1388 1475 1417
rect 1469 1328 1475 1352
rect 1501 1348 1507 1372
rect 1517 1348 1523 1492
rect 1533 1448 1539 1672
rect 1357 1248 1363 1272
rect 1453 1268 1459 1312
rect 1309 1137 1331 1143
rect 1325 1128 1331 1137
rect 1341 1128 1347 1232
rect 1469 1188 1475 1252
rect 1517 1208 1523 1332
rect 1549 1328 1555 1672
rect 1581 1628 1587 1872
rect 1629 1788 1635 1832
rect 1581 1368 1587 1612
rect 1533 1228 1539 1312
rect 1613 1308 1619 1772
rect 1645 1748 1651 2312
rect 1693 2308 1699 2472
rect 1709 2368 1715 2572
rect 1741 2528 1747 2532
rect 1709 2348 1715 2352
rect 1693 2228 1699 2292
rect 1677 2128 1683 2132
rect 1693 2048 1699 2092
rect 1661 1908 1667 2032
rect 1693 1928 1699 2032
rect 1645 1648 1651 1732
rect 1661 1708 1667 1732
rect 1645 1506 1651 1532
rect 1677 1488 1683 1852
rect 1709 1828 1715 1852
rect 1725 1788 1731 2052
rect 1741 1888 1747 2512
rect 1757 2468 1763 2512
rect 1757 2368 1763 2452
rect 1773 2308 1779 2432
rect 1773 2028 1779 2292
rect 1789 2288 1795 2592
rect 1837 2468 1843 2512
rect 1805 2348 1811 2432
rect 1789 2008 1795 2272
rect 1837 2268 1843 2292
rect 1853 2288 1859 3752
rect 1869 3748 1875 3752
rect 1901 3728 1907 3772
rect 1917 3703 1923 3712
rect 1997 3708 2003 3852
rect 2045 3708 2051 3872
rect 2061 3788 2067 3917
rect 2093 3808 2099 3972
rect 2109 3948 2115 4272
rect 2125 4148 2131 4232
rect 2141 4188 2147 4192
rect 2125 4008 2131 4112
rect 2157 3943 2163 4392
rect 2205 4328 2211 4472
rect 2205 4308 2211 4312
rect 2189 4288 2195 4292
rect 2173 4068 2179 4272
rect 2189 4048 2195 4232
rect 2205 4148 2211 4292
rect 2221 4148 2227 4432
rect 2237 4288 2243 4492
rect 2301 4188 2307 4312
rect 2333 4188 2339 4672
rect 2445 4668 2451 4932
rect 2445 4548 2451 4652
rect 2477 4648 2483 4692
rect 2413 4528 2419 4532
rect 2445 4308 2451 4532
rect 2541 4508 2547 4532
rect 2589 4488 2595 5332
rect 2637 5128 2643 5132
rect 2685 5128 2691 5332
rect 2733 5268 2739 5472
rect 2797 5263 2803 5492
rect 2829 5488 2835 5497
rect 3192 5497 3203 5503
rect 2893 5388 2899 5492
rect 2813 5288 2819 5332
rect 2781 5257 2803 5263
rect 2744 5237 2755 5243
rect 2621 5088 2627 5092
rect 2637 5088 2643 5112
rect 2669 5108 2675 5112
rect 2749 5108 2755 5237
rect 2653 4908 2659 5032
rect 2669 4908 2675 4932
rect 2685 4928 2691 5092
rect 2749 5048 2755 5092
rect 2717 4948 2723 4952
rect 2765 4848 2771 5032
rect 2781 4788 2787 5257
rect 2797 5128 2803 5232
rect 2797 5088 2803 5092
rect 2813 5088 2819 5272
rect 2845 5128 2851 5312
rect 2845 5088 2851 5092
rect 2845 5068 2851 5072
rect 2637 4708 2643 4712
rect 2621 4668 2627 4692
rect 2669 4508 2675 4512
rect 2365 4148 2371 4172
rect 2205 4108 2211 4132
rect 2157 3937 2179 3943
rect 2141 3888 2147 3912
rect 2173 3908 2179 3937
rect 2173 3888 2179 3892
rect 2093 3748 2099 3792
rect 2237 3788 2243 3952
rect 2109 3748 2115 3752
rect 2125 3728 2131 3772
rect 2173 3748 2179 3752
rect 1901 3697 1923 3703
rect 1901 3328 1907 3697
rect 2061 3568 2067 3692
rect 2125 3588 2131 3692
rect 1917 3468 1923 3492
rect 2029 3488 2035 3490
rect 2109 3468 2115 3532
rect 2253 3508 2259 4012
rect 2445 3908 2451 4292
rect 2541 4168 2547 4472
rect 2685 4288 2691 4612
rect 2717 4528 2723 4712
rect 2765 4588 2771 4692
rect 2845 4668 2851 4872
rect 2861 4728 2867 5092
rect 2877 5088 2883 5092
rect 2909 4808 2915 5312
rect 2941 5183 2947 5492
rect 2989 5388 2995 5492
rect 3117 5488 3123 5492
rect 2941 5177 2952 5183
rect 3021 5128 3027 5252
rect 3085 5128 3091 5232
rect 2893 4748 2899 4792
rect 2925 4783 2931 5092
rect 3117 5088 3123 5272
rect 3149 5148 3155 5272
rect 3144 5097 3155 5103
rect 3085 4948 3091 5072
rect 3101 4908 3107 5032
rect 3149 4988 3155 5097
rect 3165 4928 3171 5492
rect 3181 5188 3187 5472
rect 3197 5388 3203 5497
rect 3277 5497 3288 5503
rect 3245 5408 3251 5492
rect 3277 5488 3283 5497
rect 3485 5506 3491 5512
rect 3597 5508 3603 5512
rect 3757 5508 3763 5512
rect 3341 5348 3347 5432
rect 3421 5368 3427 5432
rect 3197 5208 3203 5232
rect 3213 5088 3219 5132
rect 2920 4777 2931 4783
rect 2941 4708 2947 4712
rect 2973 4708 2979 4712
rect 2781 4548 2787 4652
rect 2893 4608 2899 4692
rect 2925 4688 2931 4692
rect 3037 4688 3043 4712
rect 3069 4588 3075 4832
rect 2701 4508 2707 4512
rect 2813 4508 2819 4514
rect 2829 4388 2835 4432
rect 2861 4388 2867 4392
rect 2925 4388 2931 4392
rect 2909 4328 2915 4352
rect 3005 4328 3011 4472
rect 2589 4148 2595 4232
rect 2605 4168 2611 4252
rect 2477 4108 2483 4112
rect 2445 3888 2451 3892
rect 2381 3748 2387 3792
rect 2461 3788 2467 3892
rect 2365 3648 2371 3652
rect 2365 3508 2371 3632
rect 2429 3508 2435 3712
rect 2477 3708 2483 4092
rect 2557 3908 2563 3932
rect 2573 3863 2579 4132
rect 2653 4108 2659 4232
rect 2685 4148 2691 4272
rect 2589 3908 2595 3912
rect 2557 3857 2579 3863
rect 2541 3768 2547 3832
rect 2557 3828 2563 3857
rect 2621 3843 2627 3912
rect 2685 3906 2691 3912
rect 2653 3888 2659 3892
rect 2701 3888 2707 4272
rect 2765 4188 2771 4272
rect 2877 4208 2883 4312
rect 2893 4168 2899 4292
rect 2925 4168 2931 4172
rect 2829 4128 2835 4132
rect 2717 4108 2723 4112
rect 2749 3868 2755 4112
rect 2813 4108 2819 4112
rect 2877 4088 2883 4092
rect 2781 3948 2787 4032
rect 2941 3968 2947 4312
rect 3021 4308 3027 4552
rect 3085 4548 3091 4612
rect 3053 4283 3059 4492
rect 3117 4383 3123 4912
rect 3165 4708 3171 4872
rect 3197 4788 3203 4832
rect 3133 4528 3139 4632
rect 3213 4628 3219 4932
rect 3245 4748 3251 5312
rect 3277 5288 3283 5332
rect 3309 5308 3315 5332
rect 3437 5328 3443 5332
rect 3293 5088 3299 5092
rect 3277 4928 3283 4932
rect 3309 4928 3315 5072
rect 3341 5068 3347 5312
rect 3357 5288 3363 5312
rect 3453 4988 3459 5472
rect 3485 5268 3491 5332
rect 3645 5328 3651 5492
rect 3661 5328 3667 5472
rect 3677 5388 3683 5472
rect 3501 5128 3507 5132
rect 3469 5108 3475 5112
rect 3357 4928 3363 4952
rect 3373 4728 3379 4752
rect 3405 4748 3411 4932
rect 3437 4928 3443 4932
rect 3453 4888 3459 4972
rect 3469 4928 3475 5092
rect 3469 4908 3475 4912
rect 3437 4708 3443 4712
rect 3469 4708 3475 4892
rect 3501 4828 3507 5032
rect 3517 5008 3523 5232
rect 3565 5148 3571 5232
rect 3613 5128 3619 5192
rect 3629 5108 3635 5292
rect 3645 5128 3651 5312
rect 3645 5108 3651 5112
rect 3661 5088 3667 5312
rect 3677 5088 3683 5192
rect 3693 5108 3699 5314
rect 3773 5288 3779 5332
rect 3805 5223 3811 5657
rect 3821 5308 3827 5432
rect 3789 5217 3811 5223
rect 3789 5188 3795 5217
rect 3837 5208 3843 5312
rect 3853 5183 3859 5663
rect 3901 5488 3907 5492
rect 3933 5388 3939 5663
rect 4141 5588 4147 5663
rect 4189 5588 4195 5663
rect 4237 5588 4243 5663
rect 4573 5508 4579 5512
rect 4701 5508 4707 5512
rect 4797 5508 4803 5512
rect 5053 5508 5059 5512
rect 5181 5508 5187 5512
rect 4093 5497 4104 5503
rect 4061 5388 4067 5492
rect 4093 5488 4099 5497
rect 4157 5468 4163 5492
rect 4301 5448 4307 5452
rect 3949 5348 3955 5352
rect 3869 5323 3875 5332
rect 3869 5317 3880 5323
rect 3848 5177 3859 5183
rect 3901 5108 3907 5272
rect 3741 5097 3752 5103
rect 3533 4948 3539 4952
rect 3549 4948 3555 4992
rect 3565 4948 3571 5072
rect 3565 4928 3571 4932
rect 3149 4548 3155 4612
rect 3240 4537 3251 4543
rect 3149 4503 3155 4512
rect 3165 4508 3171 4532
rect 3245 4528 3251 4537
rect 3144 4497 3155 4503
rect 3165 4388 3171 4392
rect 3112 4377 3123 4383
rect 3165 4323 3171 4332
rect 3181 4328 3187 4412
rect 3133 4317 3171 4323
rect 3037 4277 3059 4283
rect 3037 4148 3043 4277
rect 3000 4117 3011 4123
rect 2989 4108 2995 4112
rect 2621 3837 2643 3843
rect 2493 3708 2499 3712
rect 2125 3468 2131 3492
rect 1917 3388 1923 3452
rect 1997 3328 2003 3412
rect 2029 3388 2035 3452
rect 2141 3368 2147 3492
rect 2157 3468 2163 3492
rect 2253 3488 2259 3492
rect 2269 3448 2275 3492
rect 2461 3488 2467 3572
rect 2509 3523 2515 3732
rect 2504 3517 2515 3523
rect 1917 3088 1923 3232
rect 1981 3068 1987 3072
rect 1997 2963 2003 3312
rect 1981 2957 2003 2963
rect 1869 2908 1875 2952
rect 1981 2888 1987 2957
rect 1997 2928 2003 2932
rect 2013 2928 2019 3092
rect 2029 2988 2035 3272
rect 2061 3248 2067 3312
rect 2141 3188 2147 3292
rect 2093 3108 2099 3152
rect 2077 2968 2083 3052
rect 2093 2928 2099 3072
rect 2125 2988 2131 3092
rect 2157 2988 2163 3432
rect 2285 3348 2291 3472
rect 2461 3368 2467 3472
rect 2397 3348 2403 3352
rect 2381 3328 2387 3332
rect 2301 3228 2307 3312
rect 2349 3228 2355 3292
rect 2429 3108 2435 3312
rect 2461 3268 2467 3332
rect 2477 3308 2483 3432
rect 2509 3388 2515 3492
rect 2557 3488 2563 3812
rect 2637 3788 2643 3837
rect 2749 3808 2755 3852
rect 2669 3748 2675 3792
rect 2765 3788 2771 3792
rect 2685 3748 2691 3752
rect 2781 3748 2787 3752
rect 2605 3728 2611 3732
rect 2589 3648 2595 3672
rect 2525 3348 2531 3392
rect 2605 3388 2611 3452
rect 2493 3128 2499 3312
rect 2509 3188 2515 3292
rect 2525 3148 2531 3332
rect 2621 3328 2627 3632
rect 2589 3288 2595 3312
rect 2605 3183 2611 3272
rect 2637 3228 2643 3692
rect 2669 3428 2675 3432
rect 2685 3403 2691 3732
rect 2813 3728 2819 3792
rect 2733 3628 2739 3692
rect 2701 3468 2707 3492
rect 2669 3397 2691 3403
rect 2653 3188 2659 3332
rect 2600 3177 2611 3183
rect 2477 3083 2483 3112
rect 2461 3077 2483 3083
rect 2141 2928 2147 2932
rect 2157 2928 2163 2972
rect 2173 2968 2179 3032
rect 2205 2928 2211 2992
rect 2285 2988 2291 3052
rect 2349 3048 2355 3072
rect 1965 2708 1971 2812
rect 2013 2788 2019 2912
rect 2029 2708 2035 2832
rect 1869 2628 1875 2652
rect 1869 2508 1875 2552
rect 1933 2548 1939 2632
rect 2045 2548 2051 2632
rect 1901 2388 1907 2492
rect 1885 2288 1891 2292
rect 1853 2088 1859 2272
rect 1869 2268 1875 2272
rect 1981 2108 1987 2132
rect 1997 2128 2003 2532
rect 2013 2528 2019 2532
rect 2061 2508 2067 2632
rect 2077 2508 2083 2792
rect 2093 2728 2099 2752
rect 2125 2748 2131 2832
rect 2189 2748 2195 2872
rect 2205 2868 2211 2892
rect 2173 2628 2179 2692
rect 2221 2668 2227 2972
rect 2237 2948 2243 2952
rect 2333 2928 2339 3012
rect 2397 2988 2403 3052
rect 2413 2903 2419 3072
rect 2461 2988 2467 3077
rect 2429 2928 2435 2952
rect 2477 2928 2483 3052
rect 2493 2988 2499 3112
rect 2509 3068 2515 3092
rect 2541 2948 2547 3032
rect 2413 2897 2435 2903
rect 2285 2728 2291 2852
rect 2301 2748 2307 2892
rect 2333 2743 2339 2872
rect 2328 2737 2339 2743
rect 2301 2728 2307 2732
rect 2269 2668 2275 2672
rect 2157 2568 2163 2592
rect 2125 2528 2131 2552
rect 2173 2528 2179 2612
rect 2221 2508 2227 2652
rect 2237 2608 2243 2632
rect 2317 2528 2323 2532
rect 2061 2488 2067 2492
rect 2189 2488 2195 2492
rect 2013 2448 2019 2472
rect 2269 2448 2275 2512
rect 2333 2508 2339 2737
rect 2397 2688 2403 2732
rect 2349 2508 2355 2572
rect 2397 2568 2403 2652
rect 2429 2548 2435 2897
rect 2477 2588 2483 2892
rect 2541 2743 2547 2932
rect 2573 2848 2579 3132
rect 2589 3028 2595 3092
rect 2605 3048 2611 3112
rect 2605 2808 2611 3032
rect 2653 3008 2659 3092
rect 2669 3088 2675 3397
rect 2701 3328 2707 3332
rect 2717 3308 2723 3412
rect 2765 3388 2771 3692
rect 2797 3548 2803 3712
rect 2829 3708 2835 3852
rect 2861 3788 2867 3892
rect 2941 3828 2947 3872
rect 2941 3768 2947 3772
rect 2872 3697 2883 3703
rect 2813 3588 2819 3612
rect 2877 3588 2883 3697
rect 2909 3548 2915 3632
rect 2797 3488 2803 3532
rect 2781 3388 2787 3432
rect 2733 3348 2739 3352
rect 2813 3328 2819 3332
rect 2685 3148 2691 3272
rect 2797 3188 2803 3272
rect 2621 2928 2627 2932
rect 2525 2737 2547 2743
rect 2493 2706 2499 2712
rect 2525 2688 2531 2737
rect 2605 2708 2611 2712
rect 2637 2708 2643 2712
rect 2397 2448 2403 2512
rect 2125 2408 2131 2432
rect 2061 2308 2067 2392
rect 2413 2348 2419 2532
rect 2253 2308 2259 2332
rect 2285 2308 2291 2312
rect 2525 2308 2531 2672
rect 2557 2548 2563 2632
rect 2573 2568 2579 2672
rect 2557 2528 2563 2532
rect 2589 2508 2595 2652
rect 2637 2588 2643 2672
rect 2653 2568 2659 2692
rect 2637 2388 2643 2472
rect 2669 2468 2675 2512
rect 2685 2308 2691 3112
rect 2813 3103 2819 3292
rect 2829 3288 2835 3532
rect 2845 3488 2851 3492
rect 2893 3408 2899 3532
rect 2909 3528 2915 3532
rect 2909 3488 2915 3492
rect 2941 3308 2947 3312
rect 2973 3308 2979 3552
rect 2893 3148 2899 3232
rect 2808 3097 2819 3103
rect 2717 2928 2723 3032
rect 2733 2948 2739 2952
rect 2781 2888 2787 2912
rect 2781 2648 2787 2872
rect 2797 2748 2803 3092
rect 2829 3088 2835 3112
rect 2893 3108 2899 3132
rect 2893 3088 2899 3092
rect 2925 3088 2931 3092
rect 2813 2988 2819 3052
rect 2829 3048 2835 3072
rect 2845 2963 2851 3032
rect 2829 2957 2851 2963
rect 2829 2908 2835 2957
rect 2925 2928 2931 2952
rect 2888 2897 2899 2903
rect 2829 2706 2835 2712
rect 2701 2508 2707 2552
rect 2733 2548 2739 2572
rect 2781 2528 2787 2552
rect 2813 2548 2819 2672
rect 2893 2568 2899 2897
rect 2941 2728 2947 3092
rect 3005 3088 3011 4117
rect 3021 3948 3027 4032
rect 3021 3748 3027 3752
rect 3037 3748 3043 4132
rect 3085 3868 3091 4312
rect 3133 4308 3139 4317
rect 3197 4308 3203 4492
rect 3213 4468 3219 4492
rect 3149 4203 3155 4292
rect 3133 4197 3155 4203
rect 3101 4068 3107 4092
rect 3117 3888 3123 4192
rect 3133 4188 3139 4197
rect 3149 4168 3155 4172
rect 3165 4108 3171 4292
rect 3245 4148 3251 4512
rect 3261 4508 3267 4512
rect 3261 4108 3267 4312
rect 3197 4048 3203 4072
rect 3245 4068 3251 4072
rect 3277 3948 3283 4692
rect 3517 4688 3523 4732
rect 3549 4706 3555 4712
rect 3384 4677 3395 4683
rect 3229 3928 3235 3932
rect 3277 3908 3283 3932
rect 3293 3928 3299 4632
rect 3373 4568 3379 4652
rect 3389 4628 3395 4677
rect 3405 4648 3411 4672
rect 3581 4668 3587 4912
rect 3597 4908 3603 5032
rect 3645 4948 3651 5052
rect 3645 4928 3651 4932
rect 3693 4928 3699 4932
rect 3661 4908 3667 4912
rect 3629 4868 3635 4872
rect 3661 4848 3667 4892
rect 3709 4863 3715 5092
rect 3741 5088 3747 5097
rect 3789 5097 3800 5103
rect 3789 4988 3795 5097
rect 3853 4948 3859 5032
rect 3837 4928 3843 4932
rect 3885 4928 3891 4932
rect 3901 4928 3907 5092
rect 3949 5088 3955 5132
rect 4013 5128 4019 5292
rect 4077 5268 4083 5332
rect 4093 5288 4099 5312
rect 4189 5308 4195 5312
rect 4093 5128 4099 5272
rect 4093 5108 4099 5112
rect 4061 5088 4067 5092
rect 3949 5068 3955 5072
rect 3949 4928 3955 4932
rect 3709 4857 3731 4863
rect 3645 4728 3651 4832
rect 3725 4808 3731 4857
rect 3693 4788 3699 4792
rect 3757 4768 3763 4912
rect 3869 4908 3875 4912
rect 3981 4908 3987 4932
rect 3709 4748 3715 4752
rect 3805 4728 3811 4832
rect 3725 4688 3731 4692
rect 3613 4648 3619 4652
rect 3325 4528 3331 4552
rect 3373 4528 3379 4552
rect 3309 4408 3315 4492
rect 3325 4488 3331 4492
rect 3357 4488 3363 4492
rect 3341 4477 3352 4483
rect 3309 4288 3315 4352
rect 3325 4228 3331 4312
rect 3309 4068 3315 4132
rect 3341 4048 3347 4477
rect 3373 4308 3379 4492
rect 3389 4443 3395 4612
rect 3613 4588 3619 4612
rect 3677 4588 3683 4632
rect 3709 4588 3715 4672
rect 3821 4668 3827 4872
rect 3901 4868 3907 4872
rect 3837 4708 3843 4812
rect 3901 4748 3907 4852
rect 3949 4728 3955 4832
rect 3981 4708 3987 4812
rect 4029 4703 4035 4932
rect 4093 4928 4099 5092
rect 4109 4968 4115 5072
rect 4125 5048 4131 5052
rect 4125 4968 4131 5032
rect 4173 4948 4179 4972
rect 4045 4723 4051 4832
rect 4077 4828 4083 4912
rect 4077 4788 4083 4792
rect 4205 4788 4211 5372
rect 4301 5348 4307 5432
rect 4269 5308 4275 5332
rect 4269 5106 4275 5112
rect 4333 5088 4339 5472
rect 4365 5388 4371 5492
rect 4557 5468 4563 5472
rect 4429 5388 4435 5452
rect 4669 5348 4675 5472
rect 4413 5328 4419 5332
rect 4541 5328 4547 5332
rect 4349 5288 4355 5292
rect 4397 5288 4403 5312
rect 4349 5068 4355 5072
rect 4365 4783 4371 5192
rect 4381 5108 4387 5112
rect 4413 5108 4419 5112
rect 4461 4948 4467 5232
rect 4477 5108 4483 5172
rect 4493 4943 4499 5312
rect 4477 4937 4499 4943
rect 4413 4928 4419 4932
rect 4445 4908 4451 4912
rect 4365 4777 4376 4783
rect 4477 4783 4483 4937
rect 4493 4888 4499 4912
rect 4477 4777 4488 4783
rect 4072 4737 4083 4743
rect 4045 4717 4067 4723
rect 4061 4708 4067 4717
rect 4029 4697 4051 4703
rect 3853 4668 3859 4672
rect 3757 4628 3763 4652
rect 3437 4528 3443 4552
rect 3501 4528 3507 4552
rect 3389 4437 3411 4443
rect 3389 4288 3395 4392
rect 3405 4388 3411 4437
rect 3421 4348 3427 4492
rect 3453 4488 3459 4492
rect 3453 4468 3459 4472
rect 3437 4408 3443 4432
rect 3517 4368 3523 4432
rect 3549 4388 3555 4532
rect 3405 4208 3411 4232
rect 3341 3988 3347 4032
rect 3357 3988 3363 4072
rect 3373 4008 3379 4072
rect 3133 3888 3139 3892
rect 3112 3717 3123 3723
rect 3021 3708 3027 3712
rect 3117 3708 3123 3717
rect 3149 3723 3155 3872
rect 3197 3728 3203 3732
rect 3144 3717 3155 3723
rect 3213 3708 3219 3712
rect 3096 3697 3107 3703
rect 3069 3628 3075 3692
rect 3101 3588 3107 3697
rect 3133 3588 3139 3612
rect 3037 3348 3043 3412
rect 3053 3328 3059 3512
rect 3069 3408 3075 3532
rect 3117 3528 3123 3532
rect 3149 3528 3155 3532
rect 3085 3388 3091 3492
rect 3069 3308 3075 3352
rect 3117 3328 3123 3412
rect 3053 3268 3059 3292
rect 3053 3188 3059 3252
rect 3069 3128 3075 3212
rect 3117 3188 3123 3212
rect 3133 3188 3139 3332
rect 3149 3288 3155 3512
rect 3181 3508 3187 3672
rect 3261 3568 3267 3732
rect 3277 3588 3283 3592
rect 3261 3528 3267 3552
rect 3293 3528 3299 3532
rect 3165 3148 3171 3312
rect 3181 3128 3187 3492
rect 3293 3488 3299 3512
rect 3197 3388 3203 3452
rect 3261 3388 3267 3432
rect 3309 3348 3315 3872
rect 3325 3548 3331 3712
rect 3341 3588 3347 3592
rect 3357 3588 3363 3672
rect 3373 3648 3379 3892
rect 3405 3788 3411 4112
rect 3421 4108 3427 4332
rect 3437 4188 3443 4292
rect 3469 4088 3475 4332
rect 3501 4328 3507 4332
rect 3485 4288 3491 4292
rect 3533 4288 3539 4292
rect 3533 4228 3539 4272
rect 3549 4203 3555 4332
rect 3565 4328 3571 4492
rect 3597 4388 3603 4472
rect 3613 4388 3619 4532
rect 3773 4528 3779 4572
rect 3821 4528 3827 4532
rect 3837 4528 3843 4572
rect 3853 4528 3859 4652
rect 3901 4588 3907 4692
rect 3933 4588 3939 4692
rect 4029 4648 4035 4652
rect 3901 4557 3912 4563
rect 3869 4528 3875 4532
rect 3885 4528 3891 4532
rect 3661 4388 3667 4472
rect 3741 4388 3747 4512
rect 3853 4497 3864 4503
rect 3533 4197 3555 4203
rect 3485 4128 3491 4132
rect 3501 4128 3507 4132
rect 3533 4088 3539 4197
rect 3549 4128 3555 4152
rect 3565 4108 3571 4312
rect 3421 3988 3427 4072
rect 3389 3583 3395 3732
rect 3437 3728 3443 4012
rect 3469 3928 3475 4052
rect 3501 3988 3507 4072
rect 3501 3948 3507 3972
rect 3533 3948 3539 4072
rect 3549 3988 3555 3992
rect 3453 3888 3459 3892
rect 3453 3748 3459 3752
rect 3389 3577 3400 3583
rect 3325 3468 3331 3512
rect 3341 3408 3347 3532
rect 3389 3448 3395 3512
rect 3421 3468 3427 3492
rect 3437 3428 3443 3712
rect 3469 3648 3475 3912
rect 3485 3908 3491 3932
rect 3533 3868 3539 3912
rect 3549 3908 3555 3932
rect 3581 3928 3587 4312
rect 3613 4288 3619 4292
rect 3645 4068 3651 4312
rect 3661 4288 3667 4292
rect 3501 3588 3507 3632
rect 3501 3528 3507 3572
rect 3533 3568 3539 3852
rect 3597 3788 3603 4032
rect 3661 4008 3667 4272
rect 3677 3988 3683 4332
rect 3693 4317 3704 4323
rect 3693 4263 3699 4317
rect 3741 4263 3747 4292
rect 3757 4268 3763 4272
rect 3693 4257 3715 4263
rect 3709 4188 3715 4257
rect 3725 4257 3747 4263
rect 3693 4148 3699 4152
rect 3725 4108 3731 4257
rect 3741 4128 3747 4132
rect 3725 4088 3731 4092
rect 3677 3928 3683 3972
rect 3725 3948 3731 4032
rect 3757 4028 3763 4112
rect 3773 3948 3779 4472
rect 3805 4388 3811 4492
rect 3821 4348 3827 4472
rect 3853 4388 3859 4497
rect 3821 4308 3827 4312
rect 3805 4268 3811 4292
rect 3789 4188 3795 4212
rect 3821 3983 3827 4132
rect 3816 3977 3827 3983
rect 3837 3948 3843 4272
rect 3853 4268 3859 4292
rect 3869 4188 3875 4232
rect 3901 4188 3907 4557
rect 3981 4528 3987 4532
rect 4045 4528 4051 4697
rect 4077 4703 4083 4737
rect 4077 4697 4088 4703
rect 4109 4588 4115 4712
rect 4157 4708 4163 4772
rect 4189 4728 4195 4752
rect 4125 4608 4131 4692
rect 4141 4668 4147 4672
rect 4221 4668 4227 4712
rect 4237 4708 4243 4712
rect 4285 4708 4291 4772
rect 4509 4768 4515 5072
rect 4397 4688 4403 4692
rect 4109 4557 4120 4563
rect 4093 4508 4099 4512
rect 3933 4488 3939 4492
rect 3965 4468 3971 4472
rect 3933 4388 3939 4392
rect 3997 4348 4003 4472
rect 4013 4388 4019 4412
rect 3965 4303 3971 4312
rect 3949 4297 3971 4303
rect 3853 3988 3859 4132
rect 3885 3988 3891 4072
rect 3917 3988 3923 4072
rect 3757 3908 3763 3912
rect 3693 3888 3699 3892
rect 3629 3768 3635 3772
rect 3661 3748 3667 3752
rect 3789 3743 3795 3932
rect 3869 3928 3875 3952
rect 3933 3948 3939 4032
rect 3901 3928 3907 3932
rect 3949 3928 3955 4297
rect 3981 4268 3987 4292
rect 4109 4248 4115 4557
rect 4125 4528 4131 4532
rect 3981 4148 3987 4172
rect 4045 4168 4051 4232
rect 4141 4223 4147 4612
rect 4205 4588 4211 4632
rect 4269 4588 4275 4652
rect 4413 4568 4419 4752
rect 4445 4708 4451 4712
rect 4429 4668 4435 4692
rect 4477 4648 4483 4652
rect 4189 4428 4195 4472
rect 4253 4408 4259 4472
rect 4157 4288 4163 4292
rect 4301 4268 4307 4532
rect 4525 4508 4531 5092
rect 4541 5088 4547 5252
rect 4637 5148 4643 5314
rect 4621 5108 4627 5112
rect 4637 5083 4643 5092
rect 4669 5088 4675 5332
rect 4733 5328 4739 5472
rect 4717 5288 4723 5312
rect 4632 5077 4643 5083
rect 4557 4948 4563 5032
rect 4573 4908 4579 4912
rect 4573 4708 4579 4872
rect 4605 4788 4611 5072
rect 4637 4888 4643 5012
rect 4653 4968 4659 5072
rect 4701 4908 4707 5152
rect 4717 5088 4723 5272
rect 4749 5108 4755 5292
rect 4765 5128 4771 5232
rect 4797 5168 4803 5492
rect 5181 5488 5187 5492
rect 5245 5488 5251 5512
rect 4893 5368 4899 5472
rect 5037 5388 5043 5472
rect 4893 5348 4899 5352
rect 4973 5328 4979 5332
rect 5037 5308 5043 5372
rect 5133 5328 5139 5472
rect 4829 5208 4835 5232
rect 4845 5108 4851 5292
rect 4877 5128 4883 5192
rect 4893 5108 4899 5132
rect 4925 5108 4931 5112
rect 4717 4988 4723 5012
rect 4733 4948 4739 4972
rect 4765 4928 4771 5072
rect 4845 5068 4851 5072
rect 4781 4928 4787 4972
rect 4861 4948 4867 4952
rect 4877 4928 4883 5092
rect 4925 5048 4931 5072
rect 4941 5028 4947 5112
rect 4973 5108 4979 5152
rect 4989 5088 4995 5292
rect 5085 5148 5091 5312
rect 5165 5268 5171 5472
rect 5245 5368 5251 5472
rect 5325 5348 5331 5372
rect 5229 5328 5235 5332
rect 5373 5328 5379 5472
rect 5389 5468 5395 5472
rect 5501 5348 5507 5432
rect 5597 5388 5603 5492
rect 5613 5468 5619 5472
rect 5613 5388 5619 5452
rect 5421 5328 5427 5332
rect 5197 5288 5203 5312
rect 5309 5308 5315 5312
rect 4989 4968 4995 5072
rect 5005 4988 5011 5032
rect 5149 4968 5155 5032
rect 5165 5003 5171 5232
rect 5213 5048 5219 5072
rect 5165 4997 5187 5003
rect 4957 4928 4963 4932
rect 5101 4928 5107 4932
rect 4637 4708 4643 4872
rect 4573 4628 4579 4692
rect 4541 4528 4547 4532
rect 4573 4508 4579 4512
rect 4125 4217 4147 4223
rect 4109 4148 4115 4192
rect 4045 4128 4051 4132
rect 3837 3888 3843 3892
rect 3933 3808 3939 3912
rect 3949 3868 3955 3912
rect 4045 3908 4051 4112
rect 4109 4108 4115 4132
rect 4077 3908 4083 3992
rect 3965 3848 3971 3892
rect 4029 3868 4035 3872
rect 4045 3788 4051 3892
rect 3917 3768 3923 3772
rect 3784 3737 3795 3743
rect 3549 3583 3555 3672
rect 3597 3588 3603 3732
rect 3661 3708 3667 3732
rect 3741 3708 3747 3712
rect 3677 3697 3688 3703
rect 3549 3577 3560 3583
rect 3517 3528 3523 3552
rect 3549 3488 3555 3532
rect 3597 3468 3603 3492
rect 3613 3488 3619 3532
rect 3325 3348 3331 3352
rect 3293 3248 3299 3312
rect 3357 3308 3363 3312
rect 3085 3068 3091 3072
rect 3117 3068 3123 3092
rect 3341 3088 3347 3092
rect 2957 2848 2963 3032
rect 2973 2988 2979 2992
rect 2989 2943 2995 2992
rect 3165 2968 3171 3052
rect 2984 2937 2995 2943
rect 3037 2883 3043 2932
rect 3053 2908 3059 2952
rect 3197 2948 3203 3072
rect 3277 3043 3283 3072
rect 3261 3037 3283 3043
rect 3261 2968 3267 3037
rect 3357 2968 3363 3272
rect 3069 2928 3075 2932
rect 3357 2928 3363 2952
rect 3421 2948 3427 3332
rect 3437 3108 3443 3312
rect 3501 3128 3507 3192
rect 3437 2948 3443 2992
rect 3453 2948 3459 2952
rect 3533 2928 3539 3372
rect 3549 3308 3555 3312
rect 3565 3008 3571 3072
rect 3613 2948 3619 3332
rect 3629 3188 3635 3252
rect 3645 3088 3651 3412
rect 3661 3308 3667 3492
rect 3677 3388 3683 3697
rect 3741 3508 3747 3652
rect 3837 3588 3843 3632
rect 3901 3588 3907 3672
rect 3981 3588 3987 3692
rect 3853 3528 3859 3532
rect 3917 3528 3923 3572
rect 3677 3108 3683 3232
rect 3757 3208 3763 3232
rect 3741 3108 3747 3112
rect 3773 3088 3779 3432
rect 3789 3248 3795 3312
rect 3805 3268 3811 3472
rect 3853 3388 3859 3492
rect 3917 3328 3923 3492
rect 3773 3068 3779 3072
rect 3805 2988 3811 2992
rect 3821 2968 3827 3132
rect 3837 3106 3843 3112
rect 3949 3108 3955 3112
rect 3917 3088 3923 3092
rect 3965 3088 3971 3332
rect 3997 3328 4003 3332
rect 3981 3108 3987 3112
rect 4045 3108 4051 3732
rect 4061 3588 4067 3852
rect 4093 3808 4099 3912
rect 4125 3908 4131 4217
rect 4173 4148 4179 4232
rect 4205 4148 4211 4152
rect 4237 4148 4243 4212
rect 4269 4188 4275 4232
rect 4349 4228 4355 4292
rect 4365 4188 4371 4272
rect 4477 4248 4483 4292
rect 4589 4288 4595 4532
rect 4381 4208 4387 4232
rect 4381 4168 4387 4172
rect 4397 4148 4403 4152
rect 4141 4048 4147 4092
rect 4109 3748 4115 3752
rect 4141 3748 4147 4032
rect 4205 3948 4211 4132
rect 4173 3868 4179 3872
rect 4109 3508 4115 3512
rect 4077 3388 4083 3452
rect 3821 2948 3827 2952
rect 3549 2928 3555 2932
rect 3069 2888 3075 2912
rect 3037 2877 3059 2883
rect 3053 2788 3059 2877
rect 2941 2708 2947 2712
rect 2909 2668 2915 2672
rect 3037 2668 3043 2672
rect 3069 2648 3075 2872
rect 3149 2728 3155 2772
rect 3309 2706 3315 2872
rect 3085 2668 3091 2672
rect 3117 2648 3123 2672
rect 2941 2568 2947 2572
rect 2797 2488 2803 2532
rect 2749 2308 2755 2452
rect 2061 2208 2067 2252
rect 2061 2188 2067 2192
rect 2173 2128 2179 2132
rect 1997 1968 2003 2112
rect 1757 1908 1763 1912
rect 1869 1906 1875 1912
rect 1773 1888 1779 1892
rect 1709 1488 1715 1512
rect 1725 1508 1731 1512
rect 1741 1508 1747 1532
rect 1613 1288 1619 1292
rect 1037 928 1043 1072
rect 1213 1068 1219 1072
rect 1229 968 1235 1072
rect 1149 928 1155 952
rect 957 877 968 883
rect 765 688 771 692
rect 829 668 835 692
rect 893 688 899 692
rect 797 648 803 652
rect 509 148 515 192
rect 477 128 483 132
rect 589 -43 595 292
rect 669 288 675 292
rect 685 288 691 292
rect 669 228 675 272
rect 717 128 723 272
rect 781 148 787 412
rect 829 408 835 652
rect 925 648 931 752
rect 973 748 979 872
rect 989 868 995 892
rect 1005 768 1011 892
rect 1021 748 1027 872
rect 989 723 995 732
rect 973 717 995 723
rect 957 668 963 672
rect 845 528 851 612
rect 861 528 867 632
rect 925 588 931 632
rect 845 428 851 512
rect 861 168 867 252
rect 877 188 883 252
rect 893 148 899 392
rect 973 348 979 717
rect 989 688 995 692
rect 1005 308 1011 692
rect 1021 688 1027 712
rect 1037 708 1043 912
rect 1069 748 1075 752
rect 1037 668 1043 692
rect 1053 388 1059 732
rect 1069 708 1075 712
rect 1085 688 1091 712
rect 1101 708 1107 712
rect 1149 688 1155 812
rect 1165 728 1171 732
rect 1229 723 1235 952
rect 1261 948 1267 952
rect 1293 948 1299 1072
rect 1389 948 1395 1172
rect 1469 1088 1475 1172
rect 1501 1108 1507 1132
rect 1533 1128 1539 1172
rect 1565 1108 1571 1152
rect 1581 1108 1587 1112
rect 1581 1088 1587 1092
rect 1517 1068 1523 1072
rect 1309 908 1315 912
rect 1261 897 1272 903
rect 1261 788 1267 897
rect 1341 888 1347 892
rect 1245 748 1251 772
rect 1213 717 1235 723
rect 1213 688 1219 717
rect 1261 708 1267 712
rect 1069 548 1075 612
rect 1085 563 1091 672
rect 1101 588 1107 632
rect 1213 608 1219 672
rect 1261 648 1267 692
rect 1245 568 1251 632
rect 1261 568 1267 572
rect 1085 557 1096 563
rect 1064 377 1075 383
rect 1069 348 1075 377
rect 925 248 931 290
rect 973 188 979 232
rect 893 128 899 132
rect 957 128 963 132
rect 1037 128 1043 312
rect 1069 268 1075 312
rect 1101 308 1107 332
rect 1117 128 1123 172
rect 1133 148 1139 472
rect 1149 388 1155 472
rect 1165 388 1171 492
rect 1245 448 1251 512
rect 1165 308 1171 372
rect 1181 288 1187 312
rect 1229 308 1235 312
rect 1261 268 1267 432
rect 1277 343 1283 732
rect 1293 448 1299 712
rect 1309 668 1315 692
rect 1309 388 1315 492
rect 1325 348 1331 732
rect 1357 548 1363 932
rect 1389 828 1395 932
rect 1405 728 1411 932
rect 1453 928 1459 1012
rect 1421 708 1427 892
rect 1277 337 1288 343
rect 1309 308 1315 332
rect 1197 130 1203 232
rect 1261 168 1267 252
rect 1325 168 1331 312
rect 1341 188 1347 512
rect 1357 497 1368 503
rect 1357 388 1363 497
rect 1389 208 1395 692
rect 1421 568 1427 672
rect 1421 548 1427 552
rect 1437 408 1443 912
rect 1533 788 1539 932
rect 1597 930 1603 1032
rect 1565 708 1571 872
rect 1613 748 1619 1272
rect 1629 1263 1635 1472
rect 1661 1288 1667 1412
rect 1677 1368 1683 1452
rect 1677 1328 1683 1352
rect 1677 1263 1683 1292
rect 1741 1288 1747 1432
rect 1629 1257 1651 1263
rect 1645 948 1651 1257
rect 1661 1257 1683 1263
rect 1661 1068 1667 1257
rect 1677 1088 1683 1192
rect 1725 1188 1731 1232
rect 1741 1128 1747 1192
rect 1773 1108 1779 1872
rect 1789 1808 1795 1892
rect 1837 1868 1843 1872
rect 1837 1728 1843 1812
rect 1933 1768 1939 1852
rect 2029 1788 2035 1852
rect 2013 1768 2019 1772
rect 1933 1728 1939 1752
rect 1821 1688 1827 1712
rect 1837 1708 1843 1712
rect 1885 1688 1891 1712
rect 1789 1528 1795 1532
rect 1805 1448 1811 1672
rect 1821 1528 1827 1632
rect 1837 1508 1843 1632
rect 1837 1468 1843 1492
rect 1789 1328 1795 1332
rect 1837 1328 1843 1332
rect 1853 1263 1859 1512
rect 1869 1308 1875 1672
rect 1949 1663 1955 1712
rect 1981 1708 1987 1752
rect 2045 1728 2051 1872
rect 2077 1728 2083 1832
rect 1933 1657 1955 1663
rect 1885 1528 1891 1632
rect 1901 1468 1907 1492
rect 1869 1288 1875 1292
rect 1901 1263 1907 1452
rect 1933 1368 1939 1657
rect 1949 1548 1955 1632
rect 1997 1508 2003 1552
rect 1997 1448 2003 1452
rect 2013 1428 2019 1432
rect 2077 1408 2083 1592
rect 2109 1588 2115 1892
rect 2141 1748 2147 1872
rect 2173 1748 2179 2112
rect 2189 1988 2195 2172
rect 2205 2148 2211 2272
rect 2221 2168 2227 2232
rect 2269 2168 2275 2272
rect 2429 2248 2435 2252
rect 2557 2248 2563 2272
rect 2301 2148 2307 2192
rect 2285 1908 2291 2072
rect 2317 2008 2323 2112
rect 2253 1788 2259 1832
rect 2333 1788 2339 2092
rect 2349 1988 2355 1992
rect 2381 1888 2387 2132
rect 2429 2128 2435 2232
rect 2637 2228 2643 2232
rect 2493 2108 2499 2112
rect 2557 2108 2563 2132
rect 2413 1988 2419 2092
rect 2397 1888 2403 1912
rect 2525 1908 2531 2092
rect 2141 1708 2147 1712
rect 2269 1708 2275 1752
rect 2125 1528 2131 1532
rect 2093 1508 2099 1512
rect 2109 1488 2115 1492
rect 1933 1328 1939 1352
rect 2077 1328 2083 1392
rect 1853 1257 1875 1263
rect 1901 1257 1923 1263
rect 1693 1088 1699 1092
rect 1789 1088 1795 1172
rect 1837 1128 1843 1252
rect 1853 1208 1859 1232
rect 1821 1108 1827 1112
rect 1869 1108 1875 1257
rect 1901 1108 1907 1112
rect 1805 1088 1811 1092
rect 1661 968 1667 1052
rect 1773 948 1779 1072
rect 1789 948 1795 1072
rect 1693 888 1699 912
rect 1917 788 1923 1257
rect 2093 1228 2099 1332
rect 2109 1328 2115 1352
rect 2141 1308 2147 1532
rect 2157 1508 2163 1512
rect 2189 1488 2195 1612
rect 2237 1528 2243 1552
rect 2157 1477 2168 1483
rect 1933 1188 1939 1212
rect 1997 728 2003 932
rect 2045 928 2051 1192
rect 2125 1108 2131 1292
rect 2157 1188 2163 1477
rect 2205 1468 2211 1492
rect 2253 1448 2259 1472
rect 2285 1468 2291 1712
rect 2301 1688 2307 1692
rect 2317 1568 2323 1632
rect 2173 1328 2179 1372
rect 2205 1328 2211 1332
rect 2237 1328 2243 1332
rect 2125 968 2131 1072
rect 2141 928 2147 1052
rect 2173 988 2179 1312
rect 2269 1308 2275 1352
rect 2285 1328 2291 1452
rect 2365 1348 2371 1872
rect 2381 1748 2387 1752
rect 2381 1648 2387 1732
rect 2397 1708 2403 1872
rect 2477 1748 2483 1872
rect 2397 1568 2403 1692
rect 2429 1548 2435 1632
rect 2397 1468 2403 1512
rect 2509 1508 2515 1552
rect 2477 1488 2483 1492
rect 2445 1468 2451 1472
rect 2333 1128 2339 1292
rect 2349 1168 2355 1312
rect 2509 1308 2515 1492
rect 2525 1463 2531 1872
rect 2573 1748 2579 2012
rect 2605 1948 2611 2132
rect 2557 1708 2563 1712
rect 2568 1517 2579 1523
rect 2525 1457 2547 1463
rect 2541 1348 2547 1457
rect 2573 1388 2579 1517
rect 2637 1348 2643 1692
rect 2669 1568 2675 2292
rect 2717 2208 2723 2232
rect 2685 2088 2691 2092
rect 2685 1988 2691 2072
rect 2749 1983 2755 2292
rect 2797 2288 2803 2412
rect 2877 2288 2883 2292
rect 2781 2148 2787 2192
rect 2941 2188 2947 2432
rect 3037 2328 3043 2492
rect 2957 2148 2963 2232
rect 3005 2188 3011 2312
rect 3037 2308 3043 2312
rect 3053 2308 3059 2472
rect 3069 2308 3075 2532
rect 3053 2288 3059 2292
rect 2877 2128 2883 2132
rect 2829 2103 2835 2112
rect 2829 2097 2840 2103
rect 2829 1988 2835 2097
rect 2749 1977 2760 1983
rect 2861 1908 2867 1972
rect 2893 1888 2899 2132
rect 2925 2097 2936 2103
rect 2925 1943 2931 2097
rect 2957 2043 2963 2132
rect 3037 2108 3043 2152
rect 3069 2088 3075 2212
rect 2941 2037 2963 2043
rect 2941 1968 2947 2037
rect 2925 1937 2947 1943
rect 2653 1488 2659 1492
rect 2269 1108 2275 1112
rect 2317 1108 2323 1112
rect 2493 1088 2499 1252
rect 2541 1088 2547 1332
rect 2221 968 2227 1072
rect 1773 706 1779 712
rect 1869 708 1875 712
rect 1453 628 1459 632
rect 1453 568 1459 572
rect 1453 528 1459 532
rect 1485 528 1491 532
rect 1453 383 1459 412
rect 1448 377 1459 383
rect 1453 248 1459 312
rect 1501 308 1507 312
rect 1517 288 1523 672
rect 1805 668 1811 672
rect 1741 548 1747 592
rect 1773 528 1779 632
rect 1869 548 1875 592
rect 1885 588 1891 712
rect 1997 708 2003 712
rect 1933 548 1939 552
rect 1533 468 1539 472
rect 1725 448 1731 512
rect 1853 508 1859 512
rect 1917 508 1923 512
rect 1997 508 2003 692
rect 2093 548 2099 812
rect 2237 728 2243 992
rect 2301 988 2307 1012
rect 2397 948 2403 952
rect 2205 708 2211 712
rect 2285 688 2291 912
rect 2333 888 2339 912
rect 2157 668 2163 672
rect 2285 643 2291 672
rect 2269 637 2291 643
rect 2269 588 2275 637
rect 2125 548 2131 552
rect 2269 548 2275 572
rect 2333 548 2339 652
rect 1757 403 1763 492
rect 1789 488 1795 492
rect 1741 397 1763 403
rect 1581 308 1587 372
rect 1565 288 1571 292
rect 1469 248 1475 252
rect 1581 228 1587 292
rect 1341 168 1347 172
rect 1597 148 1603 152
rect 1677 128 1683 332
rect 1741 248 1747 397
rect 1853 308 1859 492
rect 1885 428 1891 492
rect 1869 308 1875 332
rect 1933 328 1939 332
rect 1997 328 2003 492
rect 2029 428 2035 532
rect 2109 528 2115 532
rect 2045 468 2051 492
rect 2141 448 2147 512
rect 2157 508 2163 512
rect 2029 308 2035 412
rect 2141 388 2147 432
rect 1741 188 1747 232
rect 1773 168 1779 272
rect 1853 128 1859 252
rect 1933 208 1939 232
rect 1933 188 1939 192
rect 1901 148 1907 152
rect 1997 148 2003 292
rect 2029 228 2035 272
rect 2061 268 2067 312
rect 2109 268 2115 292
rect 2189 148 2195 152
rect 2221 148 2227 232
rect 1517 108 1523 112
rect 1629 108 1635 112
rect 1677 108 1683 112
rect 1821 -43 1827 12
rect 1997 -43 2003 132
rect 2237 128 2243 332
rect 2333 288 2339 532
rect 2381 528 2387 872
rect 2429 828 2435 1072
rect 2445 1008 2451 1032
rect 2445 928 2451 952
rect 2445 908 2451 912
rect 2493 648 2499 1072
rect 2541 1028 2547 1072
rect 2573 988 2579 1272
rect 2589 1108 2595 1332
rect 2621 1268 2627 1332
rect 2669 1288 2675 1552
rect 2765 1508 2771 1732
rect 2781 1508 2787 1512
rect 2733 1488 2739 1492
rect 2797 1348 2803 1572
rect 2813 1548 2819 1872
rect 2701 1308 2707 1312
rect 2605 988 2611 1152
rect 2493 528 2499 612
rect 2333 208 2339 272
rect 2333 168 2339 192
rect 2365 168 2371 392
rect 2157 108 2163 114
rect 2285 108 2291 112
rect 2397 -37 2403 432
rect 2509 428 2515 532
rect 2541 423 2547 932
rect 2573 788 2579 832
rect 2589 688 2595 812
rect 2621 708 2627 1132
rect 2669 1128 2675 1232
rect 2701 1208 2707 1292
rect 2701 988 2707 1172
rect 2717 1168 2723 1332
rect 2733 1128 2739 1312
rect 2749 1297 2760 1303
rect 2749 1188 2755 1297
rect 2733 1088 2739 1092
rect 2749 988 2755 1152
rect 2813 1148 2819 1512
rect 2845 1488 2851 1872
rect 2893 1868 2899 1872
rect 2893 1748 2899 1852
rect 2925 1848 2931 1912
rect 2941 1788 2947 1937
rect 2973 1908 2979 1952
rect 3053 1923 3059 2032
rect 3048 1917 3059 1923
rect 3069 1908 3075 1912
rect 3069 1888 3075 1892
rect 3085 1888 3091 2332
rect 3101 2148 3107 2512
rect 3149 2508 3155 2632
rect 3277 2548 3283 2672
rect 3261 2528 3267 2532
rect 3133 2128 3139 2492
rect 3149 2308 3155 2312
rect 3149 2288 3155 2292
rect 3149 2148 3155 2152
rect 3197 2128 3203 2232
rect 3213 2188 3219 2292
rect 3261 2288 3267 2512
rect 3325 2288 3331 2292
rect 3213 2148 3219 2152
rect 3117 2088 3123 2092
rect 3117 1908 3123 2032
rect 3181 1968 3187 2012
rect 3197 1988 3203 2032
rect 3165 1888 3171 1892
rect 3181 1888 3187 1952
rect 3229 1928 3235 2032
rect 3197 1908 3203 1912
rect 2989 1868 2995 1872
rect 3053 1748 3059 1832
rect 3085 1768 3091 1872
rect 3277 1808 3283 2092
rect 3325 2068 3331 2112
rect 3341 2108 3347 2752
rect 3389 2748 3395 2892
rect 3405 2888 3411 2912
rect 3421 2908 3427 2912
rect 3421 2728 3427 2892
rect 3453 2708 3459 2732
rect 3549 2728 3555 2732
rect 3597 2708 3603 2932
rect 3741 2928 3747 2932
rect 3837 2928 3843 2952
rect 3869 2948 3875 3072
rect 4013 3068 4019 3072
rect 3901 2948 3907 2992
rect 4045 2948 4051 2992
rect 3645 2728 3651 2732
rect 3517 2688 3523 2692
rect 3597 2688 3603 2692
rect 3645 2688 3651 2712
rect 3421 2648 3427 2672
rect 3501 2663 3507 2672
rect 3501 2657 3523 2663
rect 3421 2548 3427 2632
rect 3485 2508 3491 2572
rect 3501 2528 3507 2532
rect 3517 2508 3523 2657
rect 3597 2648 3603 2672
rect 3629 2663 3635 2672
rect 3629 2657 3651 2663
rect 3645 2588 3651 2657
rect 3677 2588 3683 2712
rect 3741 2688 3747 2812
rect 3533 2528 3539 2572
rect 3677 2548 3683 2552
rect 3405 2348 3411 2432
rect 3501 2328 3507 2332
rect 3549 2328 3555 2532
rect 3597 2448 3603 2472
rect 3448 2317 3459 2323
rect 3453 2243 3459 2317
rect 3469 2263 3475 2292
rect 3485 2288 3491 2312
rect 3469 2257 3491 2263
rect 3453 2237 3475 2243
rect 3421 2148 3427 2232
rect 3469 2188 3475 2237
rect 3373 2128 3379 2132
rect 3421 2128 3427 2132
rect 3485 2108 3491 2257
rect 3336 2037 3347 2043
rect 3309 1948 3315 1952
rect 3341 1888 3347 2037
rect 3357 1948 3363 2072
rect 3357 1908 3363 1912
rect 3357 1868 3363 1892
rect 3373 1828 3379 1932
rect 3373 1788 3379 1792
rect 3405 1788 3411 2032
rect 3485 1968 3491 2092
rect 3421 1928 3427 1932
rect 3501 1908 3507 2232
rect 3549 2168 3555 2292
rect 3565 2288 3571 2352
rect 3549 2148 3555 2152
rect 3597 2148 3603 2432
rect 3741 2408 3747 2672
rect 3757 2588 3763 2692
rect 3773 2528 3779 2752
rect 3853 2688 3859 2692
rect 3869 2688 3875 2932
rect 3933 2908 3939 2932
rect 3773 2388 3779 2512
rect 3821 2508 3827 2592
rect 3709 2306 3715 2332
rect 3773 2288 3779 2312
rect 3805 2308 3811 2332
rect 3837 2328 3843 2672
rect 3869 2528 3875 2592
rect 3885 2548 3891 2652
rect 3901 2588 3907 2612
rect 3933 2528 3939 2632
rect 3965 2608 3971 2932
rect 4013 2728 4019 2732
rect 3981 2648 3987 2672
rect 4045 2648 4051 2932
rect 4061 2928 4067 3152
rect 4109 3128 4115 3252
rect 4077 3088 4083 3092
rect 4125 2988 4131 3112
rect 4141 3108 4147 3452
rect 4173 3368 4179 3852
rect 4205 3748 4211 3932
rect 4221 3828 4227 3892
rect 4189 3528 4195 3712
rect 4237 3708 4243 4112
rect 4301 4108 4307 4132
rect 4461 4108 4467 4112
rect 4189 3508 4195 3512
rect 4221 3488 4227 3552
rect 4253 3388 4259 4092
rect 4301 4068 4307 4092
rect 4333 4048 4339 4092
rect 4317 3948 4323 4032
rect 4509 3888 4515 4272
rect 4589 4168 4595 4272
rect 4605 4128 4611 4132
rect 4605 3928 4611 4072
rect 4637 3963 4643 4572
rect 4669 4543 4675 4832
rect 4765 4828 4771 4912
rect 4861 4908 4867 4912
rect 4813 4788 4819 4832
rect 4685 4588 4691 4632
rect 4765 4568 4771 4652
rect 4845 4583 4851 4692
rect 4861 4648 4867 4652
rect 4845 4577 4856 4583
rect 4669 4537 4680 4543
rect 4701 4528 4707 4532
rect 4765 4508 4771 4552
rect 4813 4548 4819 4552
rect 4925 4548 4931 4752
rect 4973 4588 4979 4812
rect 4989 4688 4995 4692
rect 5069 4588 5075 4832
rect 4733 4468 4739 4492
rect 4653 4308 4659 4432
rect 4685 4308 4691 4352
rect 4781 4328 4787 4432
rect 4813 4308 4819 4512
rect 4685 4148 4691 4152
rect 4621 3957 4643 3963
rect 4605 3908 4611 3912
rect 4557 3888 4563 3892
rect 4317 3728 4323 3732
rect 4301 3488 4307 3712
rect 4317 3448 4323 3472
rect 4237 3348 4243 3352
rect 4349 3328 4355 3812
rect 4429 3748 4435 3872
rect 4605 3828 4611 3892
rect 4621 3888 4627 3957
rect 4637 3928 4643 3932
rect 4653 3908 4659 3912
rect 4669 3908 4675 4032
rect 4701 3928 4707 3972
rect 4717 3968 4723 4232
rect 4765 4148 4771 4212
rect 4749 3988 4755 4032
rect 4445 3748 4451 3812
rect 4477 3708 4483 3752
rect 4509 3748 4515 3812
rect 4621 3808 4627 3872
rect 4669 3828 4675 3892
rect 4685 3868 4691 3872
rect 4525 3788 4531 3792
rect 4573 3748 4579 3752
rect 4509 3608 4515 3732
rect 4509 3528 4515 3532
rect 4557 3528 4563 3692
rect 4637 3508 4643 3772
rect 4605 3468 4611 3492
rect 4637 3488 4643 3492
rect 4221 3308 4227 3312
rect 4221 3208 4227 3292
rect 4157 3008 4163 3092
rect 4237 3068 4243 3072
rect 4157 2968 4163 2992
rect 4205 2948 4211 3052
rect 4301 3008 4307 3312
rect 4317 3288 4323 3292
rect 4317 3128 4323 3192
rect 4317 3108 4323 3112
rect 4173 2888 4179 2892
rect 4061 2668 4067 2672
rect 4077 2588 4083 2692
rect 4109 2588 4115 2712
rect 4221 2688 4227 2692
rect 3997 2548 4003 2552
rect 3853 2448 3859 2512
rect 3645 2268 3651 2272
rect 3645 2163 3651 2252
rect 3741 2168 3747 2272
rect 3645 2157 3656 2163
rect 3869 2163 3875 2392
rect 3885 2328 3891 2512
rect 3901 2508 3907 2512
rect 3917 2388 3923 2492
rect 3949 2388 3955 2532
rect 4061 2488 4067 2532
rect 4077 2528 4083 2572
rect 4141 2548 4147 2632
rect 4173 2548 4179 2572
rect 4237 2563 4243 2992
rect 4333 2948 4339 3132
rect 4349 3068 4355 3072
rect 4269 2908 4275 2914
rect 4365 2908 4371 2912
rect 4397 2708 4403 3452
rect 4605 3348 4611 3432
rect 4653 3308 4659 3812
rect 4669 3748 4675 3792
rect 4696 3737 4707 3743
rect 4669 3708 4675 3712
rect 4685 3608 4691 3712
rect 4669 3528 4675 3532
rect 4429 3106 4435 3112
rect 4493 3108 4499 3132
rect 4669 3128 4675 3432
rect 4685 3428 4691 3592
rect 4701 3588 4707 3737
rect 4717 3508 4723 3952
rect 4749 3888 4755 3932
rect 4765 3908 4771 4132
rect 4781 4088 4787 4232
rect 4797 4148 4803 4172
rect 4781 3988 4787 4052
rect 4765 3848 4771 3892
rect 4733 3788 4739 3832
rect 4765 3788 4771 3832
rect 4813 3808 4819 4292
rect 4829 4288 4835 4532
rect 4893 4508 4899 4512
rect 4829 4228 4835 4272
rect 4845 4128 4851 4492
rect 4861 4388 4867 4452
rect 4909 4288 4915 4312
rect 4925 4143 4931 4532
rect 4989 4308 4995 4312
rect 4920 4137 4931 4143
rect 4845 3888 4851 4112
rect 4877 4108 4883 4112
rect 4861 3908 4867 3912
rect 4765 3703 4771 3752
rect 4760 3697 4771 3703
rect 4717 3408 4723 3452
rect 4749 3428 4755 3492
rect 4717 3188 4723 3272
rect 4557 2948 4563 2992
rect 4637 2968 4643 3092
rect 4669 3028 4675 3032
rect 4685 2948 4691 3112
rect 4717 2988 4723 3112
rect 4733 3088 4739 3412
rect 4749 3348 4755 3412
rect 4765 3348 4771 3352
rect 4749 3308 4755 3312
rect 4781 3308 4787 3312
rect 4781 3208 4787 3292
rect 4797 3088 4803 3412
rect 4829 3108 4835 3812
rect 4845 3728 4851 3732
rect 4861 3488 4867 3872
rect 4877 3568 4883 4092
rect 4973 3888 4979 3892
rect 4941 3868 4947 3872
rect 4893 3768 4899 3772
rect 4973 3708 4979 3712
rect 4989 3708 4995 4292
rect 5005 4288 5011 4532
rect 5085 4508 5091 4692
rect 5117 4668 5123 4772
rect 5181 4688 5187 4997
rect 5245 4988 5251 5112
rect 5309 5108 5315 5292
rect 5437 5288 5443 5312
rect 5549 5308 5555 5312
rect 5565 5283 5571 5332
rect 5549 5277 5571 5283
rect 5277 4908 5283 5092
rect 5293 5028 5299 5072
rect 5341 5048 5347 5072
rect 5341 4968 5347 5032
rect 5197 4708 5203 4712
rect 5229 4708 5235 4772
rect 5261 4668 5267 4692
rect 5309 4648 5315 4652
rect 5229 4568 5235 4612
rect 5277 4588 5283 4592
rect 5293 4528 5299 4552
rect 5325 4548 5331 4632
rect 5341 4548 5347 4632
rect 5373 4628 5379 4692
rect 5405 4608 5411 5232
rect 5485 4928 5491 5272
rect 5501 4948 5507 5032
rect 5517 4948 5523 5032
rect 5421 4708 5427 4712
rect 5437 4708 5443 4732
rect 5453 4728 5459 4732
rect 5469 4728 5475 4832
rect 5485 4708 5491 4912
rect 5501 4703 5507 4932
rect 5517 4928 5523 4932
rect 5549 4848 5555 5277
rect 5565 5268 5571 5277
rect 5565 4928 5571 5032
rect 5581 4948 5587 5012
rect 5597 4928 5603 5352
rect 5789 5348 5795 5452
rect 5853 5388 5859 5452
rect 5885 5428 5891 5472
rect 5613 5108 5619 5232
rect 5709 5148 5715 5232
rect 5757 5108 5763 5332
rect 5837 5308 5843 5312
rect 5645 4988 5651 5092
rect 5757 5088 5763 5092
rect 5773 4948 5779 5012
rect 5821 4988 5827 5292
rect 5885 5188 5891 5312
rect 5901 5308 5907 5432
rect 5917 5388 5923 5512
rect 5933 5368 5939 5452
rect 5949 5448 5955 5492
rect 5997 5488 6003 5492
rect 6093 5488 6099 5512
rect 5965 5468 5971 5472
rect 5997 5428 6003 5452
rect 5997 5388 6003 5412
rect 5901 5168 5907 5292
rect 5837 5088 5843 5092
rect 5901 4988 5907 5152
rect 5933 5088 5939 5352
rect 5949 5148 5955 5332
rect 6125 5323 6131 5472
rect 6253 5468 6259 5472
rect 6301 5348 6307 5352
rect 6205 5328 6211 5332
rect 6120 5317 6131 5323
rect 6029 5308 6035 5312
rect 5949 5108 5955 5112
rect 6093 5108 6099 5312
rect 6237 5308 6243 5312
rect 6109 5108 6115 5132
rect 6029 5088 6035 5092
rect 5949 4948 5955 4952
rect 5997 4928 6003 4932
rect 5896 4917 5907 4923
rect 5533 4748 5539 4832
rect 5613 4728 5619 4912
rect 5709 4908 5715 4912
rect 5629 4897 5640 4903
rect 5629 4788 5635 4897
rect 5565 4708 5571 4712
rect 5501 4697 5512 4703
rect 5421 4668 5427 4672
rect 5485 4583 5491 4652
rect 5613 4628 5619 4712
rect 5693 4708 5699 4732
rect 5661 4668 5667 4672
rect 5661 4648 5667 4652
rect 5677 4648 5683 4692
rect 5485 4577 5496 4583
rect 5133 4388 5139 4512
rect 5197 4508 5203 4512
rect 5005 3888 5011 3912
rect 5085 3888 5091 3892
rect 5101 3888 5107 3992
rect 5005 3748 5011 3832
rect 4877 3506 4883 3532
rect 4941 3488 4947 3512
rect 4973 3488 4979 3512
rect 4989 3503 4995 3692
rect 5005 3528 5011 3532
rect 5069 3508 5075 3532
rect 4989 3497 5011 3503
rect 4749 2948 4755 3032
rect 4413 2888 4419 2932
rect 4573 2928 4579 2932
rect 4781 2928 4787 2932
rect 4461 2908 4467 2912
rect 4669 2728 4675 2752
rect 4717 2728 4723 2892
rect 4829 2828 4835 2832
rect 4845 2803 4851 3072
rect 4861 3008 4867 3472
rect 4877 3348 4883 3392
rect 4989 3328 4995 3332
rect 4925 3188 4931 3292
rect 4973 3108 4979 3232
rect 5005 3188 5011 3497
rect 5037 3488 5043 3492
rect 5085 3488 5091 3872
rect 5133 3588 5139 4372
rect 5181 4168 5187 4272
rect 5181 4148 5187 4152
rect 5149 3748 5155 4132
rect 5277 4108 5283 4112
rect 5213 3908 5219 3912
rect 5197 3868 5203 3872
rect 5229 3748 5235 3752
rect 5261 3508 5267 3572
rect 5069 3428 5075 3432
rect 5069 3348 5075 3412
rect 5101 3343 5107 3492
rect 5197 3428 5203 3432
rect 5101 3337 5123 3343
rect 4877 3088 4883 3092
rect 4973 2988 4979 3092
rect 4989 2988 4995 3092
rect 5037 3088 5043 3092
rect 5037 3068 5043 3072
rect 4829 2797 4851 2803
rect 4749 2708 4755 2752
rect 4333 2688 4339 2692
rect 4669 2688 4675 2692
rect 4221 2557 4243 2563
rect 4109 2508 4115 2512
rect 4141 2508 4147 2532
rect 4061 2428 4067 2472
rect 4205 2448 4211 2492
rect 3885 2308 3891 2312
rect 4061 2308 4067 2312
rect 4077 2308 4083 2432
rect 4221 2388 4227 2557
rect 4269 2548 4275 2652
rect 4301 2528 4307 2672
rect 4381 2528 4387 2532
rect 4253 2488 4259 2512
rect 4237 2328 4243 2432
rect 4189 2317 4200 2323
rect 3869 2157 3891 2163
rect 3885 2148 3891 2157
rect 3965 2148 3971 2252
rect 4189 2248 4195 2317
rect 4333 2308 4339 2412
rect 4413 2328 4419 2532
rect 4429 2528 4435 2532
rect 4141 2148 4147 2192
rect 4205 2148 4211 2292
rect 4349 2288 4355 2292
rect 4285 2248 4291 2252
rect 4301 2208 4307 2232
rect 4349 2188 4355 2232
rect 4269 2148 4275 2152
rect 3517 2108 3523 2112
rect 3485 1888 3491 1892
rect 3213 1728 3219 1732
rect 2893 1708 2899 1712
rect 2893 1548 2899 1692
rect 2989 1683 2995 1692
rect 2989 1677 3011 1683
rect 3005 1588 3011 1677
rect 2845 1148 2851 1472
rect 2877 1328 2883 1532
rect 2893 1528 2899 1532
rect 2941 1508 2947 1532
rect 3133 1488 3139 1492
rect 2813 988 2819 1112
rect 2829 1068 2835 1112
rect 2637 848 2643 912
rect 2781 888 2787 912
rect 2589 668 2595 672
rect 2621 563 2627 692
rect 2653 588 2659 712
rect 2749 688 2755 832
rect 2637 563 2643 572
rect 2621 557 2643 563
rect 2557 508 2563 512
rect 2621 508 2627 532
rect 2637 508 2643 557
rect 2685 548 2691 632
rect 2749 608 2755 672
rect 2781 568 2787 692
rect 2797 688 2803 892
rect 2525 417 2547 423
rect 2509 288 2515 412
rect 2477 148 2483 272
rect 2509 148 2515 192
rect 2477 108 2483 132
rect 2397 -43 2419 -37
rect 2525 -43 2531 417
rect 2541 388 2547 392
rect 2557 328 2563 492
rect 2557 288 2563 312
rect 2637 308 2643 332
rect 2605 148 2611 152
rect 2621 128 2627 252
rect 2669 228 2675 272
rect 2685 248 2691 532
rect 2749 308 2755 312
rect 2813 288 2819 592
rect 2653 -43 2659 212
rect 2733 148 2739 272
rect 2845 148 2851 232
rect 2861 188 2867 1312
rect 2909 1108 2915 1332
rect 2941 1308 2947 1312
rect 3053 1243 3059 1332
rect 3085 1308 3091 1314
rect 3053 1237 3075 1243
rect 3053 1108 3059 1132
rect 3069 1108 3075 1237
rect 3229 1128 3235 1512
rect 3261 1388 3267 1732
rect 3341 1728 3347 1772
rect 3421 1728 3427 1832
rect 3453 1728 3459 1832
rect 3421 1668 3427 1672
rect 3437 1628 3443 1632
rect 3325 1508 3331 1592
rect 3469 1588 3475 1752
rect 3501 1728 3507 1832
rect 3533 1728 3539 1752
rect 3549 1588 3555 1712
rect 3453 1468 3459 1472
rect 3325 1457 3336 1463
rect 3293 1328 3299 1432
rect 3325 1388 3331 1457
rect 3373 1388 3379 1392
rect 3421 1388 3427 1452
rect 3325 1368 3331 1372
rect 3405 1368 3411 1372
rect 3437 1368 3443 1452
rect 3437 1328 3443 1352
rect 3453 1348 3459 1372
rect 3245 1088 3251 1092
rect 2877 948 2883 1072
rect 2893 988 2899 1052
rect 2973 1028 2979 1072
rect 3261 1063 3267 1232
rect 3245 1057 3267 1063
rect 2989 948 2995 1012
rect 3245 948 3251 1057
rect 2877 688 2883 932
rect 2909 788 2915 892
rect 2893 608 2899 652
rect 2973 588 2979 712
rect 3005 688 3011 692
rect 3037 583 3043 632
rect 3053 628 3059 712
rect 3085 688 3091 732
rect 3117 708 3123 712
rect 3149 708 3155 712
rect 3165 708 3171 932
rect 3277 928 3283 1032
rect 3293 888 3299 1312
rect 3485 1288 3491 1512
rect 3517 1408 3523 1492
rect 3501 1308 3507 1352
rect 3405 1128 3411 1132
rect 3341 1088 3347 1112
rect 3373 1088 3379 1112
rect 3421 1088 3427 1092
rect 3437 1088 3443 1132
rect 3357 988 3363 1052
rect 3389 948 3395 952
rect 3421 948 3427 1072
rect 3469 1068 3475 1072
rect 3485 1008 3491 1272
rect 3501 1108 3507 1112
rect 3421 908 3427 932
rect 3437 928 3443 932
rect 3469 928 3475 932
rect 3485 928 3491 932
rect 3261 706 3267 712
rect 3325 708 3331 872
rect 3357 728 3363 732
rect 3485 728 3491 852
rect 3501 768 3507 1092
rect 3517 888 3523 992
rect 3533 968 3539 1292
rect 3549 1108 3555 1352
rect 3565 1348 3571 2132
rect 3597 2128 3603 2132
rect 3581 2068 3587 2112
rect 3581 2048 3587 2052
rect 3613 1708 3619 1932
rect 3629 1908 3635 2032
rect 3661 1788 3667 1912
rect 3677 1908 3683 1992
rect 3709 1988 3715 2092
rect 3901 2088 3907 2112
rect 3757 1908 3763 1912
rect 3917 1908 3923 1972
rect 3629 1728 3635 1732
rect 3629 1683 3635 1712
rect 3613 1677 3635 1683
rect 3581 1508 3587 1632
rect 3597 1488 3603 1572
rect 3613 1548 3619 1677
rect 3661 1628 3667 1632
rect 3709 1588 3715 1692
rect 3613 1528 3619 1532
rect 3629 1508 3635 1512
rect 3565 1328 3571 1332
rect 3581 1108 3587 1472
rect 3613 1328 3619 1332
rect 3629 1308 3635 1492
rect 3661 1388 3667 1472
rect 3613 1288 3619 1292
rect 3613 1123 3619 1232
rect 3613 1117 3624 1123
rect 3597 1108 3603 1112
rect 3565 1088 3571 1092
rect 3581 1088 3587 1092
rect 3533 868 3539 912
rect 3549 908 3555 932
rect 3581 908 3587 972
rect 3629 928 3635 1032
rect 3645 948 3651 1312
rect 3693 1268 3699 1332
rect 3709 1288 3715 1432
rect 3725 1288 3731 1652
rect 3741 1508 3747 1552
rect 3741 1328 3747 1332
rect 3757 1328 3763 1792
rect 3773 1343 3779 1432
rect 3789 1368 3795 1832
rect 3821 1568 3827 1892
rect 3901 1708 3907 1872
rect 3965 1828 3971 1912
rect 3981 1908 3987 2132
rect 4013 2088 4019 2092
rect 4013 1928 4019 2072
rect 4045 2028 4051 2132
rect 4093 2128 4099 2132
rect 4141 2128 4147 2132
rect 4061 1988 4067 2112
rect 4141 1988 4147 2072
rect 4029 1888 4035 1892
rect 3965 1728 3971 1732
rect 3981 1708 3987 1772
rect 4045 1708 4051 1852
rect 4077 1808 4083 1832
rect 4125 1828 4131 1912
rect 3837 1488 3843 1692
rect 3997 1688 4003 1692
rect 3901 1568 3907 1632
rect 3933 1548 3939 1672
rect 3949 1668 3955 1672
rect 3997 1668 4003 1672
rect 3805 1348 3811 1432
rect 3853 1368 3859 1492
rect 3917 1448 3923 1492
rect 3965 1488 3971 1632
rect 4029 1548 4035 1632
rect 4013 1488 4019 1492
rect 3981 1437 3992 1443
rect 3981 1428 3987 1437
rect 3949 1368 3955 1412
rect 3773 1337 3795 1343
rect 3757 1308 3763 1312
rect 3789 1308 3795 1337
rect 3677 908 3683 1152
rect 3709 1148 3715 1272
rect 3725 1188 3731 1252
rect 3741 1123 3747 1232
rect 3757 1168 3763 1292
rect 3805 1288 3811 1312
rect 3837 1128 3843 1312
rect 3853 1308 3859 1352
rect 3869 1348 3875 1352
rect 3981 1348 3987 1392
rect 4045 1368 4051 1692
rect 4093 1588 4099 1692
rect 4141 1668 4147 1972
rect 4157 1888 4163 1892
rect 4173 1863 4179 1912
rect 4189 1908 4195 2012
rect 4237 1983 4243 2072
rect 4269 1988 4275 2072
rect 4237 1977 4248 1983
rect 4269 1948 4275 1972
rect 4157 1857 4179 1863
rect 4157 1728 4163 1857
rect 4173 1728 4179 1732
rect 4093 1568 4099 1572
rect 4109 1548 4115 1632
rect 4157 1488 4163 1632
rect 4173 1628 4179 1692
rect 4205 1683 4211 1932
rect 4237 1868 4243 1912
rect 4237 1788 4243 1812
rect 4253 1788 4259 1892
rect 4285 1808 4291 2092
rect 4301 2028 4307 2112
rect 4253 1728 4259 1772
rect 4200 1677 4216 1683
rect 3949 1328 3955 1332
rect 4013 1328 4019 1352
rect 3917 1308 3923 1312
rect 3997 1308 4003 1312
rect 3901 1268 3907 1272
rect 3885 1228 3891 1232
rect 3981 1128 3987 1132
rect 3741 1117 3752 1123
rect 3709 1108 3715 1112
rect 3805 1108 3811 1112
rect 3837 1088 3843 1092
rect 3789 1068 3795 1072
rect 3885 1068 3891 1092
rect 3981 1068 3987 1092
rect 4029 1088 4035 1332
rect 3757 1048 3763 1052
rect 3693 868 3699 912
rect 3709 888 3715 972
rect 3741 908 3747 932
rect 3533 728 3539 832
rect 3597 828 3603 832
rect 3629 728 3635 732
rect 3597 703 3603 712
rect 3597 697 3640 703
rect 3501 688 3507 692
rect 3021 577 3043 583
rect 3021 503 3027 577
rect 3037 548 3043 552
rect 3085 528 3091 612
rect 3133 548 3139 652
rect 3165 548 3171 632
rect 3021 497 3032 503
rect 3005 388 3011 492
rect 2861 168 2867 172
rect 2685 108 2691 112
rect 2717 108 2723 132
rect 2701 -43 2707 12
rect 2845 -43 2851 132
rect 2877 -43 2883 332
rect 2909 148 2915 272
rect 2941 108 2947 132
rect 2973 128 2979 312
rect 3005 288 3011 372
rect 3085 348 3091 512
rect 3101 388 3107 532
rect 3117 328 3123 352
rect 3165 328 3171 492
rect 3181 288 3187 672
rect 3261 583 3267 652
rect 3245 577 3267 583
rect 3197 528 3203 572
rect 2973 108 2979 112
rect 2941 -43 2947 92
rect 3005 -37 3011 192
rect 3213 148 3219 512
rect 3229 488 3235 492
rect 3245 468 3251 577
rect 3373 568 3379 592
rect 3501 548 3507 672
rect 3517 648 3523 672
rect 3565 663 3571 692
rect 3581 688 3587 692
rect 3549 657 3571 663
rect 3277 528 3283 532
rect 3245 288 3251 452
rect 3389 368 3395 432
rect 3309 308 3315 332
rect 3277 288 3283 292
rect 3341 288 3347 312
rect 3389 288 3395 352
rect 3069 128 3075 132
rect 3437 128 3443 332
rect 3485 188 3491 272
rect 3501 228 3507 272
rect 3517 128 3523 612
rect 3549 508 3555 657
rect 3565 448 3571 512
rect 3549 388 3555 392
rect 3037 108 3043 112
rect 3149 108 3155 114
rect 3325 108 3331 112
rect 2989 -43 3011 -37
rect 3341 -43 3347 32
rect 3485 -43 3491 12
rect 3533 -43 3539 172
rect 3581 148 3587 532
rect 3597 308 3603 652
rect 3661 528 3667 752
rect 3693 728 3699 832
rect 3757 728 3763 832
rect 3773 788 3779 912
rect 3837 888 3843 972
rect 3885 908 3891 932
rect 3901 928 3907 1052
rect 3933 988 3939 1052
rect 3965 888 3971 992
rect 3885 837 3896 843
rect 3821 728 3827 832
rect 3773 708 3779 712
rect 3837 708 3843 732
rect 3885 723 3891 837
rect 3917 788 3923 872
rect 3965 748 3971 872
rect 3981 788 3987 872
rect 4029 828 4035 932
rect 4045 728 4051 1352
rect 4109 1328 4115 1472
rect 4141 1328 4147 1392
rect 4173 1348 4179 1432
rect 4173 1328 4179 1332
rect 4061 1308 4067 1312
rect 4157 1308 4163 1312
rect 4077 1268 4083 1292
rect 4109 1208 4115 1272
rect 4125 1108 4131 1232
rect 4157 1123 4163 1292
rect 4189 1148 4195 1272
rect 4157 1117 4168 1123
rect 4189 1068 4195 1092
rect 4157 968 4163 1032
rect 4077 948 4083 952
rect 4125 928 4131 932
rect 4173 928 4179 932
rect 4157 908 4163 912
rect 4125 868 4131 872
rect 4061 748 4067 752
rect 3885 717 3907 723
rect 3709 688 3715 692
rect 3677 588 3683 632
rect 3709 548 3715 552
rect 3613 388 3619 432
rect 3645 408 3651 512
rect 3661 508 3667 512
rect 3645 388 3651 392
rect 3677 388 3683 432
rect 3645 288 3651 312
rect 3693 288 3699 292
rect 3709 288 3715 412
rect 3725 308 3731 652
rect 3741 508 3747 512
rect 3821 308 3827 692
rect 3869 668 3875 672
rect 3837 588 3843 652
rect 3869 468 3875 512
rect 3885 508 3891 512
rect 3901 308 3907 717
rect 3997 708 4003 712
rect 4093 688 4099 792
rect 4157 748 4163 872
rect 4173 828 4179 832
rect 4189 828 4195 852
rect 4141 688 4147 692
rect 4045 528 4051 552
rect 4077 528 4083 612
rect 4157 588 4163 632
rect 4109 528 4115 572
rect 4173 563 4179 752
rect 4189 748 4195 812
rect 4205 728 4211 1552
rect 4221 1428 4227 1672
rect 4285 1648 4291 1792
rect 4301 1728 4307 1732
rect 4349 1728 4355 2052
rect 4365 1908 4371 2272
rect 4429 2148 4435 2512
rect 4493 2328 4499 2552
rect 4589 2548 4595 2672
rect 4621 2308 4627 2532
rect 4749 2528 4755 2532
rect 4525 2268 4531 2272
rect 4509 2203 4515 2232
rect 4509 2197 4531 2203
rect 4397 1728 4403 1912
rect 4477 1888 4483 2132
rect 4525 2108 4531 2197
rect 4573 2148 4579 2232
rect 4685 2188 4691 2192
rect 4733 2148 4739 2152
rect 4765 2148 4771 2672
rect 4781 2488 4787 2592
rect 4797 2528 4803 2752
rect 4829 2708 4835 2797
rect 4797 2508 4803 2512
rect 4781 2388 4787 2472
rect 4605 2108 4611 2112
rect 4557 1908 4563 1912
rect 4301 1637 4312 1643
rect 4301 1508 4307 1637
rect 4365 1468 4371 1472
rect 4237 1388 4243 1392
rect 4221 1368 4227 1372
rect 4253 1328 4259 1452
rect 4253 1188 4259 1312
rect 4301 1308 4307 1312
rect 4317 1308 4323 1352
rect 4349 1323 4355 1432
rect 4381 1408 4387 1712
rect 4413 1708 4419 1832
rect 4445 1768 4451 1872
rect 4477 1708 4483 1712
rect 4397 1488 4403 1512
rect 4413 1468 4419 1472
rect 4429 1328 4435 1332
rect 4349 1317 4360 1323
rect 4445 1308 4451 1632
rect 4461 1528 4467 1552
rect 4461 1368 4467 1512
rect 4493 1508 4499 1532
rect 4509 1308 4515 1612
rect 4525 1408 4531 1432
rect 4253 1148 4259 1152
rect 4317 1128 4323 1292
rect 4285 1028 4291 1092
rect 4301 1088 4307 1092
rect 4333 1088 4339 1232
rect 4349 1148 4355 1232
rect 4397 1188 4403 1272
rect 4333 1048 4339 1052
rect 4349 988 4355 1032
rect 4253 968 4259 972
rect 4269 928 4275 952
rect 4221 728 4227 912
rect 4269 908 4275 912
rect 4365 903 4371 1152
rect 4360 897 4371 903
rect 4381 1137 4392 1143
rect 4205 688 4211 692
rect 4237 683 4243 892
rect 4381 888 4387 1137
rect 4429 1128 4435 1292
rect 4445 1148 4451 1272
rect 4397 1068 4403 1072
rect 4413 968 4419 1092
rect 4429 988 4435 1092
rect 4493 1088 4499 1232
rect 4509 1168 4515 1292
rect 4541 1268 4547 1272
rect 4557 1068 4563 1732
rect 4605 1728 4611 2092
rect 4765 2048 4771 2112
rect 4781 1928 4787 2232
rect 4813 2168 4819 2532
rect 4829 2268 4835 2692
rect 4845 2688 4851 2732
rect 4845 2328 4851 2532
rect 4861 2303 4867 2972
rect 4877 2948 4883 2952
rect 5069 2928 5075 3072
rect 5117 2988 5123 3337
rect 5133 3188 5139 3292
rect 5165 3148 5171 3232
rect 4877 2528 4883 2712
rect 4877 2508 4883 2512
rect 4856 2297 4867 2303
rect 4845 2288 4851 2292
rect 4877 2288 4883 2292
rect 4797 2128 4803 2132
rect 4701 1888 4707 1912
rect 4733 1908 4739 1912
rect 4749 1888 4755 1892
rect 4781 1888 4787 1892
rect 4669 1768 4675 1872
rect 4765 1868 4771 1872
rect 4813 1808 4819 2152
rect 4829 2108 4835 2232
rect 4877 2128 4883 2272
rect 4845 2028 4851 2092
rect 4877 2088 4883 2112
rect 4893 2048 4899 2832
rect 4989 2808 4995 2832
rect 5133 2768 5139 3032
rect 5149 2968 5155 2972
rect 5197 2968 5203 3392
rect 5213 3348 5219 3492
rect 5229 3488 5235 3492
rect 5229 3328 5235 3472
rect 5293 3468 5299 3872
rect 5325 3728 5331 3732
rect 5309 3648 5315 3692
rect 5341 3688 5347 4532
rect 5389 4528 5395 4532
rect 5485 4508 5491 4532
rect 5501 4508 5507 4552
rect 5453 4488 5459 4492
rect 5453 4148 5459 4232
rect 5501 4188 5507 4312
rect 5517 4308 5523 4612
rect 5709 4588 5715 4712
rect 5725 4568 5731 4672
rect 5741 4648 5747 4692
rect 5773 4628 5779 4632
rect 5789 4588 5795 4712
rect 5853 4708 5859 4852
rect 5853 4628 5859 4692
rect 5869 4588 5875 4812
rect 5885 4708 5891 4872
rect 5549 4548 5555 4552
rect 5533 4528 5539 4532
rect 5613 4508 5619 4532
rect 5581 4428 5587 4492
rect 5613 4408 5619 4492
rect 5645 4448 5651 4512
rect 5645 4308 5651 4332
rect 5661 4308 5667 4312
rect 5389 4128 5395 4132
rect 5453 4128 5459 4132
rect 5373 3848 5379 4112
rect 5581 4108 5587 4212
rect 5597 4128 5603 4132
rect 5389 3748 5395 3972
rect 5421 3948 5427 4032
rect 5357 3648 5363 3712
rect 5309 3548 5315 3632
rect 5245 3388 5251 3452
rect 5325 3448 5331 3512
rect 5341 3508 5347 3512
rect 5373 3488 5379 3572
rect 5389 3548 5395 3732
rect 5405 3588 5411 3632
rect 5421 3508 5427 3832
rect 5517 3768 5523 3852
rect 5549 3788 5555 4092
rect 5661 3928 5667 4112
rect 5693 4028 5699 4532
rect 5725 4488 5731 4492
rect 5789 4428 5795 4492
rect 5821 4388 5827 4532
rect 5901 4528 5907 4917
rect 5933 4908 5939 4912
rect 5949 4728 5955 4912
rect 5981 4897 5992 4903
rect 5981 4788 5987 4897
rect 6093 4888 6099 5092
rect 6141 4943 6147 5232
rect 6317 5108 6323 5452
rect 6349 5348 6355 5432
rect 6365 5388 6371 5432
rect 6445 5388 6451 5492
rect 6573 5488 6579 5492
rect 6637 5488 6643 5512
rect 6941 5508 6947 5512
rect 6973 5508 6979 5512
rect 7149 5508 7155 5512
rect 6461 5468 6467 5472
rect 6557 5448 6563 5472
rect 6573 5368 6579 5452
rect 6333 5288 6339 5312
rect 6461 5308 6467 5312
rect 6573 5308 6579 5314
rect 6141 4937 6163 4943
rect 5917 4588 5923 4632
rect 5773 4308 5779 4332
rect 5837 4328 5843 4332
rect 5725 4168 5731 4292
rect 5805 4288 5811 4312
rect 5741 4128 5747 4272
rect 5629 3908 5635 3912
rect 5677 3863 5683 3892
rect 5693 3888 5699 4012
rect 5741 4008 5747 4112
rect 5741 3988 5747 3992
rect 5677 3857 5699 3863
rect 5517 3728 5523 3752
rect 5645 3748 5651 3752
rect 5501 3588 5507 3632
rect 5437 3468 5443 3472
rect 5293 3128 5299 3432
rect 5357 3348 5363 3452
rect 5453 3408 5459 3492
rect 5501 3408 5507 3432
rect 5405 3328 5411 3352
rect 5501 3328 5507 3332
rect 5325 3308 5331 3312
rect 5341 3188 5347 3212
rect 5437 3188 5443 3232
rect 5517 3148 5523 3712
rect 5693 3708 5699 3857
rect 5693 3688 5699 3692
rect 5693 3568 5699 3672
rect 5549 3488 5555 3492
rect 5581 3348 5587 3432
rect 5597 3348 5603 3532
rect 5725 3508 5731 3912
rect 5741 3688 5747 3712
rect 5757 3508 5763 4272
rect 5869 4228 5875 4432
rect 5885 4308 5891 4312
rect 5901 4288 5907 4512
rect 5917 4263 5923 4572
rect 5933 4508 5939 4512
rect 5901 4257 5923 4263
rect 5773 4128 5779 4172
rect 5837 3988 5843 4132
rect 5869 4128 5875 4132
rect 5885 4008 5891 4112
rect 5901 3988 5907 4257
rect 5917 4228 5923 4232
rect 5933 4168 5939 4292
rect 5949 4288 5955 4712
rect 6013 4708 6019 4792
rect 6045 4728 6051 4832
rect 6093 4808 6099 4872
rect 6157 4788 6163 4937
rect 6013 4628 6019 4692
rect 5965 4588 5971 4612
rect 5997 4568 6003 4592
rect 5997 4548 6003 4552
rect 6029 4528 6035 4692
rect 6045 4688 6051 4712
rect 6077 4708 6083 4712
rect 6125 4628 6131 4692
rect 6157 4688 6163 4772
rect 6173 4748 6179 5072
rect 6189 4968 6195 5072
rect 6301 4988 6307 5092
rect 6349 5048 6355 5052
rect 6397 5043 6403 5292
rect 6461 5108 6467 5292
rect 6397 5037 6419 5043
rect 6349 4948 6355 5032
rect 6413 4988 6419 5037
rect 6493 4988 6499 5092
rect 6557 4948 6563 5052
rect 6605 4948 6611 5072
rect 6621 4988 6627 5092
rect 6445 4928 6451 4932
rect 6557 4928 6563 4932
rect 6269 4908 6275 4912
rect 6173 4708 6179 4712
rect 6072 4557 6099 4563
rect 6093 4548 6099 4557
rect 6141 4548 6147 4672
rect 6173 4608 6179 4692
rect 6189 4568 6195 4832
rect 6461 4828 6467 4912
rect 6589 4908 6595 4912
rect 6525 4828 6531 4892
rect 6637 4828 6643 5472
rect 6717 5468 6723 5472
rect 6813 5468 6819 5472
rect 6813 5343 6819 5452
rect 6797 5337 6819 5343
rect 6797 5328 6803 5337
rect 6861 5328 6867 5332
rect 6909 5328 6915 5472
rect 7005 5448 7011 5472
rect 6941 5348 6947 5432
rect 6685 5108 6691 5112
rect 6733 4928 6739 5032
rect 6781 4948 6787 5232
rect 6813 5068 6819 5092
rect 6813 4988 6819 5032
rect 6669 4888 6675 4912
rect 6205 4748 6211 4752
rect 6205 4708 6211 4732
rect 6237 4648 6243 4692
rect 6269 4668 6275 4732
rect 6285 4668 6291 4752
rect 6349 4728 6355 4732
rect 6237 4588 6243 4592
rect 6029 4508 6035 4512
rect 6093 4508 6099 4512
rect 6125 4508 6131 4512
rect 5965 4308 5971 4432
rect 5981 4288 5987 4292
rect 5965 4268 5971 4272
rect 5949 4148 5955 4152
rect 5965 4148 5971 4252
rect 6029 4188 6035 4292
rect 6077 4288 6083 4312
rect 6109 4308 6115 4432
rect 6141 4368 6147 4532
rect 6077 4128 6083 4152
rect 6109 4128 6115 4272
rect 5981 4008 5987 4092
rect 5613 3348 5619 3492
rect 5629 3488 5635 3492
rect 5725 3488 5731 3492
rect 5629 3468 5635 3472
rect 5645 3388 5651 3432
rect 5581 3308 5587 3312
rect 5325 3108 5331 3112
rect 5213 3088 5219 3092
rect 5149 2948 5155 2952
rect 5261 2928 5267 2992
rect 5293 2963 5299 3052
rect 5288 2957 5299 2963
rect 5309 2948 5315 3072
rect 5325 2928 5331 2992
rect 5357 2988 5363 3072
rect 5373 3068 5379 3132
rect 5373 2968 5379 3052
rect 5405 3028 5411 3092
rect 5405 2928 5411 3012
rect 5421 2928 5427 3072
rect 5469 2948 5475 3032
rect 5517 2988 5523 2992
rect 5565 2948 5571 3112
rect 5581 3008 5587 3092
rect 5613 2948 5619 3312
rect 5469 2888 5475 2912
rect 5549 2908 5555 2912
rect 4941 2708 4947 2712
rect 4957 2688 4963 2692
rect 5000 2677 5011 2683
rect 5005 2588 5011 2677
rect 4973 2468 4979 2512
rect 4989 2308 4995 2492
rect 5005 2288 5011 2432
rect 5069 2288 5075 2672
rect 5085 2508 5091 2512
rect 5085 2488 5091 2492
rect 5197 2463 5203 2832
rect 5453 2688 5459 2692
rect 5421 2668 5427 2672
rect 5245 2543 5251 2652
rect 5245 2537 5267 2543
rect 5261 2528 5267 2537
rect 5197 2457 5219 2463
rect 5197 2428 5203 2432
rect 4941 2128 4947 2252
rect 5069 2128 5075 2172
rect 5101 2148 5107 2232
rect 4877 1908 4883 1972
rect 4621 1708 4627 1712
rect 4605 1528 4611 1532
rect 4637 1508 4643 1732
rect 4781 1648 4787 1792
rect 4909 1768 4915 1872
rect 4909 1728 4915 1732
rect 4765 1508 4771 1512
rect 4781 1483 4787 1632
rect 4776 1477 4787 1483
rect 4589 1288 4595 1412
rect 4605 1308 4611 1312
rect 4621 1308 4627 1352
rect 4669 1328 4675 1392
rect 4685 1348 4691 1472
rect 4797 1468 4803 1472
rect 4765 1348 4771 1352
rect 4861 1348 4867 1672
rect 4877 1568 4883 1632
rect 4925 1588 4931 1732
rect 4941 1728 4947 2072
rect 4957 1748 4963 2112
rect 4989 1968 4995 2032
rect 5101 1908 5107 1932
rect 5117 1888 5123 2272
rect 5133 2128 5139 2292
rect 5181 2188 5187 2232
rect 5181 2148 5187 2152
rect 4989 1848 4995 1872
rect 4877 1488 4883 1532
rect 4621 1203 4627 1292
rect 4637 1288 4643 1292
rect 4605 1197 4627 1203
rect 4605 1128 4611 1197
rect 4637 1148 4643 1252
rect 4669 1148 4675 1232
rect 4557 988 4563 1052
rect 4605 988 4611 1072
rect 4269 837 4280 843
rect 4269 808 4275 837
rect 4349 808 4355 832
rect 4365 828 4371 872
rect 4397 868 4403 912
rect 4285 688 4291 792
rect 4317 708 4323 772
rect 4461 748 4467 872
rect 4525 868 4531 912
rect 4477 708 4483 832
rect 4221 677 4243 683
rect 4157 557 4179 563
rect 4157 528 4163 557
rect 3965 308 3971 312
rect 3720 277 3731 283
rect 3565 128 3571 132
rect 3629 128 3635 232
rect 3725 188 3731 277
rect 3725 148 3731 172
rect 3757 128 3763 232
rect 3789 123 3795 232
rect 3853 188 3859 272
rect 3949 168 3955 232
rect 3965 128 3971 232
rect 3981 188 3987 452
rect 4205 448 4211 672
rect 4221 528 4227 677
rect 4333 608 4339 692
rect 4269 528 4275 572
rect 4285 548 4291 552
rect 4317 508 4323 512
rect 3997 308 4003 312
rect 4013 288 4019 392
rect 4061 308 4067 432
rect 4125 308 4131 432
rect 4237 308 4243 432
rect 4253 288 4259 352
rect 3981 148 3987 172
rect 4125 148 4131 232
rect 4189 168 4195 232
rect 4205 208 4211 232
rect 4173 128 4179 152
rect 4221 128 4227 132
rect 4269 128 4275 152
rect 4285 128 4291 492
rect 4333 328 4339 452
rect 4381 368 4387 532
rect 4397 488 4403 652
rect 4429 608 4435 672
rect 4333 308 4339 312
rect 4381 288 4387 312
rect 4397 308 4403 312
rect 4429 308 4435 592
rect 4493 528 4499 532
rect 3789 117 3800 123
rect 3581 -43 3587 32
rect 3661 -43 3667 32
rect 3709 -43 3715 112
rect 4125 108 4131 112
rect 4301 108 4307 232
rect 4365 168 4371 272
rect 4333 123 4339 132
rect 4397 128 4403 192
rect 4445 188 4451 272
rect 4509 188 4515 532
rect 4525 288 4531 312
rect 4525 268 4531 272
rect 4541 208 4547 632
rect 4573 408 4579 932
rect 4621 708 4627 1092
rect 4637 828 4643 1132
rect 4669 968 4675 1032
rect 4685 928 4691 1332
rect 4797 1308 4803 1312
rect 4829 1188 4835 1272
rect 4717 1088 4723 1132
rect 4733 1128 4739 1152
rect 4797 1108 4803 1112
rect 4765 988 4771 1092
rect 4797 1088 4803 1092
rect 4669 648 4675 692
rect 4685 688 4691 912
rect 4797 728 4803 872
rect 4824 717 4835 723
rect 4765 688 4771 712
rect 4797 663 4803 712
rect 4829 668 4835 717
rect 4845 708 4851 1072
rect 4861 1068 4867 1332
rect 4877 1088 4883 1092
rect 4861 928 4867 932
rect 4893 928 4899 1512
rect 4957 1488 4963 1712
rect 4989 1708 4995 1832
rect 4973 1588 4979 1692
rect 4957 1408 4963 1472
rect 4957 1328 4963 1332
rect 4973 1308 4979 1312
rect 4909 888 4915 1112
rect 4957 1108 4963 1112
rect 4989 1088 4995 1392
rect 4973 1068 4979 1072
rect 4925 928 4931 1032
rect 4989 928 4995 1072
rect 4925 748 4931 832
rect 5005 728 5011 1752
rect 5037 1728 5043 1732
rect 5149 1688 5155 1732
rect 5165 1688 5171 1712
rect 5085 1528 5091 1532
rect 5101 1128 5107 1412
rect 5117 1348 5123 1492
rect 5133 1123 5139 1552
rect 5165 1508 5171 1672
rect 5181 1506 5187 1552
rect 5213 1528 5219 2457
rect 5229 2388 5235 2512
rect 5245 2508 5251 2512
rect 5245 2308 5251 2492
rect 5293 2208 5299 2432
rect 5341 2288 5347 2652
rect 5389 2588 5395 2632
rect 5501 2608 5507 2892
rect 5645 2788 5651 2914
rect 5549 2708 5555 2712
rect 5565 2708 5571 2772
rect 5645 2688 5651 2752
rect 5677 2728 5683 3472
rect 5693 3308 5699 3332
rect 5725 3308 5731 3392
rect 5757 3328 5763 3492
rect 5773 3448 5779 3732
rect 5805 3668 5811 3892
rect 5869 3888 5875 3932
rect 5949 3908 5955 3912
rect 5885 3828 5891 3892
rect 5997 3868 6003 3932
rect 5885 3728 5891 3772
rect 5885 3488 5891 3492
rect 5773 3328 5779 3392
rect 5789 3348 5795 3432
rect 5772 3297 5779 3303
rect 5693 3188 5699 3292
rect 5773 3108 5779 3297
rect 5741 2768 5747 2892
rect 5773 2843 5779 3032
rect 5789 2988 5795 3312
rect 5805 3268 5811 3332
rect 5869 3308 5875 3392
rect 5933 3388 5939 3512
rect 5981 3488 5987 3732
rect 5981 3448 5987 3472
rect 5949 3308 5955 3332
rect 5805 3128 5811 3252
rect 5981 3248 5987 3332
rect 6013 3108 6019 4112
rect 6157 4063 6163 4512
rect 6189 4508 6195 4552
rect 6317 4528 6323 4692
rect 6333 4588 6339 4712
rect 6381 4663 6387 4772
rect 6413 4717 6451 4723
rect 6413 4703 6419 4717
rect 6445 4708 6451 4717
rect 6408 4697 6419 4703
rect 6504 4697 6536 4703
rect 6477 4683 6483 4692
rect 6408 4677 6419 4683
rect 6477 4677 6552 4683
rect 6381 4657 6392 4663
rect 6413 4608 6419 4677
rect 6445 4648 6451 4652
rect 6477 4588 6483 4592
rect 6541 4548 6547 4632
rect 6573 4608 6579 4712
rect 6605 4688 6611 4692
rect 6621 4668 6627 4672
rect 6141 4057 6163 4063
rect 6141 3988 6147 4057
rect 6173 4008 6179 4252
rect 6205 4048 6211 4112
rect 6237 4108 6243 4252
rect 6253 4068 6259 4512
rect 6349 4428 6355 4492
rect 6301 4128 6307 4252
rect 6349 4188 6355 4412
rect 6413 4368 6419 4532
rect 6637 4528 6643 4692
rect 6669 4688 6675 4752
rect 6669 4668 6675 4672
rect 6445 4488 6451 4492
rect 6445 4328 6451 4472
rect 6525 4468 6531 4512
rect 6669 4348 6675 4432
rect 6685 4388 6691 4892
rect 6829 4888 6835 5312
rect 6957 5308 6963 5312
rect 6845 5088 6851 5092
rect 6701 4768 6707 4832
rect 6861 4808 6867 4912
rect 6701 4708 6707 4712
rect 6733 4708 6739 4732
rect 6877 4708 6883 5232
rect 6893 4988 6899 5012
rect 6941 4988 6947 5112
rect 6973 5068 6979 5092
rect 6989 5088 6995 5432
rect 7005 5328 7011 5332
rect 6909 4708 6915 4712
rect 6749 4668 6755 4672
rect 6797 4668 6803 4692
rect 6813 4688 6819 4692
rect 6877 4688 6883 4692
rect 6925 4688 6931 4932
rect 7005 4928 7011 5172
rect 7021 5048 7027 5492
rect 7229 5148 7235 5472
rect 7261 5348 7267 5472
rect 7341 5388 7347 5492
rect 7405 5388 7411 5392
rect 7261 5283 7267 5332
rect 7261 5277 7283 5283
rect 7213 5088 7219 5132
rect 7117 4948 7123 5052
rect 7261 5048 7267 5092
rect 7277 4968 7283 5277
rect 7293 5268 7299 5332
rect 7309 5308 7315 5312
rect 7293 5088 7299 5252
rect 7128 4937 7139 4943
rect 7133 4928 7139 4937
rect 7293 4928 7299 5032
rect 6941 4728 6947 4732
rect 7005 4708 7011 4892
rect 7117 4888 7123 4912
rect 7037 4728 7043 4832
rect 6941 4688 6947 4692
rect 6845 4668 6851 4672
rect 6861 4668 6867 4672
rect 6733 4568 6739 4632
rect 6781 4588 6787 4632
rect 6829 4528 6835 4552
rect 6893 4528 6899 4632
rect 6973 4588 6979 4652
rect 6973 4528 6979 4552
rect 6989 4548 6995 4672
rect 7005 4648 7011 4692
rect 6989 4528 6995 4532
rect 6413 4308 6419 4312
rect 6381 4168 6387 4272
rect 6141 3908 6147 3972
rect 6173 3908 6179 3912
rect 6045 3868 6051 3872
rect 6205 3743 6211 4032
rect 6253 3908 6259 4032
rect 6397 3928 6403 4172
rect 6429 4128 6435 4232
rect 6285 3908 6291 3912
rect 6205 3737 6227 3743
rect 6109 3728 6115 3732
rect 6221 3728 6227 3737
rect 6045 3708 6051 3712
rect 6045 3463 6051 3692
rect 6205 3528 6211 3712
rect 6093 3508 6099 3512
rect 6125 3488 6131 3512
rect 6221 3508 6227 3712
rect 6237 3708 6243 3712
rect 6029 3457 6051 3463
rect 5837 2948 5843 2972
rect 5869 2968 5875 2972
rect 5805 2888 5811 2892
rect 5885 2848 5891 3032
rect 5933 2988 5939 2992
rect 5949 2928 5955 3072
rect 5981 3068 5987 3072
rect 5981 2968 5987 3052
rect 5933 2908 5939 2912
rect 5773 2837 5795 2843
rect 5357 2488 5363 2512
rect 5421 2288 5427 2512
rect 5485 2328 5491 2332
rect 5469 2288 5475 2292
rect 5389 2268 5395 2272
rect 5501 2268 5507 2532
rect 5517 2503 5523 2672
rect 5533 2648 5539 2672
rect 5517 2497 5539 2503
rect 5517 2308 5523 2312
rect 5533 2288 5539 2497
rect 5549 2308 5555 2472
rect 5597 2388 5603 2572
rect 5629 2548 5635 2632
rect 5709 2628 5715 2632
rect 5725 2563 5731 2712
rect 5709 2557 5731 2563
rect 5645 2488 5651 2512
rect 5693 2488 5699 2492
rect 5709 2328 5715 2557
rect 5741 2528 5747 2752
rect 5773 2708 5779 2732
rect 5789 2708 5795 2837
rect 5821 2828 5827 2832
rect 5757 2668 5763 2672
rect 5725 2508 5731 2512
rect 5645 2308 5651 2312
rect 5309 2148 5315 2152
rect 5501 2148 5507 2252
rect 5533 2248 5539 2272
rect 5389 2108 5395 2112
rect 5229 1928 5235 1952
rect 5261 1908 5267 1932
rect 5277 1908 5283 1952
rect 5325 1908 5331 1932
rect 5229 1688 5235 1692
rect 5245 1488 5251 1632
rect 5277 1528 5283 1552
rect 5149 1143 5155 1232
rect 5149 1137 5171 1143
rect 5133 1117 5144 1123
rect 5101 1108 5107 1112
rect 5117 1088 5123 1092
rect 5085 788 5091 952
rect 5117 908 5123 1072
rect 5149 928 5155 932
rect 4941 708 4947 712
rect 4797 657 4819 663
rect 4653 588 4659 632
rect 4717 548 4723 592
rect 4781 588 4787 632
rect 4765 568 4771 572
rect 4621 428 4627 512
rect 4797 503 4803 632
rect 4813 528 4819 657
rect 4845 608 4851 692
rect 4909 608 4915 652
rect 4925 568 4931 672
rect 4829 548 4835 552
rect 4792 497 4803 503
rect 4557 288 4563 312
rect 4573 288 4579 352
rect 4685 348 4691 492
rect 4685 328 4691 332
rect 4813 328 4819 512
rect 4589 288 4595 292
rect 4861 288 4867 332
rect 4909 288 4915 292
rect 4813 268 4819 272
rect 4925 268 4931 512
rect 4941 468 4947 692
rect 5021 548 5027 632
rect 5101 548 5107 572
rect 4973 528 4979 532
rect 4941 308 4947 312
rect 5069 288 5075 532
rect 5005 268 5011 272
rect 4525 148 4531 172
rect 4333 117 4344 123
rect 4733 128 4739 192
rect 4749 188 4755 252
rect 4845 128 4851 232
rect 4925 148 4931 252
rect 4973 128 4979 212
rect 5005 188 5011 252
rect 5069 148 5075 272
rect 5085 188 5091 472
rect 5117 308 5123 332
rect 5165 328 5171 1137
rect 5197 1108 5203 1112
rect 5229 1088 5235 1292
rect 5293 1188 5299 1892
rect 5389 1888 5395 2092
rect 5405 1908 5411 1912
rect 5437 1888 5443 1892
rect 5533 1888 5539 2132
rect 5309 1868 5315 1872
rect 5373 1728 5379 1732
rect 5357 1703 5363 1712
rect 5357 1697 5379 1703
rect 5325 1488 5331 1532
rect 5357 1508 5363 1512
rect 5357 1488 5363 1492
rect 5213 988 5219 1052
rect 5181 928 5187 932
rect 5181 728 5187 912
rect 5181 688 5187 692
rect 5213 688 5219 832
rect 5229 568 5235 1072
rect 5309 1068 5315 1092
rect 5325 1088 5331 1092
rect 5373 1088 5379 1697
rect 5389 1548 5395 1872
rect 5549 1868 5555 2192
rect 5597 2148 5603 2232
rect 5629 1908 5635 2172
rect 5677 2148 5683 2232
rect 5693 2128 5699 2192
rect 5533 1857 5544 1863
rect 5485 1768 5491 1812
rect 5533 1748 5539 1857
rect 5613 1768 5619 1852
rect 5581 1728 5587 1752
rect 5661 1748 5667 2032
rect 5501 1668 5507 1692
rect 5549 1628 5555 1712
rect 5437 1508 5443 1512
rect 5405 1308 5411 1332
rect 5421 1328 5427 1492
rect 5549 1488 5555 1612
rect 5597 1608 5603 1732
rect 5693 1728 5699 1732
rect 5677 1668 5683 1712
rect 5725 1668 5731 2492
rect 5741 2288 5747 2312
rect 5757 2168 5763 2272
rect 5789 2188 5795 2692
rect 5821 2668 5827 2672
rect 5853 2668 5859 2692
rect 5885 2668 5891 2692
rect 5901 2688 5907 2892
rect 5949 2888 5955 2892
rect 5821 2548 5827 2652
rect 5901 2643 5907 2672
rect 5949 2668 5955 2672
rect 5901 2637 5923 2643
rect 5885 2628 5891 2632
rect 5837 2528 5843 2532
rect 5853 2528 5859 2612
rect 5837 2188 5843 2472
rect 5853 2068 5859 2432
rect 5917 2408 5923 2637
rect 5869 2128 5875 2332
rect 5885 2308 5891 2372
rect 5901 2128 5907 2212
rect 5933 2208 5939 2432
rect 5965 2348 5971 2832
rect 6013 2828 6019 3092
rect 6029 2983 6035 3457
rect 6205 3428 6211 3492
rect 6237 3468 6243 3492
rect 6125 3328 6131 3332
rect 6045 3128 6051 3132
rect 6077 3088 6083 3272
rect 6093 3188 6099 3232
rect 6141 3128 6147 3132
rect 6189 3128 6195 3132
rect 6029 2977 6040 2983
rect 5997 2708 6003 2752
rect 6045 2728 6051 2832
rect 6093 2788 6099 3032
rect 6141 2988 6147 3092
rect 6205 2928 6211 3012
rect 6237 3008 6243 3112
rect 6237 2968 6243 2992
rect 6173 2888 6179 2892
rect 6253 2808 6259 3872
rect 6269 3808 6275 3872
rect 6317 3848 6323 3872
rect 6349 3868 6355 3872
rect 6317 3828 6323 3832
rect 6269 3768 6275 3772
rect 6344 3757 6376 3763
rect 6269 3748 6275 3752
rect 6333 3708 6339 3712
rect 6397 3608 6403 3912
rect 6413 3728 6419 3972
rect 6445 3948 6451 4312
rect 6669 4308 6675 4332
rect 6781 4328 6787 4332
rect 6829 4308 6835 4332
rect 6477 4268 6483 4272
rect 6477 4248 6483 4252
rect 6509 4168 6515 4292
rect 6557 4288 6563 4292
rect 6717 4228 6723 4292
rect 6589 4128 6595 4152
rect 6733 4128 6739 4272
rect 6845 4268 6851 4272
rect 6525 4048 6531 4112
rect 6557 3948 6563 4032
rect 6461 3848 6467 3912
rect 6525 3908 6531 3932
rect 6509 3828 6515 3872
rect 6456 3757 6467 3763
rect 6461 3748 6467 3757
rect 6525 3748 6531 3752
rect 6541 3748 6547 3772
rect 6573 3768 6579 3832
rect 6589 3748 6595 3792
rect 6509 3728 6515 3732
rect 6605 3728 6611 3932
rect 6669 3788 6675 3912
rect 6701 3728 6707 3732
rect 6477 3668 6483 3712
rect 6509 3588 6515 3712
rect 6733 3708 6739 3832
rect 6749 3748 6755 4132
rect 6797 4128 6803 4232
rect 6861 4188 6867 4472
rect 6893 4388 6899 4492
rect 6909 4468 6915 4512
rect 7021 4508 7027 4512
rect 6941 4348 6947 4492
rect 7005 4328 7011 4492
rect 6941 4188 6947 4272
rect 6973 4208 6979 4312
rect 6989 4188 6995 4312
rect 7021 4303 7027 4312
rect 7037 4308 7043 4672
rect 7069 4588 7075 4712
rect 7117 4688 7123 4692
rect 7133 4608 7139 4672
rect 7149 4568 7155 4832
rect 7181 4748 7187 4912
rect 7197 4528 7203 4872
rect 7213 4548 7219 4552
rect 7309 4548 7315 5132
rect 7325 5048 7331 5112
rect 7357 5028 7363 5332
rect 7373 5128 7379 5312
rect 7421 5308 7427 5312
rect 7389 5188 7395 5292
rect 7437 5088 7443 5472
rect 7469 5348 7475 5432
rect 7565 5408 7571 5492
rect 7453 5108 7459 5332
rect 7501 5328 7507 5372
rect 7597 5348 7603 5372
rect 7549 5328 7555 5332
rect 7485 5268 7491 5312
rect 7517 5108 7523 5252
rect 7501 5088 7507 5092
rect 7373 4968 7379 5072
rect 7373 4948 7379 4952
rect 7437 4928 7443 5072
rect 7341 4688 7347 4912
rect 7453 4748 7459 5072
rect 7501 4928 7507 4932
rect 7517 4928 7523 5092
rect 7517 4888 7523 4912
rect 7533 4908 7539 5232
rect 7613 5148 7619 5452
rect 7645 5423 7651 5512
rect 7693 5468 7699 5492
rect 7725 5488 7731 5512
rect 7725 5428 7731 5432
rect 7629 5417 7651 5423
rect 7629 5388 7635 5417
rect 7645 5348 7651 5392
rect 7645 5303 7651 5332
rect 7757 5328 7763 5332
rect 7709 5308 7715 5312
rect 7773 5308 7779 5492
rect 7789 5408 7795 5472
rect 7645 5297 7667 5303
rect 7549 5048 7555 5112
rect 7629 5083 7635 5292
rect 7613 5077 7635 5083
rect 7613 5068 7619 5077
rect 7517 4708 7523 4872
rect 7533 4728 7539 4752
rect 7016 4297 7027 4303
rect 6957 4148 6963 4152
rect 7005 4148 7011 4272
rect 7037 4268 7043 4272
rect 6845 4048 6851 4132
rect 6797 3908 6803 4012
rect 6765 3748 6771 3752
rect 6781 3748 6787 3812
rect 6829 3788 6835 3992
rect 6877 3928 6883 4092
rect 6893 4088 6899 4092
rect 6909 3928 6915 4052
rect 6925 3988 6931 4072
rect 6941 4068 6947 4112
rect 6989 4068 6995 4092
rect 6845 3748 6851 3792
rect 6765 3728 6771 3732
rect 6669 3608 6675 3692
rect 6733 3628 6739 3692
rect 6797 3688 6803 3712
rect 6669 3528 6675 3552
rect 6605 3508 6611 3512
rect 6504 3497 6515 3503
rect 6317 3468 6323 3492
rect 6317 3328 6323 3452
rect 6333 3328 6339 3372
rect 6349 3368 6355 3432
rect 6365 3388 6371 3432
rect 6381 3328 6387 3492
rect 6413 3308 6419 3312
rect 6413 3148 6419 3292
rect 6429 3188 6435 3372
rect 6509 3348 6515 3497
rect 6573 3488 6579 3492
rect 6573 3468 6579 3472
rect 6605 3388 6611 3492
rect 6669 3488 6675 3512
rect 6637 3448 6643 3472
rect 6797 3468 6803 3492
rect 6749 3388 6755 3452
rect 6813 3368 6819 3732
rect 6829 3668 6835 3692
rect 6845 3548 6851 3692
rect 6861 3688 6867 3712
rect 6877 3548 6883 3892
rect 6893 3868 6899 3872
rect 6909 3808 6915 3912
rect 6941 3728 6947 4032
rect 7021 3906 7027 4092
rect 6957 3848 6963 3872
rect 6920 3697 6931 3703
rect 6605 3328 6611 3352
rect 6621 3328 6627 3332
rect 6813 3328 6819 3352
rect 6845 3328 6851 3432
rect 6669 3188 6675 3192
rect 6733 3188 6739 3192
rect 6269 3068 6275 3072
rect 6285 3028 6291 3032
rect 6301 2948 6307 2972
rect 6029 2508 6035 2692
rect 6045 2688 6051 2692
rect 6093 2608 6099 2672
rect 6109 2668 6115 2672
rect 6125 2668 6131 2692
rect 6173 2688 6179 2792
rect 6301 2768 6307 2872
rect 6205 2708 6211 2732
rect 6093 2588 6099 2592
rect 6141 2568 6147 2672
rect 6141 2388 6147 2472
rect 6173 2368 6179 2672
rect 6189 2668 6195 2692
rect 6221 2628 6227 2712
rect 6253 2688 6259 2712
rect 6301 2688 6307 2752
rect 6285 2628 6291 2672
rect 6221 2528 6227 2552
rect 6301 2548 6307 2592
rect 6317 2528 6323 2892
rect 6317 2508 6323 2512
rect 6349 2508 6355 3132
rect 6461 3108 6467 3132
rect 6509 3088 6515 3112
rect 6637 3108 6643 3132
rect 6797 3128 6803 3132
rect 6653 3108 6659 3112
rect 6701 3088 6707 3092
rect 6381 3068 6387 3072
rect 6365 2708 6371 2732
rect 6397 2728 6403 3072
rect 6477 3068 6483 3072
rect 6525 2968 6531 3052
rect 6557 3048 6563 3052
rect 6541 2948 6547 2992
rect 6557 2968 6563 3032
rect 6413 2748 6419 2912
rect 6461 2808 6467 2932
rect 6621 2928 6627 3076
rect 6669 3028 6675 3032
rect 6653 2988 6659 2992
rect 6637 2948 6643 2952
rect 6685 2948 6691 3072
rect 6749 2988 6755 3112
rect 6877 3088 6883 3532
rect 6893 3448 6899 3692
rect 6925 3588 6931 3697
rect 6909 3548 6915 3572
rect 6941 3508 6947 3712
rect 6957 3528 6963 3712
rect 6957 3508 6963 3512
rect 6941 3488 6947 3492
rect 6957 3468 6963 3472
rect 6925 3188 6931 3232
rect 6893 3108 6899 3172
rect 6957 3148 6963 3272
rect 6957 3128 6963 3132
rect 6813 3008 6819 3032
rect 6797 2983 6803 2992
rect 6797 2977 6819 2983
rect 6493 2728 6499 2892
rect 6701 2888 6707 2932
rect 6813 2928 6819 2977
rect 6925 2928 6931 3032
rect 6941 2928 6947 3012
rect 6973 2988 6979 3792
rect 6989 3748 6995 3872
rect 6989 3468 6995 3472
rect 6989 3388 6995 3432
rect 7005 3308 7011 3612
rect 7037 3608 7043 4192
rect 7053 4168 7059 4232
rect 7117 4208 7123 4492
rect 7165 4488 7171 4492
rect 7181 4308 7187 4312
rect 7197 4308 7203 4512
rect 7117 4108 7123 4112
rect 7117 3908 7123 4092
rect 7197 3888 7203 4252
rect 7229 4168 7235 4252
rect 7293 4228 7299 4292
rect 7293 4148 7299 4152
rect 7293 3948 7299 4112
rect 7277 3908 7283 3912
rect 7133 3708 7139 3712
rect 7021 3528 7027 3572
rect 7037 3308 7043 3592
rect 7069 3488 7075 3512
rect 7069 3368 7075 3472
rect 7101 3388 7107 3652
rect 7117 3508 7123 3532
rect 7133 3388 7139 3692
rect 7149 3508 7155 3832
rect 7181 3708 7187 3712
rect 7197 3688 7203 3872
rect 7261 3728 7267 3732
rect 7277 3728 7283 3892
rect 7293 3708 7299 3712
rect 7165 3588 7171 3672
rect 7197 3568 7203 3672
rect 7213 3508 7219 3632
rect 7261 3528 7267 3572
rect 7197 3368 7203 3492
rect 7213 3477 7224 3483
rect 7165 3348 7171 3352
rect 7197 3308 7203 3312
rect 6989 3188 6995 3292
rect 7005 3288 7011 3292
rect 7005 2948 7011 2992
rect 7021 2988 7027 3072
rect 7037 3068 7043 3072
rect 6717 2908 6723 2912
rect 6701 2748 6707 2792
rect 6397 2708 6403 2712
rect 6429 2708 6435 2712
rect 6573 2688 6579 2692
rect 6397 2588 6403 2672
rect 6413 2648 6419 2672
rect 6413 2548 6419 2632
rect 6429 2548 6435 2612
rect 6461 2588 6467 2592
rect 6349 2488 6355 2492
rect 5933 2123 5939 2192
rect 5965 2148 5971 2272
rect 6029 2268 6035 2272
rect 6077 2248 6083 2292
rect 6205 2288 6211 2392
rect 6429 2388 6435 2472
rect 6248 2317 6275 2323
rect 6269 2308 6275 2317
rect 6317 2308 6323 2312
rect 6013 2188 6019 2232
rect 6157 2148 6163 2252
rect 5933 2117 5944 2123
rect 5837 1908 5843 2032
rect 5869 1988 5875 2112
rect 5949 2108 5955 2112
rect 5933 1968 5939 2032
rect 5965 1948 5971 2132
rect 6157 2128 6163 2132
rect 5869 1906 5875 1932
rect 5949 1928 5955 1932
rect 5757 1728 5763 1752
rect 5773 1748 5779 1852
rect 5821 1788 5827 1872
rect 5805 1728 5811 1732
rect 5837 1703 5843 1892
rect 5933 1888 5939 1912
rect 5997 1888 6003 1932
rect 6093 1908 6099 1912
rect 5901 1848 5907 1872
rect 5949 1868 5955 1872
rect 5832 1697 5843 1703
rect 5597 1588 5603 1592
rect 5581 1508 5587 1512
rect 5645 1368 5651 1432
rect 5693 1348 5699 1652
rect 5709 1528 5715 1532
rect 5757 1508 5763 1532
rect 5805 1368 5811 1472
rect 5421 1308 5427 1312
rect 5629 1308 5635 1332
rect 5693 1328 5699 1332
rect 5533 1288 5539 1292
rect 5277 928 5283 932
rect 5309 688 5315 712
rect 5357 688 5363 932
rect 5325 548 5331 552
rect 5357 548 5363 672
rect 5373 548 5379 692
rect 5181 508 5187 512
rect 5213 288 5219 532
rect 5229 488 5235 532
rect 5229 308 5235 312
rect 5245 308 5251 332
rect 5213 268 5219 272
rect 5277 128 5283 532
rect 5309 508 5315 512
rect 5341 508 5347 532
rect 5373 388 5379 492
rect 5405 328 5411 1112
rect 5453 903 5459 1072
rect 5469 988 5475 1272
rect 5485 1128 5491 1172
rect 5533 1108 5539 1172
rect 5821 1128 5827 1532
rect 5853 1488 5859 1672
rect 5885 1548 5891 1632
rect 5885 1508 5891 1512
rect 5901 1508 5907 1712
rect 5917 1668 5923 1712
rect 5933 1488 5939 1592
rect 5853 1388 5859 1472
rect 5869 1388 5875 1472
rect 5885 1308 5891 1312
rect 5901 1268 5907 1472
rect 5821 1108 5827 1112
rect 5485 968 5491 1032
rect 5448 897 5459 903
rect 5421 708 5427 712
rect 5453 688 5459 712
rect 5469 688 5475 892
rect 5485 728 5491 732
rect 5533 708 5539 732
rect 5565 688 5571 1072
rect 5645 1068 5651 1092
rect 5885 1088 5891 1152
rect 5917 1108 5923 1312
rect 5613 928 5619 992
rect 5741 988 5747 1072
rect 5629 968 5635 972
rect 5693 848 5699 912
rect 5773 888 5779 1072
rect 5789 1048 5795 1072
rect 5837 1008 5843 1032
rect 5837 928 5843 932
rect 5565 568 5571 672
rect 5565 548 5571 552
rect 5469 388 5475 512
rect 5501 428 5507 492
rect 5484 317 5507 323
rect 5405 308 5411 312
rect 5501 308 5507 317
rect 5325 288 5331 292
rect 5405 288 5411 292
rect 5501 268 5507 272
rect 5517 268 5523 312
rect 5533 308 5539 432
rect 5549 308 5555 532
rect 5389 128 5395 152
rect 5485 148 5491 252
rect 5565 148 5571 412
rect 5597 128 5603 732
rect 5661 688 5667 692
rect 5645 588 5651 592
rect 5645 548 5651 572
rect 5693 568 5699 832
rect 5789 708 5795 912
rect 5917 868 5923 1092
rect 5933 948 5939 1472
rect 5949 1468 5955 1852
rect 6093 1828 6099 1892
rect 5981 1748 5987 1752
rect 6109 1748 6115 1832
rect 5949 1388 5955 1452
rect 5965 1363 5971 1692
rect 6013 1508 6019 1712
rect 6141 1668 6147 2112
rect 6157 1988 6163 2092
rect 6189 1968 6195 2192
rect 6205 2023 6211 2272
rect 6221 2148 6227 2292
rect 6253 2288 6259 2292
rect 6333 2268 6339 2332
rect 6429 2308 6435 2372
rect 6413 2288 6419 2292
rect 6397 2268 6403 2272
rect 6253 2188 6259 2212
rect 6285 2128 6291 2252
rect 6413 2168 6419 2272
rect 6445 2188 6451 2292
rect 6493 2248 6499 2492
rect 6525 2443 6531 2532
rect 6573 2528 6579 2632
rect 6685 2588 6691 2692
rect 6733 2548 6739 2832
rect 6829 2668 6835 2672
rect 6749 2528 6755 2532
rect 6813 2528 6819 2532
rect 6861 2528 6867 2532
rect 6877 2528 6883 2632
rect 6893 2588 6899 2692
rect 6941 2648 6947 2912
rect 7005 2888 7011 2912
rect 6973 2728 6979 2832
rect 6941 2588 6947 2592
rect 6941 2548 6947 2572
rect 6717 2508 6723 2512
rect 6797 2488 6803 2512
rect 6525 2437 6547 2443
rect 6525 2308 6531 2312
rect 6509 2228 6515 2252
rect 6541 2148 6547 2437
rect 6733 2428 6739 2432
rect 6221 2108 6227 2112
rect 6205 2017 6227 2023
rect 6061 1506 6067 1512
rect 6013 1368 6019 1412
rect 5949 1357 5971 1363
rect 5949 1188 5955 1357
rect 5949 928 5955 1052
rect 5965 948 5971 1312
rect 6013 1108 6019 1112
rect 6109 1108 6115 1212
rect 5997 948 6003 972
rect 6013 928 6019 1092
rect 6029 988 6035 1052
rect 6109 928 6115 952
rect 6141 928 6147 1612
rect 6189 1523 6195 1952
rect 6205 1708 6211 1712
rect 6189 1517 6200 1523
rect 6205 1508 6211 1512
rect 6173 1488 6179 1492
rect 6221 1488 6227 2017
rect 6285 1928 6291 2112
rect 6333 1948 6339 2032
rect 6445 1908 6451 2112
rect 6237 1888 6243 1892
rect 6317 1848 6323 1872
rect 6333 1788 6339 1812
rect 6269 1748 6275 1772
rect 6429 1763 6435 1852
rect 6429 1757 6451 1763
rect 6445 1748 6451 1757
rect 6301 1728 6307 1732
rect 6349 1728 6355 1732
rect 6429 1728 6435 1732
rect 6237 1508 6243 1512
rect 6157 1328 6163 1472
rect 6253 1428 6259 1492
rect 6285 1488 6291 1532
rect 6301 1508 6307 1612
rect 6365 1508 6371 1512
rect 6269 1468 6275 1472
rect 6173 1328 6179 1372
rect 6285 1363 6291 1472
rect 6280 1357 6291 1363
rect 6333 1363 6339 1492
rect 6397 1408 6403 1632
rect 6445 1508 6451 1732
rect 6413 1488 6419 1492
rect 6333 1357 6344 1363
rect 6157 1148 6163 1312
rect 6189 1048 6195 1052
rect 6157 948 6163 992
rect 6205 968 6211 1272
rect 6237 1108 6243 1332
rect 6301 1328 6307 1332
rect 6285 1108 6291 1192
rect 6461 1108 6467 1972
rect 6477 1728 6483 2092
rect 6589 2088 6595 2252
rect 6653 2148 6659 2372
rect 6669 2308 6675 2312
rect 6669 2208 6675 2292
rect 6733 2288 6739 2412
rect 6749 2288 6755 2352
rect 6829 2308 6835 2432
rect 6845 2308 6851 2332
rect 6861 2308 6867 2312
rect 6685 2128 6691 2232
rect 6701 2108 6707 2232
rect 6493 1906 6499 1912
rect 6493 1788 6499 1792
rect 6477 1708 6483 1712
rect 6541 1708 6547 1732
rect 6573 1728 6579 1932
rect 6541 1668 6547 1692
rect 6509 1608 6515 1652
rect 6573 1648 6579 1712
rect 6509 1508 6515 1592
rect 6541 1528 6547 1532
rect 6589 1528 6595 2072
rect 6605 1928 6611 2032
rect 6669 1948 6675 2032
rect 6701 1968 6707 2092
rect 6621 1908 6627 1932
rect 6701 1928 6707 1932
rect 6669 1908 6675 1912
rect 6717 1908 6723 2032
rect 6733 1928 6739 1932
rect 6733 1908 6739 1912
rect 6749 1888 6755 2272
rect 6781 2148 6787 2152
rect 6621 1748 6627 1832
rect 6669 1788 6675 1852
rect 6605 1508 6611 1532
rect 6573 1488 6579 1492
rect 6493 1348 6499 1352
rect 6509 1328 6515 1332
rect 6525 1128 6531 1412
rect 6541 1328 6547 1332
rect 6557 1308 6563 1432
rect 6573 1428 6579 1472
rect 6589 1468 6595 1472
rect 6589 1448 6595 1452
rect 6621 1368 6627 1732
rect 6669 1608 6675 1632
rect 6669 1508 6675 1512
rect 6637 1488 6643 1492
rect 6685 1468 6691 1872
rect 6749 1748 6755 1872
rect 6749 1708 6755 1712
rect 6765 1528 6771 1952
rect 6781 1868 6787 1892
rect 6813 1888 6819 2272
rect 6893 2248 6899 2312
rect 6845 2168 6851 2172
rect 6845 1908 6851 1912
rect 6909 1908 6915 1912
rect 6925 1888 6931 1912
rect 6941 1908 6947 2512
rect 6989 2508 6995 2712
rect 7005 2588 7011 2872
rect 7021 2708 7027 2712
rect 7037 2668 7043 2692
rect 7053 2548 7059 2572
rect 7037 2508 7043 2512
rect 6957 2288 6963 2352
rect 6989 2328 6995 2452
rect 7053 2448 7059 2532
rect 7101 2468 7107 3292
rect 7133 3188 7139 3272
rect 7197 3248 7203 3292
rect 7213 3188 7219 3477
rect 7277 3468 7283 3512
rect 7325 3508 7331 4592
rect 7421 4588 7427 4652
rect 7341 4388 7347 4512
rect 7453 4468 7459 4672
rect 7485 4668 7491 4672
rect 7501 4603 7507 4632
rect 7485 4597 7507 4603
rect 7485 4508 7491 4597
rect 7501 4548 7507 4572
rect 7341 4348 7347 4372
rect 7405 4308 7411 4352
rect 7373 4268 7379 4272
rect 7405 4188 7411 4252
rect 7421 4188 7427 4372
rect 7501 4308 7507 4532
rect 7533 4528 7539 4712
rect 7549 4568 7555 4832
rect 7565 4668 7571 4692
rect 7581 4668 7587 4672
rect 7597 4643 7603 4832
rect 7613 4768 7619 5052
rect 7645 5048 7651 5092
rect 7661 5088 7667 5297
rect 7709 5188 7715 5292
rect 7789 5288 7795 5292
rect 7661 5028 7667 5072
rect 7773 5048 7779 5232
rect 7661 4868 7667 4972
rect 7789 4948 7795 5252
rect 7805 4988 7811 5472
rect 7837 5268 7843 5472
rect 7933 5388 7939 5452
rect 7901 5328 7907 5352
rect 7981 5188 7987 5332
rect 7917 5068 7923 5072
rect 7853 4948 7859 5012
rect 7869 5008 7875 5032
rect 7949 4988 7955 5092
rect 7997 4948 8003 4952
rect 7693 4928 7699 4932
rect 7613 4708 7619 4712
rect 7661 4708 7667 4852
rect 7693 4788 7699 4912
rect 7805 4828 7811 4892
rect 7789 4708 7795 4712
rect 7581 4637 7603 4643
rect 7581 4548 7587 4637
rect 7661 4608 7667 4692
rect 7677 4548 7683 4612
rect 7725 4588 7731 4672
rect 7517 4448 7523 4512
rect 7453 4288 7459 4292
rect 7517 4288 7523 4292
rect 7501 4268 7507 4272
rect 7581 4228 7587 4532
rect 7597 4508 7603 4512
rect 7741 4508 7747 4692
rect 7805 4683 7811 4692
rect 7821 4688 7827 4712
rect 7800 4677 7811 4683
rect 7837 4568 7843 4572
rect 7789 4528 7795 4532
rect 7901 4306 7907 4872
rect 7917 4848 7923 4932
rect 8029 4908 8035 4912
rect 7949 4888 7955 4892
rect 7965 4708 7971 4892
rect 7917 4388 7923 4492
rect 7517 4168 7523 4172
rect 7613 4143 7619 4272
rect 7608 4137 7619 4143
rect 7549 4128 7555 4132
rect 7405 3908 7411 3912
rect 7453 3908 7459 3932
rect 7549 3888 7555 4112
rect 7581 4108 7587 4112
rect 7597 4108 7603 4112
rect 7581 3888 7587 3892
rect 7597 3888 7603 3892
rect 7485 3868 7491 3872
rect 7485 3768 7491 3852
rect 7549 3748 7555 3752
rect 7597 3748 7603 3872
rect 7613 3868 7619 4137
rect 7629 4108 7635 4292
rect 7725 4288 7731 4292
rect 7693 4128 7699 4212
rect 7709 4148 7715 4252
rect 7645 4108 7651 4112
rect 7693 3968 7699 4112
rect 7709 3908 7715 4132
rect 7805 4128 7811 4232
rect 7901 4148 7907 4252
rect 7933 4168 7939 4432
rect 7821 4128 7827 4132
rect 7725 3908 7731 4092
rect 7805 3908 7811 4112
rect 7901 3948 7907 4132
rect 7933 4128 7939 4132
rect 7949 4128 7955 4372
rect 7965 4368 7971 4532
rect 7981 4528 7987 4592
rect 7997 4188 8003 4692
rect 8013 4308 8019 4432
rect 8029 4388 8035 4892
rect 7981 4108 7987 4152
rect 8013 4108 8019 4112
rect 7736 3897 7747 3903
rect 7645 3748 7651 3872
rect 7709 3868 7715 3872
rect 7693 3848 7699 3852
rect 7373 3728 7379 3732
rect 7373 3708 7379 3712
rect 7453 3668 7459 3712
rect 7533 3648 7539 3712
rect 7597 3648 7603 3732
rect 7421 3528 7427 3552
rect 7485 3548 7491 3552
rect 7453 3528 7459 3532
rect 7485 3528 7491 3532
rect 7532 3517 7555 3523
rect 7293 3448 7299 3492
rect 7261 3268 7267 3332
rect 7277 3288 7283 3292
rect 7149 3128 7155 3132
rect 7213 2728 7219 3132
rect 7245 3003 7251 3072
rect 7229 2997 7251 3003
rect 7229 2928 7235 2997
rect 7213 2708 7219 2712
rect 7149 2588 7155 2672
rect 7213 2428 7219 2692
rect 7229 2668 7235 2912
rect 7293 2848 7299 3432
rect 7325 3348 7331 3492
rect 7437 3488 7443 3512
rect 7453 3508 7459 3512
rect 7549 3508 7555 3517
rect 7645 3488 7651 3732
rect 7741 3728 7747 3897
rect 7901 3888 7907 3932
rect 7949 3908 7955 4032
rect 7757 3748 7763 3852
rect 7661 3688 7667 3712
rect 7741 3628 7747 3712
rect 7757 3648 7763 3732
rect 7389 3328 7395 3472
rect 7485 3368 7491 3372
rect 7309 3288 7315 3312
rect 7437 3308 7443 3312
rect 7549 3268 7555 3332
rect 7565 3308 7571 3312
rect 7565 3288 7571 3292
rect 7309 3106 7315 3232
rect 7485 3108 7491 3112
rect 7581 3088 7587 3472
rect 7677 3388 7683 3472
rect 7741 3368 7747 3372
rect 7661 3288 7667 3332
rect 7757 3328 7763 3332
rect 7597 3108 7603 3252
rect 7693 3148 7699 3192
rect 7773 3168 7779 3832
rect 7789 3448 7795 3492
rect 7805 3388 7811 3732
rect 7853 3728 7859 3732
rect 7821 3588 7827 3632
rect 7885 3588 7891 3612
rect 7837 3288 7843 3292
rect 7805 3148 7811 3172
rect 7693 3128 7699 3132
rect 7805 3128 7811 3132
rect 7613 3108 7619 3112
rect 7677 3108 7683 3112
rect 7453 2948 7459 3072
rect 7581 3008 7587 3072
rect 7309 2908 7315 2932
rect 7293 2708 7299 2832
rect 7293 2668 7299 2692
rect 7229 2548 7235 2652
rect 7309 2508 7315 2872
rect 7325 2788 7331 2932
rect 7421 2728 7427 2892
rect 7469 2688 7475 2932
rect 7501 2708 7507 2912
rect 6989 2268 6995 2312
rect 7005 2188 7011 2272
rect 7101 2188 7107 2252
rect 7165 2248 7171 2292
rect 7197 2268 7203 2272
rect 6957 2128 6963 2132
rect 7005 2108 7011 2112
rect 7021 2108 7027 2132
rect 7133 2128 7139 2192
rect 7165 2128 7171 2132
rect 7197 2123 7203 2252
rect 7245 2228 7251 2272
rect 7261 2268 7267 2292
rect 7325 2268 7331 2312
rect 7192 2117 7203 2123
rect 6957 1908 6963 1912
rect 7021 1888 7027 2092
rect 6781 1548 6787 1632
rect 6797 1588 6803 1712
rect 6797 1508 6803 1512
rect 6733 1448 6739 1472
rect 6749 1388 6755 1412
rect 6765 1308 6771 1432
rect 6813 1363 6819 1432
rect 6813 1357 6835 1363
rect 6525 1108 6531 1112
rect 6237 1028 6243 1052
rect 6397 1048 6403 1052
rect 6397 1008 6403 1032
rect 6221 968 6227 972
rect 6269 948 6275 952
rect 6413 948 6419 1092
rect 6541 1088 6547 1252
rect 6781 1228 6787 1312
rect 6797 1308 6803 1312
rect 6813 1288 6819 1312
rect 6829 1308 6835 1357
rect 6845 1323 6851 1872
rect 6877 1768 6883 1872
rect 7021 1868 7027 1872
rect 6909 1708 6915 1832
rect 6957 1728 6963 1752
rect 7069 1728 7075 1892
rect 7101 1768 7107 2032
rect 7197 1948 7203 2032
rect 7165 1888 7171 1892
rect 7213 1748 7219 1852
rect 7245 1788 7251 2212
rect 7293 1908 7299 2192
rect 7309 2168 7315 2192
rect 7341 1928 7347 2632
rect 7357 2548 7363 2672
rect 7357 2488 7363 2532
rect 7405 2528 7411 2632
rect 7453 2568 7459 2672
rect 7485 2588 7491 2612
rect 7517 2608 7523 2692
rect 7549 2688 7555 2992
rect 7389 2368 7395 2492
rect 7421 2488 7427 2512
rect 7485 2508 7491 2512
rect 7517 2488 7523 2512
rect 7469 2308 7475 2312
rect 7341 1908 7347 1912
rect 7357 1888 7363 2252
rect 7373 2208 7379 2272
rect 7405 2188 7411 2232
rect 7405 2168 7411 2172
rect 7437 2128 7443 2272
rect 7469 2088 7475 2292
rect 7485 2288 7491 2432
rect 7533 2388 7539 2532
rect 7549 2368 7555 2672
rect 7565 2528 7571 2672
rect 7581 2588 7587 2932
rect 7613 2928 7619 2932
rect 7629 2928 7635 3092
rect 7789 3088 7795 3112
rect 7645 2948 7651 3072
rect 7709 2963 7715 3052
rect 7725 2988 7731 3032
rect 7805 3028 7811 3032
rect 7709 2957 7731 2963
rect 7645 2908 7651 2912
rect 7597 2728 7603 2872
rect 7485 2228 7491 2272
rect 7501 2268 7507 2272
rect 7533 2137 7544 2143
rect 7501 2128 7507 2132
rect 7405 1988 7411 2072
rect 7405 1908 7411 1972
rect 7485 1928 7491 2072
rect 7501 1908 7507 1912
rect 7517 1908 7523 2112
rect 7085 1688 7091 1732
rect 6909 1468 6915 1472
rect 6877 1348 6883 1452
rect 6893 1388 6899 1432
rect 6925 1368 6931 1492
rect 6941 1468 6947 1472
rect 6845 1317 6856 1323
rect 6877 1188 6883 1332
rect 6893 1288 6899 1292
rect 6909 1208 6915 1292
rect 6429 948 6435 1032
rect 6509 1008 6515 1032
rect 6541 1028 6547 1072
rect 6701 1068 6707 1072
rect 6797 1068 6803 1072
rect 6509 968 6515 972
rect 6525 948 6531 952
rect 6461 937 6499 943
rect 6285 928 6291 932
rect 5821 788 5827 832
rect 5677 548 5683 552
rect 5693 528 5699 552
rect 5677 508 5683 512
rect 5677 328 5683 492
rect 5629 168 5635 252
rect 5629 148 5635 152
rect 5661 148 5667 312
rect 5709 308 5715 652
rect 5789 548 5795 632
rect 5741 528 5747 532
rect 5853 308 5859 712
rect 5869 548 5875 692
rect 5885 648 5891 692
rect 5901 603 5907 832
rect 5933 688 5939 692
rect 5949 688 5955 912
rect 5981 908 5987 912
rect 6109 788 6115 912
rect 6141 908 6147 912
rect 6157 868 6163 912
rect 6253 903 6259 912
rect 6317 908 6323 912
rect 6253 897 6296 903
rect 6333 848 6339 932
rect 6461 928 6467 937
rect 6493 928 6499 937
rect 6541 928 6547 972
rect 6589 948 6595 1052
rect 5981 728 5987 732
rect 5901 597 5923 603
rect 5885 568 5891 572
rect 5880 537 5891 543
rect 5885 388 5891 537
rect 5885 328 5891 372
rect 5917 368 5923 597
rect 5965 508 5971 632
rect 5997 528 6003 732
rect 6029 588 6035 672
rect 6093 548 6099 692
rect 5725 148 5731 192
rect 5837 188 5843 272
rect 5837 143 5843 172
rect 5965 168 5971 312
rect 5997 228 6003 292
rect 6013 248 6019 532
rect 6157 288 6163 772
rect 6221 728 6227 732
rect 6189 648 6195 672
rect 6013 208 6019 232
rect 6109 228 6115 232
rect 5997 148 6003 152
rect 6109 148 6115 212
rect 6189 188 6195 532
rect 6205 508 6211 632
rect 6221 608 6227 712
rect 6237 708 6243 732
rect 6269 728 6275 792
rect 6285 737 6339 743
rect 6269 708 6275 712
rect 6285 708 6291 737
rect 6333 728 6339 737
rect 6317 708 6323 712
rect 6477 708 6483 912
rect 6237 688 6243 692
rect 6285 628 6291 672
rect 6301 528 6307 592
rect 6317 563 6323 632
rect 6317 557 6339 563
rect 6205 208 6211 292
rect 6317 268 6323 532
rect 6333 508 6339 557
rect 6365 528 6371 692
rect 6493 688 6499 692
rect 6509 688 6515 872
rect 6381 668 6387 672
rect 6509 548 6515 672
rect 6541 623 6547 912
rect 6573 908 6579 912
rect 6589 768 6595 932
rect 6637 903 6643 1032
rect 6653 928 6659 932
rect 6637 897 6659 903
rect 6653 788 6659 897
rect 6685 848 6691 952
rect 6733 948 6739 952
rect 6717 888 6723 912
rect 6749 908 6755 1052
rect 6765 948 6771 952
rect 6829 948 6835 1172
rect 6893 1128 6899 1132
rect 6941 1068 6947 1332
rect 6957 1128 6963 1512
rect 6973 1468 6979 1512
rect 7053 1508 7059 1512
rect 7069 1468 7075 1572
rect 6973 1328 6979 1352
rect 6989 1328 6995 1332
rect 7005 1308 7011 1432
rect 7069 1388 7075 1452
rect 6989 1088 6995 1092
rect 6893 968 6899 1052
rect 6893 948 6899 952
rect 6765 888 6771 912
rect 6877 908 6883 932
rect 6957 928 6963 932
rect 6669 808 6675 832
rect 6765 788 6771 832
rect 6749 708 6755 732
rect 6621 688 6627 692
rect 6541 617 6563 623
rect 6349 388 6355 452
rect 6397 328 6403 332
rect 6397 308 6403 312
rect 6221 148 6227 172
rect 6317 168 6323 252
rect 6317 148 6323 152
rect 6333 148 6339 292
rect 6381 208 6387 292
rect 6477 288 6483 532
rect 6557 468 6563 617
rect 6589 588 6595 632
rect 6637 608 6643 692
rect 6605 388 6611 592
rect 6653 588 6659 652
rect 6685 608 6691 692
rect 6733 688 6739 692
rect 6525 308 6531 312
rect 6365 188 6371 192
rect 6445 188 6451 272
rect 6461 188 6467 212
rect 5837 137 5848 143
rect 4557 108 4563 114
rect 5597 108 5603 112
rect 5661 108 5667 132
rect 5709 128 5715 132
rect 5965 108 5971 132
rect 6045 128 6051 132
rect 6493 128 6499 292
rect 6509 148 6515 152
rect 6589 128 6595 352
rect 6621 308 6627 512
rect 6637 308 6643 352
rect 6653 308 6659 312
rect 6621 228 6627 272
rect 6621 168 6627 192
rect 6717 163 6723 532
rect 6749 508 6755 514
rect 6733 328 6739 352
rect 6765 288 6771 752
rect 6797 688 6803 692
rect 6861 668 6867 852
rect 6909 688 6915 792
rect 6925 708 6931 912
rect 6989 848 6995 912
rect 7005 908 7011 1032
rect 7053 928 7059 1172
rect 7069 948 7075 1032
rect 7085 948 7091 1152
rect 7101 1148 7107 1492
rect 7133 1468 7139 1472
rect 7101 1128 7107 1132
rect 7053 883 7059 912
rect 7101 908 7107 912
rect 7037 877 7059 883
rect 7037 783 7043 877
rect 7037 777 7048 783
rect 7117 728 7123 992
rect 7021 708 7027 712
rect 7117 708 7123 712
rect 6813 568 6819 612
rect 6861 448 6867 652
rect 6909 528 6915 552
rect 6909 388 6915 452
rect 6845 308 6851 332
rect 6893 308 6899 332
rect 6957 308 6963 532
rect 6781 268 6787 292
rect 6829 168 6835 292
rect 6941 288 6947 292
rect 6957 188 6963 292
rect 6973 228 6979 532
rect 7037 528 7043 692
rect 7069 548 7075 592
rect 7037 508 7043 512
rect 7005 388 7011 492
rect 6989 288 6995 332
rect 7021 328 7027 472
rect 7133 328 7139 1392
rect 7165 1348 7171 1732
rect 7229 1528 7235 1752
rect 7245 1728 7251 1732
rect 7245 1528 7251 1672
rect 7261 1528 7267 1812
rect 7341 1748 7347 1792
rect 7229 1508 7235 1512
rect 7245 1488 7251 1512
rect 7293 1508 7299 1712
rect 7341 1668 7347 1712
rect 7261 1488 7267 1492
rect 7293 1488 7299 1492
rect 7277 1477 7288 1483
rect 7181 1437 7192 1443
rect 7181 1328 7187 1437
rect 7149 1088 7155 1112
rect 7149 828 7155 932
rect 7213 868 7219 932
rect 7245 908 7251 1152
rect 7261 988 7267 1452
rect 7277 1328 7283 1477
rect 7277 1188 7283 1312
rect 7293 1088 7299 1312
rect 7341 1228 7347 1312
rect 7357 1168 7363 1872
rect 7469 1828 7475 1832
rect 7437 1728 7443 1752
rect 7469 1748 7475 1792
rect 7517 1768 7523 1892
rect 7533 1868 7539 2137
rect 7565 2143 7571 2332
rect 7581 2328 7587 2512
rect 7597 2508 7603 2632
rect 7629 2548 7635 2852
rect 7645 2548 7651 2892
rect 7709 2888 7715 2892
rect 7693 2568 7699 2652
rect 7709 2588 7715 2692
rect 7613 2468 7619 2512
rect 7629 2448 7635 2532
rect 7725 2528 7731 2957
rect 7773 2948 7779 2992
rect 7757 2868 7763 2912
rect 7821 2788 7827 3232
rect 7837 3148 7843 3272
rect 7869 3128 7875 3212
rect 7885 3148 7891 3312
rect 7901 3248 7907 3872
rect 7965 3848 7971 3852
rect 8013 3788 8019 4092
rect 8029 3988 8035 4352
rect 8045 4188 8051 4232
rect 8045 4148 8051 4172
rect 8045 3668 8051 3712
rect 7917 3348 7923 3352
rect 7917 3188 7923 3272
rect 7885 3068 7891 3132
rect 7901 3108 7907 3172
rect 7789 2628 7795 2672
rect 7661 2517 7672 2523
rect 7581 2208 7587 2312
rect 7629 2308 7635 2392
rect 7661 2388 7667 2517
rect 7677 2483 7683 2492
rect 7741 2488 7747 2512
rect 7677 2477 7699 2483
rect 7645 2288 7651 2312
rect 7560 2137 7571 2143
rect 7549 2103 7555 2112
rect 7581 2103 7587 2152
rect 7661 2148 7667 2352
rect 7677 2328 7683 2412
rect 7693 2388 7699 2477
rect 7789 2428 7795 2552
rect 7821 2528 7827 2652
rect 7869 2628 7875 2912
rect 7901 2908 7907 3032
rect 7917 2708 7923 3152
rect 7933 3108 7939 3652
rect 7949 3288 7955 3492
rect 7997 3328 8003 3332
rect 7965 3208 7971 3292
rect 7981 3188 7987 3292
rect 7869 2528 7875 2532
rect 7933 2528 7939 3092
rect 7997 2688 8003 3232
rect 8013 2968 8019 3132
rect 8029 2988 8035 3332
rect 7709 2288 7715 2412
rect 7853 2348 7859 2432
rect 7949 2308 7955 2452
rect 7981 2388 7987 2612
rect 7997 2408 8003 2432
rect 7597 2108 7603 2112
rect 7661 2108 7667 2112
rect 7549 2097 7587 2103
rect 7597 2088 7603 2092
rect 7629 2088 7635 2092
rect 7629 1928 7635 1952
rect 7693 1928 7699 1952
rect 7517 1728 7523 1752
rect 7533 1748 7539 1852
rect 7549 1728 7555 1832
rect 7373 1388 7379 1452
rect 7309 1106 7315 1132
rect 7341 1008 7347 1072
rect 7277 928 7283 932
rect 7405 928 7411 1672
rect 7421 1528 7427 1692
rect 7517 1688 7523 1692
rect 7421 1488 7427 1492
rect 7469 1488 7475 1492
rect 7469 1328 7475 1332
rect 7421 1128 7427 1152
rect 7453 1108 7459 1132
rect 7469 948 7475 1312
rect 7485 1268 7491 1472
rect 7501 1348 7507 1652
rect 7517 1508 7523 1632
rect 7597 1508 7603 1872
rect 7645 1868 7651 1872
rect 7613 1528 7619 1832
rect 7693 1708 7699 1712
rect 7645 1528 7651 1692
rect 7709 1548 7715 2192
rect 7853 2148 7859 2272
rect 7725 1908 7731 1932
rect 7741 1788 7747 1892
rect 7757 1888 7763 2132
rect 7773 2088 7779 2112
rect 7789 1988 7795 2072
rect 7853 2048 7859 2132
rect 7949 2128 7955 2292
rect 7981 2188 7987 2232
rect 7917 2108 7923 2112
rect 7757 1808 7763 1872
rect 7773 1868 7779 1872
rect 7885 1728 7891 2092
rect 7933 2088 7939 2092
rect 7917 1728 7923 1872
rect 7933 1768 7939 1912
rect 7949 1908 7955 1932
rect 7709 1508 7715 1532
rect 7517 1368 7523 1492
rect 7693 1488 7699 1492
rect 7549 1448 7555 1472
rect 7629 1448 7635 1472
rect 7709 1468 7715 1472
rect 7549 1348 7555 1432
rect 7661 1348 7667 1372
rect 7485 1108 7491 1152
rect 7501 1088 7507 1332
rect 7581 1328 7587 1332
rect 7517 1308 7523 1314
rect 7613 1308 7619 1312
rect 7517 1188 7523 1212
rect 7549 988 7555 992
rect 7581 988 7587 1252
rect 7677 1188 7683 1432
rect 7709 1388 7715 1432
rect 7757 1388 7763 1512
rect 7693 1308 7699 1312
rect 7645 1106 7651 1132
rect 7741 1128 7747 1152
rect 7613 1008 7619 1072
rect 7197 728 7203 732
rect 7165 688 7171 712
rect 7213 528 7219 532
rect 7133 308 7139 312
rect 7037 288 7043 292
rect 7149 283 7155 292
rect 7144 277 7155 283
rect 6712 157 6723 163
rect 6621 148 6627 152
rect 6893 148 6899 152
rect 6957 148 6963 172
rect 7229 168 7235 252
rect 7229 148 7235 152
rect 6717 128 6723 132
rect 7101 128 7107 132
rect 7261 128 7267 692
rect 7293 548 7299 732
rect 7325 708 7331 772
rect 7469 748 7475 932
rect 7517 928 7523 932
rect 7709 928 7715 1052
rect 7341 708 7347 732
rect 7421 548 7427 672
rect 7293 288 7299 532
rect 7293 148 7299 272
rect 7325 188 7331 532
rect 7453 530 7459 532
rect 7341 488 7347 512
rect 7437 388 7443 432
rect 7485 308 7491 712
rect 7517 706 7523 812
rect 7549 688 7555 832
rect 7645 788 7651 852
rect 7709 788 7715 872
rect 7677 708 7683 712
rect 7549 568 7555 672
rect 7629 588 7635 672
rect 7549 328 7555 472
rect 7581 348 7587 432
rect 7661 388 7667 512
rect 7549 308 7555 312
rect 7709 308 7715 312
rect 7325 148 7331 172
rect 7405 168 7411 272
rect 7421 268 7427 292
rect 7517 288 7523 292
rect 7725 288 7731 432
rect 7757 308 7763 1312
rect 7773 1308 7779 1532
rect 7869 1508 7875 1512
rect 7853 1488 7859 1492
rect 7805 1368 7811 1472
rect 7805 1348 7811 1352
rect 7789 1148 7795 1152
rect 7773 1108 7779 1132
rect 7789 1108 7795 1132
rect 7773 688 7779 832
rect 7805 728 7811 1092
rect 7821 1088 7827 1332
rect 7869 1308 7875 1332
rect 7885 1288 7891 1332
rect 7901 1328 7907 1712
rect 7965 1648 7971 2112
rect 7997 1983 8003 2032
rect 7981 1977 8003 1983
rect 7981 1888 7987 1977
rect 7837 1228 7843 1232
rect 7853 1188 7859 1232
rect 7853 1108 7859 1152
rect 7869 1128 7875 1172
rect 7901 1148 7907 1312
rect 7917 1283 7923 1312
rect 7965 1308 7971 1312
rect 7917 1277 7939 1283
rect 7885 1108 7891 1112
rect 7837 988 7843 1032
rect 7773 528 7779 572
rect 7789 503 7795 632
rect 7805 588 7811 712
rect 7853 688 7859 732
rect 7917 668 7923 1072
rect 7933 708 7939 1277
rect 7949 1048 7955 1052
rect 7981 1003 7987 1872
rect 7997 1528 8003 1632
rect 7997 1108 8003 1492
rect 8029 1488 8035 1492
rect 8013 1363 8019 1432
rect 8013 1357 8035 1363
rect 7965 997 7987 1003
rect 7965 928 7971 997
rect 7981 708 7987 712
rect 7853 548 7859 552
rect 7805 528 7811 532
rect 7789 497 7800 503
rect 7901 288 7907 532
rect 7517 188 7523 272
rect 7629 268 7635 272
rect 7645 128 7651 232
rect 7757 188 7763 252
rect 7869 128 7875 232
rect 7901 168 7907 272
rect 7981 188 7987 652
rect 7997 388 8003 1052
rect 8013 968 8019 1332
rect 8029 1128 8035 1357
rect 8013 948 8019 952
rect 8013 588 8019 672
rect 7997 168 8003 232
rect 6205 108 6211 112
rect 6381 108 6387 112
rect 6589 108 6595 112
rect 6861 108 6867 112
rect 7261 108 7267 112
rect 7293 108 7299 112
rect 7421 108 7427 112
rect 3789 -43 3795 32
rect 3837 -43 3843 32
rect 4093 -43 4099 32
rect 4141 -43 4147 32
rect 4189 -43 4195 32
rect 4237 -43 4243 32
rect 4333 -43 4339 12
rect 4381 -43 4387 32
rect 4429 -43 4435 32
rect 4701 -43 4707 32
<< m3contact >>
rect 925 5602 961 5618
rect 1640 5512 1656 5528
rect 72 5472 88 5488
rect 136 5372 152 5388
rect 88 5352 104 5368
rect 376 5492 392 5508
rect 520 5492 536 5508
rect 232 5472 248 5488
rect 392 5472 408 5488
rect 344 5392 360 5408
rect 216 5352 232 5368
rect 264 5352 280 5368
rect 152 5332 168 5348
rect 248 5332 264 5348
rect 40 5312 56 5328
rect 88 5312 104 5328
rect 104 5312 120 5328
rect 248 5312 264 5328
rect 72 5232 88 5248
rect 40 5032 56 5048
rect 24 5012 40 5028
rect 88 5112 104 5128
rect 88 5072 104 5088
rect 40 4692 56 4708
rect 40 4672 56 4688
rect 88 4672 104 4688
rect 40 4552 56 4568
rect 24 4372 40 4388
rect 40 4272 56 4288
rect 56 4252 72 4268
rect 136 5092 152 5108
rect 216 5072 232 5088
rect 216 5052 232 5068
rect 248 5052 264 5068
rect 152 4952 168 4968
rect 120 4912 136 4928
rect 248 4932 264 4948
rect 168 4912 184 4928
rect 216 4912 232 4928
rect 248 4912 264 4928
rect 136 4892 152 4908
rect 136 4752 152 4768
rect 136 4732 152 4748
rect 184 4812 200 4828
rect 200 4792 216 4808
rect 168 4752 184 4768
rect 200 4732 216 4748
rect 120 4692 136 4708
rect 152 4612 168 4628
rect 120 4492 136 4508
rect 424 5372 440 5388
rect 744 5492 760 5508
rect 776 5492 792 5508
rect 824 5492 840 5508
rect 952 5492 968 5508
rect 1064 5506 1080 5508
rect 1064 5492 1080 5506
rect 648 5472 664 5488
rect 584 5452 600 5468
rect 504 5352 520 5368
rect 584 5352 600 5368
rect 760 5472 776 5488
rect 728 5392 744 5408
rect 376 5312 392 5328
rect 504 5312 520 5328
rect 552 5312 568 5328
rect 680 5312 696 5328
rect 280 5112 296 5128
rect 312 5072 328 5088
rect 440 5072 456 5088
rect 376 5032 392 5048
rect 328 5012 344 5028
rect 728 5132 744 5148
rect 584 5092 600 5108
rect 664 5092 680 5108
rect 472 4972 488 4988
rect 392 4932 408 4948
rect 424 4932 440 4948
rect 472 4932 488 4948
rect 312 4912 328 4928
rect 264 4892 280 4908
rect 344 4892 360 4908
rect 232 4872 248 4888
rect 296 4872 312 4888
rect 312 4872 328 4888
rect 360 4872 376 4888
rect 248 4772 264 4788
rect 280 4772 296 4788
rect 232 4732 248 4748
rect 232 4692 248 4708
rect 248 4692 264 4708
rect 280 4692 296 4708
rect 216 4672 232 4688
rect 184 4512 200 4528
rect 200 4492 216 4508
rect 280 4652 296 4668
rect 376 4832 392 4848
rect 344 4732 360 4748
rect 312 4692 328 4708
rect 440 4912 456 4928
rect 488 4912 504 4928
rect 488 4792 504 4808
rect 760 5012 776 5028
rect 744 4952 760 4968
rect 632 4932 648 4948
rect 536 4772 552 4788
rect 552 4752 568 4768
rect 472 4732 488 4748
rect 536 4732 552 4748
rect 552 4732 568 4748
rect 376 4712 392 4728
rect 376 4692 392 4708
rect 360 4672 376 4688
rect 344 4632 360 4648
rect 296 4592 312 4608
rect 248 4512 264 4528
rect 296 4512 312 4528
rect 360 4512 376 4528
rect 280 4492 296 4508
rect 344 4492 360 4508
rect 424 4692 440 4708
rect 408 4672 424 4688
rect 424 4612 440 4628
rect 520 4712 536 4728
rect 504 4652 520 4668
rect 792 5452 808 5468
rect 808 5352 824 5368
rect 872 5452 888 5468
rect 888 5352 904 5368
rect 840 5332 856 5348
rect 856 5312 872 5328
rect 808 5072 824 5088
rect 824 5052 840 5068
rect 824 5012 840 5028
rect 792 4992 808 5008
rect 824 4952 840 4968
rect 792 4932 808 4948
rect 776 4912 792 4928
rect 664 4772 680 4788
rect 536 4612 552 4628
rect 488 4592 504 4608
rect 424 4532 440 4548
rect 472 4512 488 4528
rect 312 4472 328 4488
rect 440 4472 456 4488
rect 248 4452 264 4468
rect 168 4372 184 4388
rect 232 4372 248 4388
rect 248 4352 264 4368
rect 312 4312 328 4328
rect 232 4292 248 4308
rect 56 4112 72 4128
rect 8 3932 24 3948
rect 8 3912 24 3928
rect 8 3512 24 3528
rect 104 3932 120 3948
rect 88 3912 104 3928
rect 40 3872 56 3888
rect 88 3892 104 3908
rect 56 3772 72 3788
rect 40 3752 56 3768
rect 88 3752 104 3768
rect 248 4272 264 4288
rect 216 4232 232 4248
rect 296 4232 312 4248
rect 248 4212 264 4228
rect 200 4112 216 4128
rect 248 4112 264 4128
rect 296 4112 312 4128
rect 184 3992 200 4008
rect 168 3952 184 3968
rect 152 3912 168 3928
rect 168 3872 184 3888
rect 184 3852 200 3868
rect 232 4092 248 4108
rect 248 4072 264 4088
rect 280 4072 296 4088
rect 296 4072 312 4088
rect 264 4032 280 4048
rect 248 3952 264 3968
rect 232 3932 248 3948
rect 216 3892 232 3908
rect 200 3772 232 3788
rect 152 3752 168 3768
rect 136 3732 152 3748
rect 344 4452 360 4468
rect 392 4432 408 4448
rect 440 4372 456 4388
rect 376 4332 392 4348
rect 424 4332 440 4348
rect 360 4272 376 4288
rect 408 4252 424 4268
rect 424 4232 440 4248
rect 360 4112 376 4128
rect 328 4072 344 4088
rect 344 4072 360 4088
rect 360 4072 376 4088
rect 360 3952 376 3968
rect 280 3892 296 3908
rect 264 3852 280 3868
rect 248 3712 264 3728
rect 184 3632 200 3648
rect 40 3492 56 3508
rect 88 3352 104 3368
rect 120 3512 136 3528
rect 200 3552 216 3568
rect 232 3532 248 3548
rect 136 3492 152 3508
rect 344 3912 360 3928
rect 568 4532 584 4548
rect 504 4512 520 4528
rect 616 4512 632 4528
rect 536 4492 552 4508
rect 504 4432 520 4448
rect 504 4412 520 4428
rect 552 4432 568 4448
rect 792 4752 808 4768
rect 808 4732 824 4748
rect 696 4692 712 4708
rect 680 4612 696 4628
rect 792 4612 808 4628
rect 600 4492 616 4508
rect 664 4492 680 4508
rect 680 4472 696 4488
rect 632 4452 648 4468
rect 568 4412 584 4428
rect 520 4392 552 4408
rect 664 4392 680 4408
rect 488 4372 504 4388
rect 488 4352 504 4368
rect 584 4372 600 4388
rect 568 4332 584 4348
rect 616 4332 632 4348
rect 648 4332 664 4348
rect 488 4312 504 4328
rect 520 4312 536 4328
rect 696 4332 712 4348
rect 472 4232 488 4248
rect 440 3932 456 3948
rect 344 3892 360 3908
rect 296 3832 312 3848
rect 296 3752 312 3768
rect 312 3712 328 3728
rect 328 3712 344 3728
rect 280 3692 296 3708
rect 296 3672 312 3688
rect 328 3532 344 3548
rect 264 3472 280 3488
rect 248 3432 264 3448
rect 312 3352 328 3368
rect 216 3332 232 3348
rect 168 3312 200 3328
rect 264 3312 280 3328
rect 184 3272 200 3288
rect 40 3132 56 3148
rect 24 3112 40 3128
rect 152 3252 168 3268
rect 72 3152 88 3168
rect 120 3152 152 3168
rect 104 3112 120 3128
rect 88 3092 104 3108
rect 40 3052 56 3068
rect 296 3292 312 3308
rect 248 3252 264 3268
rect 264 3232 280 3248
rect 136 3132 152 3148
rect 152 3132 168 3148
rect 200 3132 216 3148
rect 184 3112 200 3128
rect 168 3092 184 3108
rect 168 2992 184 3008
rect 168 2972 184 2988
rect 216 3032 232 3048
rect 200 2992 216 3008
rect 40 2932 56 2948
rect 152 2932 168 2948
rect 184 2732 200 2748
rect 88 2652 104 2668
rect 312 3252 344 3268
rect 296 3032 312 3048
rect 312 2972 328 2988
rect 232 2912 248 2928
rect 296 2912 312 2928
rect 296 2732 312 2748
rect 248 2712 264 2728
rect 216 2652 232 2668
rect 152 2632 168 2648
rect 216 2632 232 2648
rect 168 2592 184 2608
rect 120 2572 136 2588
rect 184 2512 200 2528
rect 72 2492 88 2508
rect 8 2312 24 2328
rect 136 2472 152 2488
rect 120 2312 136 2328
rect 152 2292 168 2308
rect 200 2432 216 2448
rect 280 2552 296 2568
rect 200 2292 216 2308
rect 264 2292 280 2308
rect 168 2272 184 2288
rect 88 2112 104 2128
rect 168 2112 184 2128
rect 136 2072 152 2088
rect 72 1952 88 1968
rect 40 1892 56 1908
rect 88 1872 104 1888
rect 40 1792 56 1808
rect 120 1852 136 1868
rect 40 1772 56 1788
rect 104 1772 120 1788
rect 8 1712 24 1728
rect 104 1712 120 1728
rect 104 1572 120 1588
rect 40 1352 56 1368
rect 8 1312 24 1328
rect 40 1152 56 1168
rect 24 1132 40 1148
rect 40 1092 56 1108
rect 168 1892 184 1908
rect 152 1792 168 1808
rect 184 1872 200 1888
rect 184 1772 200 1788
rect 168 1712 184 1728
rect 424 3892 440 3908
rect 376 3872 392 3888
rect 424 3872 440 3888
rect 392 3852 408 3868
rect 408 3812 424 3828
rect 504 4272 520 4288
rect 488 4092 504 4108
rect 552 4292 568 4308
rect 600 4252 616 4268
rect 616 4212 632 4228
rect 680 4212 696 4228
rect 760 4332 776 4348
rect 856 4912 872 4928
rect 1096 5472 1112 5488
rect 1304 5472 1320 5488
rect 984 5392 1000 5408
rect 984 5352 1000 5368
rect 968 5332 984 5348
rect 1128 5452 1144 5468
rect 1336 5472 1352 5488
rect 1432 5472 1448 5488
rect 1320 5372 1336 5388
rect 1224 5352 1240 5368
rect 925 5202 961 5218
rect 1016 5212 1032 5228
rect 984 5132 1000 5148
rect 952 5032 968 5048
rect 984 5032 1000 5048
rect 1240 5312 1256 5328
rect 1304 5312 1320 5328
rect 1160 5292 1176 5308
rect 1256 5292 1268 5308
rect 1268 5292 1272 5308
rect 1304 5272 1320 5288
rect 1160 5232 1176 5248
rect 1096 5132 1112 5148
rect 1080 5092 1096 5108
rect 1128 5092 1144 5108
rect 1592 5472 1608 5488
rect 1784 5472 1800 5488
rect 1560 5452 1576 5468
rect 1592 5452 1608 5468
rect 1672 5432 1688 5448
rect 1528 5372 1544 5388
rect 1400 5352 1416 5368
rect 1480 5352 1512 5368
rect 1576 5332 1592 5348
rect 1624 5332 1640 5348
rect 1464 5252 1480 5268
rect 1352 5232 1368 5248
rect 1368 5112 1384 5128
rect 1464 5112 1480 5128
rect 1448 5092 1464 5108
rect 1048 5072 1064 5088
rect 1064 5072 1080 5088
rect 1096 5072 1112 5088
rect 1128 5072 1144 5088
rect 1176 5072 1192 5088
rect 1432 5072 1448 5088
rect 1448 5072 1464 5088
rect 1016 4972 1032 4988
rect 1064 4932 1080 4948
rect 904 4912 920 4928
rect 1000 4912 1016 4928
rect 1080 4912 1096 4928
rect 1048 4872 1064 4888
rect 888 4852 904 4868
rect 1000 4852 1016 4868
rect 925 4802 961 4818
rect 872 4772 888 4788
rect 984 4752 1000 4768
rect 872 4732 888 4748
rect 1000 4732 1016 4748
rect 1400 4992 1416 5008
rect 1256 4972 1272 4988
rect 1112 4932 1128 4948
rect 1272 4952 1288 4968
rect 1144 4752 1160 4768
rect 936 4712 952 4728
rect 968 4712 984 4728
rect 1016 4712 1032 4728
rect 1096 4712 1112 4728
rect 872 4692 888 4708
rect 904 4692 920 4708
rect 984 4692 1000 4708
rect 1032 4692 1048 4708
rect 808 4332 824 4348
rect 728 4312 744 4328
rect 712 4292 728 4308
rect 728 4252 744 4268
rect 744 4212 760 4228
rect 632 4092 648 4108
rect 536 4072 552 4088
rect 664 4072 680 4088
rect 552 3992 568 4008
rect 584 3992 600 4008
rect 552 3952 568 3968
rect 488 3892 504 3908
rect 536 3892 552 3908
rect 552 3812 568 3828
rect 424 3732 440 3748
rect 488 3732 504 3748
rect 552 3732 568 3748
rect 456 3692 472 3708
rect 376 3652 392 3668
rect 360 3612 376 3628
rect 440 3612 456 3628
rect 392 3512 408 3528
rect 600 3932 616 3948
rect 728 4112 744 4128
rect 696 3912 712 3928
rect 600 3892 632 3908
rect 664 3892 680 3908
rect 616 3772 632 3788
rect 680 3872 696 3888
rect 632 3752 648 3768
rect 616 3712 632 3728
rect 648 3492 664 3508
rect 536 3472 552 3488
rect 424 3332 440 3348
rect 392 3312 408 3328
rect 360 3292 376 3308
rect 376 3292 392 3308
rect 488 3392 504 3408
rect 424 3132 440 3148
rect 456 3212 472 3228
rect 520 3252 536 3268
rect 648 3392 664 3408
rect 680 3352 696 3368
rect 664 3312 680 3328
rect 776 4312 792 4328
rect 808 4312 824 4328
rect 792 4292 808 4308
rect 808 4232 824 4248
rect 792 4212 808 4228
rect 792 4112 808 4128
rect 760 3992 776 4008
rect 776 3932 792 3948
rect 744 3892 760 3908
rect 888 4632 904 4648
rect 856 4572 872 4588
rect 872 4452 888 4468
rect 840 4432 872 4448
rect 1160 4672 1176 4688
rect 1016 4612 1032 4628
rect 1064 4592 1080 4608
rect 952 4572 968 4588
rect 1048 4572 1064 4588
rect 920 4552 936 4568
rect 920 4532 936 4548
rect 1224 4932 1240 4948
rect 1432 4912 1448 4928
rect 1288 4892 1304 4908
rect 1304 4892 1320 4908
rect 1352 4892 1368 4908
rect 1384 4892 1400 4908
rect 1320 4852 1336 4868
rect 1224 4832 1240 4848
rect 1304 4732 1320 4748
rect 1272 4692 1288 4708
rect 1240 4672 1256 4688
rect 1256 4672 1272 4688
rect 1192 4632 1208 4648
rect 1192 4572 1208 4588
rect 1224 4572 1240 4588
rect 1112 4552 1128 4568
rect 1128 4552 1144 4568
rect 1176 4552 1192 4568
rect 1336 4732 1352 4748
rect 1336 4692 1352 4708
rect 968 4532 984 4548
rect 1016 4532 1032 4548
rect 1080 4532 1096 4548
rect 1288 4532 1304 4548
rect 1304 4532 1320 4548
rect 1000 4512 1016 4528
rect 925 4402 961 4418
rect 968 4352 984 4368
rect 920 4292 936 4308
rect 984 4292 1000 4308
rect 824 4212 840 4228
rect 824 4112 840 4128
rect 872 4112 888 4128
rect 840 4092 856 4108
rect 744 3812 760 3828
rect 792 3572 808 3588
rect 776 3532 792 3548
rect 760 3512 776 3528
rect 728 3492 744 3508
rect 760 3452 776 3468
rect 712 3332 728 3348
rect 744 3332 760 3348
rect 584 3272 600 3288
rect 664 3292 680 3308
rect 696 3292 712 3308
rect 632 3232 648 3248
rect 728 3312 744 3328
rect 712 3252 728 3268
rect 728 3192 744 3208
rect 648 3152 680 3168
rect 472 3132 488 3148
rect 408 3112 424 3128
rect 440 3112 456 3128
rect 696 3112 712 3128
rect 360 3092 376 3108
rect 392 3092 408 3108
rect 536 3092 552 3108
rect 536 3052 552 3068
rect 408 2972 424 2988
rect 536 2972 552 2988
rect 440 2952 456 2968
rect 424 2932 440 2948
rect 344 2912 360 2928
rect 328 2752 344 2768
rect 360 2712 376 2728
rect 328 2672 344 2688
rect 344 2552 360 2568
rect 408 2892 424 2908
rect 376 2532 408 2548
rect 312 2492 328 2508
rect 360 2472 376 2488
rect 328 2432 344 2448
rect 312 2312 328 2328
rect 312 2132 328 2148
rect 360 2292 376 2308
rect 280 1932 296 1948
rect 328 1932 344 1948
rect 456 2912 472 2928
rect 440 2592 456 2608
rect 664 2952 680 2968
rect 872 3912 888 3928
rect 824 3892 840 3908
rect 1368 4832 1384 4848
rect 1384 4812 1400 4828
rect 1400 4732 1416 4748
rect 1384 4712 1400 4728
rect 1368 4692 1384 4708
rect 1400 4632 1416 4648
rect 1528 5292 1544 5308
rect 1496 5272 1512 5288
rect 1656 5352 1672 5368
rect 1640 5292 1656 5308
rect 1560 5212 1576 5228
rect 1544 5172 1560 5188
rect 1512 5092 1528 5108
rect 1560 5072 1576 5088
rect 1480 4952 1496 4968
rect 1464 4792 1480 4808
rect 1512 4972 1528 4988
rect 1512 4932 1528 4948
rect 1560 4932 1576 4948
rect 1640 4912 1656 4928
rect 1576 4892 1592 4908
rect 1592 4892 1608 4908
rect 1624 4872 1640 4888
rect 1560 4852 1592 4868
rect 1544 4792 1560 4808
rect 1528 4712 1544 4728
rect 1496 4692 1512 4708
rect 1512 4672 1528 4688
rect 1432 4612 1448 4628
rect 1384 4592 1400 4608
rect 1416 4592 1432 4608
rect 1384 4572 1400 4588
rect 1416 4552 1432 4568
rect 1448 4572 1464 4588
rect 1512 4532 1544 4548
rect 1432 4512 1448 4528
rect 1480 4512 1496 4528
rect 1608 4752 1624 4768
rect 1576 4712 1592 4728
rect 1608 4692 1624 4708
rect 1592 4652 1608 4668
rect 1624 4632 1640 4648
rect 1592 4592 1608 4608
rect 1624 4592 1640 4608
rect 1208 4492 1224 4508
rect 1256 4492 1272 4508
rect 1352 4492 1368 4508
rect 1464 4492 1480 4508
rect 1304 4392 1320 4408
rect 1192 4372 1208 4388
rect 1112 4352 1128 4368
rect 1048 4332 1064 4348
rect 1080 4312 1096 4328
rect 1144 4312 1160 4328
rect 1000 4252 1016 4268
rect 1096 4292 1112 4308
rect 1032 4212 1048 4228
rect 1016 4152 1032 4168
rect 920 4112 936 4128
rect 936 4092 952 4108
rect 925 4002 961 4018
rect 936 3932 952 3948
rect 968 3932 984 3948
rect 1032 3932 1048 3948
rect 1000 3912 1016 3928
rect 1048 3912 1064 3928
rect 1064 3892 1080 3908
rect 1064 3872 1080 3888
rect 920 3852 936 3868
rect 904 3832 920 3848
rect 840 3792 856 3808
rect 872 3792 888 3808
rect 856 3732 872 3748
rect 808 3532 824 3548
rect 808 3472 824 3488
rect 840 3472 856 3488
rect 888 3452 904 3468
rect 872 3392 888 3408
rect 824 3352 840 3368
rect 856 3352 872 3368
rect 1016 3852 1032 3868
rect 968 3812 1000 3828
rect 925 3602 961 3618
rect 904 3332 920 3348
rect 936 3332 952 3348
rect 920 3312 936 3328
rect 808 3272 824 3288
rect 792 3152 808 3168
rect 792 3132 808 3148
rect 712 2972 728 2988
rect 680 2912 696 2928
rect 584 2832 600 2848
rect 552 2732 568 2748
rect 472 2672 488 2688
rect 520 2672 536 2688
rect 504 2612 520 2628
rect 552 2592 568 2608
rect 456 2512 472 2528
rect 488 2512 504 2528
rect 536 2512 552 2528
rect 408 2372 424 2388
rect 408 2332 424 2348
rect 424 2292 440 2308
rect 392 2272 408 2288
rect 264 1892 280 1908
rect 376 1832 392 1848
rect 360 1812 376 1828
rect 216 1712 232 1728
rect 200 1692 216 1708
rect 248 1712 264 1728
rect 296 1712 312 1728
rect 344 1712 360 1728
rect 168 1672 184 1688
rect 152 1392 168 1408
rect 136 1352 152 1368
rect 104 1312 120 1328
rect 184 1332 200 1348
rect 168 1312 184 1328
rect 168 1292 184 1308
rect 120 1172 136 1188
rect 216 1492 232 1508
rect 328 1692 344 1708
rect 280 1672 296 1688
rect 296 1672 312 1688
rect 376 1738 392 1748
rect 376 1732 392 1738
rect 456 2132 472 2148
rect 456 2112 472 2128
rect 440 1972 456 1988
rect 568 2552 584 2568
rect 568 2272 584 2288
rect 536 2152 552 2168
rect 552 2112 568 2128
rect 632 2812 648 2828
rect 616 2706 632 2708
rect 616 2692 632 2706
rect 696 2852 712 2868
rect 680 2772 696 2788
rect 776 3072 792 3088
rect 904 3292 920 3308
rect 925 3202 961 3218
rect 872 3152 888 3168
rect 840 3112 856 3128
rect 808 3092 824 3108
rect 872 3092 888 3108
rect 1032 3572 1048 3588
rect 1016 3532 1032 3548
rect 1000 3512 1016 3528
rect 984 3392 1000 3408
rect 1016 3352 1032 3368
rect 1000 3332 1016 3348
rect 1064 3692 1080 3708
rect 1352 4372 1368 4388
rect 1448 4372 1464 4388
rect 1352 4332 1368 4348
rect 1272 4312 1288 4328
rect 1208 4292 1224 4308
rect 1432 4292 1448 4308
rect 1384 4272 1400 4288
rect 1176 4232 1192 4248
rect 1160 4212 1176 4228
rect 1160 4132 1176 4148
rect 1272 4132 1288 4148
rect 1208 4072 1224 4088
rect 1096 3972 1112 3988
rect 1144 3972 1160 3988
rect 1176 3952 1192 3968
rect 1160 3892 1176 3908
rect 1144 3872 1160 3888
rect 1192 3872 1208 3888
rect 1256 4112 1272 4128
rect 1336 4192 1352 4208
rect 1304 4152 1320 4168
rect 1352 4172 1368 4188
rect 1256 4032 1272 4048
rect 1240 3932 1256 3948
rect 1368 4152 1384 4168
rect 1400 4012 1416 4028
rect 1352 3972 1368 3988
rect 1720 5332 1736 5348
rect 1768 5252 1784 5268
rect 1752 5112 1768 5128
rect 1912 5512 1928 5528
rect 1832 5472 1848 5488
rect 1816 5314 1832 5328
rect 1816 5312 1832 5314
rect 2056 5506 2072 5508
rect 2056 5492 2072 5506
rect 2088 5472 2104 5488
rect 2008 5452 2024 5468
rect 1949 5402 1985 5418
rect 1928 5352 1944 5368
rect 1928 5332 1944 5348
rect 1896 5312 1912 5328
rect 1800 5212 1816 5228
rect 1864 5132 1880 5148
rect 1992 5272 2008 5288
rect 1944 5152 1960 5168
rect 1928 5132 1944 5148
rect 1848 5112 1860 5128
rect 1860 5112 1864 5128
rect 1912 5112 1928 5128
rect 2136 5492 2168 5508
rect 2264 5612 2280 5628
rect 2216 5512 2232 5528
rect 2232 5492 2248 5508
rect 2120 5412 2136 5428
rect 2200 5452 2216 5468
rect 2184 5432 2200 5448
rect 2136 5352 2152 5368
rect 2024 5332 2040 5348
rect 2008 5232 2024 5248
rect 1832 5092 1848 5108
rect 1992 5092 2008 5108
rect 1704 5012 1720 5028
rect 1816 5012 1832 5028
rect 1704 4932 1720 4948
rect 1656 4892 1672 4908
rect 1656 4812 1672 4828
rect 1784 4912 1800 4928
rect 1800 4872 1816 4888
rect 1736 4852 1752 4868
rect 1720 4772 1736 4788
rect 1704 4672 1720 4688
rect 1704 4652 1720 4668
rect 1752 4832 1768 4848
rect 1816 4772 1832 4788
rect 2200 5412 2216 5428
rect 2216 5332 2232 5348
rect 2184 5312 2200 5328
rect 2168 5292 2184 5308
rect 2040 5252 2072 5268
rect 2088 5252 2104 5268
rect 2024 5172 2040 5188
rect 2024 5032 2040 5048
rect 1949 5002 1985 5018
rect 1976 4932 1992 4948
rect 2168 5232 2184 5248
rect 2056 5092 2072 5108
rect 2168 5092 2184 5108
rect 2136 5052 2152 5068
rect 1992 4912 2008 4928
rect 1912 4752 1928 4768
rect 1848 4712 1864 4728
rect 1880 4712 1896 4728
rect 1944 4712 1960 4728
rect 2024 4892 2040 4908
rect 2072 4952 2088 4968
rect 2280 5472 2296 5488
rect 2296 5392 2312 5408
rect 2248 5312 2264 5328
rect 2280 5312 2296 5328
rect 2232 5292 2248 5308
rect 2280 5292 2296 5308
rect 2456 5512 2472 5528
rect 2472 5492 2488 5508
rect 2584 5506 2600 5508
rect 2584 5492 2600 5506
rect 2440 5472 2456 5488
rect 2328 5392 2344 5408
rect 2392 5392 2408 5408
rect 2328 5312 2344 5328
rect 2392 5312 2408 5328
rect 2232 5132 2248 5148
rect 2280 5112 2296 5128
rect 2296 5092 2312 5108
rect 2264 5072 2280 5088
rect 2280 5052 2296 5068
rect 2184 5032 2200 5048
rect 2264 5032 2280 5048
rect 2168 4932 2184 4948
rect 2152 4892 2168 4908
rect 2120 4872 2136 4888
rect 2216 4812 2232 4828
rect 1832 4692 1848 4708
rect 1928 4692 1944 4708
rect 2040 4692 2056 4708
rect 1752 4632 1768 4648
rect 1784 4632 1800 4648
rect 1720 4592 1736 4608
rect 1736 4572 1752 4588
rect 1768 4572 1784 4588
rect 1832 4672 1848 4688
rect 1816 4512 1832 4528
rect 1608 4472 1624 4488
rect 1640 4472 1656 4488
rect 1672 4472 1688 4488
rect 1608 4452 1624 4468
rect 1592 4352 1608 4368
rect 1480 4272 1496 4288
rect 1640 4272 1656 4288
rect 1624 4232 1640 4248
rect 1608 4192 1624 4208
rect 1592 4152 1608 4168
rect 1512 4132 1528 4148
rect 1464 4092 1480 4108
rect 1448 3992 1464 4008
rect 1352 3952 1368 3968
rect 1416 3952 1432 3968
rect 1400 3932 1416 3948
rect 1384 3912 1400 3928
rect 1336 3892 1352 3908
rect 1480 3912 1496 3928
rect 1416 3892 1432 3908
rect 1480 3892 1496 3908
rect 1464 3872 1480 3888
rect 1256 3852 1272 3868
rect 1432 3852 1448 3868
rect 1288 3832 1304 3848
rect 1416 3832 1432 3848
rect 1288 3792 1304 3808
rect 1400 3792 1416 3808
rect 1368 3732 1384 3748
rect 1208 3672 1224 3688
rect 1192 3552 1208 3568
rect 1112 3532 1128 3548
rect 1080 3512 1096 3528
rect 1096 3472 1112 3488
rect 1160 3472 1176 3488
rect 1160 3372 1176 3388
rect 1080 3352 1096 3368
rect 1064 3332 1080 3348
rect 1112 3332 1128 3348
rect 1160 3312 1176 3328
rect 1080 3292 1096 3308
rect 984 3272 1000 3288
rect 1048 3252 1064 3268
rect 1032 3092 1048 3108
rect 760 3012 776 3028
rect 728 2932 744 2948
rect 744 2852 760 2868
rect 680 2712 696 2728
rect 696 2612 712 2628
rect 744 2612 760 2628
rect 680 2552 712 2568
rect 600 2532 616 2548
rect 600 2232 616 2248
rect 776 2952 792 2968
rect 792 2892 808 2908
rect 792 2812 808 2828
rect 792 2772 808 2788
rect 792 2492 808 2508
rect 760 2472 776 2488
rect 744 2392 760 2408
rect 712 2352 728 2368
rect 744 2332 760 2348
rect 696 2312 728 2328
rect 712 2292 728 2308
rect 664 2272 680 2288
rect 632 2192 648 2208
rect 776 2172 792 2188
rect 504 2072 520 2088
rect 488 1872 504 1888
rect 600 2072 616 2088
rect 648 2072 664 2088
rect 552 1932 568 1948
rect 552 1912 568 1928
rect 536 1852 552 1868
rect 456 1832 472 1848
rect 536 1792 552 1808
rect 456 1772 472 1788
rect 424 1732 440 1748
rect 472 1732 488 1748
rect 472 1712 488 1728
rect 376 1692 392 1708
rect 408 1692 440 1708
rect 312 1652 328 1668
rect 344 1572 360 1588
rect 312 1492 328 1508
rect 328 1472 344 1488
rect 248 1452 264 1468
rect 232 1432 248 1448
rect 216 1312 232 1328
rect 264 1412 280 1428
rect 616 1872 632 1888
rect 584 1852 616 1868
rect 776 2112 792 2128
rect 680 2092 696 2108
rect 760 2092 776 2108
rect 664 1912 680 1928
rect 664 1872 680 1888
rect 568 1752 584 1768
rect 392 1652 424 1668
rect 408 1632 424 1648
rect 472 1652 488 1668
rect 376 1512 392 1528
rect 440 1512 456 1528
rect 456 1512 488 1528
rect 376 1492 392 1508
rect 408 1492 424 1508
rect 360 1372 376 1388
rect 344 1312 360 1328
rect 296 1292 312 1308
rect 328 1292 344 1308
rect 168 1192 184 1208
rect 88 1152 104 1168
rect 152 1152 184 1168
rect 232 1272 248 1288
rect 280 1272 296 1288
rect 360 1272 376 1288
rect 392 1472 408 1488
rect 392 1452 408 1468
rect 408 1332 424 1348
rect 472 1312 488 1328
rect 456 1292 472 1308
rect 584 1692 600 1708
rect 584 1652 600 1668
rect 568 1592 584 1608
rect 552 1532 568 1548
rect 696 1852 712 1868
rect 632 1832 648 1848
rect 728 1832 744 1848
rect 744 1812 760 1828
rect 824 3072 840 3088
rect 824 2952 840 2968
rect 872 2912 888 2928
rect 888 2792 904 2808
rect 824 2692 840 2708
rect 920 2992 936 3008
rect 968 2872 984 2888
rect 925 2802 961 2818
rect 1032 2912 1048 2928
rect 1016 2712 1032 2728
rect 904 2672 920 2688
rect 856 2572 872 2588
rect 840 2552 856 2568
rect 872 2532 888 2548
rect 1128 3292 1144 3308
rect 1096 3232 1112 3248
rect 1112 3132 1128 3148
rect 1064 2972 1080 2988
rect 1016 2632 1032 2648
rect 1048 2612 1064 2628
rect 968 2592 984 2608
rect 1048 2532 1064 2548
rect 920 2512 936 2528
rect 840 2492 856 2508
rect 904 2492 920 2508
rect 824 2372 856 2388
rect 808 2332 824 2348
rect 1080 2952 1096 2968
rect 1144 3112 1160 3128
rect 1144 3092 1160 3108
rect 1144 3052 1160 3068
rect 1336 3672 1352 3688
rect 1352 3652 1368 3668
rect 1352 3612 1368 3628
rect 1336 3512 1352 3528
rect 1304 3492 1320 3508
rect 1256 3452 1272 3468
rect 1256 3412 1272 3428
rect 1224 3392 1240 3408
rect 1208 3292 1224 3308
rect 1192 3272 1208 3288
rect 1384 3532 1400 3548
rect 1432 3772 1448 3788
rect 1528 4052 1544 4068
rect 1560 4012 1576 4028
rect 1592 4032 1608 4048
rect 1656 4152 1672 4168
rect 1768 4452 1784 4468
rect 1704 4432 1720 4448
rect 1784 4292 1800 4308
rect 1800 4292 1816 4308
rect 1816 4272 1832 4288
rect 1768 4252 1784 4268
rect 1672 4132 1688 4148
rect 1752 4132 1768 4148
rect 1704 4112 1720 4128
rect 1672 4092 1688 4108
rect 1656 4072 1672 4088
rect 1640 4052 1656 4068
rect 1512 3892 1528 3908
rect 1576 3892 1592 3908
rect 1592 3892 1608 3908
rect 1464 3752 1480 3768
rect 1448 3732 1464 3748
rect 1528 3732 1544 3748
rect 1592 3732 1608 3748
rect 1624 3732 1640 3748
rect 1560 3712 1576 3728
rect 1544 3652 1560 3668
rect 1496 3632 1512 3648
rect 1560 3632 1576 3648
rect 1432 3572 1448 3588
rect 1624 3692 1640 3708
rect 1688 4072 1704 4088
rect 1704 4072 1720 4088
rect 1704 4032 1720 4048
rect 1688 3772 1704 3788
rect 1800 4012 1816 4028
rect 1784 3932 1800 3948
rect 1800 3892 1816 3908
rect 1848 4652 1864 4668
rect 1896 4612 1912 4628
rect 1896 4572 1912 4588
rect 2008 4672 2024 4688
rect 1949 4602 1985 4618
rect 1896 4532 1912 4548
rect 1880 4512 1896 4528
rect 1928 4392 1944 4408
rect 1928 4352 1944 4368
rect 1912 4332 1928 4348
rect 1848 4292 1864 4308
rect 1880 4252 1896 4268
rect 1896 4232 1912 4248
rect 1864 4172 1880 4188
rect 1944 4252 1960 4268
rect 1949 4202 1985 4218
rect 1928 4132 1960 4148
rect 1832 3872 1848 3888
rect 1912 4092 1928 4108
rect 1864 4052 1880 4068
rect 1848 3792 1864 3808
rect 2008 4552 2024 4568
rect 2312 4912 2328 4928
rect 2248 4712 2264 4728
rect 2136 4706 2152 4708
rect 2136 4692 2152 4706
rect 2280 4692 2296 4708
rect 2152 4672 2168 4688
rect 2056 4492 2072 4508
rect 2024 4472 2040 4488
rect 2232 4572 2248 4588
rect 2408 5292 2424 5308
rect 2360 5092 2376 5108
rect 2392 5092 2408 5108
rect 2344 5072 2360 5088
rect 2504 5472 2520 5488
rect 2488 5392 2504 5408
rect 2632 5372 2648 5388
rect 2957 5602 2993 5618
rect 3016 5612 3032 5628
rect 3048 5612 3064 5628
rect 3176 5612 3192 5628
rect 3480 5512 3496 5528
rect 3624 5512 3628 5528
rect 3628 5512 3640 5528
rect 2808 5492 2824 5508
rect 2728 5472 2744 5488
rect 2488 5332 2504 5348
rect 2584 5332 2600 5348
rect 2568 5172 2584 5188
rect 2488 5072 2504 5088
rect 2472 5052 2488 5068
rect 2408 4972 2424 4988
rect 2392 4932 2408 4948
rect 2376 4892 2392 4908
rect 2392 4772 2408 4788
rect 2344 4712 2360 4728
rect 2360 4712 2364 4728
rect 2364 4712 2376 4728
rect 2376 4692 2392 4708
rect 2440 4952 2456 4968
rect 2536 4952 2552 4968
rect 2568 4932 2584 4948
rect 2392 4672 2408 4688
rect 2312 4572 2328 4588
rect 2296 4532 2312 4548
rect 2152 4512 2168 4528
rect 2264 4512 2280 4528
rect 2280 4512 2296 4528
rect 2232 4492 2248 4508
rect 2200 4472 2216 4488
rect 2104 4392 2120 4408
rect 2152 4392 2168 4408
rect 2104 4372 2120 4388
rect 2024 4312 2040 4328
rect 2120 4352 2136 4368
rect 2008 4272 2024 4288
rect 2088 4272 2104 4288
rect 2056 4232 2072 4248
rect 2008 4152 2024 4168
rect 2072 4152 2088 4168
rect 2040 4132 2056 4148
rect 2056 4112 2072 4128
rect 2008 4072 2024 4088
rect 1992 4052 2008 4068
rect 2008 4032 2024 4048
rect 1992 3932 2008 3948
rect 2088 3972 2104 3988
rect 2024 3912 2040 3928
rect 1960 3872 1992 3888
rect 2040 3872 2056 3888
rect 1992 3852 2008 3868
rect 1949 3802 1985 3818
rect 1880 3772 1912 3788
rect 1848 3752 1880 3768
rect 1720 3732 1736 3748
rect 1768 3732 1800 3748
rect 1816 3732 1832 3748
rect 1832 3732 1848 3748
rect 1656 3692 1672 3708
rect 1640 3652 1656 3668
rect 1576 3592 1592 3608
rect 1528 3472 1544 3488
rect 1496 3452 1512 3468
rect 1528 3412 1544 3428
rect 1256 3352 1272 3368
rect 1336 3352 1352 3368
rect 1240 3312 1256 3328
rect 1464 3312 1480 3328
rect 1256 3292 1272 3308
rect 1192 3112 1208 3128
rect 1176 3032 1192 3048
rect 1272 3272 1288 3288
rect 1224 3252 1240 3268
rect 1256 3232 1272 3248
rect 1464 3292 1480 3308
rect 1320 3252 1336 3268
rect 1448 3272 1464 3288
rect 1400 3252 1416 3268
rect 1432 3252 1448 3268
rect 1464 3252 1480 3268
rect 1368 3232 1384 3248
rect 1464 3232 1480 3248
rect 1352 3152 1368 3168
rect 1416 3152 1432 3168
rect 1320 3132 1336 3148
rect 1352 3132 1368 3148
rect 1272 3112 1288 3128
rect 1320 3112 1336 3128
rect 1256 3092 1272 3108
rect 1432 3092 1448 3108
rect 1240 3072 1256 3088
rect 1224 2992 1240 3008
rect 1304 3032 1320 3048
rect 1384 3032 1400 3048
rect 1256 2972 1272 2988
rect 1400 2972 1416 2988
rect 1336 2952 1352 2968
rect 1240 2932 1256 2948
rect 1272 2912 1288 2928
rect 1400 2914 1416 2928
rect 1400 2912 1416 2914
rect 1160 2892 1176 2908
rect 1208 2892 1224 2908
rect 1288 2852 1304 2868
rect 1240 2692 1256 2708
rect 1064 2512 1080 2528
rect 1032 2492 1048 2508
rect 1080 2472 1096 2488
rect 1000 2452 1016 2468
rect 1032 2452 1064 2468
rect 1016 2432 1032 2448
rect 925 2402 961 2418
rect 968 2412 984 2428
rect 856 2352 872 2368
rect 1064 2432 1080 2448
rect 1112 2392 1128 2408
rect 968 2332 984 2348
rect 984 2332 1000 2348
rect 984 2312 1000 2328
rect 1064 2292 1080 2308
rect 808 2192 824 2208
rect 1032 2272 1048 2288
rect 952 2232 968 2248
rect 984 2232 1000 2248
rect 872 2192 888 2208
rect 936 2172 952 2188
rect 824 2132 840 2148
rect 792 1912 808 1928
rect 888 2112 904 2128
rect 968 2172 984 2188
rect 1032 2132 1048 2148
rect 872 2032 888 2048
rect 952 2032 968 2048
rect 792 1832 808 1848
rect 776 1792 792 1808
rect 648 1752 664 1768
rect 840 1752 856 1768
rect 680 1712 696 1728
rect 744 1712 760 1728
rect 808 1712 824 1728
rect 925 2002 961 2018
rect 888 1912 904 1928
rect 872 1732 888 1748
rect 616 1692 632 1708
rect 632 1632 648 1648
rect 984 1972 1000 1988
rect 1032 1892 1048 1908
rect 1032 1732 1048 1748
rect 968 1672 984 1688
rect 1032 1672 1048 1688
rect 1048 1672 1064 1688
rect 1016 1652 1032 1668
rect 824 1612 840 1628
rect 925 1602 961 1618
rect 680 1572 696 1588
rect 584 1552 600 1568
rect 600 1532 616 1548
rect 1000 1532 1016 1548
rect 568 1492 584 1508
rect 552 1472 568 1488
rect 536 1392 552 1408
rect 552 1372 568 1388
rect 536 1312 552 1328
rect 440 1272 472 1288
rect 216 1252 232 1268
rect 360 1232 376 1248
rect 296 1152 312 1168
rect 440 1212 456 1228
rect 200 1132 216 1148
rect 232 1132 248 1148
rect 296 1132 312 1148
rect 424 1132 440 1148
rect 120 1112 136 1128
rect 200 1112 216 1128
rect 248 1112 264 1128
rect 360 1112 376 1128
rect 104 1092 120 1108
rect 88 1052 104 1068
rect 56 952 72 968
rect 88 672 104 688
rect 88 532 104 548
rect 216 1092 232 1108
rect 184 1072 200 1088
rect 232 1072 248 1088
rect 168 1052 184 1068
rect 280 1072 296 1088
rect 424 1092 440 1108
rect 392 1052 408 1068
rect 376 1032 392 1048
rect 264 952 280 968
rect 280 952 296 968
rect 152 932 168 948
rect 312 932 328 948
rect 424 1032 440 1048
rect 408 952 424 968
rect 232 912 248 928
rect 312 912 328 928
rect 376 912 392 928
rect 424 912 440 928
rect 216 892 232 908
rect 200 572 216 588
rect 248 872 264 888
rect 408 892 424 908
rect 504 1292 520 1308
rect 1128 2292 1144 2308
rect 1272 2572 1288 2588
rect 1192 2532 1208 2548
rect 1160 2352 1176 2368
rect 1144 2252 1160 2268
rect 1112 2172 1128 2188
rect 1096 2152 1112 2168
rect 1256 2492 1272 2508
rect 1496 3112 1512 3128
rect 1464 2952 1480 2968
rect 1624 3432 1640 3448
rect 1592 3352 1608 3368
rect 1640 3392 1656 3408
rect 1704 3712 1720 3728
rect 1736 3712 1752 3728
rect 1752 3712 1768 3728
rect 1752 3652 1768 3668
rect 1688 3492 1704 3508
rect 1672 3352 1688 3368
rect 1688 3352 1704 3368
rect 1608 3332 1624 3348
rect 1544 3312 1560 3328
rect 1592 3312 1608 3328
rect 1608 3252 1624 3268
rect 1640 3272 1656 3288
rect 1688 3272 1704 3288
rect 1800 3512 1816 3528
rect 1704 3232 1720 3248
rect 1528 3052 1544 3068
rect 1512 3032 1528 3048
rect 1624 3092 1640 3108
rect 1656 3112 1672 3128
rect 1640 3072 1656 3088
rect 1608 3052 1624 3068
rect 1576 3032 1592 3048
rect 1688 3092 1704 3108
rect 1672 3052 1688 3068
rect 1624 2912 1640 2928
rect 1592 2892 1608 2908
rect 1672 2892 1688 2908
rect 1496 2852 1512 2868
rect 1448 2792 1464 2808
rect 1528 2792 1544 2808
rect 1432 2772 1448 2788
rect 1496 2772 1512 2788
rect 1400 2692 1416 2708
rect 1368 2672 1384 2688
rect 1320 2652 1336 2668
rect 1480 2652 1496 2668
rect 1496 2632 1512 2648
rect 1400 2612 1416 2628
rect 1320 2592 1336 2608
rect 1384 2592 1400 2608
rect 1304 2552 1320 2568
rect 1368 2552 1384 2568
rect 1304 2532 1320 2548
rect 1192 2432 1208 2448
rect 1288 2432 1304 2448
rect 1256 2412 1272 2428
rect 1224 2332 1240 2348
rect 1240 2332 1256 2348
rect 1240 2312 1256 2328
rect 1304 2392 1320 2408
rect 1336 2432 1352 2448
rect 1176 2212 1192 2228
rect 1320 2312 1336 2328
rect 1256 2272 1272 2288
rect 1336 2272 1352 2288
rect 1368 2272 1384 2288
rect 1320 2252 1336 2268
rect 1288 2232 1304 2248
rect 1288 2132 1304 2148
rect 1192 2112 1208 2128
rect 1080 2092 1096 2108
rect 1208 2092 1224 2108
rect 1256 2072 1272 2088
rect 1128 1952 1144 1968
rect 1112 1832 1128 1848
rect 1112 1732 1128 1748
rect 1192 1852 1208 1868
rect 1240 1852 1256 1868
rect 1224 1812 1240 1828
rect 1192 1772 1208 1788
rect 1160 1652 1176 1668
rect 1144 1612 1160 1628
rect 1128 1552 1144 1568
rect 1160 1552 1176 1568
rect 712 1492 728 1508
rect 824 1492 840 1508
rect 952 1506 968 1508
rect 952 1492 968 1506
rect 1016 1492 1032 1508
rect 1144 1492 1160 1508
rect 984 1472 1000 1488
rect 616 1432 632 1448
rect 680 1432 696 1448
rect 584 1332 616 1348
rect 664 1332 680 1348
rect 648 1292 664 1308
rect 488 1272 504 1288
rect 472 1232 488 1248
rect 504 1212 520 1228
rect 552 1192 568 1208
rect 488 1132 504 1148
rect 504 1112 520 1128
rect 536 1132 552 1148
rect 568 1152 584 1168
rect 728 1312 744 1328
rect 712 1292 728 1308
rect 808 1312 824 1328
rect 1224 1752 1240 1768
rect 1368 2192 1384 2208
rect 1480 2552 1496 2568
rect 1464 2532 1480 2548
rect 1416 2512 1432 2528
rect 1400 2452 1416 2468
rect 1432 2272 1448 2288
rect 1464 2492 1480 2508
rect 1464 2452 1480 2468
rect 1448 2172 1464 2188
rect 1576 2712 1592 2728
rect 1544 2692 1560 2708
rect 1544 2512 1560 2528
rect 1816 3492 1832 3508
rect 1800 3332 1816 3348
rect 1832 3212 1848 3228
rect 1752 3192 1768 3208
rect 1736 3152 1752 3168
rect 1720 3112 1736 3128
rect 1720 3072 1736 3088
rect 1832 3132 1848 3148
rect 1784 3072 1800 3088
rect 1768 2932 1784 2948
rect 1784 2912 1800 2928
rect 1752 2832 1768 2848
rect 1704 2792 1720 2808
rect 1768 2772 1784 2788
rect 1720 2752 1736 2768
rect 1656 2692 1672 2708
rect 1800 2692 1816 2708
rect 1560 2492 1576 2508
rect 1672 2632 1688 2648
rect 1720 2632 1736 2648
rect 1640 2592 1672 2608
rect 1624 2492 1640 2508
rect 1528 2472 1544 2488
rect 1608 2472 1624 2488
rect 1512 2452 1528 2468
rect 1784 2592 1800 2608
rect 1704 2572 1720 2588
rect 1672 2512 1688 2528
rect 1688 2472 1704 2488
rect 1656 2412 1672 2428
rect 1592 2372 1624 2388
rect 1576 2352 1592 2368
rect 1496 2232 1512 2248
rect 1544 2232 1560 2248
rect 1352 2132 1368 2148
rect 1416 2132 1432 2148
rect 1464 2132 1480 2148
rect 1528 2132 1544 2148
rect 1416 2112 1432 2128
rect 1512 2112 1528 2128
rect 1560 2112 1576 2128
rect 1544 2092 1560 2108
rect 1512 1972 1528 1988
rect 1528 1932 1544 1948
rect 1272 1892 1288 1908
rect 1320 1892 1336 1908
rect 1384 1892 1400 1908
rect 1272 1872 1288 1888
rect 1480 1852 1496 1868
rect 1288 1832 1304 1848
rect 1416 1832 1432 1848
rect 1352 1812 1368 1828
rect 1384 1812 1400 1828
rect 1528 1812 1544 1828
rect 1336 1752 1352 1768
rect 1320 1732 1336 1748
rect 1240 1692 1256 1708
rect 1176 1452 1192 1468
rect 1096 1412 1112 1428
rect 1064 1372 1080 1388
rect 856 1352 872 1368
rect 824 1292 840 1308
rect 872 1332 888 1348
rect 1112 1352 1128 1368
rect 968 1332 984 1348
rect 1096 1332 1112 1348
rect 1160 1332 1176 1348
rect 936 1312 952 1328
rect 888 1292 904 1308
rect 760 1272 776 1288
rect 792 1272 808 1288
rect 888 1272 904 1288
rect 616 1252 648 1268
rect 840 1252 856 1268
rect 744 1212 760 1228
rect 728 1192 744 1208
rect 872 1212 888 1228
rect 776 1152 792 1168
rect 925 1202 961 1218
rect 1032 1312 1048 1328
rect 1096 1312 1112 1328
rect 1016 1292 1032 1308
rect 1128 1292 1144 1308
rect 1064 1272 1080 1288
rect 1320 1712 1336 1728
rect 1272 1692 1288 1708
rect 1288 1612 1304 1628
rect 1272 1572 1288 1588
rect 1256 1392 1272 1408
rect 1400 1772 1416 1788
rect 1432 1772 1448 1788
rect 1416 1712 1432 1728
rect 1512 1752 1528 1768
rect 1464 1732 1480 1748
rect 1496 1732 1512 1748
rect 1640 2312 1656 2328
rect 1608 2212 1624 2228
rect 1592 2172 1608 2188
rect 1608 2112 1624 2128
rect 1576 1992 1592 2008
rect 1560 1932 1576 1948
rect 1560 1912 1576 1928
rect 1464 1692 1484 1708
rect 1484 1692 1496 1708
rect 1480 1652 1496 1668
rect 1320 1512 1336 1528
rect 1352 1512 1368 1528
rect 1464 1512 1480 1528
rect 1256 1372 1272 1388
rect 1224 1352 1240 1368
rect 1192 1312 1208 1328
rect 1048 1172 1064 1188
rect 1176 1172 1192 1188
rect 1048 1152 1064 1168
rect 680 1132 696 1148
rect 984 1132 1000 1148
rect 1080 1132 1096 1148
rect 584 1112 600 1128
rect 616 1112 632 1128
rect 664 1112 680 1128
rect 792 1112 808 1128
rect 840 1112 856 1128
rect 520 1092 552 1108
rect 808 1092 824 1108
rect 904 1092 920 1108
rect 488 1072 504 1088
rect 616 1072 632 1088
rect 680 1072 696 1088
rect 760 1072 776 1088
rect 664 1052 680 1068
rect 536 932 552 948
rect 728 1052 744 1068
rect 488 912 504 928
rect 552 912 568 928
rect 600 912 616 928
rect 328 712 344 728
rect 392 712 408 728
rect 408 712 424 728
rect 248 692 264 708
rect 312 692 328 708
rect 392 692 408 708
rect 424 692 440 708
rect 248 672 264 688
rect 360 652 376 668
rect 360 572 376 588
rect 328 532 344 548
rect 504 692 520 708
rect 472 572 488 588
rect 440 532 472 548
rect 280 512 296 528
rect 104 412 120 428
rect 24 352 40 368
rect 40 332 56 348
rect 40 312 56 328
rect 104 312 120 328
rect 120 292 136 308
rect 104 272 120 288
rect 248 472 264 488
rect 168 392 184 408
rect 248 372 264 388
rect 184 352 200 368
rect 232 352 248 368
rect 152 332 168 348
rect 232 332 248 348
rect 200 292 216 308
rect 216 292 232 308
rect 168 272 184 288
rect 136 192 152 208
rect 56 152 72 168
rect 552 552 568 568
rect 504 532 520 548
rect 568 532 584 548
rect 488 512 504 528
rect 360 492 376 508
rect 312 452 328 468
rect 344 432 360 448
rect 296 352 312 368
rect 328 352 344 368
rect 296 332 312 348
rect 280 292 296 308
rect 696 812 712 828
rect 600 712 616 728
rect 648 612 664 628
rect 600 552 616 568
rect 664 552 680 568
rect 584 512 600 528
rect 552 492 568 508
rect 424 452 440 468
rect 440 452 456 468
rect 504 452 520 468
rect 456 432 472 448
rect 536 412 552 428
rect 488 372 504 388
rect 424 352 440 368
rect 440 332 456 348
rect 472 332 488 348
rect 360 312 376 328
rect 360 292 376 308
rect 328 272 344 288
rect 248 152 264 168
rect 264 152 280 168
rect 216 132 232 148
rect 312 132 328 148
rect 504 352 520 368
rect 536 332 552 348
rect 552 312 568 328
rect 680 512 696 528
rect 712 672 728 688
rect 696 492 712 508
rect 632 472 648 488
rect 696 452 712 468
rect 616 412 632 428
rect 600 372 616 388
rect 616 372 632 388
rect 680 352 696 368
rect 824 1052 840 1068
rect 904 992 920 1008
rect 872 912 888 928
rect 1144 1092 1160 1108
rect 1192 1092 1208 1108
rect 1240 1312 1256 1328
rect 1272 1272 1288 1288
rect 1240 1132 1256 1148
rect 1288 1192 1304 1208
rect 1336 1492 1352 1508
rect 1416 1472 1432 1488
rect 1336 1452 1352 1468
rect 1544 1712 1560 1728
rect 1560 1712 1576 1728
rect 1544 1672 1560 1688
rect 1512 1492 1528 1508
rect 1496 1372 1512 1388
rect 1528 1432 1544 1448
rect 1464 1312 1480 1328
rect 1320 1292 1336 1308
rect 1448 1252 1480 1268
rect 1352 1232 1368 1248
rect 1608 1772 1640 1788
rect 1592 1752 1608 1768
rect 1576 1612 1592 1628
rect 1560 1372 1576 1388
rect 1576 1352 1592 1368
rect 1544 1312 1560 1328
rect 1592 1312 1608 1328
rect 1736 2512 1752 2528
rect 1704 2352 1720 2368
rect 1688 2212 1704 2228
rect 1672 2132 1688 2148
rect 1688 2092 1704 2108
rect 1720 2052 1736 2068
rect 1656 2032 1672 2048
rect 1688 1912 1704 1928
rect 1672 1892 1688 1908
rect 1672 1852 1688 1868
rect 1656 1752 1672 1768
rect 1624 1712 1640 1728
rect 1656 1692 1672 1708
rect 1640 1632 1656 1648
rect 1640 1532 1656 1548
rect 1704 1812 1720 1828
rect 1752 2452 1768 2468
rect 1768 2432 1784 2448
rect 1752 2352 1768 2368
rect 1752 2272 1768 2288
rect 1832 2452 1848 2468
rect 1800 2332 1816 2348
rect 1800 2312 1816 2328
rect 1816 2292 1832 2308
rect 1768 2012 1784 2028
rect 1880 3732 1896 3748
rect 2072 3872 2088 3888
rect 2136 4192 2152 4208
rect 2120 3992 2136 4008
rect 2104 3932 2120 3948
rect 2200 4292 2216 4308
rect 2184 4272 2200 4288
rect 2168 4052 2184 4068
rect 2264 4292 2296 4308
rect 2248 4272 2264 4288
rect 2312 4272 2328 4288
rect 2472 4914 2488 4928
rect 2472 4912 2488 4914
rect 2440 4652 2456 4668
rect 2488 4672 2504 4688
rect 2472 4632 2488 4648
rect 2408 4532 2424 4548
rect 2536 4532 2552 4548
rect 2536 4492 2552 4508
rect 2632 5132 2648 5148
rect 2776 5292 2792 5308
rect 2728 5252 2744 5268
rect 3064 5492 3080 5508
rect 3112 5492 3128 5508
rect 2808 5272 2824 5288
rect 2632 5112 2648 5128
rect 2680 5112 2696 5128
rect 2616 5092 2632 5108
rect 2760 5112 2776 5128
rect 2664 5092 2696 5108
rect 2616 5072 2632 5088
rect 2632 4912 2648 4928
rect 2712 5032 2728 5048
rect 2744 5032 2760 5048
rect 2712 4952 2728 4968
rect 2744 4914 2760 4928
rect 2744 4912 2760 4914
rect 2616 4892 2632 4908
rect 2648 4892 2680 4908
rect 2760 4832 2776 4848
rect 2792 5112 2808 5128
rect 2840 5112 2856 5128
rect 2856 5092 2888 5108
rect 2792 5072 2808 5088
rect 2840 5072 2856 5088
rect 2840 5052 2856 5068
rect 2760 4732 2776 4748
rect 2632 4712 2648 4728
rect 2712 4712 2728 4728
rect 2616 4652 2632 4668
rect 2680 4612 2696 4628
rect 2632 4532 2648 4548
rect 2664 4512 2680 4528
rect 2536 4472 2552 4488
rect 2584 4472 2600 4488
rect 2456 4292 2472 4308
rect 2328 4172 2344 4188
rect 2360 4172 2376 4188
rect 2216 4132 2232 4148
rect 2280 4112 2296 4128
rect 2424 4112 2440 4128
rect 2200 4092 2216 4108
rect 2296 4092 2312 4108
rect 2392 4092 2408 4108
rect 2184 4032 2200 4048
rect 2248 4012 2264 4028
rect 2232 3952 2248 3968
rect 2104 3912 2120 3928
rect 2136 3912 2152 3928
rect 2168 3892 2184 3908
rect 2200 3906 2216 3908
rect 2200 3892 2216 3906
rect 2088 3792 2104 3808
rect 2120 3772 2136 3788
rect 2104 3752 2120 3768
rect 2168 3732 2184 3748
rect 2200 3712 2216 3728
rect 2120 3692 2136 3708
rect 2152 3692 2168 3708
rect 2056 3552 2072 3568
rect 1928 3512 1944 3528
rect 1912 3492 1928 3508
rect 1960 3492 1976 3508
rect 2024 3472 2040 3488
rect 2136 3512 2152 3528
rect 2296 3912 2312 3928
rect 2600 4432 2616 4448
rect 2824 4692 2840 4708
rect 2824 4672 2840 4688
rect 2888 4892 2904 4908
rect 3016 5332 3032 5348
rect 3096 5312 3112 5328
rect 3112 5272 3128 5288
rect 3016 5252 3032 5268
rect 2957 5202 2993 5218
rect 3080 5232 3096 5248
rect 3064 5112 3080 5128
rect 2888 4792 2920 4808
rect 3144 5132 3160 5148
rect 2984 4932 3000 4948
rect 3080 4932 3096 4948
rect 3064 4912 3080 4928
rect 3176 5472 3192 5488
rect 3592 5492 3608 5508
rect 3640 5492 3656 5508
rect 3752 5492 3768 5508
rect 3384 5472 3400 5488
rect 3560 5472 3576 5488
rect 3416 5432 3432 5448
rect 3240 5392 3256 5408
rect 3304 5332 3320 5348
rect 3336 5332 3352 5348
rect 3192 5192 3208 5208
rect 3208 5132 3224 5148
rect 3208 4932 3224 4948
rect 3160 4912 3176 4928
rect 3096 4892 3112 4908
rect 2957 4802 2993 4818
rect 2856 4712 2872 4728
rect 2968 4712 2984 4728
rect 3032 4712 3048 4728
rect 2856 4692 2872 4708
rect 2936 4692 2952 4708
rect 2952 4692 2968 4708
rect 2776 4652 2792 4668
rect 2840 4652 2856 4668
rect 2760 4572 2776 4588
rect 2920 4672 2936 4688
rect 2888 4592 2904 4608
rect 3096 4706 3112 4708
rect 3096 4692 3112 4706
rect 3096 4652 3112 4668
rect 3080 4612 3096 4628
rect 3064 4572 3080 4588
rect 3016 4552 3032 4568
rect 2744 4532 2760 4548
rect 2968 4532 2984 4548
rect 2712 4512 2728 4528
rect 2696 4492 2712 4508
rect 2808 4492 2824 4508
rect 3000 4472 3016 4488
rect 2824 4432 2840 4448
rect 2856 4392 2872 4408
rect 2920 4392 2936 4408
rect 2957 4402 2993 4418
rect 2904 4352 2920 4368
rect 2456 4132 2472 4148
rect 2584 4132 2600 4148
rect 2536 4114 2552 4128
rect 2536 4112 2552 4114
rect 2472 4092 2488 4108
rect 2440 3892 2456 3908
rect 2376 3792 2392 3808
rect 2424 3712 2440 3728
rect 2360 3652 2376 3668
rect 2312 3572 2328 3588
rect 2552 3932 2568 3948
rect 2536 3872 2552 3888
rect 2680 4132 2696 4148
rect 2648 4092 2664 4108
rect 2680 4092 2696 4108
rect 2584 3912 2600 3928
rect 2680 3912 2696 3928
rect 2648 3892 2664 3908
rect 2872 4192 2888 4208
rect 2760 4172 2776 4188
rect 2920 4172 2936 4188
rect 2728 4132 2744 4148
rect 2712 4112 2728 4128
rect 2824 4112 2840 4128
rect 2856 4112 2872 4128
rect 2696 3872 2712 3888
rect 2808 4092 2824 4108
rect 2872 4072 2888 4088
rect 2856 3972 2872 3988
rect 3048 4492 3064 4508
rect 2952 4292 2968 4308
rect 3032 4292 3048 4308
rect 3160 4892 3176 4908
rect 3160 4872 3176 4888
rect 3192 4772 3208 4788
rect 3128 4632 3144 4648
rect 3432 5312 3448 5328
rect 3272 5272 3288 5288
rect 3288 5072 3304 5088
rect 3432 5292 3448 5308
rect 3352 5272 3368 5288
rect 3416 5112 3432 5128
rect 3384 5092 3400 5108
rect 3432 5072 3448 5088
rect 3336 5052 3352 5068
rect 3544 5352 3560 5368
rect 3464 5312 3480 5328
rect 3720 5472 3736 5488
rect 3672 5372 3688 5388
rect 3720 5332 3736 5348
rect 3640 5312 3672 5328
rect 3624 5292 3640 5308
rect 3480 5252 3496 5268
rect 3496 5132 3512 5148
rect 3464 5112 3480 5128
rect 3448 4972 3464 4988
rect 3352 4952 3368 4968
rect 3272 4912 3288 4928
rect 3368 4752 3384 4768
rect 3240 4732 3256 4748
rect 3432 4912 3448 4928
rect 3480 5072 3496 5088
rect 3480 4952 3496 4968
rect 3464 4912 3480 4928
rect 3448 4872 3464 4888
rect 3400 4732 3416 4748
rect 3240 4712 3256 4728
rect 3432 4712 3448 4728
rect 3608 5192 3624 5208
rect 3560 5132 3576 5148
rect 3528 5092 3544 5108
rect 3640 5092 3656 5108
rect 3672 5192 3688 5208
rect 3768 5272 3784 5288
rect 3784 5232 3800 5248
rect 3832 5192 3848 5208
rect 3896 5472 3912 5488
rect 5021 5602 5057 5618
rect 7053 5602 7089 5618
rect 4568 5512 4584 5528
rect 4696 5512 4712 5528
rect 5048 5512 5064 5528
rect 5112 5512 5128 5528
rect 5176 5512 5192 5528
rect 6968 5512 6984 5528
rect 7144 5512 7160 5528
rect 7640 5512 7656 5528
rect 7736 5512 7752 5528
rect 3976 5472 3992 5488
rect 3997 5402 4033 5418
rect 4200 5492 4216 5508
rect 4680 5492 4696 5508
rect 4792 5492 4808 5508
rect 4904 5492 4920 5508
rect 5064 5492 5080 5508
rect 5208 5492 5224 5508
rect 4328 5472 4344 5488
rect 4152 5452 4168 5468
rect 4296 5432 4312 5448
rect 4056 5372 4072 5388
rect 4200 5372 4216 5388
rect 3944 5352 3960 5368
rect 4088 5352 4104 5368
rect 4168 5332 4184 5348
rect 4040 5292 4044 5308
rect 4044 5292 4056 5308
rect 3896 5272 3912 5288
rect 3832 5112 3848 5128
rect 3944 5132 3960 5148
rect 3688 5092 3704 5108
rect 3656 5072 3672 5088
rect 3512 4992 3528 5008
rect 3544 4992 3560 5008
rect 3528 4952 3544 4968
rect 3640 5052 3656 5068
rect 3560 4932 3576 4948
rect 3512 4912 3528 4928
rect 3496 4812 3512 4828
rect 3512 4732 3528 4748
rect 3272 4692 3288 4708
rect 3448 4692 3464 4708
rect 3464 4692 3480 4708
rect 3144 4612 3160 4628
rect 3208 4612 3224 4628
rect 3208 4552 3224 4568
rect 3160 4532 3176 4548
rect 3144 4512 3160 4528
rect 3224 4512 3240 4528
rect 3240 4512 3256 4528
rect 3160 4492 3176 4508
rect 3192 4492 3208 4508
rect 3176 4412 3192 4428
rect 3160 4392 3176 4408
rect 3144 4332 3160 4348
rect 3112 4312 3128 4328
rect 3048 4252 3064 4268
rect 2984 4092 3000 4108
rect 2957 4002 2993 4018
rect 2936 3952 2952 3968
rect 2776 3932 2792 3948
rect 2552 3812 2568 3828
rect 2456 3692 2504 3708
rect 2456 3572 2472 3588
rect 2136 3492 2152 3508
rect 2184 3492 2200 3508
rect 2248 3492 2264 3508
rect 1912 3452 1928 3468
rect 2024 3452 2040 3468
rect 2104 3452 2136 3468
rect 1949 3402 1985 3418
rect 1992 3412 2008 3428
rect 2184 3472 2200 3488
rect 2536 3512 2552 3528
rect 2152 3432 2168 3448
rect 2264 3432 2280 3448
rect 1896 3312 1912 3328
rect 1864 3092 1880 3108
rect 1976 3072 1992 3088
rect 1949 3002 1985 3018
rect 1912 2952 1928 2968
rect 2024 3272 2040 3288
rect 1912 2932 1928 2948
rect 1880 2912 1896 2928
rect 1912 2912 1928 2928
rect 1864 2892 1880 2908
rect 1992 2932 2008 2948
rect 2136 3292 2152 3308
rect 2056 3232 2072 3248
rect 2088 3152 2104 3168
rect 2104 3112 2120 3128
rect 2040 3092 2056 3108
rect 2120 3092 2136 3108
rect 2072 3052 2088 3068
rect 2072 2952 2088 2968
rect 2392 3432 2408 3448
rect 2392 3352 2408 3368
rect 2456 3352 2472 3368
rect 2264 3332 2280 3348
rect 2376 3332 2392 3348
rect 2184 3312 2200 3328
rect 2312 3312 2328 3328
rect 2296 3212 2312 3228
rect 2344 3212 2360 3228
rect 2376 3112 2392 3128
rect 2440 3292 2456 3308
rect 2664 3792 2680 3808
rect 2744 3792 2776 3808
rect 2808 3792 2824 3808
rect 2680 3752 2696 3768
rect 2600 3732 2616 3748
rect 2776 3732 2792 3748
rect 2792 3732 2808 3748
rect 2632 3712 2648 3728
rect 2568 3672 2584 3688
rect 2584 3632 2600 3648
rect 2616 3632 2632 3648
rect 2552 3452 2568 3468
rect 2600 3452 2616 3468
rect 2520 3392 2536 3408
rect 2488 3312 2504 3328
rect 2472 3292 2488 3308
rect 2456 3252 2472 3268
rect 2584 3272 2600 3288
rect 2664 3432 2680 3448
rect 2664 3412 2680 3428
rect 2696 3712 2712 3728
rect 2776 3712 2792 3728
rect 2792 3712 2808 3728
rect 2760 3692 2776 3708
rect 2728 3612 2744 3628
rect 2696 3452 2712 3468
rect 2712 3412 2728 3428
rect 2632 3212 2648 3228
rect 2568 3132 2584 3148
rect 2632 3132 2648 3148
rect 2296 3092 2312 3108
rect 2408 3092 2424 3108
rect 2456 3092 2472 3108
rect 2168 3072 2184 3088
rect 2408 3072 2424 3088
rect 2280 3052 2296 3068
rect 2152 2972 2168 2988
rect 2200 2992 2216 3008
rect 2168 2952 2184 2968
rect 2184 2952 2200 2968
rect 2376 3052 2392 3068
rect 2392 3052 2408 3068
rect 2344 3032 2360 3048
rect 2328 3012 2344 3028
rect 2216 2972 2232 2988
rect 2008 2912 2024 2928
rect 2040 2912 2056 2928
rect 2088 2912 2104 2928
rect 2136 2912 2152 2928
rect 1976 2872 1992 2888
rect 1960 2812 1976 2828
rect 2184 2872 2200 2888
rect 2120 2832 2136 2848
rect 2008 2772 2024 2788
rect 2072 2792 2088 2808
rect 2056 2732 2072 2748
rect 1864 2652 1880 2668
rect 2040 2632 2056 2648
rect 1864 2612 1880 2628
rect 1864 2552 1880 2568
rect 1912 2552 1928 2568
rect 1949 2602 1985 2618
rect 1944 2552 1960 2568
rect 1928 2532 1944 2548
rect 1992 2532 2024 2548
rect 1880 2512 1896 2528
rect 1928 2512 1944 2528
rect 1880 2432 1896 2448
rect 1896 2372 1912 2388
rect 1976 2312 1992 2328
rect 1880 2292 1912 2308
rect 1864 2272 1880 2288
rect 1832 2252 1848 2268
rect 1949 2202 1985 2218
rect 1912 2132 1928 2148
rect 1880 2114 1896 2128
rect 1880 2112 1896 2114
rect 2088 2752 2104 2768
rect 2200 2852 2216 2868
rect 2120 2732 2136 2748
rect 2152 2712 2168 2728
rect 2104 2692 2120 2708
rect 2120 2632 2136 2648
rect 2232 2952 2248 2968
rect 2472 3052 2488 3068
rect 2424 2952 2440 2968
rect 2504 3052 2520 3068
rect 2536 3032 2552 3048
rect 2488 2972 2504 2988
rect 2280 2852 2296 2868
rect 2328 2872 2344 2888
rect 2296 2732 2312 2748
rect 2296 2712 2312 2728
rect 2296 2692 2312 2708
rect 2216 2652 2232 2668
rect 2264 2652 2280 2668
rect 2312 2652 2328 2668
rect 2168 2612 2184 2628
rect 2152 2592 2168 2608
rect 2120 2552 2136 2568
rect 2088 2512 2104 2528
rect 2168 2512 2184 2528
rect 2200 2512 2216 2528
rect 2232 2592 2248 2608
rect 2232 2532 2248 2548
rect 2296 2532 2328 2548
rect 2312 2512 2328 2528
rect 2056 2492 2072 2508
rect 2184 2492 2200 2508
rect 2392 2672 2408 2688
rect 2344 2572 2360 2588
rect 2360 2552 2376 2568
rect 2392 2552 2408 2568
rect 2456 2872 2472 2888
rect 2632 3112 2648 3128
rect 2600 3032 2616 3048
rect 2584 3012 2600 3028
rect 2568 2832 2584 2848
rect 2680 3352 2696 3368
rect 2696 3332 2712 3348
rect 2936 3812 2952 3828
rect 2936 3772 2952 3788
rect 2856 3712 2872 3728
rect 2936 3712 2952 3728
rect 2824 3692 2840 3708
rect 2808 3612 2824 3628
rect 2957 3602 2993 3618
rect 2968 3552 2984 3568
rect 2792 3532 2808 3548
rect 2904 3532 2920 3548
rect 2776 3372 2792 3388
rect 2728 3352 2744 3368
rect 2808 3332 2824 3348
rect 2776 3292 2792 3308
rect 2808 3292 2824 3308
rect 2680 3132 2696 3148
rect 2776 3132 2792 3148
rect 2680 3112 2696 3128
rect 2664 3072 2680 3088
rect 2648 2992 2664 3008
rect 2616 2932 2632 2948
rect 2632 2912 2648 2928
rect 2600 2792 2616 2808
rect 2488 2712 2504 2728
rect 2632 2712 2648 2728
rect 2600 2692 2616 2708
rect 2648 2692 2664 2708
rect 2632 2672 2648 2688
rect 2472 2572 2488 2588
rect 2440 2552 2456 2568
rect 2504 2532 2520 2548
rect 2312 2472 2328 2488
rect 2008 2432 2024 2448
rect 2072 2432 2088 2448
rect 2264 2432 2280 2448
rect 2392 2432 2408 2448
rect 2056 2392 2072 2408
rect 2120 2392 2136 2408
rect 2008 2332 2024 2348
rect 2040 2312 2056 2328
rect 2488 2512 2504 2528
rect 2152 2332 2168 2348
rect 2248 2332 2264 2348
rect 2408 2332 2424 2348
rect 2280 2312 2296 2328
rect 2344 2312 2360 2328
rect 2552 2632 2568 2648
rect 2584 2652 2600 2668
rect 2568 2552 2584 2568
rect 2552 2512 2568 2528
rect 2664 2672 2680 2688
rect 2648 2552 2664 2568
rect 2632 2472 2648 2488
rect 2664 2452 2680 2468
rect 2760 3092 2776 3108
rect 2856 3512 2872 3528
rect 2840 3472 2856 3488
rect 2904 3512 2920 3528
rect 2920 3512 2936 3528
rect 2904 3472 2920 3488
rect 2888 3392 2904 3408
rect 2888 3352 2904 3368
rect 2984 3492 3000 3508
rect 2936 3292 2952 3308
rect 2824 3272 2840 3288
rect 2936 3272 2952 3288
rect 2888 3232 2904 3248
rect 2957 3202 2993 3218
rect 2888 3132 2904 3148
rect 2728 2932 2744 2948
rect 2712 2912 2728 2928
rect 2776 2872 2792 2888
rect 2760 2652 2776 2668
rect 2936 3092 2952 3108
rect 2888 3072 2904 3088
rect 2920 3072 2936 3088
rect 2808 3052 2824 3068
rect 2824 3032 2856 3048
rect 2920 2952 2936 2968
rect 2840 2932 2856 2948
rect 2888 2932 2904 2948
rect 2792 2732 2808 2748
rect 2824 2712 2840 2728
rect 2776 2632 2792 2648
rect 2728 2572 2744 2588
rect 2696 2552 2712 2568
rect 2776 2552 2792 2568
rect 3016 3932 3032 3948
rect 3016 3892 3032 3908
rect 3016 3752 3032 3768
rect 3064 4112 3080 4128
rect 3208 4452 3224 4468
rect 3096 4292 3112 4308
rect 3128 4292 3144 4308
rect 3160 4292 3176 4308
rect 3112 4192 3128 4208
rect 3096 4052 3112 4068
rect 3144 4172 3160 4188
rect 3256 4492 3272 4508
rect 3240 4132 3256 4148
rect 3176 4112 3192 4128
rect 3240 4112 3256 4128
rect 3160 4092 3176 4108
rect 3208 4092 3224 4108
rect 3256 4092 3272 4108
rect 3240 4072 3256 4088
rect 3256 4072 3272 4088
rect 3176 4052 3192 4068
rect 3192 4032 3208 4048
rect 3544 4712 3560 4728
rect 3368 4652 3384 4668
rect 3224 3932 3240 3948
rect 3272 3932 3288 3948
rect 3160 3912 3176 3928
rect 3464 4672 3480 4688
rect 3640 4932 3656 4948
rect 3688 4932 3704 4948
rect 3656 4912 3672 4928
rect 3624 4852 3640 4868
rect 3688 4872 3704 4888
rect 3832 4932 3864 4948
rect 3880 4932 3896 4948
rect 4184 5292 4200 5308
rect 4088 5272 4104 5288
rect 4072 5252 4088 5268
rect 4008 5112 4024 5128
rect 4088 5112 4104 5128
rect 4056 5092 4072 5108
rect 3997 5002 4033 5018
rect 3976 4932 3992 4948
rect 3864 4912 3880 4928
rect 3896 4912 3912 4928
rect 3944 4912 3960 4928
rect 3736 4892 3752 4908
rect 3656 4832 3672 4848
rect 3704 4832 3720 4848
rect 3688 4792 3704 4808
rect 3720 4792 3736 4808
rect 3848 4892 3864 4908
rect 3816 4872 3832 4888
rect 3800 4832 3816 4848
rect 3704 4752 3720 4768
rect 3752 4752 3768 4768
rect 3640 4712 3656 4728
rect 3752 4692 3768 4708
rect 3704 4672 3736 4688
rect 3768 4672 3784 4688
rect 3576 4652 3592 4668
rect 3400 4632 3416 4648
rect 3608 4632 3624 4648
rect 3672 4632 3688 4648
rect 3384 4612 3400 4628
rect 3608 4612 3624 4628
rect 3320 4552 3336 4568
rect 3368 4552 3384 4568
rect 3320 4492 3336 4508
rect 3352 4492 3368 4508
rect 3304 4392 3320 4408
rect 3304 4352 3320 4368
rect 3304 4252 3320 4268
rect 3320 4212 3336 4228
rect 3320 4172 3336 4188
rect 3304 4052 3320 4068
rect 3896 4852 3912 4868
rect 3832 4832 3848 4848
rect 3832 4812 3848 4828
rect 3864 4752 3880 4768
rect 3912 4832 3928 4848
rect 3944 4832 3960 4848
rect 3880 4732 3896 4748
rect 3896 4732 3912 4748
rect 3976 4812 3992 4828
rect 3928 4712 3944 4728
rect 4104 5072 4120 5088
rect 4120 5052 4136 5068
rect 4168 4972 4184 4988
rect 4104 4952 4120 4968
rect 4072 4912 4088 4928
rect 4088 4912 4104 4928
rect 4040 4832 4056 4848
rect 4072 4812 4088 4828
rect 4072 4792 4088 4808
rect 4264 5292 4280 5308
rect 4264 5112 4280 5128
rect 4648 5472 4664 5488
rect 4728 5472 4744 5488
rect 4744 5472 4760 5488
rect 4424 5452 4440 5468
rect 4552 5452 4568 5468
rect 4632 5352 4648 5368
rect 4408 5332 4424 5348
rect 4664 5332 4680 5348
rect 4408 5312 4424 5328
rect 4536 5312 4552 5328
rect 4344 5272 4360 5288
rect 4392 5272 4408 5288
rect 4456 5232 4472 5248
rect 4360 5192 4376 5208
rect 4344 5052 4360 5068
rect 4296 4932 4312 4948
rect 4248 4912 4264 4928
rect 4152 4772 4168 4788
rect 4280 4772 4296 4788
rect 4408 5112 4424 5128
rect 4376 5092 4392 5108
rect 4424 5092 4440 5108
rect 4440 5072 4456 5088
rect 4472 5172 4488 5188
rect 4536 5252 4552 5268
rect 4520 5092 4536 5108
rect 4504 5072 4520 5088
rect 4408 4912 4424 4928
rect 4392 4892 4408 4908
rect 4440 4892 4456 4908
rect 4488 4872 4504 4888
rect 3816 4652 3832 4668
rect 3848 4652 3864 4668
rect 3752 4612 3768 4628
rect 3768 4572 3784 4588
rect 3832 4572 3848 4588
rect 3432 4552 3448 4568
rect 3496 4552 3512 4568
rect 3752 4532 3768 4548
rect 3448 4492 3464 4508
rect 3400 4452 3416 4468
rect 3384 4392 3400 4408
rect 3368 4292 3384 4308
rect 3496 4472 3512 4488
rect 3448 4452 3464 4468
rect 3432 4392 3448 4408
rect 3480 4372 3496 4388
rect 3560 4492 3576 4508
rect 3512 4352 3528 4368
rect 3416 4332 3432 4348
rect 3496 4332 3512 4348
rect 3400 4192 3416 4208
rect 3368 4172 3384 4188
rect 3400 4132 3416 4148
rect 3400 4112 3416 4128
rect 3336 4032 3352 4048
rect 3368 3992 3384 4008
rect 3352 3972 3368 3988
rect 3288 3912 3304 3928
rect 3256 3892 3272 3908
rect 3368 3892 3384 3908
rect 3128 3872 3144 3888
rect 3192 3872 3208 3888
rect 3080 3852 3096 3868
rect 3032 3732 3048 3748
rect 3128 3732 3144 3748
rect 3032 3712 3048 3728
rect 3128 3712 3144 3728
rect 3160 3772 3176 3788
rect 3240 3752 3256 3768
rect 3192 3732 3208 3748
rect 3176 3712 3192 3728
rect 3224 3712 3240 3728
rect 3016 3692 3032 3708
rect 3048 3692 3060 3708
rect 3060 3692 3064 3708
rect 3064 3612 3080 3628
rect 3112 3692 3128 3708
rect 3208 3692 3224 3708
rect 3160 3672 3176 3688
rect 3176 3672 3192 3688
rect 3128 3612 3144 3628
rect 3112 3532 3128 3548
rect 3016 3512 3032 3528
rect 3032 3412 3048 3428
rect 3144 3512 3160 3528
rect 3080 3492 3096 3508
rect 3128 3492 3144 3508
rect 3064 3392 3080 3408
rect 3112 3412 3128 3428
rect 3064 3352 3080 3368
rect 3048 3312 3064 3328
rect 3048 3292 3064 3308
rect 3048 3252 3064 3268
rect 3064 3212 3080 3228
rect 3112 3212 3128 3228
rect 3272 3592 3288 3608
rect 3256 3552 3272 3568
rect 3224 3512 3240 3528
rect 3288 3512 3304 3528
rect 3272 3492 3288 3508
rect 3144 3272 3160 3288
rect 3160 3132 3176 3148
rect 3288 3472 3304 3488
rect 3192 3452 3208 3468
rect 3256 3432 3272 3448
rect 3336 3752 3352 3768
rect 3336 3592 3352 3608
rect 3432 4172 3448 4188
rect 3432 4112 3448 4128
rect 3432 4092 3448 4108
rect 3480 4272 3496 4288
rect 3528 4272 3544 4288
rect 3528 4212 3544 4228
rect 3800 4532 3816 4548
rect 3976 4672 3992 4688
rect 4024 4632 4040 4648
rect 3997 4602 4033 4618
rect 3928 4572 3944 4588
rect 3880 4532 3896 4548
rect 3816 4512 3832 4528
rect 3848 4512 3880 4528
rect 3768 4472 3784 4488
rect 3608 4372 3624 4388
rect 3736 4372 3752 4388
rect 3672 4332 3688 4348
rect 3480 4132 3512 4148
rect 3496 4112 3512 4128
rect 3544 4152 3560 4168
rect 3544 4092 3560 4108
rect 3560 4092 3576 4108
rect 3416 4072 3432 4088
rect 3448 4072 3464 4088
rect 3464 4072 3480 4088
rect 3496 4072 3512 4088
rect 3432 4052 3448 4068
rect 3464 4052 3480 4068
rect 3432 4012 3448 4028
rect 3368 3632 3384 3648
rect 3352 3572 3368 3588
rect 3480 3972 3496 3988
rect 3496 3972 3512 3988
rect 3544 3992 3560 4008
rect 3480 3932 3496 3948
rect 3544 3932 3560 3948
rect 3560 3932 3576 3948
rect 3448 3872 3464 3888
rect 3448 3752 3464 3768
rect 3400 3692 3416 3708
rect 3320 3532 3336 3548
rect 3336 3532 3352 3548
rect 3416 3532 3432 3548
rect 3320 3512 3336 3528
rect 3320 3452 3336 3468
rect 3352 3492 3368 3508
rect 3416 3452 3432 3468
rect 3384 3432 3400 3448
rect 3528 3912 3544 3928
rect 3608 4272 3624 4288
rect 3656 4272 3672 4288
rect 3640 4052 3656 4068
rect 3576 3912 3592 3928
rect 3528 3852 3544 3868
rect 3480 3692 3496 3708
rect 3512 3692 3528 3708
rect 3464 3632 3480 3648
rect 3496 3632 3512 3648
rect 3448 3572 3464 3588
rect 3496 3572 3512 3588
rect 3464 3532 3480 3548
rect 3656 3992 3672 4008
rect 3704 4272 3720 4288
rect 3688 4152 3704 4168
rect 3688 4112 3704 4128
rect 3752 4252 3768 4268
rect 3736 4112 3752 4128
rect 3752 4112 3768 4128
rect 3720 4072 3736 4088
rect 3720 4032 3736 4048
rect 3640 3972 3656 3988
rect 3672 3972 3688 3988
rect 3752 4012 3768 4028
rect 3816 4472 3832 4488
rect 3784 4332 3800 4348
rect 3832 4312 3848 4328
rect 3816 4292 3832 4308
rect 3832 4272 3848 4288
rect 3800 4252 3816 4268
rect 3784 4212 3800 4228
rect 3800 4092 3816 4108
rect 3848 4252 3864 4268
rect 3864 4232 3880 4248
rect 3976 4532 3992 4548
rect 4088 4712 4104 4728
rect 4104 4712 4120 4728
rect 4184 4752 4200 4768
rect 4232 4712 4248 4728
rect 4200 4692 4216 4708
rect 4408 4752 4424 4768
rect 4504 4752 4520 4768
rect 4312 4712 4328 4728
rect 4392 4712 4408 4728
rect 4264 4692 4280 4708
rect 4264 4672 4280 4688
rect 4344 4672 4360 4688
rect 4392 4672 4408 4688
rect 4136 4652 4152 4668
rect 4216 4652 4232 4668
rect 4264 4652 4280 4668
rect 4360 4652 4376 4668
rect 4200 4632 4216 4648
rect 4136 4612 4152 4628
rect 4120 4592 4136 4608
rect 3944 4512 3960 4528
rect 4040 4512 4056 4528
rect 4072 4512 4088 4528
rect 3992 4492 4008 4508
rect 4088 4492 4104 4508
rect 3928 4472 3944 4488
rect 3960 4452 3976 4468
rect 3928 4392 3944 4408
rect 4008 4412 4024 4428
rect 3912 4332 3928 4348
rect 3960 4332 3976 4348
rect 3944 4312 3960 4328
rect 3928 4292 3944 4308
rect 3928 4132 3944 4148
rect 3928 4092 3944 4108
rect 3928 4032 3944 4048
rect 3880 3972 3896 3988
rect 3864 3952 3880 3968
rect 3720 3932 3736 3948
rect 3784 3932 3800 3948
rect 3672 3912 3688 3928
rect 3608 3892 3624 3908
rect 3752 3892 3768 3908
rect 3768 3892 3784 3908
rect 3688 3872 3704 3888
rect 3544 3772 3560 3788
rect 3592 3772 3608 3788
rect 3624 3772 3640 3788
rect 3592 3752 3608 3768
rect 3656 3752 3672 3768
rect 3768 3752 3784 3768
rect 3976 4292 3992 4308
rect 3976 4252 3992 4268
rect 4120 4512 4136 4528
rect 4104 4232 4120 4248
rect 3997 4202 4033 4218
rect 3976 4172 3992 4188
rect 4504 4732 4520 4748
rect 4440 4712 4456 4728
rect 4456 4692 4472 4708
rect 4504 4692 4520 4708
rect 4424 4652 4440 4668
rect 4472 4632 4488 4648
rect 4184 4532 4200 4548
rect 4296 4532 4312 4548
rect 4488 4532 4504 4548
rect 4184 4412 4200 4428
rect 4248 4392 4264 4408
rect 4152 4272 4168 4288
rect 4232 4272 4248 4288
rect 4408 4514 4424 4528
rect 4408 4512 4424 4514
rect 4632 5132 4648 5148
rect 4616 5092 4648 5108
rect 4600 5072 4616 5088
rect 4776 5312 4792 5328
rect 4744 5292 4760 5308
rect 4712 5272 4728 5288
rect 4696 5152 4712 5168
rect 4664 5072 4680 5088
rect 4552 5032 4568 5048
rect 4568 4892 4584 4908
rect 4568 4872 4584 4888
rect 4632 5012 4648 5028
rect 4648 4932 4664 4948
rect 5368 5492 5384 5508
rect 5848 5506 5864 5508
rect 5848 5492 5864 5506
rect 5016 5472 5032 5488
rect 5128 5472 5144 5488
rect 5144 5472 5160 5488
rect 5176 5472 5192 5488
rect 5240 5472 5256 5488
rect 5272 5472 5288 5488
rect 5368 5472 5384 5488
rect 5448 5472 5464 5488
rect 5032 5372 5048 5388
rect 4888 5352 4904 5368
rect 4968 5332 4984 5348
rect 4984 5312 5000 5328
rect 5080 5312 5096 5328
rect 5112 5312 5128 5328
rect 4984 5292 5000 5308
rect 5032 5292 5048 5308
rect 4824 5192 4840 5208
rect 4792 5152 4808 5168
rect 4760 5112 4776 5128
rect 4872 5192 4888 5208
rect 4968 5152 4984 5168
rect 4888 5132 4904 5148
rect 4920 5112 4936 5128
rect 4760 5092 4776 5108
rect 4840 5092 4856 5108
rect 4872 5092 4888 5108
rect 4920 5092 4936 5108
rect 4712 5072 4728 5088
rect 4760 5072 4776 5088
rect 4712 5012 4728 5028
rect 4728 4972 4744 4988
rect 4840 5052 4856 5068
rect 4776 4972 4792 4988
rect 4856 4952 4872 4968
rect 4856 4932 4872 4948
rect 4920 5032 4936 5048
rect 4952 5092 4968 5108
rect 5021 5202 5057 5218
rect 5320 5372 5336 5388
rect 5240 5352 5256 5368
rect 5272 5332 5288 5348
rect 5384 5452 5400 5468
rect 5608 5452 5624 5468
rect 5848 5452 5864 5468
rect 5512 5372 5528 5388
rect 5592 5372 5608 5388
rect 5592 5352 5608 5368
rect 5416 5332 5432 5348
rect 5464 5332 5480 5348
rect 5496 5332 5512 5348
rect 5176 5312 5192 5328
rect 5224 5312 5240 5328
rect 5256 5292 5272 5308
rect 5304 5292 5320 5308
rect 5192 5272 5208 5288
rect 5160 5252 5176 5268
rect 5128 5092 5144 5108
rect 4936 5012 4952 5028
rect 5144 5032 5160 5048
rect 5000 4972 5016 4988
rect 5208 5032 5224 5048
rect 4984 4952 5000 4968
rect 4904 4932 4920 4948
rect 5096 4932 5112 4948
rect 4824 4912 4840 4928
rect 4952 4912 4968 4928
rect 4632 4872 4648 4888
rect 4552 4692 4568 4708
rect 4568 4612 4584 4628
rect 4632 4572 4648 4588
rect 4536 4512 4552 4528
rect 4520 4492 4536 4508
rect 4568 4492 4584 4508
rect 4312 4312 4328 4328
rect 4312 4252 4328 4268
rect 4168 4232 4184 4248
rect 4104 4192 4120 4208
rect 4040 4152 4056 4168
rect 4040 4112 4056 4128
rect 3992 4092 4008 4108
rect 3960 3972 3976 3988
rect 3896 3912 3912 3928
rect 3928 3912 3944 3928
rect 3832 3892 3848 3908
rect 3912 3892 3928 3908
rect 3832 3872 3848 3888
rect 4072 3992 4088 4008
rect 3960 3892 3976 3908
rect 4040 3892 4056 3908
rect 3944 3852 3960 3868
rect 4024 3852 4040 3868
rect 3960 3832 3976 3848
rect 3928 3792 3944 3808
rect 3997 3802 4033 3818
rect 4056 3852 4072 3868
rect 3912 3772 3928 3788
rect 4040 3732 4056 3748
rect 3720 3712 3736 3728
rect 3864 3712 3880 3728
rect 3656 3692 3672 3708
rect 3512 3552 3544 3568
rect 3496 3512 3512 3528
rect 3480 3492 3496 3508
rect 3528 3492 3544 3508
rect 3576 3512 3592 3528
rect 3544 3472 3560 3488
rect 3608 3472 3624 3488
rect 3592 3452 3608 3468
rect 3432 3412 3448 3428
rect 3640 3412 3656 3428
rect 3336 3392 3352 3408
rect 3528 3372 3544 3388
rect 3320 3352 3336 3368
rect 3432 3352 3448 3368
rect 3304 3332 3320 3348
rect 3416 3332 3432 3348
rect 3352 3312 3368 3328
rect 3384 3292 3388 3308
rect 3388 3292 3400 3308
rect 3352 3272 3368 3288
rect 3288 3232 3304 3248
rect 3176 3112 3192 3128
rect 3224 3112 3240 3128
rect 3000 3072 3032 3088
rect 3080 3072 3096 3088
rect 3336 3072 3352 3088
rect 3112 3052 3128 3068
rect 2968 2992 3000 3008
rect 3048 2952 3064 2968
rect 3000 2892 3016 2908
rect 3208 3032 3224 3048
rect 3400 3112 3416 3128
rect 3352 2952 3368 2968
rect 3064 2932 3080 2948
rect 3192 2932 3208 2948
rect 3432 3312 3448 3328
rect 3496 3192 3512 3208
rect 3432 3092 3448 3108
rect 3512 3072 3528 3088
rect 3432 2992 3448 3008
rect 3448 2952 3464 2968
rect 3368 2932 3384 2948
rect 3416 2932 3432 2948
rect 3448 2932 3464 2948
rect 3544 3292 3560 3308
rect 3544 3092 3560 3108
rect 3560 3072 3576 3088
rect 3576 3052 3592 3068
rect 3560 2992 3576 3008
rect 3624 3252 3640 3268
rect 3688 3692 3704 3708
rect 3736 3692 3752 3708
rect 3976 3692 3992 3708
rect 3896 3672 3912 3688
rect 3736 3652 3752 3668
rect 3688 3512 3704 3528
rect 3832 3632 3848 3648
rect 3912 3572 3928 3588
rect 3848 3532 3864 3548
rect 3848 3492 3864 3508
rect 3800 3472 3816 3488
rect 3736 3312 3752 3328
rect 3656 3292 3672 3308
rect 3752 3192 3768 3208
rect 3672 3092 3688 3108
rect 3736 3092 3752 3108
rect 3784 3312 3800 3328
rect 3880 3472 3896 3488
rect 3997 3402 4033 3418
rect 3992 3332 4008 3348
rect 3816 3312 3832 3328
rect 3912 3312 3928 3328
rect 3848 3272 3864 3288
rect 3800 3252 3816 3268
rect 3784 3232 3800 3248
rect 3816 3132 3832 3148
rect 3768 3072 3784 3088
rect 3768 3052 3784 3068
rect 3656 3032 3672 3048
rect 3800 2992 3816 3008
rect 3832 3112 3848 3128
rect 3912 3092 3928 3108
rect 3944 3092 3960 3108
rect 3976 3112 3992 3128
rect 4232 4212 4248 4228
rect 4200 4152 4216 4168
rect 4344 4212 4360 4228
rect 4504 4272 4520 4288
rect 4472 4232 4488 4248
rect 4376 4192 4392 4208
rect 4264 4172 4280 4188
rect 4376 4172 4392 4188
rect 4392 4152 4408 4168
rect 4248 4132 4264 4148
rect 4440 4132 4456 4148
rect 4136 4032 4152 4048
rect 4088 3792 4104 3808
rect 4104 3752 4120 3768
rect 4232 4112 4248 4128
rect 4200 3932 4216 3948
rect 4168 3912 4184 3928
rect 4184 3872 4200 3888
rect 4168 3852 4184 3868
rect 4136 3732 4152 3748
rect 4152 3732 4168 3748
rect 4072 3712 4088 3728
rect 4136 3692 4152 3708
rect 4104 3512 4120 3528
rect 4104 3492 4120 3508
rect 4152 3492 4168 3508
rect 4136 3472 4152 3488
rect 4136 3452 4152 3468
rect 4104 3252 4120 3268
rect 4056 3152 4072 3168
rect 4040 3092 4056 3108
rect 3864 3072 3880 3088
rect 3960 3072 3976 3088
rect 3816 2952 3848 2968
rect 3544 2932 3560 2948
rect 3736 2932 3752 2948
rect 3192 2912 3208 2928
rect 3256 2914 3272 2928
rect 3256 2912 3272 2914
rect 3336 2912 3352 2928
rect 3112 2892 3128 2908
rect 3320 2892 3336 2908
rect 2952 2832 2968 2848
rect 2957 2802 2993 2818
rect 3064 2872 3080 2888
rect 3304 2872 3320 2888
rect 3000 2712 3004 2728
rect 3004 2712 3016 2728
rect 2936 2692 2952 2708
rect 3016 2692 3032 2708
rect 3032 2672 3048 2688
rect 2904 2652 2920 2668
rect 3032 2652 3048 2668
rect 3144 2772 3160 2788
rect 3336 2752 3352 2768
rect 3080 2672 3096 2688
rect 3144 2672 3160 2688
rect 3064 2632 3080 2648
rect 3112 2632 3128 2648
rect 2936 2572 2952 2588
rect 2888 2552 2904 2568
rect 3064 2532 3080 2548
rect 2760 2512 2776 2528
rect 2872 2514 2888 2528
rect 2872 2512 2888 2514
rect 2936 2512 2952 2528
rect 3032 2492 3048 2508
rect 2792 2472 2808 2488
rect 2744 2452 2760 2468
rect 2712 2352 2728 2368
rect 2936 2432 2952 2448
rect 2792 2412 2808 2428
rect 2104 2292 2120 2308
rect 2312 2292 2328 2308
rect 2472 2292 2488 2308
rect 2376 2272 2392 2288
rect 2552 2272 2568 2288
rect 2056 2252 2072 2268
rect 2056 2192 2072 2208
rect 2184 2172 2200 2188
rect 2168 2132 2184 2148
rect 2008 2112 2024 2128
rect 1976 2092 1992 2108
rect 1848 2072 1864 2088
rect 1784 1992 1800 2008
rect 2024 2092 2040 2108
rect 1992 1952 2008 1968
rect 1752 1912 1768 1928
rect 1864 1912 1880 1928
rect 1768 1892 1784 1908
rect 1784 1892 1800 1908
rect 1736 1872 1752 1888
rect 1688 1712 1704 1728
rect 1736 1532 1752 1548
rect 1704 1512 1736 1528
rect 1624 1472 1640 1488
rect 1576 1292 1592 1308
rect 1608 1292 1624 1308
rect 1528 1212 1544 1228
rect 1512 1192 1528 1208
rect 1384 1172 1400 1188
rect 1464 1172 1480 1188
rect 1528 1172 1544 1188
rect 1320 1092 1336 1108
rect 968 1072 984 1088
rect 1032 1072 1048 1088
rect 1208 1072 1224 1088
rect 1256 1072 1272 1088
rect 1192 1032 1208 1048
rect 1176 972 1192 988
rect 1144 952 1160 968
rect 1224 952 1240 968
rect 1256 952 1272 968
rect 1192 932 1208 948
rect 984 912 1000 928
rect 984 892 1000 908
rect 925 802 961 818
rect 920 752 936 768
rect 760 672 776 688
rect 808 672 824 688
rect 888 672 904 688
rect 824 652 840 668
rect 792 632 808 648
rect 744 612 760 628
rect 728 512 744 528
rect 792 514 808 528
rect 792 512 808 514
rect 776 412 792 428
rect 408 292 424 308
rect 600 292 616 308
rect 680 292 696 308
rect 712 292 728 308
rect 504 192 520 208
rect 376 152 392 168
rect 440 132 456 148
rect 472 132 488 148
rect 152 114 168 128
rect 152 112 168 114
rect 248 112 264 128
rect 424 112 440 128
rect 536 114 552 128
rect 536 112 552 114
rect 664 272 680 288
rect 664 212 680 228
rect 600 152 616 168
rect 760 252 776 268
rect 1000 752 1016 768
rect 968 732 984 748
rect 952 672 968 688
rect 920 632 936 648
rect 840 612 856 628
rect 856 512 872 528
rect 840 412 856 428
rect 824 392 840 408
rect 888 392 904 408
rect 925 402 961 418
rect 872 252 888 268
rect 856 152 872 168
rect 984 692 1000 708
rect 1000 692 1016 708
rect 968 332 984 348
rect 1208 892 1224 908
rect 1064 872 1080 888
rect 1144 812 1160 828
rect 1048 732 1064 748
rect 1064 732 1080 748
rect 1032 692 1048 708
rect 1016 672 1032 688
rect 1032 652 1048 668
rect 1032 514 1048 528
rect 1032 512 1048 514
rect 1064 712 1080 728
rect 1096 692 1112 708
rect 1128 692 1144 708
rect 1160 732 1176 748
rect 1336 952 1352 968
rect 1416 1092 1432 1108
rect 1496 1132 1512 1148
rect 1560 1152 1576 1168
rect 1576 1112 1592 1128
rect 1576 1092 1592 1108
rect 1448 1072 1464 1088
rect 1464 1052 1480 1068
rect 1512 1052 1528 1068
rect 1448 1032 1464 1048
rect 1448 1012 1464 1028
rect 1400 952 1416 968
rect 1272 932 1288 948
rect 1288 932 1304 948
rect 1320 932 1336 948
rect 1352 932 1368 948
rect 1240 912 1256 928
rect 1304 892 1320 908
rect 1336 872 1352 888
rect 1240 772 1256 788
rect 1320 732 1336 748
rect 1192 692 1208 708
rect 1256 712 1272 728
rect 1080 672 1096 688
rect 1064 612 1080 628
rect 1160 632 1176 648
rect 1240 632 1272 648
rect 1208 592 1224 608
rect 1096 572 1112 588
rect 1256 552 1272 568
rect 1160 492 1176 508
rect 1144 472 1160 488
rect 1048 372 1064 388
rect 1048 352 1064 368
rect 1032 332 1048 348
rect 1096 332 1112 348
rect 1032 312 1048 328
rect 1000 292 1016 308
rect 952 272 968 288
rect 920 232 936 248
rect 968 232 984 248
rect 1000 152 1016 168
rect 888 132 904 148
rect 1048 292 1064 308
rect 1064 252 1080 268
rect 1112 172 1128 188
rect 1080 132 1096 148
rect 1240 432 1272 448
rect 1160 372 1176 388
rect 1176 312 1192 328
rect 1224 312 1240 328
rect 1304 652 1320 668
rect 1288 432 1304 448
rect 1384 812 1400 828
rect 1432 912 1448 928
rect 1416 892 1432 908
rect 1368 712 1372 728
rect 1372 712 1384 728
rect 1400 712 1416 728
rect 1368 552 1384 568
rect 1336 512 1352 528
rect 1304 332 1320 348
rect 1320 332 1336 348
rect 1352 292 1368 308
rect 1400 672 1416 688
rect 1416 672 1432 688
rect 1416 552 1432 568
rect 1400 512 1416 528
rect 1496 892 1512 908
rect 1560 872 1576 888
rect 1672 1452 1688 1468
rect 1656 1412 1672 1428
rect 1736 1432 1752 1448
rect 1672 1352 1688 1368
rect 1720 1312 1736 1328
rect 1640 1272 1656 1288
rect 1624 1092 1640 1108
rect 1672 1192 1688 1208
rect 1736 1192 1752 1208
rect 1720 1172 1736 1188
rect 2104 1892 2120 1908
rect 2040 1872 2056 1888
rect 2088 1872 2104 1888
rect 1832 1852 1848 1868
rect 1832 1812 1848 1828
rect 1784 1792 1800 1808
rect 1949 1802 1985 1818
rect 2008 1772 2024 1788
rect 1928 1752 1944 1768
rect 1832 1712 1848 1728
rect 1928 1712 1944 1728
rect 1896 1692 1912 1708
rect 1816 1672 1832 1688
rect 1880 1672 1896 1688
rect 1912 1672 1928 1688
rect 1784 1532 1800 1548
rect 1832 1632 1848 1648
rect 1848 1512 1864 1528
rect 1832 1452 1848 1468
rect 1800 1432 1816 1448
rect 1832 1432 1848 1448
rect 1784 1332 1800 1348
rect 1832 1312 1848 1328
rect 1832 1252 1848 1268
rect 2056 1772 2072 1788
rect 2072 1712 2088 1728
rect 1976 1692 1992 1708
rect 1880 1512 1896 1528
rect 1880 1472 1896 1488
rect 1896 1452 1912 1468
rect 1880 1312 1896 1328
rect 1864 1292 1880 1308
rect 2072 1592 2088 1608
rect 1992 1552 2008 1568
rect 1944 1532 1960 1548
rect 2056 1512 2072 1528
rect 1992 1432 2008 1448
rect 1949 1402 1985 1418
rect 2008 1412 2024 1428
rect 2424 2252 2440 2268
rect 2424 2232 2440 2248
rect 2552 2232 2568 2248
rect 2296 2192 2312 2208
rect 2216 2152 2232 2168
rect 2264 2152 2280 2168
rect 2200 2132 2216 2148
rect 2216 2112 2232 2128
rect 2328 2112 2344 2128
rect 2280 2072 2296 2088
rect 2184 1972 2200 1988
rect 2328 2092 2344 2108
rect 2344 2092 2360 2108
rect 2312 1992 2328 2008
rect 2344 1992 2360 2008
rect 2632 2212 2648 2228
rect 2456 2132 2472 2148
rect 2488 2112 2504 2128
rect 2536 2112 2552 2128
rect 2408 2092 2424 2108
rect 2488 2092 2504 2108
rect 2552 2092 2568 2108
rect 2568 2012 2584 2028
rect 2360 1872 2392 1888
rect 2424 1872 2440 1888
rect 2472 1872 2488 1888
rect 2248 1772 2264 1788
rect 2264 1752 2280 1768
rect 2136 1732 2152 1748
rect 2168 1712 2184 1728
rect 2136 1692 2152 1708
rect 2184 1612 2200 1628
rect 2104 1572 2120 1588
rect 2120 1532 2152 1548
rect 2088 1512 2104 1528
rect 2104 1492 2120 1508
rect 2120 1432 2136 1448
rect 2072 1392 2088 1408
rect 1928 1352 1944 1368
rect 2104 1352 2120 1368
rect 1928 1312 1944 1328
rect 1912 1292 1928 1308
rect 1944 1272 1960 1288
rect 2040 1272 2056 1288
rect 1784 1172 1800 1188
rect 1768 1092 1784 1108
rect 1848 1192 1864 1208
rect 1816 1112 1832 1128
rect 1896 1092 1912 1108
rect 1688 1072 1704 1088
rect 1800 1072 1816 1088
rect 1848 1072 1864 1088
rect 1720 1052 1736 1068
rect 1880 1032 1896 1048
rect 1784 932 1800 948
rect 1688 912 1704 928
rect 1816 912 1832 928
rect 1880 914 1896 928
rect 1880 912 1896 914
rect 1928 1252 1944 1268
rect 2152 1512 2168 1528
rect 2232 1552 2248 1568
rect 1928 1212 1944 1228
rect 2088 1212 2104 1228
rect 2040 1192 2056 1208
rect 1949 1002 1985 1018
rect 1608 732 1624 748
rect 2184 1472 2200 1488
rect 2200 1452 2216 1468
rect 2296 1692 2312 1708
rect 2344 1692 2360 1708
rect 2312 1552 2328 1568
rect 2312 1492 2328 1508
rect 2344 1472 2360 1488
rect 2280 1452 2296 1468
rect 2248 1432 2264 1448
rect 2168 1372 2184 1388
rect 2264 1352 2280 1368
rect 2232 1332 2248 1348
rect 2200 1312 2216 1328
rect 2152 1172 2168 1188
rect 2120 1072 2136 1088
rect 2136 1052 2152 1068
rect 2312 1432 2328 1448
rect 2376 1752 2392 1768
rect 2440 1732 2456 1748
rect 2504 1692 2520 1708
rect 2376 1632 2392 1648
rect 2392 1552 2408 1568
rect 2504 1552 2520 1568
rect 2424 1532 2440 1548
rect 2424 1512 2440 1528
rect 2472 1492 2488 1508
rect 2392 1452 2408 1468
rect 2440 1452 2456 1468
rect 2376 1352 2392 1368
rect 2360 1332 2376 1348
rect 2280 1312 2296 1328
rect 2312 1312 2328 1328
rect 2488 1312 2504 1328
rect 2264 1292 2280 1308
rect 2328 1292 2344 1308
rect 2232 1132 2248 1148
rect 2536 1712 2552 1728
rect 2552 1692 2568 1708
rect 2632 1692 2648 1708
rect 2536 1492 2552 1508
rect 2536 1472 2552 1488
rect 2712 2192 2728 2208
rect 2680 2112 2696 2128
rect 2680 2092 2696 2108
rect 2680 2072 2696 2088
rect 2872 2272 2888 2288
rect 2776 2192 2792 2208
rect 2957 2402 2993 2418
rect 3048 2472 3064 2488
rect 3032 2312 3048 2328
rect 2984 2272 3000 2288
rect 3080 2332 3096 2348
rect 3048 2292 3064 2308
rect 3064 2212 3080 2228
rect 3032 2152 3048 2168
rect 2760 2132 2776 2148
rect 2872 2132 2904 2148
rect 2792 2112 2808 2128
rect 2824 2112 2840 2128
rect 2808 2092 2820 2108
rect 2820 2092 2824 2108
rect 2856 1972 2872 1988
rect 3048 2112 3064 2128
rect 2984 2092 3000 2108
rect 2957 2002 2993 2018
rect 2936 1952 2952 1968
rect 2968 1952 2984 1968
rect 2776 1872 2792 1888
rect 2840 1872 2856 1888
rect 2728 1712 2744 1728
rect 2664 1552 2680 1568
rect 2648 1472 2664 1488
rect 2584 1332 2600 1348
rect 2504 1292 2520 1308
rect 2488 1252 2504 1268
rect 2344 1152 2360 1168
rect 2264 1112 2280 1128
rect 2392 1112 2408 1128
rect 2456 1112 2472 1128
rect 2296 1092 2312 1108
rect 2312 1092 2328 1108
rect 2360 1092 2376 1108
rect 2568 1292 2584 1308
rect 2568 1272 2584 1288
rect 2360 1072 2376 1088
rect 2424 1072 2440 1088
rect 2168 972 2184 988
rect 2296 1052 2312 1068
rect 2296 1012 2312 1028
rect 2232 992 2248 1008
rect 2184 912 2200 928
rect 2088 812 2104 828
rect 1768 712 1784 728
rect 1864 712 1880 728
rect 1992 712 2008 728
rect 1480 692 1496 708
rect 1560 692 1576 708
rect 1848 692 1864 708
rect 1592 672 1608 688
rect 1832 672 1848 688
rect 1448 612 1464 628
rect 1448 572 1464 588
rect 1480 532 1496 548
rect 1448 512 1464 528
rect 1448 412 1464 428
rect 1432 392 1448 408
rect 1416 332 1432 348
rect 1496 312 1512 328
rect 1432 292 1448 308
rect 1496 292 1512 308
rect 1800 652 1816 668
rect 1768 632 1784 648
rect 1736 592 1752 608
rect 1656 572 1672 588
rect 1672 532 1688 548
rect 1864 592 1880 608
rect 1992 692 2008 708
rect 1912 672 1928 688
rect 1949 602 1985 618
rect 1880 572 1896 588
rect 1944 572 1960 588
rect 1928 552 1944 568
rect 1816 532 1832 548
rect 1608 512 1624 528
rect 1896 512 1912 528
rect 1688 492 1704 508
rect 1528 472 1544 488
rect 2360 972 2376 988
rect 2408 952 2424 968
rect 2392 932 2408 948
rect 2280 912 2296 928
rect 2344 912 2360 928
rect 2200 712 2216 728
rect 2120 706 2136 708
rect 2120 692 2136 706
rect 2216 692 2232 708
rect 2328 872 2344 888
rect 2376 872 2392 888
rect 2360 692 2376 708
rect 2184 672 2200 688
rect 2152 652 2168 668
rect 2328 652 2344 668
rect 2056 532 2072 548
rect 2120 532 2136 548
rect 2264 532 2280 548
rect 1784 492 1800 508
rect 1848 492 1864 508
rect 1912 492 1928 508
rect 1720 432 1736 448
rect 1576 372 1592 388
rect 1672 332 1688 348
rect 1560 292 1576 308
rect 1512 272 1528 288
rect 1544 252 1560 268
rect 1448 232 1480 248
rect 1640 272 1656 288
rect 1576 212 1592 228
rect 1384 192 1400 208
rect 1320 152 1352 168
rect 1592 152 1608 168
rect 1256 132 1272 148
rect 1496 132 1512 148
rect 712 112 728 128
rect 744 114 760 128
rect 744 112 760 114
rect 952 112 968 128
rect 1032 112 1048 128
rect 1720 292 1736 308
rect 1880 412 1896 428
rect 1864 332 1880 348
rect 1928 332 1944 348
rect 2104 512 2120 528
rect 2296 512 2312 528
rect 2040 452 2056 468
rect 2152 492 2168 508
rect 2216 472 2232 488
rect 2136 432 2152 448
rect 2024 412 2040 428
rect 1992 312 2008 328
rect 2232 332 2248 348
rect 2056 312 2072 328
rect 1880 292 1896 308
rect 1992 292 2008 308
rect 2024 292 2040 308
rect 1816 272 1832 288
rect 1736 232 1752 248
rect 1848 252 1864 268
rect 1768 152 1784 168
rect 1704 132 1720 148
rect 1928 232 1944 248
rect 1928 192 1944 208
rect 1949 202 1985 218
rect 1896 152 1912 168
rect 2088 292 2104 308
rect 2056 252 2072 268
rect 2104 252 2120 268
rect 2216 232 2232 248
rect 2024 212 2040 228
rect 2184 152 2200 168
rect 1992 132 2008 148
rect 1608 112 1624 128
rect 1672 112 1688 128
rect 1512 92 1528 108
rect 1624 92 1640 108
rect 925 2 961 18
rect 1816 12 1832 28
rect 2280 292 2296 308
rect 2440 992 2456 1008
rect 2456 912 2472 928
rect 2440 892 2456 908
rect 2424 812 2440 828
rect 2536 1012 2552 1028
rect 2792 1572 2808 1588
rect 2776 1512 2792 1528
rect 2728 1492 2744 1508
rect 2760 1492 2776 1508
rect 2808 1532 2824 1548
rect 2808 1512 2824 1528
rect 2744 1332 2760 1348
rect 2792 1332 2808 1348
rect 2696 1292 2712 1308
rect 2664 1272 2680 1288
rect 2616 1252 2632 1268
rect 2600 1152 2616 1168
rect 2616 1132 2632 1148
rect 2520 944 2552 948
rect 2520 932 2536 944
rect 2536 932 2552 944
rect 2520 672 2536 688
rect 2488 632 2504 648
rect 2488 612 2504 628
rect 2376 512 2392 528
rect 2360 392 2376 408
rect 2328 192 2344 208
rect 2328 152 2344 168
rect 2360 152 2376 168
rect 2328 132 2344 148
rect 2232 112 2248 128
rect 2280 112 2296 128
rect 2152 92 2168 108
rect 2248 92 2260 108
rect 2260 92 2264 108
rect 2504 412 2520 428
rect 2568 832 2584 848
rect 2584 812 2600 828
rect 2696 1192 2712 1208
rect 2696 1172 2712 1188
rect 2664 1112 2680 1128
rect 2728 1312 2744 1328
rect 2712 1152 2728 1168
rect 2744 1152 2760 1168
rect 2728 1112 2744 1128
rect 2728 1092 2744 1108
rect 2888 1852 2904 1868
rect 2920 1832 2936 1848
rect 3064 1912 3080 1928
rect 3048 1892 3064 1908
rect 3256 2512 3272 2528
rect 3272 2512 3288 2528
rect 3112 2272 3128 2288
rect 3096 2132 3112 2148
rect 3144 2312 3160 2328
rect 3144 2292 3160 2308
rect 3192 2232 3208 2248
rect 3144 2152 3160 2168
rect 3144 2132 3160 2148
rect 3256 2272 3272 2288
rect 3320 2272 3336 2288
rect 3208 2172 3224 2188
rect 3208 2152 3224 2168
rect 3128 2112 3144 2128
rect 3256 2112 3272 2128
rect 3112 2072 3128 2088
rect 3240 2072 3256 2088
rect 3112 2032 3128 2048
rect 3176 2012 3192 2028
rect 3192 1972 3208 1988
rect 3176 1952 3192 1968
rect 3160 1892 3176 1908
rect 3192 1912 3208 1928
rect 2952 1872 2968 1888
rect 3064 1872 3080 1888
rect 2984 1852 3000 1868
rect 3048 1832 3064 1848
rect 3256 1832 3272 1848
rect 3416 2892 3432 2908
rect 3400 2872 3416 2888
rect 3448 2732 3464 2748
rect 3544 2732 3560 2748
rect 3432 2712 3448 2728
rect 3496 2712 3512 2728
rect 3560 2712 3576 2728
rect 4008 3052 4024 3068
rect 3896 2992 3912 3008
rect 3997 3002 4033 3018
rect 4040 2992 4056 3008
rect 3864 2932 3880 2948
rect 3896 2932 3912 2948
rect 3720 2912 3736 2928
rect 3848 2912 3864 2928
rect 3736 2812 3752 2828
rect 3640 2732 3656 2748
rect 3640 2712 3656 2728
rect 3576 2692 3592 2708
rect 3384 2672 3400 2688
rect 3416 2672 3432 2688
rect 3512 2672 3528 2688
rect 3592 2672 3608 2688
rect 3416 2632 3432 2648
rect 3480 2572 3496 2588
rect 3384 2532 3400 2548
rect 3448 2532 3464 2548
rect 3496 2512 3512 2528
rect 3592 2632 3608 2648
rect 3768 2752 3784 2768
rect 3752 2712 3768 2728
rect 3704 2672 3720 2688
rect 3528 2572 3544 2588
rect 3672 2572 3688 2588
rect 3720 2552 3736 2568
rect 3672 2532 3688 2548
rect 3512 2492 3528 2508
rect 3400 2332 3416 2348
rect 3496 2332 3512 2348
rect 3624 2512 3640 2528
rect 3592 2472 3608 2488
rect 3560 2352 3576 2368
rect 3352 2292 3368 2308
rect 3432 2272 3448 2288
rect 3480 2312 3496 2328
rect 3544 2312 3560 2328
rect 3368 2132 3384 2148
rect 3416 2112 3432 2128
rect 3352 2072 3368 2088
rect 3320 2052 3336 2068
rect 3304 1952 3320 1968
rect 3368 1952 3384 1968
rect 3352 1892 3368 1908
rect 3352 1852 3368 1868
rect 3384 1892 3400 1908
rect 3368 1812 3384 1828
rect 3272 1792 3288 1808
rect 3368 1792 3384 1808
rect 3480 1952 3496 1968
rect 3416 1932 3432 1948
rect 3448 1932 3464 1948
rect 3464 1912 3480 1928
rect 3544 2152 3560 2168
rect 3752 2572 3768 2588
rect 3928 2892 3944 2908
rect 3848 2672 3864 2688
rect 3816 2592 3832 2608
rect 3784 2532 3800 2548
rect 3736 2392 3752 2408
rect 3768 2372 3784 2388
rect 3704 2332 3720 2348
rect 3800 2332 3816 2348
rect 3640 2292 3656 2308
rect 3768 2312 3784 2328
rect 3880 2652 3896 2668
rect 3864 2592 3880 2608
rect 3928 2632 3944 2648
rect 3896 2612 3912 2628
rect 4008 2732 4024 2748
rect 3976 2692 3992 2708
rect 4072 3092 4088 3108
rect 4104 3032 4120 3048
rect 4216 3892 4232 3908
rect 4216 3812 4232 3828
rect 4216 3752 4232 3768
rect 4408 4112 4424 4128
rect 4456 4112 4472 4128
rect 4248 4092 4264 4108
rect 4232 3692 4248 3708
rect 4216 3552 4232 3568
rect 4184 3512 4200 3528
rect 4296 4052 4312 4068
rect 4328 4032 4344 4048
rect 4312 3932 4328 3948
rect 4440 3906 4456 3908
rect 4440 3892 4456 3906
rect 4584 4152 4600 4168
rect 4600 4132 4616 4148
rect 4552 4092 4568 4108
rect 4600 4072 4616 4088
rect 4856 4892 4872 4908
rect 4920 4892 4936 4908
rect 5064 4832 5080 4848
rect 4760 4812 4776 4828
rect 4968 4812 4984 4828
rect 4808 4772 4824 4788
rect 4920 4752 4936 4768
rect 4680 4572 4696 4588
rect 4856 4632 4872 4648
rect 4728 4552 4744 4568
rect 4760 4552 4776 4568
rect 4808 4552 4824 4568
rect 4696 4532 4712 4548
rect 4664 4512 4680 4528
rect 4952 4712 4968 4728
rect 5021 4802 5057 4818
rect 4984 4672 5000 4688
rect 5000 4672 5016 4688
rect 5112 4772 5128 4788
rect 4792 4532 4808 4548
rect 4824 4532 4840 4548
rect 4808 4512 4824 4528
rect 4728 4452 4744 4468
rect 4648 4432 4664 4448
rect 4680 4352 4696 4368
rect 4776 4312 4792 4328
rect 4680 4152 4696 4168
rect 4664 4032 4680 4048
rect 4552 3912 4568 3928
rect 4600 3912 4616 3928
rect 4552 3892 4568 3908
rect 4344 3872 4360 3888
rect 4520 3872 4536 3888
rect 4344 3812 4360 3828
rect 4312 3732 4328 3748
rect 4280 3506 4296 3508
rect 4280 3492 4296 3506
rect 4312 3432 4328 3448
rect 4168 3352 4184 3368
rect 4232 3352 4248 3368
rect 4184 3332 4200 3348
rect 4296 3332 4312 3348
rect 4632 3932 4648 3948
rect 4648 3912 4664 3928
rect 4696 3972 4712 3988
rect 4760 4212 4776 4228
rect 4728 4092 4744 4108
rect 4744 3972 4760 3988
rect 4712 3952 4728 3968
rect 4680 3892 4696 3908
rect 4440 3812 4456 3828
rect 4504 3812 4520 3828
rect 4600 3812 4616 3828
rect 4456 3772 4472 3788
rect 4472 3752 4488 3768
rect 4680 3852 4696 3868
rect 4648 3812 4680 3828
rect 4520 3792 4536 3808
rect 4616 3792 4632 3808
rect 4632 3772 4648 3788
rect 4568 3752 4584 3768
rect 4616 3732 4632 3748
rect 4600 3692 4616 3708
rect 4504 3592 4520 3608
rect 4504 3532 4520 3548
rect 4536 3512 4568 3528
rect 4488 3492 4504 3508
rect 4632 3492 4648 3508
rect 4376 3472 4392 3488
rect 4568 3472 4584 3488
rect 4392 3452 4408 3468
rect 4600 3452 4616 3468
rect 4168 3292 4184 3308
rect 4216 3292 4232 3308
rect 4216 3192 4232 3208
rect 4264 3112 4276 3128
rect 4276 3112 4280 3128
rect 4248 3092 4264 3108
rect 4232 3052 4248 3068
rect 4152 2992 4168 3008
rect 4152 2952 4168 2968
rect 4312 3272 4328 3288
rect 4312 3192 4328 3208
rect 4328 3132 4344 3148
rect 4312 3092 4328 3108
rect 4232 2992 4248 3008
rect 4296 2992 4312 3008
rect 4200 2932 4216 2948
rect 4168 2872 4184 2888
rect 4072 2692 4088 2708
rect 4056 2652 4072 2668
rect 3976 2632 3992 2648
rect 4040 2632 4056 2648
rect 3960 2592 3976 2608
rect 3997 2602 4033 2618
rect 4120 2672 4136 2688
rect 4216 2672 4232 2688
rect 4072 2572 4088 2588
rect 3944 2532 3960 2548
rect 3992 2532 4008 2548
rect 3896 2512 3912 2528
rect 3848 2432 3864 2448
rect 3864 2392 3880 2408
rect 3832 2312 3848 2328
rect 3784 2292 3800 2308
rect 3640 2272 3656 2288
rect 3848 2272 3864 2288
rect 3912 2492 3928 2508
rect 3992 2512 4008 2528
rect 4168 2572 4184 2588
rect 4360 3072 4376 3088
rect 4344 3052 4360 3068
rect 4296 2932 4312 2948
rect 4344 2912 4360 2928
rect 4264 2892 4280 2908
rect 4360 2892 4376 2908
rect 4600 3432 4616 3448
rect 4472 3332 4488 3348
rect 4568 3314 4584 3328
rect 4568 3312 4584 3314
rect 4664 3792 4680 3808
rect 4664 3692 4680 3708
rect 4680 3592 4696 3608
rect 4664 3532 4680 3548
rect 4648 3292 4664 3308
rect 4488 3132 4504 3148
rect 4424 3112 4440 3128
rect 4744 3932 4760 3948
rect 4792 4172 4808 4188
rect 4776 4072 4792 4088
rect 4776 4052 4792 4068
rect 4728 3832 4744 3848
rect 4760 3832 4776 3848
rect 4840 4492 4856 4508
rect 4888 4492 4904 4508
rect 4824 4212 4840 4228
rect 4856 4452 4872 4468
rect 4904 4272 4920 4288
rect 4904 4172 4920 4188
rect 4936 4512 4952 4528
rect 4936 4312 4952 4328
rect 4984 4312 5000 4328
rect 4968 4292 4984 4308
rect 4840 4112 4856 4128
rect 4856 4112 4872 4128
rect 4824 4092 4840 4108
rect 4872 4092 4888 4108
rect 4856 3912 4872 3928
rect 4840 3872 4856 3888
rect 4824 3812 4840 3828
rect 4808 3792 4824 3808
rect 4760 3772 4776 3788
rect 4744 3752 4760 3768
rect 4760 3752 4776 3768
rect 4776 3512 4792 3528
rect 4712 3492 4728 3508
rect 4744 3492 4760 3508
rect 4680 3412 4696 3428
rect 4728 3412 4760 3428
rect 4792 3412 4808 3428
rect 4712 3392 4728 3408
rect 4680 3332 4696 3348
rect 4696 3312 4712 3328
rect 4712 3272 4728 3288
rect 4712 3112 4728 3128
rect 4488 3052 4504 3068
rect 4552 2992 4568 3008
rect 4664 3012 4680 3028
rect 4632 2952 4648 2968
rect 4760 3352 4776 3368
rect 4744 3292 4760 3308
rect 4776 3292 4792 3308
rect 4776 3192 4792 3208
rect 4744 3112 4760 3128
rect 4808 3332 4824 3348
rect 4840 3732 4856 3748
rect 4968 3892 4984 3908
rect 4936 3852 4952 3868
rect 4888 3772 4904 3788
rect 4952 3752 4968 3768
rect 4968 3712 4984 3728
rect 5128 4692 5144 4708
rect 5496 5292 5512 5308
rect 5544 5292 5560 5308
rect 5432 5272 5448 5288
rect 5480 5272 5496 5288
rect 5256 5092 5272 5108
rect 5368 5106 5384 5108
rect 5368 5092 5384 5106
rect 5224 4932 5240 4948
rect 5336 5032 5352 5048
rect 5288 5012 5304 5028
rect 5384 4912 5400 4928
rect 5224 4772 5240 4788
rect 5192 4712 5208 4728
rect 5256 4732 5272 4748
rect 5384 4732 5400 4748
rect 5304 4692 5320 4708
rect 5128 4672 5144 4688
rect 5240 4672 5256 4688
rect 5352 4672 5368 4688
rect 5224 4652 5240 4668
rect 5256 4652 5272 4668
rect 5336 4652 5352 4668
rect 5304 4632 5320 4648
rect 5336 4632 5352 4648
rect 5224 4612 5240 4628
rect 5272 4592 5288 4608
rect 5224 4552 5240 4568
rect 5288 4552 5304 4568
rect 5112 4532 5128 4548
rect 5272 4532 5288 4548
rect 5368 4612 5384 4628
rect 5432 5092 5448 5108
rect 5496 4932 5528 4948
rect 5432 4732 5464 4748
rect 5416 4712 5432 4728
rect 5464 4712 5480 4728
rect 5560 5252 5576 5268
rect 5560 5032 5576 5048
rect 5576 5012 5592 5028
rect 5896 5432 5912 5448
rect 5880 5412 5896 5428
rect 5784 5332 5800 5348
rect 5672 5312 5688 5328
rect 5704 5132 5720 5148
rect 5832 5312 5848 5328
rect 5816 5292 5848 5308
rect 5752 5092 5768 5108
rect 5768 5012 5784 5028
rect 5640 4972 5656 4988
rect 5720 4972 5736 4988
rect 5848 5232 5864 5248
rect 5928 5492 5944 5508
rect 6008 5492 6024 5508
rect 5928 5452 5944 5468
rect 6232 5492 6248 5508
rect 6584 5492 6600 5508
rect 5992 5472 6008 5488
rect 6088 5472 6104 5488
rect 5960 5452 5976 5468
rect 5992 5452 6008 5468
rect 5944 5432 5960 5448
rect 5992 5412 6008 5428
rect 6045 5402 6081 5418
rect 5928 5352 5944 5368
rect 5880 5172 5896 5188
rect 5896 5152 5912 5168
rect 5832 5072 5848 5088
rect 5912 5092 5928 5108
rect 5944 5332 5960 5348
rect 6248 5452 6264 5468
rect 6312 5452 6328 5468
rect 6248 5372 6264 5388
rect 6296 5352 6312 5368
rect 6200 5332 6216 5348
rect 6232 5312 6248 5328
rect 6280 5312 6296 5328
rect 6024 5292 6040 5308
rect 5944 5132 5960 5148
rect 5944 5112 5960 5128
rect 5992 5112 6008 5128
rect 6104 5132 6120 5148
rect 6024 5092 6040 5108
rect 5960 5072 5976 5088
rect 6045 5002 6081 5018
rect 5944 4952 5960 4968
rect 5672 4932 5688 4948
rect 5768 4932 5784 4948
rect 5624 4912 5640 4928
rect 5704 4912 5720 4928
rect 5752 4912 5768 4928
rect 5544 4832 5560 4848
rect 5528 4732 5544 4748
rect 5880 4872 5896 4888
rect 5848 4852 5864 4868
rect 5688 4732 5704 4748
rect 5560 4712 5576 4728
rect 5608 4712 5624 4728
rect 5640 4712 5656 4728
rect 5416 4652 5432 4668
rect 5528 4652 5544 4668
rect 5400 4592 5416 4608
rect 5816 4712 5832 4728
rect 5656 4652 5672 4668
rect 5656 4632 5688 4648
rect 5512 4612 5528 4628
rect 5608 4612 5624 4628
rect 5416 4552 5432 4568
rect 5496 4552 5512 4568
rect 5320 4532 5336 4548
rect 5384 4532 5400 4548
rect 5176 4512 5192 4528
rect 5080 4492 5096 4508
rect 5021 4402 5057 4418
rect 5192 4492 5208 4508
rect 5128 4372 5144 4388
rect 5016 4272 5032 4288
rect 5000 4112 5016 4128
rect 5021 4002 5057 4018
rect 5096 3992 5112 4008
rect 5064 3912 5068 3928
rect 5068 3912 5080 3928
rect 5112 3892 5128 3908
rect 5000 3872 5016 3888
rect 5080 3872 5096 3888
rect 5000 3832 5016 3848
rect 5000 3712 5016 3728
rect 4984 3692 5000 3708
rect 4872 3552 4888 3568
rect 4872 3532 4888 3548
rect 4936 3512 4952 3528
rect 5021 3602 5057 3618
rect 5000 3532 5016 3548
rect 5064 3532 5080 3548
rect 4968 3472 4984 3488
rect 4840 3292 4856 3308
rect 4840 3072 4856 3088
rect 4728 2972 4744 2988
rect 4440 2932 4456 2948
rect 4568 2932 4584 2948
rect 4744 2932 4760 2948
rect 4776 2932 4792 2948
rect 4456 2912 4472 2928
rect 4808 2912 4824 2928
rect 4456 2892 4472 2908
rect 4712 2892 4728 2908
rect 4408 2872 4424 2888
rect 4408 2772 4424 2788
rect 4664 2752 4680 2768
rect 4824 2812 4840 2828
rect 4872 3392 4888 3408
rect 4984 3332 5000 3348
rect 4920 3292 4936 3308
rect 4968 3232 4984 3248
rect 5032 3492 5048 3508
rect 5096 3732 5112 3748
rect 5144 4292 5160 4308
rect 5176 4152 5192 4168
rect 5256 4112 5272 4128
rect 5272 4092 5288 4108
rect 5320 3932 5336 3948
rect 5208 3912 5224 3928
rect 5192 3852 5208 3868
rect 5224 3752 5240 3768
rect 5272 3732 5288 3748
rect 5176 3712 5192 3728
rect 5128 3572 5144 3588
rect 5256 3572 5272 3588
rect 5128 3552 5144 3568
rect 5208 3492 5224 3508
rect 5080 3472 5096 3488
rect 5064 3432 5080 3448
rect 5064 3412 5080 3428
rect 5192 3412 5208 3428
rect 5192 3392 5208 3408
rect 5021 3202 5057 3218
rect 4968 3092 4984 3108
rect 5096 3092 5112 3108
rect 4872 3072 4888 3088
rect 4856 2992 4872 3008
rect 5032 3072 5048 3088
rect 5064 3072 5080 3088
rect 5032 3052 5048 3068
rect 4856 2972 4872 2988
rect 4984 2972 5000 2988
rect 4744 2752 4760 2768
rect 4792 2752 4808 2768
rect 4712 2712 4728 2728
rect 4776 2712 4792 2728
rect 4328 2692 4344 2708
rect 4552 2706 4568 2708
rect 4552 2692 4568 2706
rect 4664 2692 4680 2708
rect 4456 2672 4472 2688
rect 4632 2672 4648 2688
rect 4264 2652 4280 2668
rect 4168 2532 4184 2548
rect 4072 2512 4088 2528
rect 4104 2512 4120 2528
rect 4088 2492 4104 2508
rect 4136 2492 4152 2508
rect 4056 2472 4072 2488
rect 4072 2432 4088 2448
rect 4200 2432 4216 2448
rect 4056 2412 4072 2428
rect 4056 2312 4072 2328
rect 4280 2572 4296 2588
rect 4232 2532 4248 2548
rect 4488 2552 4504 2568
rect 4376 2532 4392 2548
rect 4408 2532 4424 2548
rect 4296 2512 4312 2528
rect 4248 2472 4264 2488
rect 4232 2432 4248 2448
rect 4328 2412 4344 2428
rect 4248 2352 4264 2368
rect 3880 2292 3896 2308
rect 4296 2312 4312 2328
rect 4424 2512 4440 2528
rect 4360 2312 4376 2328
rect 4344 2292 4360 2308
rect 4408 2292 4424 2308
rect 4184 2232 4200 2248
rect 3997 2202 4033 2218
rect 4136 2192 4152 2208
rect 4360 2272 4376 2288
rect 4280 2232 4296 2248
rect 4344 2232 4360 2248
rect 4296 2192 4312 2208
rect 4264 2152 4280 2168
rect 4312 2152 4328 2168
rect 3544 2132 3560 2148
rect 3560 2132 3576 2148
rect 3592 2132 3608 2148
rect 3864 2132 3880 2148
rect 3960 2132 3976 2148
rect 3976 2132 3992 2148
rect 4136 2132 4152 2148
rect 3512 2112 3528 2128
rect 3528 1912 3544 1928
rect 3432 1892 3448 1908
rect 3496 1892 3512 1908
rect 3480 1872 3496 1888
rect 3416 1832 3432 1848
rect 3448 1832 3464 1848
rect 3336 1772 3352 1788
rect 3400 1772 3416 1788
rect 3080 1752 3096 1768
rect 2856 1732 2872 1748
rect 3016 1732 3032 1748
rect 3208 1732 3224 1748
rect 2888 1712 2904 1728
rect 3032 1712 3048 1728
rect 2872 1692 2888 1708
rect 3000 1692 3016 1708
rect 2957 1602 2993 1618
rect 2872 1532 2904 1548
rect 2936 1532 2952 1548
rect 2856 1332 2872 1348
rect 2888 1512 2904 1528
rect 3224 1512 3240 1528
rect 2920 1492 2936 1508
rect 3144 1492 3160 1508
rect 3128 1472 3144 1488
rect 2904 1332 2920 1348
rect 2968 1332 2984 1348
rect 3176 1332 3192 1348
rect 2872 1312 2888 1328
rect 2808 1132 2824 1148
rect 2840 1132 2856 1148
rect 2760 1112 2776 1128
rect 2808 1112 2824 1128
rect 2840 1112 2856 1128
rect 2792 1092 2808 1108
rect 2776 1072 2792 1088
rect 2840 1092 2856 1108
rect 2824 1052 2840 1068
rect 2664 932 2680 948
rect 2696 892 2712 908
rect 2776 872 2792 888
rect 2632 832 2648 848
rect 2632 692 2648 708
rect 2600 672 2616 688
rect 2584 652 2600 668
rect 2680 632 2696 648
rect 2632 572 2648 588
rect 2552 512 2568 528
rect 2600 512 2616 528
rect 2744 592 2760 608
rect 2792 672 2808 688
rect 2808 592 2824 608
rect 2776 552 2792 568
rect 2728 532 2744 548
rect 2584 492 2588 508
rect 2588 492 2600 508
rect 2616 492 2632 508
rect 2424 352 2440 368
rect 2504 272 2520 288
rect 2504 192 2520 208
rect 2472 132 2488 148
rect 2472 92 2488 108
rect 2536 392 2552 408
rect 2632 332 2648 348
rect 2552 312 2568 328
rect 2616 252 2632 268
rect 2600 152 2616 168
rect 2760 514 2776 528
rect 2760 512 2776 514
rect 2696 312 2712 328
rect 2744 312 2760 328
rect 2728 292 2744 308
rect 2840 306 2856 308
rect 2840 292 2856 306
rect 2728 272 2744 288
rect 2760 272 2776 288
rect 2680 232 2696 248
rect 2648 212 2680 228
rect 2632 132 2648 148
rect 2536 114 2552 128
rect 2536 112 2552 114
rect 2616 112 2632 128
rect 2840 232 2856 248
rect 2792 172 2808 188
rect 2888 1292 2900 1308
rect 2900 1292 2904 1308
rect 2872 1112 2888 1128
rect 2936 1312 2952 1328
rect 3080 1292 3096 1308
rect 2957 1202 2993 1218
rect 3048 1132 3064 1148
rect 3464 1752 3480 1768
rect 3416 1652 3432 1668
rect 3432 1612 3448 1628
rect 3320 1592 3336 1608
rect 3528 1752 3544 1768
rect 3480 1672 3496 1688
rect 3496 1632 3512 1648
rect 3368 1572 3384 1588
rect 3544 1572 3560 1588
rect 3416 1452 3432 1468
rect 3448 1452 3464 1468
rect 3368 1392 3384 1408
rect 3320 1372 3336 1388
rect 3400 1372 3416 1388
rect 3448 1372 3464 1388
rect 3384 1352 3400 1368
rect 3432 1352 3448 1368
rect 3160 1112 3176 1128
rect 3192 1112 3208 1128
rect 2872 1072 2888 1088
rect 3160 1072 3176 1088
rect 3240 1072 3256 1088
rect 2888 1052 2904 1068
rect 2968 1012 3000 1028
rect 3160 952 3176 968
rect 3272 1032 3288 1048
rect 3160 932 3176 948
rect 3064 912 3080 928
rect 2957 802 2993 818
rect 3080 732 3096 748
rect 3048 712 3064 728
rect 2888 692 2904 708
rect 2936 692 2952 708
rect 2872 672 2888 688
rect 2920 672 2936 688
rect 2904 632 2920 648
rect 2888 592 2904 608
rect 3000 692 3016 708
rect 3016 692 3032 708
rect 3144 712 3160 728
rect 3496 1472 3512 1488
rect 3512 1392 3528 1408
rect 3496 1372 3512 1388
rect 3496 1352 3512 1368
rect 3544 1352 3560 1368
rect 3480 1272 3496 1288
rect 3400 1132 3416 1148
rect 3432 1132 3448 1148
rect 3336 1112 3352 1128
rect 3368 1072 3384 1088
rect 3416 1072 3432 1088
rect 3304 1052 3320 1068
rect 3352 1052 3368 1068
rect 3384 952 3400 968
rect 3464 1052 3480 1068
rect 3496 1092 3512 1108
rect 3480 992 3496 1008
rect 3416 932 3432 948
rect 3464 932 3480 948
rect 3432 912 3448 928
rect 3480 912 3496 928
rect 3288 872 3304 888
rect 3256 712 3272 728
rect 3112 692 3128 708
rect 3160 692 3176 708
rect 3480 852 3496 868
rect 3352 732 3368 748
rect 3512 1032 3528 1048
rect 3512 992 3528 1008
rect 3784 2112 3800 2128
rect 3912 2112 3928 2128
rect 3704 2092 3720 2108
rect 3576 2052 3592 2068
rect 3576 2032 3592 2048
rect 3624 2032 3640 2048
rect 3608 1932 3624 1948
rect 3672 1992 3688 2008
rect 3896 2072 3912 2088
rect 3912 1972 3928 1988
rect 3864 1932 3880 1948
rect 3752 1912 3768 1928
rect 3752 1792 3768 1808
rect 3624 1732 3640 1748
rect 3704 1712 3720 1728
rect 3608 1692 3624 1708
rect 3704 1692 3720 1708
rect 3592 1572 3608 1588
rect 3576 1492 3592 1508
rect 3656 1612 3672 1628
rect 3720 1652 3736 1668
rect 3736 1652 3752 1668
rect 3608 1512 3640 1528
rect 3624 1492 3640 1508
rect 3576 1472 3592 1488
rect 3560 1312 3576 1328
rect 3560 1292 3576 1308
rect 3608 1332 3624 1348
rect 3656 1372 3672 1388
rect 3640 1332 3656 1348
rect 3672 1312 3688 1328
rect 3608 1292 3624 1308
rect 3592 1272 3608 1288
rect 3592 1112 3608 1128
rect 3544 1092 3560 1108
rect 3560 1092 3592 1108
rect 3576 972 3592 988
rect 3528 952 3544 968
rect 3544 932 3560 948
rect 3512 872 3528 888
rect 3736 1552 3752 1568
rect 3736 1332 3752 1348
rect 3768 1432 3784 1448
rect 3800 1672 3816 1688
rect 3944 1872 3960 1888
rect 3832 1712 3848 1728
rect 4008 2072 4024 2088
rect 3992 1932 4008 1948
rect 4088 2112 4104 2128
rect 4168 2112 4184 2128
rect 4040 2012 4056 2028
rect 4104 2092 4120 2108
rect 4184 2012 4200 2028
rect 4056 1972 4072 1988
rect 4136 1972 4152 1988
rect 4008 1912 4024 1928
rect 4024 1872 4040 1888
rect 4040 1852 4056 1868
rect 3960 1812 3976 1828
rect 3997 1802 4033 1818
rect 3976 1772 3992 1788
rect 3960 1732 3976 1748
rect 4120 1812 4136 1828
rect 4072 1792 4088 1808
rect 4056 1712 4072 1728
rect 4104 1712 4120 1728
rect 3832 1692 3848 1708
rect 3896 1692 3912 1708
rect 3992 1692 4008 1708
rect 4088 1692 4104 1708
rect 3816 1552 3832 1568
rect 3928 1672 3944 1688
rect 3896 1552 3912 1568
rect 3944 1652 3960 1668
rect 3992 1652 4008 1668
rect 4024 1632 4040 1648
rect 3896 1512 3912 1528
rect 3832 1472 3848 1488
rect 3784 1352 3800 1368
rect 3880 1472 3896 1488
rect 4008 1472 4024 1488
rect 3912 1432 3928 1448
rect 3944 1412 3960 1428
rect 3976 1412 3992 1428
rect 3976 1392 3992 1408
rect 3997 1402 4033 1418
rect 3848 1352 3864 1368
rect 3752 1312 3768 1328
rect 3800 1332 3816 1348
rect 3704 1272 3720 1288
rect 3720 1272 3736 1288
rect 3688 1252 3704 1268
rect 3672 1152 3688 1168
rect 3656 1072 3672 1088
rect 3656 952 3672 968
rect 3640 932 3656 948
rect 3592 912 3608 928
rect 3640 912 3656 928
rect 3720 1252 3736 1268
rect 3704 1132 3720 1148
rect 3704 1112 3720 1128
rect 3816 1292 3832 1308
rect 3800 1232 3816 1248
rect 3752 1152 3768 1168
rect 4072 1632 4088 1648
rect 4120 1672 4136 1688
rect 4152 1892 4168 1908
rect 4264 1972 4280 1988
rect 4200 1932 4216 1948
rect 4168 1732 4184 1748
rect 4136 1652 4152 1668
rect 4152 1632 4168 1648
rect 4088 1572 4104 1588
rect 4088 1552 4104 1568
rect 4184 1672 4200 1688
rect 4216 1892 4232 1908
rect 4232 1852 4248 1868
rect 4232 1812 4248 1828
rect 4344 2052 4360 2068
rect 4296 2012 4312 2028
rect 4328 1912 4344 1928
rect 4280 1792 4296 1808
rect 4248 1772 4264 1788
rect 4216 1692 4232 1708
rect 4200 1632 4216 1648
rect 4168 1612 4184 1628
rect 4200 1572 4216 1588
rect 4200 1552 4216 1568
rect 4184 1512 4200 1528
rect 4008 1352 4024 1368
rect 4040 1352 4056 1368
rect 3864 1332 3880 1348
rect 3944 1332 3960 1348
rect 3848 1292 3864 1308
rect 3912 1292 3928 1308
rect 3960 1292 3976 1308
rect 3992 1292 4008 1308
rect 3896 1252 3912 1268
rect 3880 1212 3896 1228
rect 3960 1132 3976 1148
rect 3976 1132 3992 1148
rect 3800 1112 3816 1128
rect 3832 1112 3848 1128
rect 3864 1112 3876 1128
rect 3876 1112 3880 1128
rect 3880 1112 3896 1128
rect 3944 1112 3960 1128
rect 3832 1092 3848 1108
rect 3864 1092 3880 1108
rect 3816 1072 3832 1088
rect 4024 1072 4040 1088
rect 3784 1052 3800 1068
rect 3880 1052 3896 1068
rect 3976 1052 3992 1068
rect 3752 1032 3768 1048
rect 3704 972 3720 988
rect 3832 972 3848 988
rect 3608 892 3624 908
rect 3672 892 3688 908
rect 3736 932 3752 948
rect 3768 912 3784 928
rect 3816 912 3832 928
rect 3752 872 3768 888
rect 3528 852 3544 868
rect 3688 852 3704 868
rect 3496 752 3512 768
rect 3592 812 3608 828
rect 3656 752 3672 768
rect 3624 732 3640 748
rect 3544 712 3548 728
rect 3548 712 3560 728
rect 3592 712 3608 728
rect 3640 712 3656 728
rect 3576 692 3592 708
rect 3448 672 3464 688
rect 3496 672 3512 688
rect 3128 652 3144 668
rect 3048 612 3064 628
rect 3080 612 3096 628
rect 2904 492 2920 508
rect 3032 552 3048 568
rect 3064 552 3080 568
rect 3160 632 3176 648
rect 2957 402 2993 418
rect 2872 332 2888 348
rect 2856 152 2872 168
rect 2680 112 2696 128
rect 2712 92 2728 108
rect 2696 12 2712 28
rect 2968 312 2984 328
rect 2904 132 2920 148
rect 3144 472 3160 488
rect 3096 372 3112 388
rect 3112 352 3128 368
rect 3080 332 3096 348
rect 3160 312 3176 328
rect 3192 572 3208 588
rect 3368 592 3384 608
rect 3224 532 3240 548
rect 3208 512 3224 528
rect 3192 292 3208 308
rect 3000 272 3016 288
rect 3176 272 3192 288
rect 3016 252 3032 268
rect 3048 252 3064 268
rect 3000 192 3016 208
rect 2968 112 2984 128
rect 2936 92 2952 108
rect 2957 2 2993 18
rect 3224 472 3240 488
rect 3592 672 3608 688
rect 3512 632 3528 648
rect 3512 612 3528 628
rect 3496 532 3512 548
rect 3272 512 3288 528
rect 3304 514 3320 528
rect 3304 512 3320 514
rect 3464 492 3480 508
rect 3240 452 3256 468
rect 3384 432 3400 448
rect 3384 352 3400 368
rect 3432 352 3448 368
rect 3304 332 3320 348
rect 3272 312 3288 328
rect 3336 312 3352 328
rect 3352 312 3368 328
rect 3272 292 3288 308
rect 3432 332 3448 348
rect 3320 272 3336 288
rect 3400 272 3416 288
rect 3112 132 3128 148
rect 3048 112 3064 128
rect 3064 112 3080 128
rect 3480 292 3496 308
rect 3480 272 3496 288
rect 3496 212 3512 228
rect 3496 132 3512 148
rect 3592 652 3608 668
rect 3576 532 3592 548
rect 3560 432 3576 448
rect 3544 392 3560 408
rect 3528 172 3544 188
rect 3320 112 3336 128
rect 3032 92 3048 108
rect 3144 92 3160 108
rect 3320 92 3336 108
rect 3464 92 3480 108
rect 3480 12 3496 28
rect 3800 892 3816 908
rect 3880 932 3896 948
rect 3960 992 3976 1008
rect 3997 1002 4033 1018
rect 3944 912 3960 928
rect 3992 952 4008 968
rect 3960 872 3976 888
rect 3768 772 3784 788
rect 3832 732 3848 748
rect 3688 712 3704 728
rect 3768 712 3784 728
rect 4024 812 4040 828
rect 3896 732 3912 748
rect 4168 1432 4184 1448
rect 4136 1392 4152 1408
rect 4168 1332 4184 1348
rect 4152 1312 4168 1328
rect 4056 1292 4072 1308
rect 4072 1252 4088 1268
rect 4104 1192 4120 1208
rect 4088 1112 4104 1128
rect 4184 1272 4200 1288
rect 4168 1252 4184 1268
rect 4056 1092 4072 1108
rect 4088 1072 4104 1088
rect 4184 1052 4200 1068
rect 4072 952 4088 968
rect 4120 952 4136 968
rect 4152 952 4168 968
rect 4120 932 4136 948
rect 4168 932 4184 948
rect 4152 912 4168 928
rect 4088 892 4104 908
rect 4120 872 4136 888
rect 4152 872 4168 888
rect 4120 852 4136 868
rect 4088 792 4104 808
rect 4056 752 4072 768
rect 3704 692 3720 708
rect 3736 692 3752 708
rect 3784 692 3800 708
rect 3816 692 3832 708
rect 3784 672 3800 688
rect 3704 652 3736 668
rect 3672 572 3688 588
rect 3704 552 3720 568
rect 3656 512 3672 528
rect 3672 432 3688 448
rect 3640 392 3656 408
rect 3704 412 3720 428
rect 3608 372 3624 388
rect 3640 372 3656 388
rect 3784 552 3800 568
rect 3784 532 3800 548
rect 3752 512 3768 528
rect 3736 492 3752 508
rect 3848 672 3880 688
rect 3832 572 3848 588
rect 3880 492 3896 508
rect 3864 452 3880 468
rect 3880 312 3896 328
rect 3928 712 3944 728
rect 4040 712 4056 728
rect 3912 692 3928 708
rect 3960 692 3976 708
rect 3992 692 4008 708
rect 4120 752 4136 768
rect 4184 852 4200 868
rect 4168 812 4200 828
rect 4168 752 4184 768
rect 4136 732 4152 748
rect 4152 732 4168 748
rect 4104 712 4120 728
rect 4008 672 4024 688
rect 4136 672 4152 688
rect 4152 632 4168 648
rect 3997 602 4033 618
rect 4072 612 4088 628
rect 4040 552 4056 568
rect 4104 572 4120 588
rect 4296 1732 4312 1748
rect 4536 2532 4552 2548
rect 4712 2532 4728 2548
rect 4568 2512 4584 2528
rect 4632 2514 4648 2528
rect 4632 2512 4648 2514
rect 4744 2512 4760 2528
rect 4744 2492 4760 2508
rect 4664 2292 4680 2308
rect 4456 2252 4472 2268
rect 4520 2252 4536 2268
rect 4568 2232 4584 2248
rect 4392 1912 4408 1928
rect 4488 2114 4504 2128
rect 4488 2112 4504 2114
rect 4680 2192 4696 2208
rect 4728 2152 4744 2168
rect 4776 2592 4792 2608
rect 4840 2732 4856 2748
rect 4808 2532 4824 2548
rect 4792 2492 4808 2508
rect 4776 2472 4792 2488
rect 4616 2132 4632 2148
rect 4664 2132 4680 2148
rect 4760 2132 4776 2148
rect 4600 2112 4616 2128
rect 4648 2112 4664 2128
rect 4712 2112 4728 2128
rect 4520 2092 4536 2108
rect 4680 2092 4696 2108
rect 4552 1912 4568 1928
rect 4568 1892 4584 1908
rect 4360 1712 4376 1728
rect 4392 1712 4408 1728
rect 4296 1692 4312 1708
rect 4360 1692 4376 1708
rect 4280 1632 4296 1648
rect 4280 1512 4296 1528
rect 4360 1452 4376 1468
rect 4216 1412 4232 1428
rect 4232 1392 4248 1408
rect 4216 1372 4232 1388
rect 4312 1352 4328 1368
rect 4440 1752 4456 1768
rect 4520 1752 4536 1768
rect 4504 1732 4520 1748
rect 4552 1732 4568 1748
rect 4488 1712 4504 1728
rect 4408 1692 4424 1708
rect 4456 1692 4472 1708
rect 4472 1692 4488 1708
rect 4440 1632 4456 1648
rect 4392 1512 4408 1528
rect 4408 1472 4424 1488
rect 4376 1392 4392 1408
rect 4376 1352 4392 1368
rect 4424 1312 4440 1328
rect 4504 1612 4520 1628
rect 4456 1552 4472 1568
rect 4488 1532 4504 1548
rect 4472 1432 4488 1448
rect 4456 1352 4472 1368
rect 4472 1312 4488 1328
rect 4520 1392 4536 1408
rect 4520 1312 4536 1328
rect 4296 1292 4312 1308
rect 4280 1272 4296 1288
rect 4296 1232 4312 1248
rect 4248 1172 4264 1188
rect 4248 1152 4264 1168
rect 4344 1232 4360 1248
rect 4216 1112 4232 1128
rect 4312 1112 4328 1128
rect 4264 1092 4280 1108
rect 4312 1092 4328 1108
rect 4264 1032 4280 1048
rect 4392 1172 4408 1188
rect 4360 1152 4376 1168
rect 4296 1072 4312 1088
rect 4328 1072 4344 1088
rect 4328 1032 4344 1048
rect 4280 1012 4296 1028
rect 4248 972 4264 988
rect 4344 972 4360 988
rect 4264 952 4280 968
rect 4264 912 4280 928
rect 4296 912 4312 928
rect 4344 912 4360 928
rect 4344 892 4360 908
rect 4216 712 4232 728
rect 4216 692 4232 708
rect 4200 672 4216 688
rect 4440 1132 4456 1148
rect 4392 1052 4408 1068
rect 4520 1252 4536 1268
rect 4536 1252 4552 1268
rect 4504 1152 4520 1168
rect 4536 1112 4552 1128
rect 4760 2032 4776 2048
rect 4840 2672 4856 2688
rect 4840 2312 4856 2328
rect 4872 2952 4888 2968
rect 4936 2932 4952 2948
rect 5128 3292 5144 3308
rect 5160 3132 5176 3148
rect 5160 3112 5176 3128
rect 5112 2972 5128 2988
rect 4936 2892 4952 2908
rect 4968 2892 4984 2908
rect 5112 2892 5128 2908
rect 4872 2712 4888 2728
rect 4872 2512 4888 2528
rect 4872 2312 4888 2328
rect 4872 2292 4888 2308
rect 4840 2272 4856 2288
rect 4824 2252 4840 2268
rect 4808 2152 4824 2168
rect 4792 2112 4808 2128
rect 4728 1912 4744 1928
rect 4776 1912 4792 1928
rect 4776 1892 4792 1908
rect 4696 1872 4712 1888
rect 4744 1872 4760 1888
rect 4760 1852 4776 1868
rect 4872 2072 4888 2088
rect 4984 2792 5000 2808
rect 5021 2802 5057 2818
rect 5144 2972 5160 2988
rect 5224 3472 5240 3488
rect 5320 3712 5336 3728
rect 5480 4492 5496 4508
rect 5448 4472 5464 4488
rect 5464 4312 5480 4328
rect 5496 4312 5512 4328
rect 5368 4292 5384 4308
rect 5464 4292 5480 4308
rect 5560 4572 5576 4588
rect 5736 4632 5752 4648
rect 5768 4612 5784 4628
rect 5864 4812 5880 4828
rect 5848 4612 5864 4628
rect 5544 4552 5560 4568
rect 5720 4552 5736 4568
rect 5528 4532 5544 4548
rect 5784 4532 5800 4548
rect 5816 4532 5832 4548
rect 5608 4492 5624 4508
rect 5576 4412 5592 4428
rect 5640 4432 5656 4448
rect 5608 4392 5624 4408
rect 5640 4332 5656 4348
rect 5656 4312 5672 4328
rect 5512 4272 5528 4288
rect 5576 4212 5592 4228
rect 5352 4132 5368 4148
rect 5384 4132 5400 4148
rect 5544 4132 5560 4148
rect 5640 4132 5656 4148
rect 5592 4112 5608 4128
rect 5384 3972 5400 3988
rect 5368 3832 5384 3848
rect 5416 3932 5432 3948
rect 5512 3906 5528 3908
rect 5512 3892 5528 3906
rect 5416 3872 5432 3888
rect 5416 3832 5432 3848
rect 5336 3672 5352 3688
rect 5304 3632 5320 3648
rect 5352 3632 5368 3648
rect 5368 3572 5384 3588
rect 5304 3532 5320 3548
rect 5336 3512 5352 3528
rect 5240 3452 5256 3468
rect 5288 3452 5304 3468
rect 5352 3492 5368 3508
rect 5400 3572 5416 3588
rect 5384 3532 5400 3548
rect 5384 3512 5400 3528
rect 5720 4472 5736 4488
rect 5784 4412 5800 4428
rect 5944 4912 5960 4928
rect 5992 4912 6008 4928
rect 5928 4892 5944 4908
rect 6360 5432 6376 5448
rect 6744 5506 6760 5508
rect 6744 5492 6760 5506
rect 6936 5492 6952 5508
rect 7016 5492 7032 5508
rect 6568 5472 6584 5488
rect 6632 5472 6648 5488
rect 6664 5472 6680 5488
rect 6808 5472 6824 5488
rect 6904 5472 6920 5488
rect 6456 5452 6472 5468
rect 6568 5452 6584 5468
rect 6552 5432 6568 5448
rect 6440 5372 6456 5388
rect 6344 5332 6360 5348
rect 6488 5332 6504 5348
rect 6408 5312 6424 5328
rect 6456 5312 6472 5328
rect 6392 5292 6408 5308
rect 6424 5292 6436 5308
rect 6436 5292 6440 5308
rect 6568 5292 6584 5308
rect 6328 5272 6344 5288
rect 6152 5092 6168 5108
rect 6136 4912 6152 4928
rect 6088 4872 6104 4888
rect 6008 4792 6024 4808
rect 5912 4572 5928 4588
rect 5816 4372 5832 4388
rect 5768 4332 5784 4348
rect 5832 4332 5848 4348
rect 5720 4312 5736 4328
rect 5800 4312 5816 4328
rect 5720 4292 5736 4308
rect 5752 4292 5768 4308
rect 5736 4272 5752 4288
rect 5752 4272 5768 4288
rect 5736 4112 5752 4128
rect 5688 4012 5704 4028
rect 5656 3912 5672 3928
rect 5624 3892 5640 3908
rect 5672 3892 5688 3908
rect 5592 3872 5608 3888
rect 5640 3872 5656 3888
rect 5736 3992 5752 4008
rect 5720 3912 5736 3928
rect 5544 3772 5560 3788
rect 5512 3752 5528 3768
rect 5640 3752 5656 3768
rect 5480 3732 5496 3748
rect 5656 3732 5672 3748
rect 5576 3714 5592 3728
rect 5576 3712 5592 3714
rect 5496 3632 5512 3648
rect 5416 3492 5432 3508
rect 5352 3452 5384 3468
rect 5432 3452 5448 3468
rect 5320 3432 5336 3448
rect 5448 3392 5464 3408
rect 5496 3392 5512 3408
rect 5400 3352 5416 3368
rect 5448 3332 5464 3348
rect 5320 3312 5336 3328
rect 5496 3312 5512 3328
rect 5432 3232 5448 3248
rect 5336 3212 5352 3228
rect 5704 3712 5720 3728
rect 5672 3692 5688 3708
rect 5704 3692 5720 3708
rect 5688 3672 5704 3688
rect 5688 3552 5704 3568
rect 5592 3532 5608 3548
rect 5544 3472 5560 3488
rect 5544 3352 5560 3368
rect 5736 3672 5752 3688
rect 5880 4312 5896 4328
rect 5896 4272 5912 4288
rect 5928 4492 5944 4508
rect 5864 4212 5880 4228
rect 5768 4172 5784 4188
rect 5848 4152 5864 4168
rect 5832 4132 5848 4148
rect 5864 4112 5880 4128
rect 5880 3992 5896 4008
rect 5912 4212 5928 4228
rect 5912 4172 5928 4188
rect 6088 4792 6104 4808
rect 6152 4772 6168 4788
rect 6040 4712 6056 4728
rect 6072 4712 6088 4728
rect 6024 4692 6040 4708
rect 5960 4612 5976 4628
rect 6008 4612 6024 4628
rect 5992 4592 6008 4608
rect 5992 4532 6008 4548
rect 6088 4632 6104 4648
rect 6344 5032 6360 5048
rect 6456 5092 6472 5108
rect 6616 5092 6632 5108
rect 6456 5052 6472 5068
rect 6248 4932 6264 4948
rect 6600 4932 6616 4948
rect 6328 4912 6344 4928
rect 6440 4912 6456 4928
rect 6552 4912 6568 4928
rect 6264 4892 6280 4908
rect 6328 4892 6344 4908
rect 6408 4852 6424 4868
rect 6184 4832 6200 4848
rect 6168 4732 6184 4748
rect 6168 4712 6184 4728
rect 6136 4672 6152 4688
rect 6045 4602 6081 4618
rect 6120 4612 6136 4628
rect 6168 4592 6184 4608
rect 6584 4892 6600 4908
rect 6712 5452 6728 5468
rect 6664 5332 6680 5348
rect 6856 5332 6872 5348
rect 6936 5432 6952 5448
rect 6984 5432 7016 5448
rect 6824 5312 6840 5328
rect 6920 5312 6936 5328
rect 6680 5092 6696 5108
rect 6648 5072 6664 5088
rect 6808 5052 6824 5068
rect 6808 5032 6824 5048
rect 6776 4932 6792 4948
rect 6680 4912 6696 4928
rect 6760 4912 6776 4928
rect 6680 4892 6696 4908
rect 6664 4872 6680 4888
rect 6456 4812 6472 4828
rect 6520 4812 6536 4828
rect 6632 4812 6648 4828
rect 6376 4772 6392 4788
rect 6200 4752 6216 4768
rect 6280 4752 6296 4768
rect 6200 4732 6232 4748
rect 6264 4732 6280 4748
rect 6216 4672 6232 4688
rect 6344 4732 6360 4748
rect 6200 4632 6216 4648
rect 6232 4632 6248 4648
rect 6296 4632 6312 4648
rect 6232 4592 6248 4608
rect 6072 4532 6088 4548
rect 6088 4532 6104 4548
rect 6024 4492 6040 4508
rect 6088 4492 6104 4508
rect 6120 4492 6136 4508
rect 6024 4292 6040 4308
rect 6040 4292 6056 4308
rect 5944 4272 5960 4288
rect 5976 4272 5992 4288
rect 5960 4252 5976 4268
rect 5928 4152 5960 4168
rect 6152 4512 6168 4528
rect 6136 4352 6152 4368
rect 6120 4312 6136 4328
rect 6072 4272 6088 4288
rect 6045 4202 6081 4218
rect 6072 4152 6088 4168
rect 5960 4132 5976 4148
rect 6008 4112 6024 4128
rect 6088 4112 6104 4128
rect 6104 4112 6120 4128
rect 5976 3992 5992 4008
rect 5896 3972 5912 3988
rect 5864 3932 5880 3948
rect 5992 3932 6008 3948
rect 5608 3492 5624 3508
rect 5720 3492 5736 3508
rect 5624 3472 5640 3488
rect 5656 3472 5672 3488
rect 5624 3452 5640 3468
rect 5640 3432 5656 3448
rect 5576 3332 5592 3348
rect 5608 3312 5624 3328
rect 5528 3292 5544 3308
rect 5576 3292 5592 3308
rect 5368 3132 5384 3148
rect 5288 3112 5304 3128
rect 5256 3092 5272 3108
rect 5320 3092 5336 3108
rect 5208 3072 5224 3088
rect 5272 3052 5288 3068
rect 5288 3052 5304 3068
rect 5256 2992 5272 3008
rect 5144 2952 5160 2968
rect 5224 2952 5240 2968
rect 5176 2932 5192 2948
rect 5272 2952 5288 2968
rect 5320 2992 5336 3008
rect 5304 2932 5320 2948
rect 5560 3112 5576 3128
rect 5384 3092 5400 3108
rect 5352 2972 5368 2988
rect 5416 3072 5432 3088
rect 5400 3012 5416 3028
rect 5512 2992 5528 3008
rect 5576 2992 5592 3008
rect 5640 3072 5656 3088
rect 5208 2912 5224 2928
rect 5304 2912 5320 2928
rect 5400 2912 5416 2928
rect 5416 2912 5432 2928
rect 5208 2892 5224 2908
rect 5288 2892 5304 2908
rect 5320 2892 5336 2908
rect 5496 2892 5512 2908
rect 5544 2892 5560 2908
rect 5464 2872 5480 2888
rect 5368 2852 5384 2868
rect 5128 2752 5144 2768
rect 4936 2712 4952 2728
rect 4904 2692 4920 2708
rect 5080 2692 5096 2708
rect 4952 2672 4968 2688
rect 5160 2672 5176 2688
rect 4936 2532 4952 2548
rect 4920 2512 4936 2528
rect 4968 2512 4984 2528
rect 4904 2492 4908 2508
rect 4908 2492 4920 2508
rect 4984 2492 5000 2508
rect 4968 2452 4984 2468
rect 5021 2402 5057 2418
rect 5112 2532 5128 2548
rect 5128 2512 5144 2528
rect 5080 2492 5096 2508
rect 5080 2472 5096 2488
rect 5448 2712 5464 2728
rect 5336 2706 5352 2708
rect 5336 2692 5352 2706
rect 5448 2692 5464 2708
rect 5272 2672 5288 2688
rect 5240 2652 5256 2668
rect 5416 2652 5432 2668
rect 5224 2512 5240 2528
rect 5304 2512 5320 2528
rect 5192 2412 5208 2428
rect 5000 2272 5016 2288
rect 4936 2252 4952 2268
rect 4920 2152 4936 2168
rect 5096 2232 5112 2248
rect 5064 2172 5080 2188
rect 5096 2132 5112 2148
rect 5064 2112 5080 2128
rect 4936 2072 4952 2088
rect 4888 2032 4904 2048
rect 4840 2012 4856 2028
rect 4872 1972 4888 1988
rect 4840 1892 4856 1908
rect 4904 1872 4920 1888
rect 4776 1792 4792 1808
rect 4808 1792 4824 1808
rect 4664 1752 4680 1768
rect 4744 1752 4760 1768
rect 4600 1712 4616 1728
rect 4616 1692 4632 1708
rect 4600 1532 4616 1548
rect 4904 1752 4920 1768
rect 4792 1732 4808 1748
rect 4904 1732 4920 1748
rect 4792 1712 4808 1728
rect 4824 1692 4840 1708
rect 4856 1672 4872 1688
rect 4776 1632 4792 1648
rect 4760 1512 4776 1528
rect 4680 1492 4696 1508
rect 4840 1512 4856 1528
rect 4584 1412 4600 1428
rect 4664 1392 4680 1408
rect 4616 1352 4632 1368
rect 4632 1332 4648 1348
rect 4792 1452 4808 1468
rect 4760 1352 4776 1368
rect 5021 2002 5057 2018
rect 4984 1952 5000 1968
rect 5096 1932 5112 1948
rect 5176 2172 5192 2188
rect 5176 2152 5192 2168
rect 5176 2132 5192 2148
rect 5128 2112 5144 2128
rect 4984 1872 5000 1888
rect 5192 1872 5208 1888
rect 4968 1772 4984 1788
rect 4952 1732 4968 1748
rect 4952 1712 4968 1728
rect 4872 1552 4888 1568
rect 4872 1532 4888 1548
rect 4888 1512 4904 1528
rect 4872 1352 4888 1368
rect 4680 1332 4696 1348
rect 4600 1292 4616 1308
rect 4600 1232 4616 1248
rect 4632 1272 4648 1288
rect 4632 1252 4648 1268
rect 4568 1132 4584 1148
rect 4616 1172 4632 1188
rect 4664 1232 4680 1248
rect 4632 1132 4648 1148
rect 4568 1092 4584 1108
rect 4616 1092 4632 1108
rect 4600 1072 4616 1088
rect 4440 1052 4456 1068
rect 4552 1052 4568 1068
rect 4504 1032 4520 1048
rect 4424 972 4440 988
rect 4408 952 4424 968
rect 4424 952 4440 968
rect 4408 912 4424 928
rect 4456 912 4472 928
rect 4504 912 4520 928
rect 4296 872 4312 888
rect 4376 872 4392 888
rect 4392 852 4408 868
rect 4360 812 4376 828
rect 4264 792 4296 808
rect 4344 792 4360 808
rect 4312 772 4328 788
rect 4296 712 4312 728
rect 4520 852 4536 868
rect 4456 732 4472 748
rect 4392 712 4408 728
rect 4456 712 4472 728
rect 4536 712 4552 728
rect 4184 552 4200 568
rect 4040 492 4056 508
rect 4104 472 4120 488
rect 3976 452 3992 468
rect 3880 292 3896 308
rect 3960 292 3976 308
rect 3640 272 3656 288
rect 3688 272 3704 288
rect 3576 132 3592 148
rect 3848 272 3864 288
rect 3720 132 3736 148
rect 3560 112 3576 128
rect 3608 112 3624 128
rect 3688 112 3704 128
rect 3704 112 3720 128
rect 3944 152 3960 168
rect 4232 652 4248 668
rect 4328 592 4344 608
rect 4264 572 4280 588
rect 4280 552 4296 568
rect 4344 532 4360 548
rect 4312 512 4328 528
rect 4360 512 4376 528
rect 4280 492 4296 508
rect 4216 472 4232 488
rect 4200 432 4216 448
rect 4008 392 4024 408
rect 3992 312 4008 328
rect 4248 352 4264 368
rect 4264 292 4280 308
rect 3997 202 4033 218
rect 3976 172 3992 188
rect 4200 192 4216 208
rect 4168 152 4200 168
rect 4264 152 4280 168
rect 4120 132 4136 148
rect 4216 132 4232 148
rect 4328 452 4344 468
rect 4424 592 4440 608
rect 4408 552 4424 568
rect 4392 472 4408 488
rect 4376 352 4392 368
rect 4392 312 4408 328
rect 4328 292 4344 308
rect 4488 532 4504 548
rect 4376 272 4392 288
rect 4472 272 4488 288
rect 4392 192 4408 208
rect 4360 152 4376 168
rect 4520 252 4536 268
rect 4664 952 4680 968
rect 4792 1312 4808 1328
rect 4840 1312 4856 1328
rect 4824 1292 4828 1308
rect 4828 1292 4840 1308
rect 4824 1272 4840 1288
rect 4728 1152 4744 1168
rect 4760 1132 4776 1148
rect 4792 1092 4808 1108
rect 4792 1072 4808 1088
rect 4840 1072 4856 1088
rect 4760 972 4776 988
rect 4728 914 4744 928
rect 4728 912 4744 914
rect 4632 812 4648 828
rect 4616 692 4632 708
rect 4792 872 4808 888
rect 4760 712 4776 728
rect 4808 672 4824 688
rect 4872 1092 4888 1108
rect 4856 1052 4872 1068
rect 4856 932 4872 948
rect 5000 1752 5016 1768
rect 4952 1392 4968 1408
rect 4984 1392 5000 1408
rect 4952 1332 4968 1348
rect 4968 1292 4984 1308
rect 4904 1112 4920 1128
rect 4952 1112 4968 1128
rect 4984 1072 5000 1088
rect 4968 1052 4984 1068
rect 4952 972 4968 988
rect 4920 912 4936 928
rect 4952 892 4968 908
rect 4904 872 4920 888
rect 4920 732 4936 748
rect 5192 1732 5208 1748
rect 5032 1712 5048 1728
rect 5016 1692 5032 1708
rect 5048 1692 5064 1708
rect 5128 1692 5144 1708
rect 5144 1672 5176 1688
rect 5021 1602 5057 1618
rect 5128 1552 5144 1568
rect 5080 1532 5096 1548
rect 5096 1412 5112 1428
rect 5021 1202 5057 1218
rect 5112 1332 5128 1348
rect 5096 1112 5112 1128
rect 5176 1552 5192 1568
rect 5160 1492 5176 1508
rect 5240 2492 5256 2508
rect 5240 2292 5256 2308
rect 5384 2632 5400 2648
rect 5560 2772 5576 2788
rect 5640 2772 5656 2788
rect 5544 2712 5560 2728
rect 5640 2752 5656 2768
rect 5608 2712 5624 2728
rect 5720 3392 5736 3408
rect 5896 3912 5912 3928
rect 5944 3912 5960 3928
rect 5928 3892 5944 3908
rect 5928 3872 5944 3888
rect 5976 3852 5992 3868
rect 5944 3832 5960 3848
rect 5880 3812 5896 3828
rect 5880 3772 5896 3788
rect 5832 3752 5848 3768
rect 5960 3732 5976 3748
rect 5800 3652 5816 3668
rect 5928 3512 5944 3528
rect 5960 3512 5976 3528
rect 5800 3472 5816 3488
rect 5880 3472 5896 3488
rect 5768 3432 5800 3448
rect 5768 3392 5784 3408
rect 5864 3392 5880 3408
rect 5848 3332 5864 3348
rect 5752 3312 5768 3328
rect 5784 3312 5800 3328
rect 5768 3032 5784 3048
rect 5992 3712 6008 3728
rect 5992 3492 6008 3508
rect 5976 3432 5992 3448
rect 5944 3292 5960 3308
rect 5800 3252 5816 3268
rect 5992 3292 6008 3308
rect 5976 3232 5992 3248
rect 5800 3112 5816 3128
rect 6232 4532 6248 4548
rect 6664 4752 6680 4768
rect 6424 4692 6440 4708
rect 6552 4672 6568 4688
rect 6440 4632 6472 4648
rect 6536 4632 6552 4648
rect 6408 4592 6424 4608
rect 6472 4592 6488 4608
rect 6632 4692 6648 4708
rect 6600 4672 6616 4688
rect 6616 4652 6632 4668
rect 6568 4592 6584 4608
rect 6616 4552 6632 4568
rect 6312 4512 6328 4528
rect 6184 4492 6200 4508
rect 6232 4306 6248 4308
rect 6232 4292 6248 4306
rect 6216 4112 6232 4128
rect 6232 4092 6248 4108
rect 6344 4412 6360 4428
rect 6648 4632 6664 4648
rect 6664 4552 6680 4568
rect 6536 4512 6552 4528
rect 6440 4472 6456 4488
rect 6408 4352 6424 4368
rect 6520 4452 6536 4468
rect 6456 4432 6472 4448
rect 6664 4432 6680 4448
rect 6952 5292 6968 5308
rect 6840 5072 6856 5088
rect 6824 4872 6840 4888
rect 6856 4792 6872 4808
rect 6696 4752 6712 4768
rect 6728 4732 6744 4748
rect 6696 4712 6712 4728
rect 6888 5012 6904 5028
rect 6952 5092 6968 5108
rect 7000 5312 7016 5328
rect 7000 5292 7016 5308
rect 7000 5172 7016 5188
rect 6968 5052 6984 5068
rect 6920 4932 6936 4948
rect 6968 4932 6984 4948
rect 6904 4712 6920 4728
rect 6712 4692 6728 4708
rect 6760 4692 6776 4708
rect 6792 4692 6808 4708
rect 7032 5472 7048 5488
rect 7032 5332 7048 5348
rect 7176 5312 7192 5328
rect 7053 5202 7089 5218
rect 7400 5392 7416 5408
rect 7208 5132 7240 5148
rect 7128 5092 7144 5108
rect 7240 5072 7256 5088
rect 7016 5032 7032 5048
rect 7256 5032 7272 5048
rect 7304 5312 7320 5328
rect 7304 5292 7320 5308
rect 7336 5292 7352 5308
rect 7288 5252 7304 5268
rect 7304 5132 7320 5148
rect 7288 5072 7304 5088
rect 7112 4932 7128 4948
rect 6936 4892 6952 4908
rect 7000 4892 7016 4908
rect 6936 4712 6952 4728
rect 7112 4872 7128 4888
rect 7053 4802 7089 4818
rect 7032 4712 7048 4728
rect 7080 4712 7096 4728
rect 7016 4692 7032 4708
rect 6808 4672 6824 4688
rect 6840 4672 6856 4688
rect 6872 4672 6888 4688
rect 6888 4672 6904 4688
rect 6936 4672 6952 4688
rect 6744 4652 6760 4668
rect 6856 4652 6872 4668
rect 6728 4632 6744 4648
rect 6824 4632 6840 4648
rect 6888 4632 6904 4648
rect 6696 4572 6712 4588
rect 6776 4572 6792 4588
rect 6824 4552 6840 4568
rect 6808 4532 6824 4548
rect 6872 4532 6888 4548
rect 6936 4572 6952 4588
rect 6968 4572 6984 4588
rect 6968 4552 6984 4568
rect 7032 4672 7048 4688
rect 7000 4632 7016 4648
rect 6728 4512 6744 4528
rect 6840 4512 6856 4528
rect 6984 4512 7000 4528
rect 6856 4492 6872 4508
rect 6888 4492 6904 4508
rect 6856 4472 6872 4488
rect 6536 4332 6552 4348
rect 6664 4332 6680 4348
rect 6776 4332 6792 4348
rect 6824 4332 6840 4348
rect 6440 4312 6456 4328
rect 6408 4292 6424 4308
rect 6344 4172 6360 4188
rect 6392 4172 6408 4188
rect 6296 4112 6312 4128
rect 6248 4052 6264 4068
rect 6200 4032 6216 4048
rect 6168 3992 6184 4008
rect 6136 3972 6152 3988
rect 6168 3912 6184 3928
rect 6024 3892 6040 3908
rect 6040 3872 6056 3888
rect 6072 3872 6088 3888
rect 6104 3872 6120 3888
rect 6136 3832 6152 3848
rect 6045 3802 6081 3818
rect 6024 3772 6040 3788
rect 6184 3772 6200 3788
rect 6104 3732 6120 3748
rect 6408 3972 6424 3988
rect 6280 3912 6296 3928
rect 6296 3912 6312 3928
rect 6248 3892 6264 3908
rect 6328 3892 6344 3908
rect 6264 3872 6280 3888
rect 6040 3712 6056 3728
rect 6024 3472 6040 3488
rect 6120 3512 6136 3528
rect 6200 3512 6216 3528
rect 6088 3492 6104 3508
rect 6232 3692 6248 3708
rect 6216 3492 6232 3508
rect 5928 3092 5944 3108
rect 5848 3072 5864 3088
rect 5832 2972 5848 2988
rect 5864 2952 5880 2968
rect 5800 2872 5816 2888
rect 5928 2992 5944 3008
rect 5976 3052 5992 3068
rect 5976 2952 5992 2968
rect 5976 2932 5992 2948
rect 5896 2912 5912 2928
rect 5944 2912 5960 2928
rect 5896 2892 5912 2908
rect 5928 2892 5944 2908
rect 5736 2752 5752 2768
rect 5672 2712 5688 2728
rect 5720 2712 5736 2728
rect 5496 2592 5512 2608
rect 5416 2512 5432 2528
rect 5352 2472 5368 2488
rect 5352 2306 5368 2308
rect 5352 2292 5368 2306
rect 5448 2332 5464 2348
rect 5480 2332 5496 2348
rect 5464 2312 5480 2328
rect 5464 2292 5480 2308
rect 5528 2632 5544 2648
rect 5624 2632 5640 2648
rect 5592 2572 5608 2588
rect 5528 2512 5544 2528
rect 5512 2312 5528 2328
rect 5544 2472 5560 2488
rect 5704 2612 5720 2628
rect 5608 2532 5624 2548
rect 5656 2512 5672 2528
rect 5640 2472 5656 2488
rect 5688 2472 5704 2488
rect 5720 2532 5736 2548
rect 5768 2732 5784 2748
rect 5880 2832 5896 2848
rect 5816 2812 5832 2828
rect 5752 2672 5768 2688
rect 5736 2512 5752 2528
rect 5768 2512 5784 2528
rect 5720 2492 5736 2508
rect 5640 2312 5656 2328
rect 5704 2312 5720 2328
rect 5656 2292 5672 2308
rect 5624 2272 5640 2288
rect 5384 2252 5400 2268
rect 5496 2252 5512 2268
rect 5288 2192 5304 2208
rect 5304 2152 5320 2168
rect 5528 2232 5544 2248
rect 5672 2232 5688 2248
rect 5544 2192 5560 2208
rect 5352 2132 5368 2148
rect 5400 2132 5416 2148
rect 5448 2132 5464 2148
rect 5272 2114 5288 2128
rect 5272 2112 5288 2114
rect 5384 2112 5400 2128
rect 5432 2112 5448 2128
rect 5224 1952 5240 1968
rect 5272 1952 5288 1968
rect 5256 1932 5272 1948
rect 5320 1932 5336 1948
rect 5256 1692 5272 1708
rect 5224 1672 5240 1688
rect 5240 1632 5256 1648
rect 5208 1512 5224 1528
rect 5272 1552 5288 1568
rect 5256 1492 5272 1508
rect 5224 1332 5240 1348
rect 5176 1312 5192 1328
rect 5224 1292 5240 1308
rect 5144 1112 5160 1128
rect 5112 1092 5128 1108
rect 5021 802 5057 818
rect 5144 912 5160 928
rect 5128 892 5144 908
rect 4936 712 4952 728
rect 5000 712 5016 728
rect 4648 632 4680 648
rect 4776 632 4792 648
rect 4712 592 4728 608
rect 4760 572 4776 588
rect 4600 532 4616 548
rect 4728 532 4744 548
rect 4824 652 4840 668
rect 4840 592 4856 608
rect 4904 592 4920 608
rect 4840 572 4856 588
rect 4824 552 4840 568
rect 4920 552 4936 568
rect 4616 412 4632 428
rect 4568 392 4584 408
rect 4568 352 4584 368
rect 4552 312 4568 328
rect 4680 332 4696 348
rect 4856 332 4872 348
rect 4616 312 4632 328
rect 4808 312 4824 328
rect 4760 292 4776 308
rect 4888 312 4904 328
rect 4904 292 4920 308
rect 4584 272 4600 288
rect 4968 672 4984 688
rect 5016 632 5032 648
rect 5096 572 5112 588
rect 4968 532 4984 548
rect 5144 532 5160 548
rect 4936 452 4952 468
rect 5021 402 5057 418
rect 4936 312 4952 328
rect 5128 492 5144 508
rect 5080 472 5096 488
rect 4744 252 4760 268
rect 4808 252 4824 268
rect 4920 252 4936 268
rect 5000 252 5016 268
rect 4616 232 4632 248
rect 4536 192 4552 208
rect 4728 192 4744 208
rect 4504 172 4536 188
rect 4472 152 4488 168
rect 4616 152 4632 168
rect 4840 232 4856 248
rect 4968 212 4984 228
rect 5112 332 5128 348
rect 5192 1112 5208 1128
rect 5208 1092 5224 1108
rect 5400 1912 5416 1928
rect 5432 1892 5448 1908
rect 5304 1852 5320 1868
rect 5368 1732 5384 1748
rect 5320 1532 5336 1548
rect 5352 1492 5368 1508
rect 5304 1312 5320 1328
rect 5288 1172 5304 1188
rect 5176 1072 5192 1088
rect 5208 1052 5224 1068
rect 5176 932 5192 948
rect 5176 712 5192 728
rect 5176 672 5192 688
rect 5624 2172 5640 2188
rect 5592 2132 5608 2148
rect 5576 2112 5592 2128
rect 5688 2192 5704 2208
rect 5656 2132 5672 2148
rect 5704 2112 5720 2128
rect 5640 1892 5656 1908
rect 5480 1812 5496 1828
rect 5624 1832 5640 1848
rect 5576 1752 5592 1768
rect 5640 1752 5656 1768
rect 5704 1752 5720 1768
rect 5656 1732 5672 1748
rect 5688 1732 5704 1748
rect 5528 1712 5544 1728
rect 5560 1712 5576 1728
rect 5496 1652 5512 1668
rect 5544 1612 5560 1628
rect 5384 1532 5400 1548
rect 5432 1512 5448 1528
rect 5416 1492 5432 1508
rect 5384 1332 5400 1348
rect 5608 1712 5624 1728
rect 5736 2312 5752 2328
rect 5944 2872 5960 2888
rect 5944 2692 5960 2708
rect 5912 2672 5928 2688
rect 5848 2652 5864 2668
rect 5880 2652 5896 2668
rect 5912 2652 5928 2668
rect 5944 2652 5960 2668
rect 5848 2612 5864 2628
rect 5880 2612 5896 2628
rect 5832 2532 5848 2548
rect 5896 2552 5912 2568
rect 5832 2472 5848 2488
rect 5816 2306 5832 2308
rect 5816 2292 5832 2306
rect 5784 2172 5800 2188
rect 5752 2152 5768 2168
rect 5784 2132 5800 2148
rect 5752 2092 5768 2108
rect 5912 2392 5928 2408
rect 5880 2372 5896 2388
rect 5864 2332 5880 2348
rect 5912 2312 5928 2328
rect 5896 2212 5912 2228
rect 6168 3452 6184 3468
rect 6232 3452 6248 3468
rect 6045 3402 6081 3418
rect 6200 3412 6216 3428
rect 6120 3332 6136 3348
rect 6040 3132 6056 3148
rect 6040 3112 6056 3128
rect 6088 3232 6104 3248
rect 6136 3132 6152 3148
rect 6184 3132 6200 3148
rect 6232 3112 6248 3128
rect 6136 3092 6152 3108
rect 6072 3072 6088 3088
rect 6120 3032 6136 3048
rect 6045 3002 6081 3018
rect 6008 2812 6024 2828
rect 5992 2752 6008 2768
rect 6168 3072 6184 3088
rect 6184 3032 6200 3048
rect 6200 3012 6216 3028
rect 6152 2952 6168 2968
rect 6104 2932 6120 2948
rect 6232 2992 6248 3008
rect 6136 2892 6152 2908
rect 6216 2892 6232 2908
rect 6168 2872 6184 2888
rect 6344 3852 6360 3868
rect 6312 3832 6328 3848
rect 6312 3812 6328 3828
rect 6264 3792 6280 3808
rect 6264 3772 6280 3788
rect 6296 3772 6312 3788
rect 6264 3732 6280 3748
rect 6328 3692 6344 3708
rect 6456 4292 6472 4308
rect 6552 4292 6568 4308
rect 6472 4252 6488 4268
rect 6472 4232 6488 4248
rect 6664 4272 6680 4288
rect 6712 4212 6728 4228
rect 6504 4152 6520 4168
rect 6584 4152 6600 4168
rect 6472 4132 6488 4148
rect 6840 4252 6856 4268
rect 6744 4132 6760 4148
rect 6536 4112 6552 4128
rect 6600 4112 6616 4128
rect 6728 4112 6744 4128
rect 6520 4032 6536 4048
rect 6520 3932 6536 3948
rect 6552 3932 6568 3948
rect 6600 3932 6616 3948
rect 6472 3912 6488 3928
rect 6424 3872 6440 3888
rect 6552 3912 6568 3928
rect 6488 3872 6504 3888
rect 6456 3832 6472 3848
rect 6504 3812 6520 3828
rect 6504 3772 6520 3788
rect 6536 3772 6552 3788
rect 6520 3752 6536 3768
rect 6584 3792 6600 3808
rect 6440 3732 6456 3748
rect 6456 3732 6472 3748
rect 6504 3732 6520 3748
rect 6664 3912 6680 3928
rect 6648 3852 6664 3868
rect 6680 3892 6696 3908
rect 6728 3832 6744 3848
rect 6536 3712 6552 3728
rect 6696 3712 6712 3728
rect 6472 3652 6488 3668
rect 6392 3592 6408 3608
rect 6920 4492 6936 4508
rect 7016 4492 7032 4508
rect 6904 4452 6920 4468
rect 6872 4312 6888 4328
rect 7000 4312 7032 4328
rect 6968 4192 6984 4208
rect 7096 4692 7112 4708
rect 7112 4672 7128 4688
rect 7128 4592 7144 4608
rect 7192 4872 7208 4888
rect 7160 4712 7176 4728
rect 7144 4552 7160 4568
rect 7112 4532 7128 4548
rect 7144 4532 7160 4548
rect 7288 4692 7304 4708
rect 7208 4552 7224 4568
rect 7320 5032 7336 5048
rect 7368 5312 7384 5328
rect 7416 5312 7432 5328
rect 7384 5292 7400 5308
rect 7560 5392 7576 5408
rect 7496 5372 7512 5388
rect 7592 5372 7608 5388
rect 7544 5332 7560 5348
rect 7480 5252 7496 5268
rect 7512 5252 7528 5268
rect 7496 5072 7512 5088
rect 7352 5012 7368 5028
rect 7368 4932 7384 4948
rect 7336 4912 7352 4928
rect 7496 4932 7512 4948
rect 7672 5472 7688 5488
rect 7752 5492 7768 5508
rect 7864 5506 7880 5508
rect 7864 5492 7880 5506
rect 7720 5472 7736 5488
rect 7688 5452 7704 5468
rect 7720 5412 7736 5428
rect 7640 5392 7656 5408
rect 7688 5352 7704 5368
rect 7736 5332 7752 5348
rect 7624 5292 7640 5308
rect 7656 5312 7672 5328
rect 7704 5312 7720 5328
rect 7752 5312 7768 5328
rect 7800 5472 7816 5488
rect 7784 5392 7800 5408
rect 7784 5332 7800 5348
rect 7608 5132 7624 5148
rect 7608 5092 7624 5108
rect 7576 5072 7592 5088
rect 7608 5052 7624 5068
rect 7544 5032 7560 5048
rect 7528 4892 7544 4908
rect 7512 4872 7528 4888
rect 7464 4832 7480 4848
rect 7448 4732 7464 4748
rect 7400 4712 7416 4728
rect 7592 4832 7608 4848
rect 7528 4752 7544 4768
rect 7432 4692 7448 4708
rect 7416 4652 7432 4668
rect 7384 4632 7400 4648
rect 7320 4592 7336 4608
rect 7304 4512 7320 4528
rect 7053 4402 7089 4418
rect 7032 4292 7048 4308
rect 7000 4272 7016 4288
rect 6936 4172 6952 4188
rect 6952 4152 6968 4168
rect 7032 4252 7048 4268
rect 7032 4192 7048 4208
rect 6936 4132 6952 4148
rect 6760 4114 6776 4128
rect 6760 4112 6776 4114
rect 6792 4112 6808 4128
rect 7016 4112 7032 4128
rect 6904 4092 6908 4108
rect 6908 4092 6920 4108
rect 6840 4032 6856 4048
rect 6792 4012 6808 4028
rect 6760 3912 6776 3928
rect 6824 3992 6840 4008
rect 6808 3892 6824 3908
rect 6776 3872 6792 3888
rect 6776 3812 6792 3828
rect 6760 3752 6776 3768
rect 6888 4072 6904 4088
rect 6920 4072 6936 4088
rect 6904 4052 6920 4068
rect 7016 4092 7032 4108
rect 6936 4052 6952 4068
rect 6984 4052 7000 4068
rect 6936 4032 6952 4048
rect 6840 3912 6856 3928
rect 6872 3912 6888 3928
rect 6840 3792 6856 3808
rect 6744 3732 6760 3748
rect 6808 3732 6824 3748
rect 6760 3712 6776 3728
rect 6616 3692 6628 3708
rect 6628 3692 6632 3708
rect 6632 3692 6648 3708
rect 6744 3692 6760 3708
rect 6792 3672 6808 3688
rect 6728 3612 6744 3628
rect 6664 3592 6680 3608
rect 6664 3552 6680 3568
rect 6424 3512 6440 3528
rect 6664 3512 6680 3528
rect 6472 3492 6488 3508
rect 6296 3472 6312 3488
rect 6312 3452 6328 3468
rect 6360 3432 6376 3448
rect 6328 3372 6344 3388
rect 6344 3352 6360 3368
rect 6424 3372 6440 3388
rect 6328 3312 6344 3328
rect 6376 3312 6392 3328
rect 6408 3292 6424 3308
rect 6600 3492 6616 3508
rect 6648 3492 6664 3508
rect 6568 3452 6584 3468
rect 6712 3472 6728 3488
rect 6744 3452 6760 3468
rect 6792 3452 6808 3468
rect 6632 3432 6648 3448
rect 6600 3372 6616 3388
rect 6840 3692 6856 3708
rect 6824 3652 6840 3668
rect 6856 3672 6872 3688
rect 6888 3852 6904 3868
rect 6904 3792 6920 3808
rect 6888 3772 6904 3788
rect 6920 3772 6936 3788
rect 6952 3832 6968 3848
rect 6968 3792 6984 3808
rect 6952 3712 6968 3728
rect 6872 3532 6888 3548
rect 6840 3432 6856 3448
rect 6600 3352 6616 3368
rect 6808 3352 6824 3368
rect 6440 3332 6456 3348
rect 6616 3332 6632 3348
rect 6472 3292 6488 3308
rect 6664 3192 6680 3208
rect 6728 3192 6744 3208
rect 6568 3172 6584 3188
rect 6328 3132 6344 3148
rect 6344 3132 6360 3148
rect 6408 3132 6424 3148
rect 6456 3132 6472 3148
rect 6632 3132 6648 3148
rect 6792 3132 6808 3148
rect 6264 3072 6280 3088
rect 6328 3072 6344 3088
rect 6264 3052 6280 3068
rect 6280 3012 6296 3028
rect 6296 2972 6312 2988
rect 6168 2792 6184 2808
rect 6248 2792 6264 2808
rect 6088 2772 6104 2788
rect 6040 2712 6056 2728
rect 6152 2712 6168 2728
rect 6024 2692 6040 2708
rect 6056 2692 6072 2708
rect 5992 2512 6008 2528
rect 6040 2672 6056 2688
rect 6088 2672 6104 2688
rect 6045 2602 6081 2618
rect 6296 2752 6312 2768
rect 6200 2732 6216 2748
rect 6264 2712 6280 2728
rect 6104 2652 6136 2668
rect 6088 2592 6104 2608
rect 6136 2552 6152 2568
rect 6040 2512 6056 2528
rect 6024 2492 6040 2508
rect 6008 2472 6024 2488
rect 6136 2372 6152 2388
rect 6184 2652 6200 2668
rect 6248 2672 6264 2688
rect 6216 2612 6232 2628
rect 6280 2612 6296 2628
rect 6296 2592 6312 2608
rect 6216 2552 6232 2568
rect 6264 2532 6280 2548
rect 6328 2712 6344 2728
rect 6312 2512 6328 2528
rect 6504 3112 6520 3128
rect 6456 3092 6472 3108
rect 6520 3092 6536 3108
rect 6648 3092 6664 3108
rect 6696 3092 6712 3108
rect 6376 3072 6392 3088
rect 6504 3072 6520 3088
rect 6360 2732 6376 2748
rect 6472 3052 6488 3068
rect 6552 3032 6568 3048
rect 6536 2992 6552 3008
rect 6552 2952 6568 2968
rect 6680 3072 6696 3088
rect 6664 3012 6680 3028
rect 6648 2992 6664 3008
rect 6632 2952 6648 2968
rect 6904 3572 6920 3588
rect 6952 3512 6968 3528
rect 6936 3492 6952 3508
rect 6952 3452 6968 3468
rect 6888 3432 6904 3448
rect 6952 3352 6968 3368
rect 6920 3232 6936 3248
rect 6888 3172 6904 3188
rect 6952 3132 6968 3148
rect 6760 3072 6776 3088
rect 6840 3072 6856 3088
rect 6792 2992 6824 3008
rect 6744 2972 6760 2988
rect 6712 2952 6728 2968
rect 6680 2932 6696 2948
rect 6616 2912 6632 2928
rect 6488 2892 6504 2908
rect 6600 2892 6616 2908
rect 6456 2792 6472 2808
rect 6408 2732 6424 2748
rect 6888 2932 6904 2948
rect 6936 3012 6952 3028
rect 6984 3732 7000 3748
rect 7000 3612 7016 3628
rect 6984 3452 7000 3468
rect 6984 3432 7000 3448
rect 7160 4472 7176 4488
rect 7176 4312 7192 4328
rect 7192 4292 7208 4308
rect 7192 4252 7208 4268
rect 7112 4192 7128 4208
rect 7048 4152 7064 4168
rect 7048 4132 7064 4148
rect 7144 4132 7160 4148
rect 7112 4112 7128 4128
rect 7053 4002 7089 4018
rect 7112 3892 7128 3908
rect 7288 4212 7304 4228
rect 7288 4132 7304 4148
rect 7224 4114 7240 4128
rect 7224 4112 7240 4114
rect 7288 3932 7304 3948
rect 7224 3912 7236 3928
rect 7236 3912 7240 3928
rect 7208 3892 7224 3908
rect 7272 3892 7288 3908
rect 7144 3832 7160 3848
rect 7096 3732 7112 3748
rect 7128 3692 7144 3708
rect 7096 3652 7112 3668
rect 7032 3592 7048 3608
rect 7053 3602 7089 3618
rect 7016 3572 7032 3588
rect 7064 3512 7080 3528
rect 7112 3532 7128 3548
rect 7176 3692 7192 3708
rect 7304 3872 7320 3888
rect 7256 3712 7272 3728
rect 7272 3712 7288 3728
rect 7288 3692 7304 3708
rect 7160 3672 7176 3688
rect 7192 3672 7208 3688
rect 7208 3632 7224 3648
rect 7192 3552 7208 3568
rect 7256 3572 7272 3588
rect 7208 3492 7224 3508
rect 7128 3372 7144 3388
rect 7064 3352 7080 3368
rect 7160 3352 7176 3368
rect 7192 3352 7208 3368
rect 7096 3332 7112 3348
rect 7128 3332 7144 3348
rect 7192 3312 7208 3328
rect 6984 3292 7000 3308
rect 7000 3272 7016 3288
rect 7053 3202 7089 3218
rect 7080 3172 7096 3188
rect 7032 3072 7048 3088
rect 7000 2992 7016 3008
rect 7016 2972 7032 2988
rect 7064 2932 7080 2948
rect 6712 2912 6728 2928
rect 6920 2912 6936 2928
rect 7064 2912 7080 2928
rect 6712 2892 6728 2908
rect 6696 2872 6712 2888
rect 6568 2832 6584 2848
rect 6696 2792 6712 2808
rect 6392 2712 6408 2728
rect 6424 2712 6440 2728
rect 6488 2712 6504 2728
rect 6552 2692 6584 2708
rect 6680 2692 6696 2708
rect 6520 2672 6536 2688
rect 6568 2672 6584 2688
rect 6584 2652 6600 2668
rect 6408 2632 6424 2648
rect 6472 2632 6488 2648
rect 6568 2632 6584 2648
rect 6392 2572 6408 2588
rect 6360 2552 6376 2568
rect 6424 2612 6440 2628
rect 6456 2592 6472 2608
rect 6520 2532 6536 2548
rect 6392 2512 6408 2528
rect 6312 2492 6328 2508
rect 6344 2472 6360 2488
rect 6424 2472 6440 2488
rect 6200 2392 6216 2408
rect 6168 2352 6184 2368
rect 5960 2332 5976 2348
rect 5960 2272 5976 2288
rect 5928 2192 5944 2208
rect 6024 2252 6040 2268
rect 6424 2372 6440 2388
rect 6328 2332 6344 2348
rect 6312 2312 6328 2328
rect 6280 2292 6296 2308
rect 6008 2232 6024 2248
rect 6072 2232 6088 2248
rect 6045 2202 6081 2218
rect 6184 2192 6200 2208
rect 6104 2132 6120 2148
rect 6152 2132 6168 2148
rect 5848 2052 5864 2068
rect 5944 2092 5960 2108
rect 5864 1972 5880 1988
rect 5928 1952 5944 1968
rect 6072 2092 6088 2108
rect 5864 1932 5880 1948
rect 5944 1932 5976 1948
rect 5992 1932 6008 1948
rect 5832 1892 5848 1908
rect 5816 1872 5832 1888
rect 5752 1752 5768 1768
rect 5768 1732 5784 1748
rect 5800 1732 5816 1748
rect 5960 1892 5976 1908
rect 6008 1892 6024 1908
rect 6088 1892 6104 1908
rect 5928 1872 5960 1888
rect 5976 1872 5992 1888
rect 6040 1872 6056 1888
rect 5944 1852 5960 1868
rect 5896 1832 5912 1848
rect 5848 1672 5864 1688
rect 5672 1652 5704 1668
rect 5720 1652 5736 1668
rect 5592 1592 5608 1608
rect 5592 1572 5608 1588
rect 5576 1512 5592 1528
rect 5560 1492 5576 1508
rect 5544 1472 5560 1488
rect 5704 1532 5720 1548
rect 5752 1532 5768 1548
rect 5816 1532 5832 1548
rect 5736 1492 5752 1508
rect 5768 1472 5784 1488
rect 5800 1352 5816 1368
rect 5512 1332 5528 1348
rect 5624 1332 5640 1348
rect 5720 1332 5736 1348
rect 5432 1312 5448 1328
rect 5512 1312 5528 1328
rect 5560 1312 5576 1328
rect 5688 1312 5704 1328
rect 5736 1312 5752 1328
rect 5400 1292 5432 1308
rect 5480 1292 5496 1308
rect 5464 1272 5480 1288
rect 5528 1272 5544 1288
rect 5400 1112 5416 1128
rect 5320 1072 5336 1088
rect 5304 1052 5320 1068
rect 5240 952 5256 968
rect 5336 952 5352 968
rect 5272 932 5288 948
rect 5352 932 5368 948
rect 5272 912 5288 928
rect 5240 892 5256 908
rect 5336 892 5352 908
rect 5368 692 5384 708
rect 5304 672 5320 688
rect 5288 652 5304 668
rect 5224 552 5240 568
rect 5320 552 5336 568
rect 5384 632 5400 648
rect 5352 532 5368 548
rect 5176 492 5192 508
rect 5160 312 5176 328
rect 5192 292 5208 308
rect 5256 492 5272 508
rect 5224 472 5240 488
rect 5240 332 5256 348
rect 5224 312 5240 328
rect 5208 252 5224 268
rect 5064 132 5080 148
rect 5176 132 5192 148
rect 5352 512 5368 528
rect 5304 492 5320 508
rect 5336 492 5352 508
rect 5368 492 5384 508
rect 5384 492 5400 508
rect 5448 1072 5464 1088
rect 5432 932 5448 948
rect 5480 1172 5496 1188
rect 5528 1172 5544 1188
rect 5832 1512 5848 1528
rect 5880 1532 5896 1548
rect 5880 1512 5896 1528
rect 5912 1652 5928 1668
rect 5928 1592 5944 1608
rect 5896 1492 5912 1508
rect 5848 1472 5864 1488
rect 5928 1472 5944 1488
rect 5864 1372 5880 1388
rect 5880 1292 5896 1308
rect 5896 1252 5912 1268
rect 5880 1152 5896 1168
rect 5512 1092 5528 1108
rect 5656 1092 5672 1108
rect 5816 1092 5832 1108
rect 5864 1092 5880 1108
rect 5576 1072 5592 1088
rect 5480 1032 5496 1048
rect 5480 952 5496 968
rect 5416 712 5432 728
rect 5448 712 5464 728
rect 5416 692 5432 708
rect 5480 732 5496 748
rect 5528 732 5544 748
rect 5736 1072 5752 1088
rect 5880 1072 5896 1088
rect 5640 1052 5656 1068
rect 5608 992 5624 1008
rect 5624 972 5640 988
rect 5784 1032 5800 1048
rect 5832 992 5848 1008
rect 5832 932 5848 948
rect 5768 872 5784 888
rect 5688 832 5704 848
rect 5592 732 5608 748
rect 5576 712 5592 728
rect 5448 672 5464 688
rect 5464 672 5480 688
rect 5512 672 5528 688
rect 5432 552 5448 568
rect 5560 552 5576 568
rect 5528 532 5544 548
rect 5544 532 5560 548
rect 5512 492 5528 508
rect 5528 432 5544 448
rect 5496 412 5512 428
rect 5464 372 5480 388
rect 5288 312 5304 328
rect 5320 292 5336 308
rect 5400 292 5416 308
rect 5480 292 5496 308
rect 5496 292 5512 308
rect 5400 272 5416 288
rect 5432 272 5448 288
rect 5560 412 5576 428
rect 5480 252 5528 268
rect 5384 152 5400 168
rect 5528 152 5544 168
rect 5464 132 5480 148
rect 5560 132 5576 148
rect 5656 672 5672 688
rect 5640 592 5656 608
rect 5640 572 5656 588
rect 6104 1832 6120 1848
rect 6045 1802 6081 1818
rect 6088 1812 6104 1828
rect 5976 1752 5992 1768
rect 5976 1732 5992 1748
rect 6072 1714 6088 1728
rect 6072 1712 6088 1714
rect 5960 1692 5976 1708
rect 5944 1452 5960 1468
rect 6152 2092 6168 2108
rect 6248 2272 6264 2288
rect 6264 2272 6280 2288
rect 6392 2272 6424 2288
rect 6280 2252 6296 2268
rect 6392 2252 6408 2268
rect 6248 2212 6264 2228
rect 6472 2252 6488 2268
rect 6696 2672 6712 2688
rect 6888 2712 6904 2728
rect 6792 2706 6808 2708
rect 6792 2692 6808 2706
rect 6888 2692 6904 2708
rect 6856 2672 6872 2688
rect 6824 2652 6840 2668
rect 6728 2532 6744 2548
rect 6808 2532 6824 2548
rect 6856 2532 6872 2548
rect 7048 2892 7064 2908
rect 7000 2872 7016 2888
rect 6968 2712 7000 2728
rect 6936 2632 6952 2648
rect 6936 2592 6952 2608
rect 6936 2572 6952 2588
rect 6952 2532 6968 2548
rect 6744 2512 6760 2528
rect 6712 2492 6728 2508
rect 6792 2472 6808 2488
rect 6520 2312 6536 2328
rect 6488 2232 6504 2248
rect 6504 2212 6520 2228
rect 6440 2172 6456 2188
rect 6728 2432 6744 2448
rect 6728 2412 6744 2428
rect 6568 2372 6584 2388
rect 6648 2372 6664 2388
rect 6632 2272 6648 2288
rect 6584 2252 6600 2268
rect 6264 2112 6280 2128
rect 6504 2114 6520 2128
rect 6504 2112 6520 2114
rect 6216 2092 6232 2108
rect 6184 1952 6200 1968
rect 6168 1732 6184 1748
rect 6136 1652 6152 1668
rect 6136 1612 6152 1628
rect 6056 1512 6072 1528
rect 6008 1412 6024 1428
rect 6045 1402 6081 1418
rect 6024 1352 6040 1368
rect 5944 1052 5960 1068
rect 5928 932 5944 948
rect 5976 1292 5992 1308
rect 6104 1212 6120 1228
rect 6008 1112 6024 1128
rect 5976 1052 5992 1068
rect 5992 972 6008 988
rect 6088 1072 6104 1088
rect 6024 1052 6040 1068
rect 6088 1032 6104 1048
rect 6045 1002 6081 1018
rect 6040 952 6056 968
rect 6104 952 6120 968
rect 6088 932 6104 948
rect 6200 1732 6216 1748
rect 6200 1712 6216 1728
rect 6168 1492 6184 1508
rect 6200 1492 6216 1508
rect 6328 1932 6344 1948
rect 6280 1912 6296 1928
rect 6472 2092 6488 2108
rect 6456 1972 6472 1988
rect 6232 1872 6248 1888
rect 6312 1832 6328 1848
rect 6328 1812 6344 1828
rect 6264 1772 6280 1788
rect 6296 1732 6312 1748
rect 6424 1732 6440 1748
rect 6248 1712 6264 1728
rect 6344 1712 6360 1728
rect 6424 1712 6440 1728
rect 6296 1612 6312 1628
rect 6280 1532 6296 1548
rect 6232 1512 6248 1528
rect 6248 1492 6264 1508
rect 6216 1472 6232 1488
rect 6312 1512 6328 1528
rect 6360 1512 6376 1528
rect 6328 1492 6344 1508
rect 6264 1452 6280 1468
rect 6248 1412 6264 1428
rect 6168 1372 6184 1388
rect 6344 1472 6360 1488
rect 6360 1452 6376 1468
rect 6408 1492 6424 1508
rect 6408 1452 6424 1468
rect 6392 1392 6408 1408
rect 6376 1372 6392 1388
rect 6232 1332 6248 1348
rect 6296 1332 6312 1348
rect 6312 1332 6328 1348
rect 6392 1332 6408 1348
rect 6200 1272 6216 1288
rect 6152 1132 6168 1148
rect 6152 1072 6168 1088
rect 6184 1032 6200 1048
rect 6152 992 6168 1008
rect 6312 1312 6328 1328
rect 6408 1312 6424 1328
rect 6280 1192 6296 1208
rect 6664 2292 6680 2308
rect 6712 2292 6728 2308
rect 6744 2352 6760 2368
rect 6776 2312 6788 2328
rect 6788 2312 6792 2328
rect 6792 2312 6808 2328
rect 6840 2332 6856 2348
rect 6904 2312 6920 2328
rect 6760 2292 6776 2308
rect 6824 2292 6840 2308
rect 6856 2292 6872 2308
rect 6696 2232 6712 2248
rect 6664 2192 6680 2208
rect 6680 2112 6696 2128
rect 6568 1932 6584 1948
rect 6488 1912 6504 1928
rect 6488 1792 6504 1808
rect 6472 1712 6488 1728
rect 6520 1712 6536 1728
rect 6536 1692 6552 1708
rect 6504 1652 6520 1668
rect 6536 1652 6552 1668
rect 6568 1632 6584 1648
rect 6504 1592 6520 1608
rect 6536 1532 6552 1548
rect 6696 1952 6712 1968
rect 6616 1932 6632 1948
rect 6664 1932 6680 1948
rect 6696 1932 6712 1948
rect 6600 1912 6616 1928
rect 6632 1912 6648 1928
rect 6664 1912 6680 1928
rect 6728 1932 6744 1948
rect 6728 1912 6744 1928
rect 6680 1892 6696 1908
rect 6712 1892 6728 1908
rect 6776 2132 6792 2148
rect 6760 1952 6776 1968
rect 6680 1872 6696 1888
rect 6632 1852 6648 1868
rect 6664 1852 6680 1868
rect 6616 1832 6632 1848
rect 6600 1532 6616 1548
rect 6584 1512 6600 1528
rect 6488 1492 6504 1508
rect 6568 1492 6584 1508
rect 6520 1412 6536 1428
rect 6488 1352 6504 1368
rect 6504 1332 6520 1348
rect 6536 1312 6552 1328
rect 6584 1452 6600 1468
rect 6584 1432 6600 1448
rect 6568 1412 6584 1428
rect 6664 1592 6680 1608
rect 6664 1512 6680 1528
rect 6632 1492 6648 1508
rect 6664 1492 6680 1508
rect 6744 1732 6760 1748
rect 6696 1712 6712 1728
rect 6744 1692 6760 1708
rect 6792 1892 6808 1908
rect 6920 2292 6936 2308
rect 6888 2232 6904 2248
rect 6840 2172 6856 2188
rect 6920 2132 6936 2148
rect 6840 2114 6856 2128
rect 6840 2112 6856 2114
rect 6840 1912 6856 1928
rect 6920 1912 6936 1928
rect 6904 1892 6920 1908
rect 7053 2802 7089 2818
rect 7016 2712 7032 2728
rect 7032 2652 7048 2668
rect 7000 2572 7016 2588
rect 7048 2572 7064 2588
rect 7064 2532 7080 2548
rect 7016 2512 7032 2528
rect 6984 2492 7000 2508
rect 7032 2492 7048 2508
rect 6984 2452 7000 2468
rect 6952 2352 6968 2368
rect 7128 3272 7144 3288
rect 7192 3232 7208 3248
rect 7432 4532 7448 4548
rect 7336 4512 7352 4528
rect 7432 4492 7448 4508
rect 7480 4652 7496 4668
rect 7464 4512 7480 4528
rect 7496 4572 7512 4588
rect 7480 4492 7496 4508
rect 7448 4452 7464 4468
rect 7416 4372 7432 4388
rect 7400 4352 7416 4368
rect 7336 4332 7352 4348
rect 7368 4292 7384 4308
rect 7368 4252 7384 4268
rect 7400 4252 7416 4268
rect 7480 4312 7496 4328
rect 7576 4672 7592 4688
rect 7560 4652 7576 4668
rect 7768 5292 7784 5308
rect 7784 5272 7800 5288
rect 7784 5252 7800 5268
rect 7704 5172 7720 5188
rect 7704 5132 7720 5148
rect 7752 5092 7768 5108
rect 7672 5072 7688 5088
rect 7640 5032 7656 5048
rect 7768 5032 7784 5048
rect 7656 5012 7672 5028
rect 7656 4972 7672 4988
rect 7624 4952 7640 4968
rect 7928 5372 7944 5388
rect 7896 5352 7912 5368
rect 7832 5252 7848 5268
rect 7880 5112 7896 5128
rect 7832 5072 7848 5088
rect 7912 5052 7928 5068
rect 7848 5012 7864 5028
rect 7864 4992 7880 5008
rect 7976 5072 7992 5088
rect 7944 4972 7960 4988
rect 7992 4952 8008 4968
rect 7832 4932 7848 4948
rect 7896 4932 7912 4948
rect 7688 4912 7704 4928
rect 7720 4914 7736 4928
rect 7720 4912 7736 4914
rect 7864 4912 7880 4928
rect 7656 4852 7672 4868
rect 7608 4752 7624 4768
rect 7608 4712 7624 4728
rect 7896 4892 7912 4908
rect 7896 4872 7912 4888
rect 7800 4812 7816 4828
rect 7816 4712 7832 4728
rect 7736 4692 7752 4708
rect 7784 4692 7816 4708
rect 7544 4552 7560 4568
rect 7704 4672 7720 4688
rect 7672 4612 7688 4628
rect 7656 4592 7672 4608
rect 7720 4572 7736 4588
rect 7624 4532 7640 4548
rect 7528 4512 7544 4528
rect 7512 4432 7528 4448
rect 7560 4312 7576 4328
rect 7448 4292 7464 4308
rect 7512 4272 7528 4288
rect 7544 4272 7560 4288
rect 7496 4252 7512 4268
rect 7864 4672 7880 4688
rect 7832 4572 7848 4588
rect 7784 4532 7800 4548
rect 7592 4492 7608 4508
rect 7640 4492 7656 4508
rect 7736 4492 7752 4508
rect 7624 4312 7640 4328
rect 7928 4912 7944 4928
rect 8024 4912 8040 4928
rect 7976 4892 7992 4908
rect 7944 4872 7960 4888
rect 7912 4832 7928 4848
rect 7992 4712 8008 4728
rect 7912 4692 7928 4708
rect 7960 4692 7976 4708
rect 7992 4692 8008 4708
rect 7976 4592 7992 4608
rect 7912 4372 7928 4388
rect 7576 4212 7592 4228
rect 7512 4172 7528 4188
rect 7464 4112 7480 4128
rect 7544 4112 7560 4128
rect 7576 4112 7592 4128
rect 7416 4092 7432 4108
rect 7512 4092 7528 4108
rect 7448 3932 7464 3948
rect 7400 3912 7416 3928
rect 7528 3912 7544 3928
rect 7592 4092 7608 4108
rect 7592 3912 7608 3928
rect 7576 3892 7592 3908
rect 7480 3872 7496 3888
rect 7512 3872 7528 3888
rect 7544 3872 7560 3888
rect 7592 3872 7608 3888
rect 7544 3752 7560 3768
rect 7720 4272 7736 4288
rect 7704 4252 7720 4268
rect 7688 4212 7704 4228
rect 7672 4132 7688 4148
rect 7800 4232 7816 4248
rect 7640 4112 7656 4128
rect 7624 4092 7640 4108
rect 7688 3952 7704 3968
rect 7640 3912 7656 3928
rect 7944 4372 7960 4388
rect 7928 4152 7944 4168
rect 7816 4132 7832 4148
rect 7720 4112 7736 4128
rect 7800 4112 7816 4128
rect 7720 4092 7736 4108
rect 7768 3912 7784 3928
rect 7960 4352 7976 4368
rect 7960 4292 7976 4308
rect 8024 4372 8040 4388
rect 8024 4352 8040 4368
rect 8008 4292 8024 4308
rect 7976 4152 7992 4168
rect 7928 4112 7944 4128
rect 7944 4112 7960 4128
rect 8008 4112 8024 4128
rect 7896 3932 7912 3948
rect 7640 3892 7656 3908
rect 7704 3892 7720 3908
rect 7640 3872 7656 3888
rect 7608 3852 7624 3868
rect 7704 3852 7720 3868
rect 7688 3832 7704 3848
rect 7336 3732 7352 3748
rect 7688 3732 7704 3748
rect 7368 3712 7384 3728
rect 7448 3652 7464 3668
rect 7624 3692 7640 3708
rect 7528 3632 7544 3648
rect 7592 3632 7608 3648
rect 7416 3552 7432 3568
rect 7480 3552 7496 3568
rect 7448 3532 7464 3548
rect 7480 3532 7496 3548
rect 7560 3532 7576 3548
rect 7336 3512 7352 3528
rect 7432 3512 7464 3528
rect 7320 3492 7336 3508
rect 7272 3452 7288 3468
rect 7288 3432 7304 3448
rect 7240 3312 7256 3328
rect 7224 3292 7228 3308
rect 7228 3292 7240 3308
rect 7272 3272 7288 3288
rect 7256 3252 7272 3268
rect 7208 3172 7224 3188
rect 7144 3132 7160 3148
rect 7208 3132 7224 3148
rect 7112 3072 7128 3088
rect 7144 3072 7160 3088
rect 7160 2914 7176 2928
rect 7160 2912 7176 2914
rect 7176 2712 7188 2728
rect 7188 2712 7192 2728
rect 7160 2692 7176 2708
rect 7208 2692 7224 2708
rect 7128 2672 7144 2688
rect 7144 2572 7160 2588
rect 7192 2512 7208 2528
rect 7096 2452 7112 2468
rect 7048 2432 7064 2448
rect 7528 3492 7544 3508
rect 7544 3492 7560 3508
rect 7816 3872 7832 3888
rect 7752 3852 7768 3868
rect 7704 3692 7720 3708
rect 7656 3672 7672 3688
rect 7752 3632 7768 3648
rect 7736 3612 7752 3628
rect 7656 3492 7672 3508
rect 7544 3472 7560 3488
rect 7576 3472 7592 3488
rect 7640 3472 7656 3488
rect 7336 3352 7352 3368
rect 7400 3452 7416 3468
rect 7480 3372 7496 3388
rect 7384 3312 7400 3328
rect 7432 3292 7448 3308
rect 7304 3272 7320 3288
rect 7560 3292 7576 3308
rect 7560 3272 7576 3288
rect 7544 3252 7560 3268
rect 7560 3132 7576 3148
rect 7480 3112 7496 3128
rect 7672 3372 7688 3388
rect 7736 3372 7752 3388
rect 7608 3332 7624 3348
rect 7752 3332 7768 3348
rect 7624 3292 7640 3308
rect 7656 3272 7672 3288
rect 7592 3252 7608 3268
rect 7688 3192 7704 3208
rect 7848 3732 7864 3748
rect 7784 3432 7800 3448
rect 7816 3632 7832 3648
rect 7880 3612 7896 3628
rect 7800 3372 7816 3388
rect 7880 3332 7896 3348
rect 7880 3312 7896 3328
rect 7832 3272 7848 3288
rect 7816 3232 7832 3248
rect 7800 3172 7816 3188
rect 7768 3152 7784 3168
rect 7688 3132 7704 3148
rect 7752 3132 7768 3148
rect 7800 3132 7816 3148
rect 7608 3112 7624 3128
rect 7624 3112 7640 3128
rect 7672 3112 7688 3128
rect 7784 3112 7800 3128
rect 7544 2992 7560 3008
rect 7576 2992 7592 3008
rect 7320 2932 7336 2948
rect 7352 2932 7368 2948
rect 7464 2932 7480 2948
rect 7304 2892 7320 2908
rect 7288 2832 7304 2848
rect 7256 2672 7272 2688
rect 7224 2652 7240 2668
rect 7288 2652 7304 2668
rect 7336 2912 7352 2928
rect 7448 2712 7464 2728
rect 7432 2692 7448 2708
rect 7480 2712 7496 2728
rect 7448 2672 7464 2688
rect 7336 2632 7352 2648
rect 7053 2402 7089 2418
rect 7208 2412 7224 2428
rect 7144 2292 7160 2308
rect 7272 2292 7288 2308
rect 6984 2252 7000 2268
rect 7096 2252 7112 2268
rect 7192 2272 7208 2288
rect 7160 2232 7176 2248
rect 7128 2192 7144 2208
rect 7000 2172 7016 2188
rect 6952 2112 6968 2128
rect 7160 2132 7176 2148
rect 7256 2252 7272 2268
rect 7320 2252 7336 2268
rect 7240 2212 7256 2228
rect 6952 2092 6968 2108
rect 7000 2092 7032 2108
rect 6936 1892 6968 1908
rect 7000 1892 7016 1908
rect 7053 2002 7089 2018
rect 7032 1912 7048 1928
rect 7064 1892 7080 1908
rect 6808 1872 6824 1888
rect 7000 1872 7016 1888
rect 6776 1852 6792 1868
rect 6808 1712 6824 1728
rect 6824 1692 6840 1708
rect 6792 1572 6808 1588
rect 6776 1532 6792 1548
rect 6760 1512 6776 1528
rect 6792 1492 6808 1508
rect 6680 1452 6696 1468
rect 6728 1432 6744 1448
rect 6744 1412 6760 1428
rect 6616 1314 6632 1328
rect 6616 1312 6632 1314
rect 6792 1332 6808 1348
rect 6536 1252 6552 1268
rect 6520 1112 6536 1128
rect 6232 1092 6248 1108
rect 6360 1092 6376 1108
rect 6408 1092 6424 1108
rect 6264 1072 6280 1088
rect 6328 1072 6344 1088
rect 6248 1032 6264 1048
rect 6392 1032 6408 1048
rect 6232 1012 6248 1028
rect 6392 992 6408 1008
rect 6216 972 6232 988
rect 6248 952 6280 968
rect 6792 1292 6808 1308
rect 7016 1852 7032 1868
rect 6952 1752 6968 1768
rect 7032 1752 7048 1768
rect 7000 1732 7016 1748
rect 7192 1932 7208 1948
rect 7160 1872 7176 1888
rect 7096 1752 7112 1768
rect 7288 2192 7320 2208
rect 7480 2612 7496 2628
rect 7512 2592 7528 2608
rect 7400 2512 7416 2528
rect 7480 2512 7496 2528
rect 7352 2472 7368 2488
rect 7416 2472 7432 2488
rect 7512 2472 7528 2488
rect 7480 2432 7496 2448
rect 7384 2352 7400 2368
rect 7400 2312 7416 2328
rect 7464 2312 7480 2328
rect 7352 2272 7368 2288
rect 7352 2252 7368 2268
rect 7336 1912 7352 1928
rect 7400 2232 7416 2248
rect 7368 2192 7384 2208
rect 7400 2172 7416 2188
rect 7400 2114 7416 2128
rect 7400 2112 7416 2114
rect 7432 2112 7448 2128
rect 7704 3052 7720 3068
rect 7800 3012 7816 3028
rect 7768 2992 7784 3008
rect 7720 2972 7736 2988
rect 7640 2932 7656 2948
rect 7656 2932 7672 2948
rect 7608 2912 7640 2928
rect 7672 2912 7688 2928
rect 7640 2892 7656 2908
rect 7592 2872 7608 2888
rect 7624 2852 7640 2868
rect 7576 2512 7592 2528
rect 7544 2352 7560 2368
rect 7560 2332 7576 2348
rect 7496 2272 7512 2288
rect 7544 2272 7560 2288
rect 7480 2212 7496 2228
rect 7496 2112 7528 2128
rect 7400 2072 7416 2088
rect 7464 2072 7496 2088
rect 7496 1912 7512 1928
rect 7400 1892 7416 1908
rect 7512 1892 7528 1908
rect 7448 1872 7464 1888
rect 7256 1812 7272 1828
rect 7240 1772 7256 1788
rect 7224 1752 7240 1768
rect 7160 1732 7176 1748
rect 6904 1692 6920 1708
rect 7032 1692 7048 1708
rect 7080 1672 7096 1688
rect 7053 1602 7089 1618
rect 7064 1572 7080 1588
rect 6888 1512 6904 1528
rect 6952 1512 6968 1528
rect 6984 1512 7000 1528
rect 6856 1472 6872 1488
rect 6872 1452 6888 1468
rect 6904 1452 6920 1468
rect 6888 1372 6904 1388
rect 6936 1452 6952 1468
rect 6920 1352 6936 1368
rect 6936 1332 6952 1348
rect 6856 1312 6872 1328
rect 6808 1272 6824 1288
rect 6776 1212 6792 1228
rect 6920 1312 6936 1328
rect 6888 1272 6904 1288
rect 6904 1192 6920 1208
rect 6824 1172 6840 1188
rect 6872 1172 6888 1188
rect 6616 1112 6632 1128
rect 6568 1092 6584 1108
rect 6728 1106 6744 1108
rect 6728 1092 6744 1106
rect 6648 1072 6664 1088
rect 6792 1072 6808 1088
rect 6440 1052 6456 1068
rect 6584 1052 6600 1068
rect 6696 1052 6712 1068
rect 6744 1052 6760 1068
rect 6536 1012 6552 1028
rect 6504 992 6520 1008
rect 6504 972 6520 988
rect 6536 972 6552 988
rect 6520 952 6536 968
rect 6264 932 6280 948
rect 6280 932 6296 948
rect 6376 932 6392 948
rect 6408 932 6424 948
rect 6008 912 6024 928
rect 5912 852 5928 868
rect 5816 772 5832 788
rect 5848 712 5864 728
rect 5784 692 5800 708
rect 5736 672 5752 688
rect 5816 672 5832 688
rect 5672 552 5704 568
rect 5608 512 5624 528
rect 5688 512 5704 528
rect 5656 492 5672 508
rect 5656 312 5688 328
rect 5608 272 5624 288
rect 5624 152 5640 168
rect 5784 632 5800 648
rect 5736 512 5752 528
rect 5816 514 5832 528
rect 5816 512 5832 514
rect 5736 492 5752 508
rect 5864 692 5880 708
rect 5880 632 5896 648
rect 5976 892 5992 908
rect 6136 892 6152 908
rect 6312 892 6328 908
rect 6120 852 6136 868
rect 6152 852 6168 868
rect 6632 1032 6648 1048
rect 6472 912 6488 928
rect 6488 912 6504 928
rect 6552 912 6568 928
rect 6168 832 6184 848
rect 6328 832 6344 848
rect 6264 792 6280 808
rect 6152 772 6168 788
rect 5976 732 6008 748
rect 5928 672 5944 688
rect 5880 572 5896 588
rect 5864 532 5880 548
rect 6072 692 6088 708
rect 6136 692 6152 708
rect 6045 602 6081 618
rect 5976 512 5992 528
rect 5912 352 5928 368
rect 5880 312 5896 328
rect 5720 292 5736 308
rect 5720 192 5736 208
rect 5944 252 5960 268
rect 5832 172 5848 188
rect 5736 152 5752 168
rect 5656 132 5672 148
rect 5704 132 5720 148
rect 6216 732 6248 748
rect 6184 632 6200 648
rect 6168 512 6184 528
rect 6024 252 6040 268
rect 6008 232 6024 248
rect 6104 232 6120 248
rect 5992 212 6008 228
rect 6008 192 6024 208
rect 6045 202 6081 218
rect 6104 212 6120 228
rect 5960 152 5976 168
rect 5992 152 6008 168
rect 6072 152 6088 168
rect 6392 732 6408 748
rect 6504 872 6520 888
rect 6232 692 6248 708
rect 6264 692 6280 708
rect 6312 692 6328 708
rect 6360 692 6376 708
rect 6472 692 6488 708
rect 6280 672 6296 688
rect 6344 672 6360 688
rect 6280 612 6296 628
rect 6216 592 6232 608
rect 6296 592 6312 608
rect 6312 532 6328 548
rect 6280 512 6296 528
rect 6200 492 6216 508
rect 6264 492 6280 508
rect 6488 672 6504 688
rect 6376 652 6392 668
rect 6568 892 6584 908
rect 6600 912 6616 928
rect 6600 892 6616 908
rect 6648 952 6664 968
rect 6728 952 6744 968
rect 6648 932 6664 948
rect 6696 932 6712 948
rect 6760 952 6776 968
rect 6888 1132 6904 1148
rect 6920 1072 6936 1088
rect 7048 1492 7064 1508
rect 7048 1472 7064 1488
rect 7096 1492 7112 1508
rect 7080 1472 7096 1488
rect 6968 1452 6984 1468
rect 7032 1452 7048 1468
rect 7064 1452 7080 1468
rect 6968 1352 6984 1368
rect 6984 1332 7000 1348
rect 7053 1202 7089 1218
rect 7048 1172 7064 1188
rect 6952 1112 6968 1128
rect 7016 1112 7032 1128
rect 6984 1092 7000 1108
rect 6984 1072 7000 1088
rect 6872 1052 6888 1068
rect 6888 1052 6904 1068
rect 6936 1052 6952 1068
rect 6856 972 6872 988
rect 6936 1032 6952 1048
rect 6888 952 6904 968
rect 6824 932 6840 948
rect 6872 932 6888 948
rect 6776 912 6792 928
rect 6840 912 6856 928
rect 6904 912 6920 928
rect 6952 912 6968 928
rect 6824 892 6840 908
rect 6712 872 6728 888
rect 6760 872 6776 888
rect 6856 852 6872 868
rect 6680 832 6696 848
rect 6760 832 6776 848
rect 6664 792 6680 808
rect 6584 752 6600 768
rect 6760 752 6776 768
rect 6744 732 6760 748
rect 6616 672 6632 688
rect 6584 632 6600 648
rect 6376 532 6392 548
rect 6504 532 6520 548
rect 6456 514 6472 528
rect 6456 512 6472 514
rect 6344 492 6348 508
rect 6348 492 6360 508
rect 6344 452 6360 468
rect 6392 332 6408 348
rect 6392 312 6408 328
rect 6312 252 6328 268
rect 6200 192 6216 208
rect 6184 172 6200 188
rect 6216 172 6232 188
rect 6312 152 6328 168
rect 6648 652 6664 668
rect 6600 592 6616 608
rect 6632 592 6648 608
rect 6552 452 6568 468
rect 6728 672 6744 688
rect 6680 592 6696 608
rect 6712 532 6728 548
rect 6584 352 6600 368
rect 6520 312 6536 328
rect 6488 292 6504 308
rect 6360 192 6392 208
rect 6456 212 6472 228
rect 6440 172 6456 188
rect 5960 132 5976 148
rect 6040 132 6056 148
rect 6328 132 6344 148
rect 6408 132 6424 148
rect 4968 112 4984 128
rect 5208 114 5224 128
rect 5208 112 5224 114
rect 5272 112 5288 128
rect 5496 112 5512 128
rect 5592 112 5608 128
rect 5688 112 5704 128
rect 5832 112 5848 128
rect 6504 152 6520 168
rect 6568 132 6584 148
rect 6632 352 6648 368
rect 6648 312 6664 328
rect 6616 292 6632 308
rect 6600 272 6616 288
rect 6696 272 6712 288
rect 6616 212 6632 228
rect 6616 192 6632 208
rect 6616 152 6632 168
rect 6744 492 6760 508
rect 6728 352 6744 368
rect 6824 692 6840 708
rect 6792 672 6808 688
rect 6904 792 6920 808
rect 6936 892 6952 908
rect 7080 1152 7096 1168
rect 7128 1452 7144 1468
rect 7128 1392 7144 1408
rect 7096 1132 7112 1148
rect 7112 1072 7128 1088
rect 7112 992 7128 1008
rect 7064 932 7080 948
rect 7032 912 7048 928
rect 7000 892 7016 908
rect 7096 892 7112 908
rect 6984 832 7000 848
rect 7053 802 7089 818
rect 7016 712 7032 728
rect 7032 692 7048 708
rect 7112 692 7128 708
rect 6808 612 6824 628
rect 6888 632 6904 648
rect 6904 552 6920 568
rect 7016 532 7032 548
rect 6904 452 6920 468
rect 6856 432 6872 448
rect 6840 332 6856 348
rect 6888 332 6904 348
rect 6952 292 6968 308
rect 6776 252 6792 268
rect 6936 272 6952 288
rect 7064 592 7080 608
rect 6984 512 7000 528
rect 7032 512 7048 528
rect 7000 492 7016 508
rect 7016 472 7032 488
rect 6984 332 7000 348
rect 7053 402 7089 418
rect 7240 1732 7256 1748
rect 7240 1672 7256 1688
rect 7336 1792 7352 1808
rect 7288 1712 7304 1728
rect 7176 1512 7192 1528
rect 7224 1512 7256 1528
rect 7320 1692 7336 1708
rect 7336 1652 7352 1668
rect 7256 1492 7272 1508
rect 7256 1452 7272 1468
rect 7224 1332 7240 1348
rect 7240 1152 7256 1168
rect 7144 1112 7160 1128
rect 7144 1072 7160 1088
rect 7208 1072 7224 1088
rect 7176 892 7192 908
rect 7288 1472 7304 1488
rect 7304 1352 7320 1368
rect 7272 1172 7288 1188
rect 7336 1212 7352 1228
rect 7464 1812 7480 1828
rect 7464 1792 7480 1808
rect 7432 1752 7448 1768
rect 7368 1732 7384 1748
rect 7704 2872 7720 2888
rect 7672 2572 7688 2588
rect 7704 2572 7720 2588
rect 7688 2552 7704 2568
rect 7640 2532 7656 2548
rect 7592 2492 7608 2508
rect 7608 2452 7624 2468
rect 7736 2912 7752 2928
rect 7784 2872 7800 2888
rect 7752 2852 7768 2868
rect 7864 3212 7880 3228
rect 7832 3132 7848 3148
rect 7960 3832 7976 3848
rect 8040 4172 8056 4188
rect 7928 3692 7944 3708
rect 7928 3652 7944 3668
rect 8040 3652 8056 3668
rect 7912 3352 7928 3368
rect 7912 3272 7928 3288
rect 7896 3232 7912 3248
rect 7896 3172 7912 3188
rect 7864 3112 7880 3128
rect 7832 3092 7848 3108
rect 7848 3072 7864 3088
rect 7912 3152 7928 3168
rect 7880 3052 7896 3068
rect 7880 2912 7896 2928
rect 7816 2652 7832 2668
rect 7784 2612 7800 2628
rect 7784 2552 7800 2568
rect 7640 2512 7656 2528
rect 7624 2432 7640 2448
rect 7624 2392 7640 2408
rect 7688 2492 7704 2508
rect 7672 2412 7688 2428
rect 7656 2372 7672 2388
rect 7656 2352 7672 2368
rect 7640 2312 7656 2328
rect 7608 2292 7624 2308
rect 7576 2192 7592 2208
rect 7576 2152 7592 2168
rect 7560 2112 7576 2128
rect 7736 2472 7752 2488
rect 7896 2892 7912 2908
rect 7976 3512 7992 3528
rect 8024 3332 8040 3348
rect 7992 3312 8008 3328
rect 7976 3292 7992 3308
rect 7944 3272 7960 3288
rect 7960 3192 7976 3208
rect 7992 3232 8008 3248
rect 7864 2612 7880 2628
rect 8008 3132 8024 3148
rect 7976 2612 7992 2628
rect 7864 2512 7880 2528
rect 7928 2512 7944 2528
rect 7944 2512 7960 2528
rect 7944 2452 7960 2468
rect 7704 2412 7720 2428
rect 7784 2412 7800 2428
rect 7848 2332 7864 2348
rect 8024 2512 8040 2528
rect 7992 2392 8008 2408
rect 7816 2292 7832 2308
rect 7720 2272 7736 2288
rect 7704 2192 7720 2208
rect 7656 2132 7672 2148
rect 7592 2112 7608 2128
rect 7672 2112 7688 2128
rect 7656 2092 7672 2108
rect 7592 2072 7608 2088
rect 7624 2072 7640 2088
rect 7624 1952 7640 1968
rect 7688 1952 7704 1968
rect 7656 1892 7672 1908
rect 7592 1872 7608 1888
rect 7528 1852 7544 1868
rect 7512 1752 7528 1768
rect 7448 1732 7464 1748
rect 7528 1732 7544 1748
rect 7496 1712 7512 1728
rect 7544 1712 7560 1728
rect 7400 1692 7416 1708
rect 7416 1692 7432 1708
rect 7496 1692 7508 1708
rect 7508 1692 7512 1708
rect 7400 1672 7416 1688
rect 7384 1472 7400 1488
rect 7368 1372 7384 1388
rect 7352 1152 7368 1168
rect 7304 1132 7320 1148
rect 7288 1072 7304 1088
rect 7384 1072 7400 1088
rect 7336 992 7352 1008
rect 7512 1672 7528 1688
rect 7544 1672 7560 1688
rect 7496 1652 7512 1668
rect 7416 1492 7432 1508
rect 7464 1492 7480 1508
rect 7464 1472 7480 1488
rect 7464 1332 7480 1348
rect 7416 1152 7432 1168
rect 7448 1132 7464 1148
rect 7512 1632 7528 1648
rect 7576 1512 7592 1528
rect 7640 1852 7656 1868
rect 7688 1692 7704 1708
rect 7752 2132 7768 2148
rect 7880 2132 7896 2148
rect 7720 1932 7736 1948
rect 7768 2072 7800 2088
rect 7976 2172 7992 2188
rect 7880 2112 7896 2128
rect 7880 2092 7896 2108
rect 7912 2092 7928 2108
rect 7848 2032 7864 2048
rect 7832 1952 7848 1968
rect 7816 1912 7832 1928
rect 7784 1892 7800 1908
rect 7768 1852 7784 1868
rect 7752 1792 7768 1808
rect 7736 1772 7752 1788
rect 7928 2072 7944 2088
rect 7944 1932 7960 1948
rect 7928 1912 7944 1928
rect 7896 1712 7912 1728
rect 7704 1532 7720 1548
rect 7768 1532 7784 1548
rect 7608 1512 7624 1528
rect 7736 1512 7748 1528
rect 7748 1512 7752 1528
rect 7592 1492 7608 1508
rect 7608 1492 7624 1508
rect 7688 1492 7704 1508
rect 7544 1472 7560 1488
rect 7704 1452 7720 1468
rect 7576 1432 7592 1448
rect 7624 1432 7640 1448
rect 7704 1432 7720 1448
rect 7512 1352 7528 1368
rect 7656 1372 7672 1388
rect 7496 1332 7512 1348
rect 7480 1252 7496 1268
rect 7480 1152 7496 1168
rect 7576 1312 7592 1328
rect 7592 1312 7608 1328
rect 7512 1292 7528 1308
rect 7608 1292 7624 1308
rect 7576 1252 7592 1268
rect 7512 1212 7528 1228
rect 7544 1072 7560 1088
rect 7544 992 7560 1008
rect 7736 1352 7752 1368
rect 7688 1312 7704 1328
rect 7752 1312 7768 1328
rect 7688 1292 7704 1308
rect 7672 1172 7688 1188
rect 7736 1152 7752 1168
rect 7640 1132 7656 1148
rect 7704 1072 7720 1088
rect 7704 1052 7720 1068
rect 7608 992 7624 1008
rect 7608 952 7624 968
rect 7512 932 7528 948
rect 7272 912 7288 928
rect 7240 892 7256 908
rect 7208 852 7224 868
rect 7144 812 7160 828
rect 7320 772 7336 788
rect 7192 732 7208 748
rect 7160 712 7176 728
rect 7240 712 7256 728
rect 7208 692 7224 708
rect 7256 692 7272 708
rect 7160 672 7176 688
rect 7224 672 7240 688
rect 7208 532 7224 548
rect 7016 312 7032 328
rect 7128 312 7144 328
rect 7032 292 7048 308
rect 7048 292 7064 308
rect 7128 292 7160 308
rect 7160 272 7176 288
rect 7224 252 7240 268
rect 6968 212 6984 228
rect 6952 172 6968 188
rect 6760 152 6776 168
rect 6824 152 6840 168
rect 6888 152 6904 168
rect 6968 152 6984 168
rect 7224 152 7240 168
rect 6712 132 6728 148
rect 6920 132 6936 148
rect 7096 132 7112 148
rect 7176 132 7192 148
rect 7720 932 7736 948
rect 7704 872 7720 888
rect 7640 852 7656 868
rect 7512 812 7528 828
rect 7336 732 7352 748
rect 7464 732 7480 748
rect 7480 712 7496 728
rect 7368 532 7384 548
rect 7448 532 7464 548
rect 7272 292 7288 308
rect 7368 492 7384 508
rect 7336 472 7352 488
rect 7432 432 7448 448
rect 7672 712 7688 728
rect 7656 692 7672 708
rect 7688 692 7704 708
rect 7736 692 7752 708
rect 7624 672 7640 688
rect 7544 552 7560 568
rect 7544 472 7560 488
rect 7656 372 7672 388
rect 7576 332 7592 348
rect 7656 312 7672 328
rect 7704 312 7720 328
rect 7464 292 7480 308
rect 7512 292 7528 308
rect 7544 292 7560 308
rect 7592 292 7608 308
rect 7320 172 7336 188
rect 7864 1512 7880 1528
rect 7848 1472 7864 1488
rect 7800 1352 7816 1368
rect 7816 1332 7832 1348
rect 7864 1332 7880 1348
rect 7768 1292 7784 1308
rect 7784 1152 7800 1168
rect 7768 1132 7800 1148
rect 7768 832 7784 848
rect 7832 1312 7848 1328
rect 7992 2032 8008 2048
rect 7960 1632 7976 1648
rect 7944 1332 7960 1348
rect 7960 1312 7976 1328
rect 7880 1272 7896 1288
rect 7848 1232 7864 1248
rect 7832 1212 7848 1228
rect 7864 1172 7880 1188
rect 7848 1152 7864 1168
rect 7944 1292 7960 1308
rect 7896 1132 7912 1148
rect 7880 1112 7896 1128
rect 7912 1092 7928 1108
rect 7832 1052 7848 1068
rect 7832 1032 7848 1048
rect 7832 932 7848 948
rect 7896 914 7912 928
rect 7896 912 7912 914
rect 7848 732 7864 748
rect 7768 672 7784 688
rect 7768 572 7784 588
rect 7944 1032 7960 1048
rect 7992 1492 8008 1508
rect 8024 1492 8040 1508
rect 7992 1092 8008 1108
rect 7992 1052 8008 1068
rect 7976 692 7992 708
rect 7912 652 7928 668
rect 7976 652 7992 668
rect 7800 572 7816 588
rect 7848 552 7864 568
rect 7800 512 7816 528
rect 7880 514 7896 528
rect 7880 512 7896 514
rect 7784 312 7800 328
rect 7768 292 7784 308
rect 7864 306 7880 308
rect 7864 292 7880 306
rect 7608 272 7624 288
rect 7720 272 7736 288
rect 7416 252 7432 268
rect 7624 252 7640 268
rect 7752 252 7768 268
rect 7560 232 7576 248
rect 7640 232 7656 248
rect 7672 232 7688 248
rect 7512 172 7528 188
rect 7544 172 7560 188
rect 7464 152 7480 168
rect 7288 132 7304 148
rect 7864 232 7880 248
rect 7720 132 7736 148
rect 7832 132 7848 148
rect 8024 1072 8040 1088
rect 8008 952 8024 968
rect 8008 672 8024 688
rect 6328 112 6344 128
rect 6376 112 6392 128
rect 6520 112 6536 128
rect 6584 112 6600 128
rect 6856 112 6872 128
rect 6936 112 6952 128
rect 7256 112 7272 128
rect 7304 112 7320 128
rect 4120 92 4136 108
rect 4296 92 4312 108
rect 4552 92 4568 108
rect 5592 92 5608 108
rect 5960 92 5976 108
rect 6024 92 6028 108
rect 6028 92 6040 108
rect 6200 92 6216 108
rect 7288 92 7304 108
rect 7416 92 7432 108
rect 4328 12 4344 28
rect 5021 2 5057 18
rect 7053 2 7089 18
<< metal3 >>
rect 3032 5617 3048 5623
rect 1656 5517 1912 5523
rect 2232 5517 2456 5523
rect 3496 5517 3624 5523
rect 4584 5517 4696 5523
rect 5064 5517 5112 5523
rect 5128 5517 5176 5523
rect 6984 5517 7144 5523
rect 7656 5517 7736 5523
rect 392 5497 520 5503
rect 760 5497 776 5503
rect 792 5497 824 5503
rect 968 5497 1064 5503
rect 2072 5497 2136 5503
rect 2168 5497 2232 5503
rect 2488 5497 2584 5503
rect 3080 5497 3112 5503
rect 3608 5497 3640 5503
rect 3656 5497 3752 5503
rect 4696 5497 4792 5503
rect 4920 5497 5064 5503
rect 5224 5497 5368 5503
rect 5864 5497 5928 5503
rect 6024 5497 6232 5503
rect 6600 5497 6744 5503
rect 6952 5497 7016 5503
rect 7768 5497 7864 5503
rect 77 5488 83 5492
rect 248 5477 392 5483
rect 664 5477 760 5483
rect 1112 5477 1304 5483
rect 1320 5477 1336 5483
rect 1352 5477 1432 5483
rect 1608 5477 1784 5483
rect 1848 5477 2072 5483
rect 2104 5477 2280 5483
rect 2296 5477 2440 5483
rect 2520 5477 2728 5483
rect 3400 5477 3560 5483
rect 3736 5477 3896 5483
rect 3992 5477 4328 5483
rect 4664 5477 4728 5483
rect 5032 5477 5128 5483
rect 5192 5477 5240 5483
rect 5288 5477 5368 5483
rect 5384 5477 5448 5483
rect 6008 5477 6088 5483
rect 6104 5477 6568 5483
rect 6584 5477 6632 5483
rect 6680 5477 6808 5483
rect 6920 5477 7032 5483
rect 7736 5477 7800 5483
rect 600 5457 792 5463
rect 888 5457 1080 5463
rect 1096 5457 1128 5463
rect 1576 5457 1592 5463
rect 2024 5457 2200 5463
rect 4168 5457 4424 5463
rect 4568 5457 5384 5463
rect 5400 5457 5608 5463
rect 5864 5457 5928 5463
rect 5944 5457 5960 5463
rect 6008 5457 6248 5463
rect 6264 5457 6312 5463
rect 6328 5457 6456 5463
rect 6472 5457 6568 5463
rect 6584 5457 6712 5463
rect 7704 5457 7800 5463
rect 1688 5437 2184 5443
rect 3432 5437 4296 5443
rect 5912 5437 5944 5443
rect 6376 5437 6552 5443
rect 6568 5437 6936 5443
rect 6952 5437 6984 5443
rect 7725 5428 7731 5432
rect 360 5397 728 5403
rect 744 5397 984 5403
rect 1000 5397 1939 5403
rect 2136 5417 2200 5423
rect 152 5377 328 5383
rect 344 5377 424 5383
rect 1336 5377 1528 5383
rect 1933 5383 1939 5397
rect 2312 5397 2328 5403
rect 2408 5397 2488 5403
rect 3256 5397 3688 5403
rect 5896 5417 5992 5423
rect 7416 5397 7560 5403
rect 7656 5397 7784 5403
rect 1933 5377 2632 5383
rect 2648 5377 3672 5383
rect 4072 5377 4200 5383
rect 5048 5377 5320 5383
rect 5528 5377 5592 5383
rect 6264 5377 6440 5383
rect 7512 5377 7592 5383
rect 7608 5377 7928 5383
rect 104 5357 216 5363
rect 232 5357 264 5363
rect 536 5357 584 5363
rect 824 5357 888 5363
rect 1000 5357 1096 5363
rect 1112 5357 1224 5363
rect 1416 5357 1480 5363
rect 1512 5357 1656 5363
rect 1944 5357 2136 5363
rect 3560 5357 3944 5363
rect 3960 5357 4088 5363
rect 4648 5357 4888 5363
rect 5256 5357 5592 5363
rect 5944 5357 6296 5363
rect 7704 5357 7896 5363
rect 168 5337 248 5343
rect 856 5337 968 5343
rect 984 5337 1576 5343
rect 1592 5337 1624 5343
rect 1736 5337 1784 5343
rect 1800 5337 1928 5343
rect 2040 5337 2216 5343
rect 2232 5337 2264 5343
rect 2280 5337 2488 5343
rect 2600 5337 3016 5343
rect 3320 5337 3336 5343
rect 3736 5337 4168 5343
rect 4424 5337 4664 5343
rect 4984 5337 5272 5343
rect 5432 5337 5464 5343
rect 5480 5337 5496 5343
rect 5800 5337 5944 5343
rect 6216 5337 6344 5343
rect 6504 5337 6664 5343
rect 6872 5337 7032 5343
rect 7560 5337 7736 5343
rect 7752 5337 7784 5343
rect 56 5317 88 5323
rect 120 5317 248 5323
rect 264 5317 376 5323
rect 392 5317 504 5323
rect 520 5317 552 5323
rect 696 5317 856 5323
rect 1256 5317 1304 5323
rect 1832 5317 1896 5323
rect 2200 5317 2248 5323
rect 2296 5317 2328 5323
rect 2344 5317 2392 5323
rect 3112 5317 3432 5323
rect 3480 5317 3640 5323
rect 3672 5317 4408 5323
rect 4552 5317 4776 5323
rect 5000 5317 5080 5323
rect 5128 5317 5176 5323
rect 5192 5317 5224 5323
rect 5688 5317 5832 5323
rect 6248 5317 6280 5323
rect 6296 5317 6408 5323
rect 6424 5317 6456 5323
rect 6840 5317 6920 5323
rect 7016 5317 7176 5323
rect 7320 5317 7368 5323
rect 7384 5317 7416 5323
rect 7672 5317 7704 5323
rect 7768 5317 7784 5323
rect 1176 5297 1256 5303
rect 1544 5297 1640 5303
rect 2184 5297 2232 5303
rect 2248 5297 2280 5303
rect 2424 5297 2776 5303
rect 3448 5297 3624 5303
rect 4056 5297 4184 5303
rect 4280 5297 4408 5303
rect 4424 5297 4744 5303
rect 5000 5297 5032 5303
rect 5272 5297 5304 5303
rect 5320 5297 5496 5303
rect 5512 5297 5544 5303
rect 5560 5297 5816 5303
rect 5848 5297 6024 5303
rect 6040 5297 6392 5303
rect 6440 5297 6568 5303
rect 6632 5297 6952 5303
rect 6968 5297 7000 5303
rect 7016 5297 7304 5303
rect 7352 5297 7384 5303
rect 7640 5297 7768 5303
rect 1320 5277 1496 5283
rect 1512 5277 1992 5283
rect 2824 5277 3112 5283
rect 3128 5277 3272 5283
rect 3288 5277 3352 5283
rect 3368 5277 3768 5283
rect 3784 5277 3896 5283
rect 4104 5277 4344 5283
rect 4360 5277 4392 5283
rect 4728 5277 5192 5283
rect 5208 5277 5432 5283
rect 5448 5277 5480 5283
rect 6040 5277 6328 5283
rect 88 5257 1272 5263
rect 1288 5257 1464 5263
rect 1480 5257 1768 5263
rect 1784 5257 2040 5263
rect 2072 5257 2088 5263
rect 2744 5257 3016 5263
rect 3496 5257 4072 5263
rect 4088 5257 4536 5263
rect 4552 5257 5160 5263
rect 5576 5257 6920 5263
rect 6936 5257 7288 5263
rect 7496 5257 7512 5263
rect 7800 5257 7832 5263
rect 1176 5237 1352 5243
rect 1368 5237 2008 5243
rect 2184 5237 3080 5243
rect 3800 5237 3848 5243
rect 4472 5237 5848 5243
rect 1032 5217 1560 5223
rect 1816 5217 2616 5223
rect 3208 5197 3608 5203
rect 3624 5197 3672 5203
rect 3848 5197 4360 5203
rect 4840 5197 4872 5203
rect 1560 5177 2024 5183
rect 2584 5177 4472 5183
rect 4488 5177 5880 5183
rect 5896 5177 7000 5183
rect 1432 5157 1944 5163
rect 1960 5157 4056 5163
rect 4712 5157 4792 5163
rect 4808 5157 4968 5163
rect 4984 5157 5896 5163
rect 744 5137 984 5143
rect 1000 5137 1096 5143
rect 1880 5137 1928 5143
rect 2248 5137 2632 5143
rect 3160 5137 3208 5143
rect 3405 5137 3496 5143
rect 104 5117 280 5123
rect 1384 5117 1464 5123
rect 1768 5117 1848 5123
rect 1928 5117 2264 5123
rect 2648 5117 2680 5123
rect 2776 5117 2792 5123
rect 3405 5123 3411 5137
rect 3576 5137 3944 5143
rect 4648 5137 4888 5143
rect 5672 5137 5704 5143
rect 5960 5137 6104 5143
rect 7240 5137 7304 5143
rect 7320 5137 7608 5143
rect 7624 5137 7704 5143
rect 3080 5117 3411 5123
rect 3432 5117 3464 5123
rect 4024 5117 4088 5123
rect 4280 5117 4408 5123
rect 4776 5117 4872 5123
rect 4936 5117 5944 5123
rect 5960 5117 5976 5123
rect 7816 5117 7880 5123
rect 3645 5108 3651 5112
rect 152 5097 584 5103
rect 680 5097 1080 5103
rect 1144 5097 1448 5103
rect 1464 5097 1512 5103
rect 1848 5097 1992 5103
rect 2072 5097 2168 5103
rect 2312 5097 2360 5103
rect 2408 5097 2616 5103
rect 2696 5097 2856 5103
rect 3400 5097 3528 5103
rect 3704 5097 4056 5103
rect 4392 5097 4424 5103
rect 4440 5097 4520 5103
rect 4536 5097 4616 5103
rect 4648 5097 4760 5103
rect 4856 5097 4872 5103
rect 4888 5097 4920 5103
rect 4968 5097 5128 5103
rect 5272 5097 5368 5103
rect 5448 5097 5752 5103
rect 5928 5097 6024 5103
rect 6040 5097 6152 5103
rect 6472 5097 6616 5103
rect 6632 5097 6680 5103
rect 6968 5097 7128 5103
rect 7624 5097 7752 5103
rect 104 5077 216 5083
rect 232 5077 312 5083
rect 328 5077 440 5083
rect 824 5077 1016 5083
rect 1032 5077 1048 5083
rect 1080 5077 1096 5083
rect 1112 5077 1128 5083
rect 1192 5077 1432 5083
rect 1576 5077 2264 5083
rect 2360 5077 2488 5083
rect 2632 5077 2792 5083
rect 2856 5077 2904 5083
rect 3304 5077 3432 5083
rect 3496 5077 3656 5083
rect 3672 5077 3752 5083
rect 4120 5077 4440 5083
rect 4456 5077 4504 5083
rect 4616 5077 4664 5083
rect 4728 5077 4760 5083
rect 5848 5077 5960 5083
rect 6664 5077 6840 5083
rect 7256 5077 7288 5083
rect 7512 5077 7576 5083
rect 7592 5077 7672 5083
rect 7848 5077 7976 5083
rect 232 5057 248 5063
rect 840 5057 2136 5063
rect 2152 5057 2280 5063
rect 2488 5057 2840 5063
rect 3352 5057 3640 5063
rect 4136 5057 4344 5063
rect 4856 5057 4888 5063
rect 4904 5057 5656 5063
rect 6472 5057 6488 5063
rect 6504 5057 6808 5063
rect 6984 5057 7608 5063
rect 56 5037 376 5043
rect 968 5037 984 5043
rect 2040 5037 2184 5043
rect 2280 5037 2712 5043
rect 2760 5037 4115 5043
rect 40 5017 328 5023
rect 344 5017 760 5023
rect 776 5017 824 5023
rect 1720 5017 1816 5023
rect 4109 5023 4115 5037
rect 4568 5037 4920 5043
rect 4936 5037 5139 5043
rect 808 4997 1400 5003
rect 3528 4997 3544 5003
rect 4109 5017 4632 5023
rect 4728 5017 4936 5023
rect 5133 5023 5139 5037
rect 5160 5037 5208 5043
rect 5224 5037 5336 5043
rect 5576 5037 6344 5043
rect 6824 5037 7016 5043
rect 7032 5037 7256 5043
rect 7272 5037 7320 5043
rect 7336 5037 7544 5043
rect 7560 5037 7640 5043
rect 7784 5037 7928 5043
rect 5133 5017 5288 5023
rect 5304 5017 5576 5023
rect 5592 5017 5768 5023
rect 6904 5017 7352 5023
rect 7368 5017 7656 5023
rect 7672 5017 7848 5023
rect 7832 4997 7864 5003
rect 488 4977 1016 4983
rect 1245 4977 1256 4983
rect 1528 4977 2408 4983
rect 3464 4977 4168 4983
rect 4744 4977 4776 4983
rect 4792 4977 5000 4983
rect 5656 4977 5720 4983
rect 7672 4977 7944 4983
rect 168 4957 328 4963
rect 760 4957 824 4963
rect 1288 4957 1480 4963
rect 2088 4957 2440 4963
rect 2552 4957 2712 4963
rect 3368 4957 3480 4963
rect 3544 4957 4104 4963
rect 4872 4957 4984 4963
rect 5000 4957 5944 4963
rect 7640 4957 7992 4963
rect 264 4937 392 4943
rect 440 4937 472 4943
rect 648 4937 792 4943
rect 1080 4937 1107 4943
rect 136 4917 168 4923
rect 232 4917 248 4923
rect 264 4917 312 4923
rect 456 4917 472 4923
rect 744 4917 776 4923
rect 792 4917 856 4923
rect 872 4917 904 4923
rect 920 4917 1000 4923
rect 1101 4923 1107 4937
rect 1128 4937 1224 4943
rect 1528 4937 1560 4943
rect 1576 4937 1704 4943
rect 1992 4937 2168 4943
rect 2408 4937 2568 4943
rect 2584 4937 2979 4943
rect 1101 4917 1432 4923
rect 1448 4917 1640 4923
rect 1800 4917 1992 4923
rect 2328 4917 2472 4923
rect 2648 4917 2744 4923
rect 2973 4923 2979 4937
rect 3000 4937 3080 4943
rect 3096 4937 3208 4943
rect 3224 4937 3560 4943
rect 3656 4937 3688 4943
rect 3864 4937 3880 4943
rect 3992 4937 4296 4943
rect 4664 4937 4856 4943
rect 4920 4937 5096 4943
rect 5240 4937 5496 4943
rect 5528 4937 5672 4943
rect 5784 4937 6248 4943
rect 6456 4937 6600 4943
rect 6696 4937 6776 4943
rect 6792 4937 6920 4943
rect 6984 4937 7112 4943
rect 7384 4937 7496 4943
rect 7848 4937 7864 4943
rect 7885 4937 7896 4943
rect 6445 4928 6451 4932
rect 2973 4917 3064 4923
rect 3288 4917 3432 4923
rect 3480 4917 3512 4923
rect 3672 4917 3864 4923
rect 3912 4917 3944 4923
rect 3960 4917 4072 4923
rect 4264 4917 4408 4923
rect 4840 4917 4952 4923
rect 5400 4917 5624 4923
rect 5720 4917 5752 4923
rect 5768 4917 5944 4923
rect 6008 4917 6136 4923
rect 6568 4917 6680 4923
rect 7352 4917 7688 4923
rect 7736 4917 7848 4923
rect 7880 4917 7928 4923
rect 7944 4917 8024 4923
rect 1085 4908 1091 4912
rect 4573 4908 4579 4912
rect 152 4897 264 4903
rect 1096 4897 1288 4903
rect 1320 4897 1352 4903
rect 1368 4897 1384 4903
rect 1400 4897 1576 4903
rect 1608 4897 1656 4903
rect 2040 4897 2152 4903
rect 2632 4897 2648 4903
rect 2680 4897 2888 4903
rect 3112 4897 3160 4903
rect 3752 4897 3848 4903
rect 4360 4897 4392 4903
rect 4408 4897 4440 4903
rect 4872 4897 4920 4903
rect 6280 4897 6312 4903
rect 6408 4897 6584 4903
rect 6696 4897 6936 4903
rect 7016 4897 7528 4903
rect 7912 4897 7976 4903
rect 248 4877 296 4883
rect 328 4877 360 4883
rect 1064 4877 1528 4883
rect 1544 4877 1624 4883
rect 1816 4877 2120 4883
rect 3176 4877 3448 4883
rect 3704 4877 3816 4883
rect 4504 4877 4568 4883
rect 4648 4877 5880 4883
rect 5896 4877 6024 4883
rect 6104 4877 6664 4883
rect 6680 4877 6824 4883
rect 6840 4877 7112 4883
rect 7128 4877 7192 4883
rect 7208 4877 7512 4883
rect 7912 4877 7944 4883
rect 904 4857 1000 4863
rect 1336 4857 1560 4863
rect 1592 4857 1736 4863
rect 3640 4857 3896 4863
rect 5864 4857 6392 4863
rect 6424 4857 7656 4863
rect 392 4837 1224 4843
rect 1384 4837 1752 4843
rect 3720 4837 3800 4843
rect 3848 4837 3896 4843
rect 3960 4837 4040 4843
rect 5080 4837 5544 4843
rect 6200 4837 7464 4843
rect 7608 4837 7912 4843
rect 200 4817 632 4823
rect 216 4797 488 4803
rect 1400 4817 1656 4823
rect 2232 4817 2936 4823
rect 984 4797 1464 4803
rect 1560 4797 2888 4803
rect 3512 4817 3832 4823
rect 3848 4817 3976 4823
rect 4088 4817 4760 4823
rect 4776 4817 4968 4823
rect 3736 4797 4072 4803
rect 5880 4817 6456 4823
rect 6472 4817 6520 4823
rect 6536 4817 6632 4823
rect 6024 4797 6088 4803
rect 6440 4797 6856 4803
rect 264 4777 280 4783
rect 552 4777 664 4783
rect 888 4777 1720 4783
rect 1832 4777 2392 4783
rect 3208 4777 4152 4783
rect 4168 4777 4280 4783
rect 4824 4777 5112 4783
rect 5128 4777 5224 4783
rect 6168 4777 6376 4783
rect -51 4757 136 4763
rect 184 4757 552 4763
rect 808 4757 968 4763
rect 1000 4757 1144 4763
rect 1624 4757 1912 4763
rect 2376 4757 3368 4763
rect 3400 4757 3704 4763
rect 3768 4757 3864 4763
rect 3912 4757 4184 4763
rect 4520 4757 4920 4763
rect 6216 4757 6280 4763
rect 6680 4757 6696 4763
rect 7544 4757 7608 4763
rect 152 4737 200 4743
rect 248 4737 344 4743
rect 488 4737 536 4743
rect 568 4737 808 4743
rect 1016 4737 1304 4743
rect 1352 4737 1400 4743
rect 1448 4737 2760 4743
rect 3192 4737 3240 4743
rect 3416 4737 3512 4743
rect 3544 4737 3880 4743
rect 3928 4737 4504 4743
rect 5096 4737 5256 4743
rect 5400 4737 5432 4743
rect 6184 4737 6200 4743
rect 6232 4737 6243 4743
rect 6280 4737 6344 4743
rect 6648 4737 6728 4743
rect 6744 4737 7448 4743
rect 973 4728 979 4732
rect 5453 4728 5459 4732
rect -51 4717 376 4723
rect 392 4717 520 4723
rect 1032 4717 1096 4723
rect 1336 4717 1347 4723
rect 1341 4708 1347 4717
rect 1400 4717 1528 4723
rect 1592 4717 1848 4723
rect 1896 4717 1944 4723
rect 2264 4717 2344 4723
rect 2376 4717 2632 4723
rect 2728 4717 2856 4723
rect 2872 4717 2968 4723
rect 3048 4717 3240 4723
rect 3448 4717 3544 4723
rect 3656 4717 3928 4723
rect 3960 4717 4088 4723
rect 4120 4717 4232 4723
rect 4253 4717 4280 4723
rect 136 4697 232 4703
rect 264 4697 280 4703
rect 328 4697 376 4703
rect 712 4697 856 4703
rect 888 4697 904 4703
rect 920 4697 984 4703
rect 1048 4697 1059 4703
rect 1149 4697 1272 4703
rect 56 4677 88 4683
rect 232 4677 360 4683
rect 376 4677 408 4683
rect 1149 4683 1155 4697
rect 1384 4697 1496 4703
rect 1528 4697 1608 4703
rect 1848 4697 1928 4703
rect 2056 4697 2136 4703
rect 2296 4697 2376 4703
rect 2872 4697 2936 4703
rect 2968 4697 3096 4703
rect 3288 4697 3448 4703
rect 3768 4697 4184 4703
rect 4253 4703 4259 4717
rect 4344 4717 4392 4723
rect 4424 4717 4440 4723
rect 5208 4717 5416 4723
rect 5480 4717 5560 4723
rect 5624 4717 5640 4723
rect 5656 4717 5816 4723
rect 6056 4717 6072 4723
rect 6184 4717 6696 4723
rect 6712 4717 6904 4723
rect 7096 4717 7160 4723
rect 7624 4717 7816 4723
rect 7832 4717 7992 4723
rect 4216 4697 4259 4703
rect 4280 4697 4440 4703
rect 4472 4697 4504 4703
rect 4568 4697 5112 4703
rect 5144 4697 5304 4703
rect 5320 4697 6024 4703
rect 6040 4697 6424 4703
rect 6440 4697 6632 4703
rect 6728 4697 6760 4703
rect 6808 4697 7016 4703
rect 7112 4697 7288 4703
rect 7720 4697 7736 4703
rect 7752 4697 7784 4703
rect 7816 4697 7912 4703
rect 7976 4697 7992 4703
rect 493 4677 1155 4683
rect 493 4663 499 4677
rect 1176 4677 1240 4683
rect 1272 4677 1432 4683
rect 1528 4677 1704 4683
rect 1720 4677 1832 4683
rect 2024 4677 2152 4683
rect 2408 4677 2488 4683
rect 2936 4677 3448 4683
rect 3496 4677 3704 4683
rect 3736 4677 3768 4683
rect 3800 4677 3976 4683
rect 3992 4677 4264 4683
rect 4296 4677 4312 4683
rect 4360 4677 4392 4683
rect 5016 4677 5128 4683
rect 5256 4677 5352 4683
rect 5368 4677 6136 4683
rect 6152 4677 6216 4683
rect 6232 4677 6536 4683
rect 6568 4677 6584 4683
rect 6680 4677 6808 4683
rect 6856 4677 6872 4683
rect 6904 4677 6936 4683
rect 7048 4677 7112 4683
rect 7144 4677 7576 4683
rect 7720 4677 7864 4683
rect 296 4657 499 4663
rect 520 4657 1592 4663
rect 1720 4657 1848 4663
rect 2456 4657 2616 4663
rect 2632 4657 2776 4663
rect 2856 4657 3096 4663
rect 3384 4657 3576 4663
rect 3864 4657 4136 4663
rect 4168 4657 4216 4663
rect 4280 4657 4360 4663
rect 4440 4657 5208 4663
rect 5240 4657 5256 4663
rect 5352 4657 5416 4663
rect 5432 4657 5528 4663
rect 5672 4657 6248 4663
rect 6264 4657 6616 4663
rect 6632 4657 6648 4663
rect 6760 4657 6856 4663
rect 7432 4657 7480 4663
rect 7496 4657 7560 4663
rect 904 4637 1192 4643
rect 1416 4637 1512 4643
rect 1613 4637 1624 4643
rect 1768 4637 1784 4643
rect 2280 4637 2472 4643
rect 3144 4637 3400 4643
rect 3416 4637 3608 4643
rect 3688 4637 4024 4643
rect 4216 4637 4472 4643
rect 5352 4637 5656 4643
rect 5688 4637 5736 4643
rect 5752 4637 6088 4643
rect 6216 4637 6232 4643
rect 6312 4637 6440 4643
rect 6552 4637 6648 4643
rect 6744 4637 6824 4643
rect 6904 4637 7000 4643
rect 168 4617 424 4623
rect 440 4617 536 4623
rect 552 4617 680 4623
rect 808 4617 904 4623
rect 920 4617 1016 4623
rect 1448 4617 1896 4623
rect 1912 4617 1928 4623
rect 312 4597 488 4603
rect 1080 4597 1384 4603
rect 1432 4597 1592 4603
rect 1640 4597 1720 4603
rect 2696 4617 3080 4623
rect 3096 4617 3144 4623
rect 3160 4617 3208 4623
rect 3224 4617 3384 4623
rect 3624 4617 3752 4623
rect 4072 4617 4136 4623
rect 4152 4617 4568 4623
rect 5240 4617 5368 4623
rect 5528 4617 5608 4623
rect 5976 4617 6008 4623
rect 4136 4597 5272 4603
rect 5416 4597 5992 4603
rect 6136 4617 7672 4623
rect 6104 4597 6168 4603
rect 6488 4597 6568 4603
rect 6685 4597 7128 4603
rect 968 4577 1016 4583
rect 1064 4577 1192 4583
rect 1400 4577 1448 4583
rect 1784 4577 1832 4583
rect 2248 4577 2312 4583
rect 3080 4577 3768 4583
rect 3784 4577 3832 4583
rect 3944 4577 4616 4583
rect 4648 4577 4680 4583
rect 5501 4577 5560 4583
rect 5501 4568 5507 4577
rect 6685 4583 6691 4597
rect 7144 4597 7320 4603
rect 7672 4597 7976 4603
rect 5928 4577 6691 4583
rect 6952 4577 6968 4583
rect 7512 4577 7720 4583
rect 7837 4568 7843 4572
rect 936 4557 1112 4563
rect 1192 4557 1416 4563
rect 1432 4557 2008 4563
rect 3032 4557 3208 4563
rect 3336 4557 3368 4563
rect 3448 4557 3496 4563
rect 3512 4557 4728 4563
rect 4776 4557 4808 4563
rect 4888 4557 5224 4563
rect 5304 4557 5416 4563
rect 5560 4557 5720 4563
rect 5736 4557 6408 4563
rect 6840 4557 6968 4563
rect 6984 4557 7144 4563
rect 7224 4557 7544 4563
rect 45 4548 51 4552
rect 328 4537 424 4543
rect 584 4537 872 4543
rect 936 4537 968 4543
rect 1112 4537 1288 4543
rect 1320 4537 1512 4543
rect 1544 4537 1816 4543
rect 1848 4537 1896 4543
rect 2312 4537 2408 4543
rect 2552 4537 2632 4543
rect 2760 4537 2968 4543
rect 3176 4537 3752 4543
rect 3768 4537 3784 4543
rect 3816 4537 3880 4543
rect 3992 4537 4184 4543
rect 4312 4537 4488 4543
rect 4712 4537 4792 4543
rect 4808 4537 4824 4543
rect 4840 4537 5112 4543
rect 5288 4537 5320 4543
rect 5400 4537 5528 4543
rect 5800 4537 5816 4543
rect 6008 4537 6072 4543
rect 6104 4537 6232 4543
rect 6664 4537 6808 4543
rect 6824 4537 6872 4543
rect 7128 4537 7144 4543
rect 7325 4537 7432 4543
rect 1821 4528 1827 4532
rect 200 4517 248 4523
rect 488 4517 504 4523
rect 520 4517 616 4523
rect 1016 4517 1400 4523
rect 1416 4517 1432 4523
rect 1496 4517 1507 4523
rect 2168 4517 2264 4523
rect 2680 4517 2712 4523
rect 3160 4517 3224 4523
rect 3256 4517 3816 4523
rect 3832 4517 3848 4523
rect 3880 4517 3912 4523
rect 3960 4517 4040 4523
rect 4088 4517 4120 4523
rect 4424 4517 4536 4523
rect 4680 4517 4808 4523
rect 4840 4517 4936 4523
rect 4952 4517 5176 4523
rect 5208 4517 6152 4523
rect 6168 4517 6312 4523
rect 6328 4517 6536 4523
rect 6552 4517 6664 4523
rect 6744 4517 6840 4523
rect 7325 4523 7331 4537
rect 7640 4537 7784 4543
rect 7320 4517 7331 4523
rect 7352 4517 7464 4523
rect 7480 4517 7528 4523
rect 2061 4508 2067 4512
rect 5197 4508 5203 4512
rect 136 4497 200 4503
rect 216 4497 280 4503
rect 296 4497 344 4503
rect 616 4497 664 4503
rect 1224 4497 1256 4503
rect 1368 4497 1464 4503
rect 2088 4497 2232 4503
rect 2248 4497 2536 4503
rect 2712 4497 2808 4503
rect 3064 4497 3160 4503
rect 3208 4497 3256 4503
rect 3368 4497 3448 4503
rect 3576 4497 3992 4503
rect 4024 4497 4088 4503
rect 4536 4497 4568 4503
rect 4856 4497 4888 4503
rect 5096 4497 5192 4503
rect 5496 4497 5608 4503
rect 6008 4497 6024 4503
rect 6136 4497 6184 4503
rect 6872 4497 6888 4503
rect 6936 4497 7016 4503
rect 7448 4497 7480 4503
rect 7608 4497 7640 4503
rect 7656 4497 7736 4503
rect 3325 4488 3331 4492
rect 328 4477 440 4483
rect 456 4477 680 4483
rect 1624 4477 1640 4483
rect 1656 4477 1672 4483
rect 2040 4477 2200 4483
rect 2552 4477 2584 4483
rect 3016 4477 3304 4483
rect 3336 4477 3496 4483
rect 3512 4477 3768 4483
rect 3784 4477 3816 4483
rect 4216 4477 5448 4483
rect 5464 4477 5720 4483
rect 5736 4477 6440 4483
rect 6872 4477 7160 4483
rect 264 4457 328 4463
rect 360 4457 424 4463
rect 440 4457 632 4463
rect 648 4457 872 4463
rect 1624 4457 1768 4463
rect 3224 4457 3400 4463
rect 3464 4457 3896 4463
rect 3912 4457 3960 4463
rect 4744 4457 4856 4463
rect 6536 4457 6904 4463
rect 7464 4457 7480 4463
rect 408 4437 488 4443
rect 520 4437 552 4443
rect 872 4437 1704 4443
rect 2840 4437 4648 4443
rect 4664 4437 5640 4443
rect 5656 4437 6424 4443
rect 6472 4437 6483 4443
rect 6680 4437 7512 4443
rect 520 4417 568 4423
rect -51 4397 520 4403
rect 552 4397 664 4403
rect 1320 4397 1928 4403
rect 2120 4397 2152 4403
rect 3192 4417 3992 4423
rect 4024 4417 4184 4423
rect 3240 4397 3304 4403
rect 3400 4397 3432 4403
rect 3944 4397 4248 4403
rect 5592 4417 5784 4423
rect 5800 4417 6344 4423
rect 5624 4397 6904 4403
rect 2861 4388 2867 4392
rect 2925 4388 2931 4392
rect 3165 4388 3171 4392
rect 40 4377 168 4383
rect 184 4377 232 4383
rect 456 4377 488 4383
rect 600 4377 1192 4383
rect 1368 4377 1448 4383
rect 1944 4377 2104 4383
rect 3496 4377 3608 4383
rect 3640 4377 3736 4383
rect 3752 4377 5128 4383
rect 5832 4377 7416 4383
rect 7928 4377 7944 4383
rect 7960 4377 8024 4383
rect -51 4357 248 4363
rect 504 4357 968 4363
rect 1128 4357 1592 4363
rect 1944 4357 2120 4363
rect 2920 4357 3288 4363
rect 3320 4357 3512 4363
rect 3688 4357 4568 4363
rect 4584 4357 4680 4363
rect 6152 4357 6168 4363
rect 6424 4357 7400 4363
rect 7976 4357 8024 4363
rect 392 4337 424 4343
rect 584 4337 616 4343
rect 664 4337 696 4343
rect 776 4337 808 4343
rect 1064 4337 1352 4343
rect 1544 4337 1912 4343
rect 2056 4337 3144 4343
rect 3432 4337 3496 4343
rect 3688 4337 3784 4343
rect 3800 4337 3912 4343
rect 5656 4337 5768 4343
rect 5848 4337 6536 4343
rect 6552 4337 6616 4343
rect 6792 4337 6824 4343
rect 6840 4337 7336 4343
rect 2029 4328 2035 4332
rect -51 4303 -45 4323
rect 328 4317 344 4323
rect 360 4317 488 4323
rect 536 4317 728 4323
rect 792 4317 808 4323
rect 1096 4317 1144 4323
rect 3128 4317 3192 4323
rect 3240 4317 3720 4323
rect 3736 4317 3832 4323
rect 3928 4317 3944 4323
rect 4328 4317 4776 4323
rect 4952 4317 4984 4323
rect 5480 4317 5496 4323
rect 5736 4317 5800 4323
rect 5816 4317 5880 4323
rect 6136 4317 6147 4323
rect 6456 4317 6872 4323
rect 6888 4317 7000 4323
rect 7032 4317 7176 4323
rect 7496 4317 7560 4323
rect 7576 4317 7624 4323
rect 5661 4308 5667 4312
rect -51 4297 8 4303
rect 248 4297 552 4303
rect 728 4297 792 4303
rect 936 4297 984 4303
rect 1000 4297 1096 4303
rect 1224 4297 1432 4303
rect 1816 4297 1848 4303
rect 2216 4297 2264 4303
rect 2296 4297 2456 4303
rect 2968 4297 3032 4303
rect 3112 4297 3128 4303
rect 3176 4297 3368 4303
rect 3384 4297 3656 4303
rect 3672 4297 3816 4303
rect 3832 4297 3848 4303
rect 3944 4297 3976 4303
rect 4984 4297 5144 4303
rect 5384 4297 5464 4303
rect 5672 4297 5720 4303
rect 5768 4297 5976 4303
rect 5992 4297 6024 4303
rect 6056 4297 6232 4303
rect 6328 4297 6408 4303
rect 6424 4297 6456 4303
rect 6472 4297 6552 4303
rect 6568 4297 7032 4303
rect 7208 4297 7368 4303
rect 7384 4297 7448 4303
rect 7976 4297 8008 4303
rect 2013 4288 2019 4292
rect 56 4277 248 4283
rect 392 4277 504 4283
rect 1400 4277 1480 4283
rect 1656 4277 1816 4283
rect 2104 4277 2184 4283
rect 2200 4277 2248 4283
rect 2264 4277 2312 4283
rect 3496 4277 3528 4283
rect 3624 4277 3656 4283
rect 3720 4277 3736 4283
rect 3848 4277 3896 4283
rect 3960 4277 4152 4283
rect 4248 4277 4504 4283
rect 4920 4277 5016 4283
rect 5528 4277 5736 4283
rect 5768 4277 5896 4283
rect 5960 4277 5976 4283
rect 5992 4277 6072 4283
rect 6088 4277 6664 4283
rect 7032 4277 7512 4283
rect 7560 4277 7720 4283
rect 3757 4268 3763 4272
rect 72 4257 408 4263
rect 424 4257 600 4263
rect 744 4257 1000 4263
rect 1784 4257 1880 4263
rect 1896 4257 1944 4263
rect 3064 4257 3304 4263
rect 3816 4257 3848 4263
rect 3864 4257 3896 4263
rect 3992 4257 4312 4263
rect 5976 4257 6472 4263
rect 6856 4257 7032 4263
rect 7048 4257 7192 4263
rect 7384 4257 7400 4263
rect 7512 4257 7704 4263
rect 232 4237 296 4243
rect 312 4237 424 4243
rect 440 4237 472 4243
rect 824 4237 1176 4243
rect 1192 4237 1368 4243
rect 1384 4237 1624 4243
rect 1912 4237 2056 4243
rect 3880 4237 4104 4243
rect 4184 4237 4472 4243
rect 6488 4237 7800 4243
rect 264 4217 616 4223
rect 632 4217 680 4223
rect 696 4217 744 4223
rect 808 4217 824 4223
rect 840 4217 1032 4223
rect 1048 4217 1160 4223
rect 1352 4197 1576 4203
rect 1592 4197 1608 4203
rect 3544 4217 3784 4223
rect 2152 4197 2872 4203
rect 3128 4197 3400 4203
rect 4248 4217 4344 4223
rect 4360 4217 4760 4223
rect 4776 4217 4824 4223
rect 5592 4217 5864 4223
rect 4120 4197 4376 4203
rect 6744 4217 7288 4223
rect 7592 4217 7688 4223
rect 6984 4197 7032 4203
rect 7048 4197 7112 4203
rect 24 4177 1352 4183
rect 1880 4177 2040 4183
rect 2344 4177 2360 4183
rect 2376 4177 2760 4183
rect 3160 4177 3320 4183
rect 3448 4177 3544 4183
rect 3560 4177 3880 4183
rect 3992 4177 4264 4183
rect 4392 4177 4792 4183
rect 4808 4177 4904 4183
rect 5784 4177 5912 4183
rect 6360 4177 6392 4183
rect 6952 4177 7160 4183
rect 7528 4177 8040 4183
rect 1032 4157 1304 4163
rect 1320 4157 1368 4163
rect 1608 4157 1656 4163
rect 2024 4157 2072 4163
rect 2925 4157 2931 4172
rect 2952 4157 3544 4163
rect 3560 4157 3672 4163
rect 3704 4157 4040 4163
rect 4216 4157 4392 4163
rect 4408 4157 4584 4163
rect 4696 4157 4856 4163
rect 4872 4157 5176 4163
rect 5864 4157 5928 4163
rect 6088 4157 6456 4163
rect 6472 4157 6504 4163
rect 6600 4157 6952 4163
rect 6968 4157 7048 4163
rect 7944 4157 7976 4163
rect 1176 4137 1272 4143
rect 1528 4137 1672 4143
rect 1688 4137 1752 4143
rect 1768 4137 1928 4143
rect 1960 4137 2040 4143
rect 2056 4137 2216 4143
rect 2472 4137 2584 4143
rect 2616 4137 2680 4143
rect 2696 4137 2728 4143
rect 2840 4137 3240 4143
rect 3416 4137 3480 4143
rect 3512 4137 3928 4143
rect 3960 4137 4248 4143
rect 4456 4137 4600 4143
rect 5368 4137 5384 4143
rect 5400 4137 5544 4143
rect 5656 4137 5832 4143
rect 5848 4137 5960 4143
rect 6504 4137 6744 4143
rect 7064 4137 7139 4143
rect 2829 4128 2835 4132
rect -51 4117 56 4123
rect 72 4117 200 4123
rect 264 4117 296 4123
rect 744 4117 776 4123
rect 840 4117 872 4123
rect 888 4117 920 4123
rect 1112 4117 1256 4123
rect 1277 4117 1672 4123
rect 248 4097 488 4103
rect 504 4097 632 4103
rect 648 4097 840 4103
rect 856 4097 888 4103
rect 1277 4103 1283 4117
rect 1688 4117 1704 4123
rect 1752 4117 1816 4123
rect 1832 4117 2056 4123
rect 2440 4117 2536 4123
rect 2728 4117 2792 4123
rect 2845 4117 2856 4123
rect 2872 4117 3064 4123
rect 3192 4117 3240 4123
rect 3256 4117 3400 4123
rect 3448 4117 3496 4123
rect 3704 4117 3736 4123
rect 3768 4117 4040 4123
rect 4248 4117 4344 4123
rect 4424 4117 4456 4123
rect 4472 4117 4840 4123
rect 4872 4117 5000 4123
rect 5272 4117 5592 4123
rect 5752 4117 5864 4123
rect 5944 4117 6008 4123
rect 6024 4117 6088 4123
rect 6120 4117 6216 4123
rect 6232 4117 6296 4123
rect 6552 4117 6600 4123
rect 6616 4117 6728 4123
rect 6776 4117 6792 4123
rect 7032 4117 7112 4123
rect 7133 4123 7139 4137
rect 7160 4137 7288 4143
rect 7688 4137 7816 4143
rect 7133 4117 7224 4123
rect 7480 4117 7544 4123
rect 7592 4117 7640 4123
rect 7656 4117 7720 4123
rect 7816 4117 7928 4123
rect 7960 4117 8008 4123
rect 952 4097 1283 4103
rect 1480 4097 1672 4103
rect 1864 4097 1912 4103
rect 2216 4097 2296 4103
rect 2408 4097 2472 4103
rect 2664 4097 2680 4103
rect 2824 4097 2984 4103
rect 3144 4097 3160 4103
rect 3576 4097 3720 4103
rect 3789 4097 3800 4103
rect 3944 4097 3992 4103
rect 4232 4097 4248 4103
rect 4568 4097 4728 4103
rect 4840 4097 4872 4103
rect 5288 4097 5640 4103
rect 5656 4097 6232 4103
rect 6920 4097 7016 4103
rect 7432 4097 7512 4103
rect 7608 4097 7624 4103
rect 7640 4097 7720 4103
rect 264 4077 280 4083
rect 312 4077 328 4083
rect 376 4077 536 4083
rect 680 4077 1208 4083
rect 1672 4077 1688 4083
rect 1720 4077 2008 4083
rect 2888 4077 3240 4083
rect 3272 4077 3320 4083
rect 3336 4077 3416 4083
rect 3480 4077 3496 4083
rect 3736 4077 3832 4083
rect 3848 4077 4600 4083
rect 4616 4077 4776 4083
rect 6904 4077 6920 4083
rect 1533 4068 1539 4072
rect 1656 4057 1848 4063
rect 1880 4057 1992 4063
rect 2008 4057 2168 4063
rect 3112 4057 3176 4063
rect 3320 4057 3432 4063
rect 3480 4057 3640 4063
rect 4312 4057 4776 4063
rect 6264 4057 6840 4063
rect 6920 4057 6936 4063
rect 6952 4057 6984 4063
rect 280 4037 1256 4043
rect 1608 4037 1704 4043
rect 2024 4037 2184 4043
rect 3208 4037 3336 4043
rect 3736 4037 3928 4043
rect 3944 4037 3976 4043
rect 4152 4037 4328 4043
rect 4344 4037 4664 4043
rect 6216 4037 6520 4043
rect 6536 4037 6840 4043
rect 6856 4037 6936 4043
rect 200 3997 552 4003
rect 600 3997 760 4003
rect 1416 4017 1560 4023
rect 1576 4017 1800 4023
rect 1816 4017 2248 4023
rect 1464 3997 2024 4003
rect 2104 3997 2120 4003
rect 3448 4017 3752 4023
rect 3384 3997 3544 4003
rect 3672 3997 4072 4003
rect 5704 4017 6440 4023
rect 6456 4017 6792 4023
rect 5112 3997 5736 4003
rect 5896 3997 5976 4003
rect 5992 3997 6024 4003
rect 6184 3997 6824 4003
rect 1112 3977 1144 3983
rect 1368 3977 2088 3983
rect 3368 3977 3480 3983
rect 3512 3977 3640 3983
rect 3656 3977 3672 3983
rect 3896 3977 3960 3983
rect 4712 3977 4744 3983
rect 5400 3977 5896 3983
rect 6024 3977 6136 3983
rect 6152 3977 6408 3983
rect 184 3957 248 3963
rect 328 3957 360 3963
rect 568 3957 1176 3963
rect 1192 3957 1352 3963
rect 1368 3957 1416 3963
rect 2248 3957 2936 3963
rect 3432 3957 3864 3963
rect 3880 3957 3928 3963
rect 4728 3957 7688 3963
rect 24 3937 104 3943
rect 248 3937 440 3943
rect 456 3937 600 3943
rect 792 3937 936 3943
rect 984 3937 1032 3943
rect 1048 3937 1240 3943
rect 1416 3937 1448 3943
rect 1800 3937 1992 3943
rect 2376 3937 2552 3943
rect 2568 3937 2776 3943
rect 3032 3937 3224 3943
rect 3240 3937 3272 3943
rect 3496 3937 3528 3943
rect 3576 3937 3720 3943
rect 3800 3937 4200 3943
rect 4328 3937 4632 3943
rect 4760 3937 5320 3943
rect 5432 3937 5864 3943
rect 5880 3937 5992 3943
rect 6536 3937 6552 3943
rect 6568 3937 6600 3943
rect 7304 3937 7448 3943
rect 7464 3937 7896 3943
rect 24 3917 88 3923
rect 168 3917 344 3923
rect 376 3917 696 3923
rect 888 3917 1000 3923
rect 1400 3917 1416 3923
rect 1496 3917 2024 3923
rect 2040 3917 2104 3923
rect 2152 3917 2296 3923
rect 2600 3917 2680 3923
rect 3176 3917 3288 3923
rect 3544 3917 3576 3923
rect 3688 3917 3896 3923
rect 4568 3917 4600 3923
rect 4664 3917 4856 3923
rect 5080 3917 5208 3923
rect 5672 3917 5720 3923
rect 5912 3917 5944 3923
rect 6184 3917 6280 3923
rect 6312 3917 6472 3923
rect 6568 3917 6664 3923
rect 6776 3917 6840 3923
rect 6856 3917 6872 3923
rect 7240 3917 7400 3923
rect 7544 3917 7592 3923
rect 7656 3917 7752 3923
rect 104 3897 200 3903
rect 232 3897 280 3903
rect 360 3897 424 3903
rect 440 3897 488 3903
rect 504 3897 536 3903
rect 552 3897 600 3903
rect 632 3897 664 3903
rect 840 3897 851 3903
rect 1080 3897 1160 3903
rect 1352 3897 1400 3903
rect 1432 3897 1480 3903
rect 1816 3897 2168 3903
rect 2189 3897 2200 3903
rect 56 3877 168 3883
rect 392 3877 424 3883
rect 696 3877 728 3883
rect 744 3877 1064 3883
rect 1160 3877 1192 3883
rect 1256 3877 1464 3883
rect 1517 3883 1523 3892
rect 1512 3877 1523 3883
rect 1816 3877 1832 3883
rect 1848 3877 1960 3883
rect 1992 3877 2040 3883
rect 2189 3883 2195 3897
rect 2456 3897 2648 3903
rect 3032 3897 3256 3903
rect 3384 3897 3608 3903
rect 3624 3897 3688 3903
rect 3736 3897 3752 3903
rect 3784 3897 3832 3903
rect 3928 3897 3960 3903
rect 4056 3897 4216 3903
rect 4456 3897 4552 3903
rect 4696 3897 4707 3903
rect 4728 3897 4968 3903
rect 4984 3897 5112 3903
rect 5528 3897 5619 3903
rect 2088 3877 2195 3883
rect 2552 3877 2696 3883
rect 3144 3877 3192 3883
rect 3464 3877 3688 3883
rect 3848 3877 4184 3883
rect 4360 3877 4520 3883
rect 4856 3877 5000 3883
rect 5016 3877 5080 3883
rect 5432 3877 5592 3883
rect 5613 3883 5619 3897
rect 5640 3897 5672 3903
rect 5944 3897 5987 3903
rect 5613 3877 5640 3883
rect 5981 3883 5987 3897
rect 6008 3897 6024 3903
rect 6264 3897 6328 3903
rect 6696 3897 6808 3903
rect 7128 3897 7208 3903
rect 7224 3897 7272 3903
rect 7592 3897 7640 3903
rect 5981 3877 6040 3883
rect 6088 3877 6104 3883
rect 6440 3877 6488 3883
rect 6504 3877 6760 3883
rect 6792 3877 6952 3883
rect 7320 3877 7480 3883
rect 7528 3877 7539 3883
rect 7560 3877 7592 3883
rect 7709 3883 7715 3892
rect 7656 3877 7816 3883
rect 200 3857 264 3863
rect 280 3857 392 3863
rect 936 3857 1000 3863
rect 1032 3857 1256 3863
rect 2008 3857 3080 3863
rect 3544 3857 3944 3863
rect 4040 3857 4056 3863
rect 4184 3857 4680 3863
rect 4696 3857 4856 3863
rect 4952 3857 5192 3863
rect 5992 3857 6344 3863
rect 6904 3857 6968 3863
rect 7624 3857 7704 3863
rect 7720 3857 7752 3863
rect 312 3837 392 3843
rect 920 3837 1240 3843
rect 1432 3837 3944 3843
rect 3976 3837 4728 3843
rect 4776 3837 5000 3843
rect 5016 3837 5368 3843
rect 5384 3837 5416 3843
rect 6152 3837 6163 3843
rect 6248 3837 6312 3843
rect 6472 3837 6728 3843
rect 6968 3837 7144 3843
rect 7704 3837 7960 3843
rect 424 3817 552 3823
rect 760 3817 968 3823
rect 1000 3817 1800 3823
rect 24 3797 840 3803
rect 888 3797 1288 3803
rect 1416 3797 1848 3803
rect 2568 3817 2936 3823
rect 2104 3797 2376 3803
rect 2680 3797 2744 3803
rect 2792 3797 2808 3803
rect 4232 3817 4344 3823
rect 4360 3817 4440 3823
rect 4456 3817 4504 3823
rect 4616 3817 4648 3823
rect 4680 3817 4824 3823
rect 4104 3797 4520 3803
rect 4632 3797 4664 3803
rect 4680 3797 4760 3803
rect 4824 3797 5064 3803
rect 6328 3817 6408 3823
rect 6424 3817 6504 3823
rect 6520 3817 6776 3823
rect 6792 3817 6984 3823
rect 6280 3797 6584 3803
rect 6600 3797 6840 3803
rect 6920 3797 6968 3803
rect 2765 3788 2771 3792
rect 72 3777 200 3783
rect 632 3777 1432 3783
rect 1704 3777 1880 3783
rect 1912 3777 2120 3783
rect 3208 3777 3544 3783
rect 3640 3777 3795 3783
rect 56 3757 88 3763
rect 168 3757 296 3763
rect 648 3757 1016 3763
rect 1480 3757 1848 3763
rect 2696 3757 2824 3763
rect 2840 3757 3016 3763
rect 3256 3757 3336 3763
rect 3464 3757 3592 3763
rect 3672 3757 3768 3763
rect 3789 3763 3795 3777
rect 3928 3777 4040 3783
rect 4200 3777 4456 3783
rect 4648 3777 4760 3783
rect 5560 3777 5720 3783
rect 5896 3777 6024 3783
rect 6200 3777 6264 3783
rect 6312 3777 6323 3783
rect 6520 3777 6536 3783
rect 6856 3777 6888 3783
rect 3789 3757 4104 3763
rect 4120 3757 4216 3763
rect 4488 3757 4568 3763
rect 4584 3757 4744 3763
rect 4776 3757 4952 3763
rect 5240 3757 5512 3763
rect 5656 3757 5832 3763
rect 5928 3757 6168 3763
rect 6184 3757 6520 3763
rect 6776 3757 7544 3763
rect 2109 3748 2115 3752
rect 152 3737 312 3743
rect 328 3737 424 3743
rect 504 3737 552 3743
rect 872 3737 1368 3743
rect 1464 3737 1528 3743
rect 1640 3737 1720 3743
rect 1848 3737 1880 3743
rect 2136 3737 2168 3743
rect 2616 3737 2760 3743
rect 2808 3737 3032 3743
rect 3048 3737 3096 3743
rect 3112 3737 3128 3743
rect 3208 3737 4024 3743
rect 4056 3737 4136 3743
rect 4168 3737 4312 3743
rect 4632 3737 4840 3743
rect 5112 3737 5272 3743
rect 5496 3737 5656 3743
rect 5976 3737 6104 3743
rect 6280 3737 6440 3743
rect 6472 3737 6504 3743
rect 6760 3737 6808 3743
rect 6824 3737 6984 3743
rect 7112 3737 7336 3743
rect 7704 3737 7848 3743
rect 1741 3728 1747 3732
rect 1789 3728 1795 3732
rect -51 3717 8 3723
rect 264 3717 312 3723
rect 344 3717 616 3723
rect 1288 3717 1560 3723
rect 1768 3717 1784 3723
rect 2109 3717 2200 3723
rect 1629 3708 1635 3712
rect 296 3697 456 3703
rect 1080 3697 1624 3703
rect 2109 3703 2115 3717
rect 2440 3717 2584 3723
rect 2648 3717 2680 3723
rect 2712 3717 2776 3723
rect 3048 3717 3128 3723
rect 3192 3717 3224 3723
rect 3736 3717 3864 3723
rect 3896 3717 4072 3723
rect 4088 3717 4824 3723
rect 4984 3717 5000 3723
rect 5192 3717 5320 3723
rect 5592 3717 5704 3723
rect 5736 3717 5992 3723
rect 6008 3717 6040 3723
rect 6552 3717 6563 3723
rect 6712 3717 6760 3723
rect 6968 3717 7256 3723
rect 7288 3717 7368 3723
rect 1672 3697 2115 3703
rect 2136 3697 2152 3703
rect 2776 3697 2824 3703
rect 3032 3697 3048 3703
rect 3128 3697 3208 3703
rect 3416 3697 3480 3703
rect 3528 3697 3656 3703
rect 3704 3697 3736 3703
rect 3992 3697 4088 3703
rect 4104 3697 4136 3703
rect 4248 3697 4600 3703
rect 4616 3697 4664 3703
rect 4680 3697 4984 3703
rect 5688 3697 5704 3703
rect 6008 3697 6232 3703
rect 6344 3697 6616 3703
rect 6648 3697 6744 3703
rect 6856 3697 7128 3703
rect 7192 3697 7288 3703
rect 7640 3697 7704 3703
rect 7720 3697 7928 3703
rect 312 3677 344 3683
rect 1224 3677 1320 3683
rect 1352 3677 2568 3683
rect 2600 3677 3160 3683
rect 3192 3677 3448 3683
rect 3912 3677 5336 3683
rect 5704 3677 5736 3683
rect 6808 3677 6856 3683
rect 6872 3677 7160 3683
rect 7208 3677 7656 3683
rect 392 3657 1352 3663
rect 1485 3657 1544 3663
rect 1485 3643 1491 3657
rect 1656 3657 1752 3663
rect 1768 3657 2008 3663
rect 2376 3657 3736 3663
rect 3752 3657 5800 3663
rect 5880 3657 6088 3663
rect 6104 3657 6472 3663
rect 6840 3657 7096 3663
rect 7192 3657 7448 3663
rect 7464 3657 7928 3663
rect 7944 3657 8040 3663
rect 200 3637 1491 3643
rect 1512 3637 1560 3643
rect 1592 3637 2584 3643
rect 2632 3637 3368 3643
rect 3480 3637 3496 3643
rect 3848 3637 5192 3643
rect 5320 3637 5352 3643
rect 5368 3637 5496 3643
rect 7224 3637 7528 3643
rect 7544 3637 7592 3643
rect 7768 3637 7816 3643
rect 376 3617 440 3623
rect 1368 3617 2088 3623
rect 2744 3617 2808 3623
rect 1592 3597 2392 3603
rect 3080 3617 3128 3623
rect 4520 3597 4680 3603
rect 6744 3617 7000 3623
rect 6408 3597 6664 3603
rect 6680 3597 7032 3603
rect 7752 3617 7880 3623
rect 3277 3588 3283 3592
rect 3341 3588 3347 3592
rect 808 3577 1032 3583
rect 1448 3577 2312 3583
rect 2472 3577 2600 3583
rect 3368 3577 3448 3583
rect 3512 3577 3912 3583
rect 5144 3577 5256 3583
rect 5384 3577 5400 3583
rect 6920 3577 7016 3583
rect 7176 3577 7256 3583
rect -51 3557 200 3563
rect 1144 3557 1192 3563
rect 1208 3557 1731 3563
rect 248 3537 328 3543
rect 792 3537 808 3543
rect 1032 3537 1112 3543
rect 1400 3537 1704 3543
rect 1725 3543 1731 3557
rect 1800 3557 2056 3563
rect 2984 3557 3256 3563
rect 3272 3557 3512 3563
rect 4232 3557 4760 3563
rect 4888 3557 5128 3563
rect 5144 3557 5688 3563
rect 6680 3557 7192 3563
rect 7432 3557 7480 3563
rect 1725 3537 2792 3543
rect 2920 3537 3112 3543
rect 3128 3537 3224 3543
rect 3352 3537 3416 3543
rect 3432 3537 3464 3543
rect 3912 3537 4504 3543
rect 4680 3537 4712 3543
rect 4888 3537 5000 3543
rect 5080 3537 5304 3543
rect 5400 3537 5592 3543
rect 6888 3537 7112 3543
rect 7128 3537 7448 3543
rect 7496 3537 7560 3543
rect -51 3517 8 3523
rect 136 3517 392 3523
rect 408 3517 424 3523
rect 776 3517 1000 3523
rect 1016 3517 1080 3523
rect 1352 3517 1528 3523
rect 1544 3517 1800 3523
rect 1944 3517 2136 3523
rect 2520 3517 2536 3523
rect 2872 3517 2904 3523
rect 2936 3517 3016 3523
rect 3032 3517 3128 3523
rect 3160 3517 3224 3523
rect 3240 3517 3288 3523
rect 3336 3517 3496 3523
rect 3592 3517 3688 3523
rect 3704 3517 3720 3523
rect 4120 3517 4184 3523
rect 4525 3517 4536 3523
rect 4568 3517 4776 3523
rect 4792 3517 4936 3523
rect 5400 3517 5928 3523
rect 5976 3517 6120 3523
rect 6136 3517 6200 3523
rect 6440 3517 6664 3523
rect 6712 3517 6952 3523
rect 6984 3517 7064 3523
rect 7080 3517 7336 3523
rect 7352 3517 7432 3523
rect 7464 3517 7976 3523
rect 56 3497 136 3503
rect 184 3497 648 3503
rect 664 3497 728 3503
rect 744 3497 968 3503
rect 1032 3497 1304 3503
rect 1704 3497 1816 3503
rect 1928 3497 1960 3503
rect 1976 3497 2136 3503
rect 2200 3497 2248 3503
rect 2568 3497 2984 3503
rect 3096 3497 3128 3503
rect 3288 3497 3352 3503
rect 3368 3497 3432 3503
rect 3496 3497 3528 3503
rect 3544 3497 3800 3503
rect 3864 3497 4104 3503
rect 4168 3497 4280 3503
rect 4504 3497 4632 3503
rect 4728 3497 4744 3503
rect 4872 3497 5032 3503
rect 5048 3497 5192 3503
rect 5224 3497 5352 3503
rect 5368 3497 5416 3503
rect 5432 3497 5608 3503
rect 5736 3497 5992 3503
rect 6008 3497 6088 3503
rect 6232 3497 6472 3503
rect 6616 3497 6648 3503
rect 6952 3497 7208 3503
rect 7336 3497 7528 3503
rect 7560 3497 7656 3503
rect 280 3477 536 3483
rect 824 3477 840 3483
rect 1112 3477 1160 3483
rect 1544 3477 1688 3483
rect 2040 3477 2184 3483
rect 2856 3477 2904 3483
rect 3304 3477 3544 3483
rect 3560 3477 3608 3483
rect 3816 3477 3880 3483
rect 4152 3477 4376 3483
rect 4584 3477 4968 3483
rect 4984 3477 5080 3483
rect 5240 3477 5544 3483
rect 5560 3477 5624 3483
rect 5672 3477 5800 3483
rect 5896 3477 6024 3483
rect 6312 3477 6632 3483
rect 6648 3477 6712 3483
rect 6968 3477 7544 3483
rect 7560 3477 7576 3483
rect 7592 3477 7640 3483
rect 6957 3468 6963 3472
rect 776 3457 888 3463
rect 1272 3457 1400 3463
rect 1416 3457 1496 3463
rect 1512 3457 1912 3463
rect 2040 3457 2104 3463
rect 2568 3457 2600 3463
rect 2632 3457 2696 3463
rect 2712 3457 3128 3463
rect 3208 3457 3320 3463
rect 3432 3457 3592 3463
rect 3608 3457 4136 3463
rect 4408 3457 4600 3463
rect 4616 3457 4888 3463
rect 4920 3457 5240 3463
rect 5304 3457 5352 3463
rect 5384 3457 5395 3463
rect 5640 3457 6168 3463
rect 6184 3457 6232 3463
rect 6248 3457 6312 3463
rect 6584 3457 6744 3463
rect 6808 3457 6936 3463
rect 7288 3457 7400 3463
rect 1576 3437 1624 3443
rect 2168 3437 2264 3443
rect 2280 3437 2392 3443
rect 2680 3437 2744 3443
rect 2765 3437 3256 3443
rect 1272 3417 1528 3423
rect 888 3397 984 3403
rect 1240 3397 1640 3403
rect 1656 3397 1768 3403
rect 1784 3397 1928 3403
rect 2008 3417 2664 3423
rect 2765 3423 2771 3437
rect 3272 3437 3384 3443
rect 3400 3437 3416 3443
rect 4328 3437 4600 3443
rect 4616 3437 5064 3443
rect 5336 3437 5640 3443
rect 5800 3437 5976 3443
rect 5992 3437 6360 3443
rect 6648 3437 6840 3443
rect 6904 3437 6984 3443
rect 7304 3437 7784 3443
rect 2728 3417 2771 3423
rect 3048 3417 3112 3423
rect 3128 3417 3432 3423
rect 3448 3417 3640 3423
rect 2536 3397 2888 3403
rect 2904 3397 3064 3403
rect 3080 3397 3336 3403
rect 4696 3417 4728 3423
rect 4760 3417 4792 3423
rect 5080 3417 5192 3423
rect 4728 3397 4872 3403
rect 4904 3397 5192 3403
rect 5208 3397 5448 3403
rect 5512 3397 5720 3403
rect 5736 3397 5768 3403
rect 5784 3397 5864 3403
rect 6232 3417 6344 3423
rect -51 3377 1160 3383
rect 1192 3377 2776 3383
rect 2792 3377 3528 3383
rect 3544 3377 6328 3383
rect 6440 3377 6600 3383
rect 7144 3377 7480 3383
rect 7496 3377 7672 3383
rect 7688 3377 7736 3383
rect 7752 3377 7800 3383
rect 104 3357 312 3363
rect 696 3357 824 3363
rect 872 3357 1016 3363
rect 1032 3357 1080 3363
rect 1224 3357 1256 3363
rect 1352 3357 1368 3363
rect 1608 3357 1672 3363
rect 2408 3357 2456 3363
rect 2696 3357 2728 3363
rect 2792 3357 2888 3363
rect 3080 3357 3320 3363
rect 3336 3357 3432 3363
rect 4184 3357 4232 3363
rect 5416 3357 5544 3363
rect 6360 3357 6600 3363
rect 6616 3357 6808 3363
rect 6968 3357 7064 3363
rect 7176 3357 7192 3363
rect 7208 3357 7336 3363
rect 7549 3357 7912 3363
rect 4765 3348 4771 3352
rect -51 3337 216 3343
rect 232 3337 424 3343
rect 728 3337 744 3343
rect 920 3337 936 3343
rect 1016 3337 1064 3343
rect 1128 3337 1576 3343
rect 1624 3337 1800 3343
rect 2280 3337 2376 3343
rect 2712 3337 2808 3343
rect 2824 3337 3176 3343
rect 3320 3337 3416 3343
rect 4008 3337 4184 3343
rect 4312 3337 4323 3343
rect 4488 3337 4680 3343
rect 4824 3337 4984 3343
rect 5464 3337 5576 3343
rect 5592 3337 5619 3343
rect 5613 3328 5619 3337
rect 5864 3337 6120 3343
rect 6456 3337 6616 3343
rect 7112 3337 7128 3343
rect 7549 3343 7555 3357
rect 7144 3337 7555 3343
rect 7624 3337 7752 3343
rect 7896 3337 8024 3343
rect 200 3317 264 3323
rect 408 3317 664 3323
rect 744 3317 904 3323
rect 1176 3317 1240 3323
rect 1272 3317 1464 3323
rect 1608 3317 1896 3323
rect 2200 3317 2312 3323
rect 2504 3317 3048 3323
rect 3368 3317 3432 3323
rect 3752 3317 3784 3323
rect 3832 3317 3912 3323
rect 4584 3317 4696 3323
rect 5336 3317 5496 3323
rect 5768 3317 5784 3323
rect 6344 3317 6376 3323
rect 7208 3317 7240 3323
rect 7400 3317 7880 3323
rect 7896 3317 7992 3323
rect 381 3308 387 3312
rect 1261 3308 1267 3312
rect -51 3297 8 3303
rect 312 3297 360 3303
rect 680 3297 696 3303
rect 920 3297 1080 3303
rect 1144 3297 1208 3303
rect 1400 3297 1464 3303
rect 1816 3297 2136 3303
rect 2456 3297 2472 3303
rect 2824 3297 2936 3303
rect 3064 3297 3096 3303
rect 3400 3297 3544 3303
rect 4184 3297 4216 3303
rect 4664 3297 4744 3303
rect 4792 3297 4840 3303
rect 4856 3297 4920 3303
rect 5144 3297 5528 3303
rect 5544 3297 5576 3303
rect 5960 3297 5992 3303
rect 6040 3297 6408 3303
rect 6424 3297 6472 3303
rect 7000 3297 7176 3303
rect 7240 3297 7432 3303
rect 7576 3297 7624 3303
rect 7640 3297 7976 3303
rect 200 3277 584 3283
rect 824 3277 984 3283
rect 1288 3277 1448 3283
rect 1656 3277 1688 3283
rect 2040 3277 2584 3283
rect 2840 3277 2936 3283
rect 2952 3277 3144 3283
rect 3368 3277 3848 3283
rect 4328 3277 4712 3283
rect 7144 3277 7272 3283
rect 7320 3277 7560 3283
rect 7672 3277 7832 3283
rect 7928 3277 7944 3283
rect 168 3257 248 3263
rect 344 3257 360 3263
rect 376 3257 520 3263
rect 728 3257 1048 3263
rect 1240 3257 1320 3263
rect 1416 3257 1432 3263
rect 1480 3257 1608 3263
rect 2296 3257 2456 3263
rect 2472 3257 3048 3263
rect 3640 3257 3800 3263
rect 3816 3257 4104 3263
rect 5816 3257 7256 3263
rect 7272 3257 7544 3263
rect 7560 3257 7592 3263
rect 280 3237 632 3243
rect 909 3237 1096 3243
rect 909 3223 915 3237
rect 1272 3237 1368 3243
rect 1480 3237 1704 3243
rect 2072 3237 2888 3243
rect 2952 3237 3288 3243
rect 3304 3237 3368 3243
rect 3800 3237 4968 3243
rect 5992 3237 6088 3243
rect 6936 3237 7192 3243
rect 7768 3237 7816 3243
rect 7912 3237 7992 3243
rect 472 3217 915 3223
rect 984 3217 1832 3223
rect 2312 3217 2344 3223
rect 2360 3217 2632 3223
rect 1768 3197 2936 3203
rect 3128 3217 4200 3223
rect 3512 3197 3640 3203
rect 3656 3197 3752 3203
rect 4232 3197 4312 3203
rect 4328 3197 4776 3203
rect 5080 3217 5288 3223
rect 5304 3217 5336 3223
rect 7880 3217 8115 3223
rect 7704 3197 7960 3203
rect 733 3188 739 3192
rect 6669 3188 6675 3192
rect 6733 3188 6739 3192
rect 2280 3177 6568 3183
rect 6744 3177 6888 3183
rect 6904 3177 6920 3183
rect 7096 3177 7208 3183
rect 7816 3177 7896 3183
rect 7912 3177 8115 3183
rect -51 3157 72 3163
rect 88 3157 120 3163
rect 152 3157 632 3163
rect 680 3157 792 3163
rect 888 3157 1352 3163
rect 1432 3157 1736 3163
rect 1944 3157 2088 3163
rect 4072 3157 5064 3163
rect 7784 3157 7912 3163
rect 56 3137 136 3143
rect 168 3137 200 3143
rect 488 3137 792 3143
rect 1128 3137 1320 3143
rect 1848 3137 2552 3143
rect 2584 3137 2632 3143
rect 2648 3137 2680 3143
rect 2696 3137 2776 3143
rect 2904 3137 3160 3143
rect 3832 3137 4328 3143
rect 4504 3137 5160 3143
rect 5384 3137 6040 3143
rect 6152 3137 6184 3143
rect 6200 3137 6328 3143
rect 6360 3137 6408 3143
rect 6648 3137 6792 3143
rect 6808 3137 6952 3143
rect 7160 3137 7208 3143
rect 7224 3137 7288 3143
rect 7576 3137 7688 3143
rect 7768 3137 7800 3143
rect 7848 3137 8008 3143
rect 8072 3137 8115 3143
rect -51 3117 24 3123
rect 40 3117 104 3123
rect 120 3117 184 3123
rect 424 3117 440 3123
rect 712 3117 840 3123
rect 1160 3117 1192 3123
rect 1208 3117 1272 3123
rect 1336 3117 1496 3123
rect 1672 3117 1720 3123
rect 1736 3117 2104 3123
rect 2696 3117 3176 3123
rect 3240 3117 3400 3123
rect 3848 3117 3976 3123
rect 4280 3117 4424 3123
rect 4728 3117 4744 3123
rect 4776 3117 5160 3123
rect 5304 3117 5560 3123
rect 5576 3117 5800 3123
rect 6056 3117 6232 3123
rect 6520 3117 7075 3123
rect 184 3097 360 3103
rect 408 3097 520 3103
rect 824 3097 872 3103
rect 1048 3097 1144 3103
rect 1272 3097 1432 3103
rect 1448 3097 1624 3103
rect 1640 3097 1688 3103
rect 1880 3097 2040 3103
rect 2136 3097 2296 3103
rect 2424 3097 2456 3103
rect 2952 3097 3432 3103
rect 3448 3097 3544 3103
rect 3560 3097 3672 3103
rect 3752 3097 3912 3103
rect 3960 3097 4040 3103
rect 4264 3097 4312 3103
rect 4984 3097 5096 3103
rect 5272 3097 5320 3103
rect 5336 3097 5384 3103
rect 5944 3097 6120 3103
rect 6152 3097 6456 3103
rect 6536 3097 6648 3103
rect 6664 3097 6696 3103
rect 7069 3103 7075 3117
rect 7496 3117 7608 3123
rect 7640 3117 7672 3123
rect 7800 3117 7816 3123
rect 7832 3117 7864 3123
rect 7069 3097 7832 3103
rect 7848 3097 8056 3103
rect 93 3083 99 3092
rect 93 3077 104 3083
rect 792 3077 824 3083
rect 984 3077 1240 3083
rect 1256 3077 1640 3083
rect 1656 3077 1720 3083
rect 1800 3077 1976 3083
rect 2008 3077 2168 3083
rect 2184 3077 2392 3083
rect 2424 3077 2664 3083
rect 2952 3077 3000 3083
rect 3032 3077 3043 3083
rect 3352 3077 3512 3083
rect 3576 3077 3768 3083
rect 3880 3077 3960 3083
rect 3976 3077 4360 3083
rect 4856 3077 4872 3083
rect 4888 3077 5032 3083
rect 5080 3077 5208 3083
rect 5224 3077 5416 3083
rect 5656 3077 5848 3083
rect 5864 3077 6072 3083
rect 6184 3077 6264 3083
rect 6344 3077 6376 3083
rect 6392 3077 6504 3083
rect 6696 3077 6760 3083
rect 6776 3077 6840 3083
rect 7048 3077 7112 3083
rect 7128 3077 7144 3083
rect 7309 3077 7848 3083
rect 56 3057 536 3063
rect 552 3057 872 3063
rect 1160 3057 1528 3063
rect 1544 3057 1608 3063
rect 1688 3057 2072 3063
rect 2296 3057 2376 3063
rect 2408 3057 2440 3063
rect 2488 3057 2504 3063
rect 2520 3057 2808 3063
rect 2840 3057 3112 3063
rect 3128 3057 3576 3063
rect 3784 3057 4008 3063
rect 4024 3057 4232 3063
rect 4360 3057 4488 3063
rect 5048 3057 5272 3063
rect 5304 3057 5976 3063
rect 6280 3057 6472 3063
rect 7309 3063 7315 3077
rect 8109 3083 8115 3103
rect 7864 3077 8115 3083
rect 6488 3057 7315 3063
rect 7720 3057 7880 3063
rect 232 3037 296 3043
rect 920 3037 1176 3043
rect 1192 3037 1304 3043
rect 1320 3037 1384 3043
rect 1400 3037 1512 3043
rect 1528 3037 1576 3043
rect 2360 3037 2536 3043
rect 2616 3037 2824 3043
rect 2856 3037 3208 3043
rect 3240 3037 3656 3043
rect 3981 3037 4099 3043
rect 776 3017 1432 3023
rect 184 2997 200 3003
rect 936 2997 1224 3003
rect 1240 2997 1427 3003
rect 2344 3017 2584 3023
rect 3981 3023 3987 3037
rect 2600 3017 3987 3023
rect 4093 3023 4099 3037
rect 4120 3037 5768 3043
rect 5784 3037 5992 3043
rect 6013 3037 6120 3043
rect 328 2977 408 2983
rect 552 2977 712 2983
rect 1080 2977 1256 2983
rect 1421 2983 1427 2997
rect 2216 2997 2648 3003
rect 2664 2997 2968 3003
rect 3000 2997 3432 3003
rect 3448 2997 3560 3003
rect 3816 2997 3896 3003
rect 4093 3017 4664 3023
rect 6013 3023 6019 3037
rect 6152 3037 6184 3043
rect 8109 3043 8115 3063
rect 6568 3037 8115 3043
rect 5416 3017 6019 3023
rect 4056 2997 4152 3003
rect 4248 2997 4296 3003
rect 4568 2997 4856 3003
rect 5272 2997 5320 3003
rect 5528 2997 5576 3003
rect 5864 2997 5928 3003
rect 6216 3017 6280 3023
rect 6680 3017 6936 3023
rect 7816 3017 7832 3023
rect 6248 2997 6536 3003
rect 6664 2997 6792 3003
rect 6824 2997 6952 3003
rect 6968 2997 7000 3003
rect 7560 2997 7576 3003
rect 7592 2997 7768 3003
rect 1421 2977 2152 2983
rect 2232 2977 2488 2983
rect 2509 2977 2776 2983
rect 1405 2968 1411 2972
rect -51 2957 440 2963
rect 456 2957 648 2963
rect 680 2957 776 2963
rect 840 2957 1080 2963
rect 1325 2957 1336 2963
rect 1432 2957 1464 2963
rect 1901 2957 1912 2963
rect 2088 2957 2168 2963
rect 2200 2957 2232 2963
rect 2509 2963 2515 2977
rect 2792 2977 2904 2983
rect 2920 2977 4728 2983
rect 4872 2977 4984 2983
rect 5000 2977 5112 2983
rect 5160 2977 5352 2983
rect 5368 2977 5832 2983
rect 5848 2977 6296 2983
rect 6312 2977 6744 2983
rect 6760 2977 7016 2983
rect 7032 2977 7720 2983
rect 2440 2957 2515 2963
rect 2936 2957 3048 2963
rect 3064 2957 3352 2963
rect 3464 2957 3816 2963
rect 4168 2957 4632 2963
rect 4888 2957 5144 2963
rect 5240 2957 5272 2963
rect 5320 2957 5864 2963
rect 5992 2957 6152 2963
rect 6168 2957 6552 2963
rect 6648 2957 6712 2963
rect 56 2937 152 2943
rect 744 2937 1240 2943
rect 1256 2937 1560 2943
rect 1592 2937 1768 2943
rect 1784 2937 1912 2943
rect 1928 2937 1992 2943
rect 2632 2937 2712 2943
rect 2744 2937 2840 2943
rect 3080 2937 3192 2943
rect 3384 2937 3416 2943
rect 3432 2937 3448 2943
rect 3752 2937 3864 2943
rect 3912 2937 4200 2943
rect 4312 2937 4440 2943
rect 4584 2937 4744 2943
rect 4792 2937 4936 2943
rect 4952 2937 5176 2943
rect 5192 2937 5304 2943
rect 5320 2937 5976 2943
rect 5992 2937 6104 2943
rect 6120 2937 6680 2943
rect 6904 2937 7064 2943
rect 7336 2937 7352 2943
rect 7368 2937 7464 2943
rect 7480 2937 7640 2943
rect 3549 2928 3555 2932
rect -51 2903 -45 2923
rect 264 2917 296 2923
rect 360 2917 456 2923
rect 472 2917 680 2923
rect 888 2917 1032 2923
rect 1288 2917 1400 2923
rect 1640 2917 1656 2923
rect 1672 2917 1784 2923
rect 1896 2917 1912 2923
rect 2024 2917 2040 2923
rect 2056 2917 2088 2923
rect 2104 2917 2136 2923
rect 2648 2917 2712 2923
rect 2728 2917 3192 2923
rect 3272 2917 3336 2923
rect 3736 2917 3848 2923
rect 4360 2917 4456 2923
rect 4824 2917 5208 2923
rect 5320 2917 5400 2923
rect 5432 2917 5896 2923
rect 5912 2917 5944 2923
rect 5960 2917 6616 2923
rect 6632 2917 6664 2923
rect 6728 2917 6920 2923
rect 7080 2917 7160 2923
rect 7352 2917 7448 2923
rect 7464 2917 7608 2923
rect 7640 2917 7672 2923
rect 7752 2917 7880 2923
rect -51 2897 408 2903
rect 808 2897 1160 2903
rect 1176 2897 1208 2903
rect 1608 2897 1672 2903
rect 1736 2897 1864 2903
rect 2989 2897 3000 2903
rect 3128 2897 3320 2903
rect 3432 2897 3928 2903
rect 4280 2897 4360 2903
rect 4472 2897 4712 2903
rect 4952 2897 4968 2903
rect 4984 2897 5080 2903
rect 5128 2897 5208 2903
rect 5224 2897 5288 2903
rect 5336 2897 5347 2903
rect 5512 2897 5544 2903
rect 5944 2897 6136 2903
rect 6152 2897 6216 2903
rect 6504 2897 6600 2903
rect 6616 2897 6712 2903
rect 7064 2897 7304 2903
rect 7656 2897 7896 2903
rect 984 2877 1976 2883
rect 2200 2877 2328 2883
rect 2344 2877 2456 2883
rect 2792 2877 3064 2883
rect 3320 2877 3400 2883
rect 4184 2877 4408 2883
rect 5480 2877 5800 2883
rect 5816 2877 5944 2883
rect 5960 2877 6168 2883
rect 6712 2877 7000 2883
rect 7608 2877 7704 2883
rect 7720 2877 7784 2883
rect 712 2857 744 2863
rect 760 2857 1288 2863
rect 1512 2857 2200 2863
rect 2216 2857 2280 2863
rect 2296 2857 2792 2863
rect 2824 2857 5368 2863
rect 7640 2857 7752 2863
rect 600 2837 1752 2843
rect 2136 2837 2568 2843
rect 2968 2837 3032 2843
rect 3784 2837 5880 2843
rect 6584 2837 7288 2843
rect 648 2817 792 2823
rect 840 2797 888 2803
rect 1976 2817 2056 2823
rect 2072 2817 2696 2823
rect 2712 2817 2808 2823
rect 1464 2797 1528 2803
rect 1544 2797 1704 2803
rect 1720 2797 2072 2803
rect 2088 2797 2600 2803
rect 3608 2817 3736 2823
rect 3005 2797 4984 2803
rect 696 2777 792 2783
rect 1448 2777 1496 2783
rect 1512 2777 1768 2783
rect 1784 2777 2008 2783
rect 3005 2783 3011 2797
rect 6024 2817 6552 2823
rect 6184 2797 6248 2803
rect 6472 2797 6696 2803
rect 2040 2777 3011 2783
rect 3160 2777 4408 2783
rect 5576 2777 5640 2783
rect 6104 2777 6344 2783
rect 168 2757 328 2763
rect 344 2757 1688 2763
rect 1736 2757 2088 2763
rect 2104 2757 2648 2763
rect 2664 2757 3336 2763
rect 3784 2757 3816 2763
rect 4680 2757 4744 2763
rect 4760 2757 4792 2763
rect 4808 2757 5128 2763
rect 5656 2757 5736 2763
rect 6008 2757 6296 2763
rect 200 2737 296 2743
rect 312 2737 552 2743
rect 2072 2737 2120 2743
rect 2312 2737 2488 2743
rect 2808 2737 3448 2743
rect 3560 2737 3640 2743
rect 4024 2737 4840 2743
rect 5784 2737 6200 2743
rect 6376 2737 6408 2743
rect 264 2717 360 2723
rect 696 2717 1016 2723
rect 1592 2717 2152 2723
rect 2168 2717 2296 2723
rect 2504 2717 2632 2723
rect 2840 2717 3000 2723
rect 3448 2717 3496 2723
rect 3576 2717 3603 2723
rect 840 2697 1176 2703
rect 1256 2697 1400 2703
rect 1560 2697 1656 2703
rect 1704 2697 1800 2703
rect 1816 2697 2024 2703
rect 2120 2697 2296 2703
rect 2312 2697 2472 2703
rect 2616 2697 2648 2703
rect 2952 2697 3016 2703
rect 3096 2697 3576 2703
rect 3597 2703 3603 2717
rect 3656 2717 3752 2723
rect 4728 2717 4776 2723
rect 4792 2717 4872 2723
rect 4888 2717 4936 2723
rect 5464 2717 5544 2723
rect 5560 2717 5608 2723
rect 5624 2717 5672 2723
rect 5736 2717 6040 2723
rect 6168 2717 6264 2723
rect 6344 2717 6392 2723
rect 6440 2717 6488 2723
rect 6904 2717 6968 2723
rect 7032 2717 7176 2723
rect 7464 2717 7480 2723
rect 3597 2697 3976 2703
rect 4088 2697 4328 2703
rect 4568 2697 4664 2703
rect 4920 2697 5080 2703
rect 5352 2697 5448 2703
rect 5960 2697 6008 2703
rect 6040 2697 6056 2703
rect 6072 2697 6552 2703
rect 6584 2697 6680 2703
rect 6808 2697 6888 2703
rect 7176 2697 7208 2703
rect 344 2677 472 2683
rect 536 2677 904 2683
rect 1384 2677 2392 2683
rect 2648 2677 2664 2683
rect 2680 2677 3032 2683
rect 3096 2677 3144 2683
rect 3160 2677 3384 2683
rect 3432 2677 3512 2683
rect 3528 2677 3592 2683
rect 3720 2677 3848 2683
rect 4136 2677 4216 2683
rect 4472 2677 4632 2683
rect 4856 2677 4952 2683
rect 5176 2677 5272 2683
rect 5768 2677 5912 2683
rect 6056 2677 6088 2683
rect 6120 2677 6232 2683
rect 6264 2677 6488 2683
rect 6536 2677 6568 2683
rect 6712 2677 6856 2683
rect 7144 2677 7256 2683
rect 7272 2677 7448 2683
rect 6109 2668 6115 2672
rect 104 2657 216 2663
rect 1336 2657 1480 2663
rect 1880 2657 2216 2663
rect 2280 2657 2312 2663
rect 2600 2657 2760 2663
rect 2776 2657 2904 2663
rect 3048 2657 3880 2663
rect 3896 2657 4056 2663
rect 4072 2657 4264 2663
rect 5256 2657 5416 2663
rect 5896 2657 5912 2663
rect 5928 2657 5944 2663
rect 6136 2657 6184 2663
rect 6200 2657 6584 2663
rect 7048 2657 7224 2663
rect 7304 2657 7816 2663
rect 168 2637 216 2643
rect 1032 2637 1496 2643
rect 1688 2637 1720 2643
rect 2056 2637 2120 2643
rect 2568 2637 2776 2643
rect 3080 2637 3112 2643
rect 3128 2637 3416 2643
rect 3608 2637 3928 2643
rect 3944 2637 3976 2643
rect 3992 2637 4040 2643
rect 5400 2637 5528 2643
rect 5544 2637 5624 2643
rect 5640 2637 6408 2643
rect 6488 2637 6568 2643
rect 6952 2637 7336 2643
rect 520 2617 600 2623
rect 712 2617 744 2623
rect 824 2617 1048 2623
rect 1416 2617 1464 2623
rect 1480 2617 1864 2623
rect 184 2597 264 2603
rect 456 2597 552 2603
rect 568 2597 968 2603
rect 1000 2597 1320 2603
rect 1400 2597 1640 2603
rect 1752 2597 1784 2603
rect 2184 2617 3896 2623
rect 2168 2597 2232 2603
rect 3832 2597 3864 2603
rect 3880 2597 3960 2603
rect 5864 2617 5880 2623
rect 4792 2597 5496 2603
rect 6232 2617 6264 2623
rect 6296 2617 6424 2623
rect 6440 2617 7480 2623
rect 7800 2617 7864 2623
rect 7880 2617 7976 2623
rect 6104 2597 6296 2603
rect 6328 2597 6456 2603
rect 6952 2597 7512 2603
rect 7528 2597 7624 2603
rect 136 2577 376 2583
rect 392 2577 856 2583
rect 872 2577 904 2583
rect 1288 2577 1507 2583
rect 296 2557 328 2563
rect 584 2557 680 2563
rect 712 2557 840 2563
rect 1320 2557 1368 2563
rect 1437 2557 1480 2563
rect 408 2537 600 2543
rect 888 2537 1048 2543
rect 1064 2537 1192 2543
rect 1437 2543 1443 2557
rect 1501 2563 1507 2577
rect 1720 2577 2312 2583
rect 2328 2577 2344 2583
rect 2360 2577 2472 2583
rect 2744 2577 2936 2583
rect 3496 2577 3528 2583
rect 3544 2577 3672 2583
rect 3688 2577 3752 2583
rect 3768 2577 4072 2583
rect 4184 2577 4280 2583
rect 5608 2577 6392 2583
rect 6408 2577 6936 2583
rect 7016 2577 7048 2583
rect 7064 2577 7144 2583
rect 7688 2577 7704 2583
rect 1501 2557 1864 2563
rect 1928 2557 1944 2563
rect 2136 2557 2360 2563
rect 2408 2557 2440 2563
rect 2456 2557 2568 2563
rect 2664 2557 2696 2563
rect 2712 2557 2776 2563
rect 2792 2557 2888 2563
rect 2904 2557 3720 2563
rect 3736 2557 4488 2563
rect 5912 2557 6136 2563
rect 6232 2557 6360 2563
rect 7704 2557 7784 2563
rect 1320 2537 1443 2543
rect 1944 2537 1992 2543
rect 2024 2537 2232 2543
rect 2328 2537 2504 2543
rect 2760 2537 3064 2543
rect 3400 2537 3448 2543
rect 3688 2537 3784 2543
rect 3800 2537 3944 2543
rect 4008 2537 4168 2543
rect 4248 2537 4376 2543
rect 4424 2537 4536 2543
rect 4552 2537 4712 2543
rect 4824 2537 4936 2543
rect 4952 2537 5112 2543
rect 5624 2537 5720 2543
rect 5736 2537 5832 2543
rect 6280 2537 6520 2543
rect 6744 2537 6808 2543
rect 6872 2537 6952 2543
rect 6968 2537 7064 2543
rect 200 2517 456 2523
rect 504 2517 536 2523
rect 936 2517 1064 2523
rect 1432 2517 1544 2523
rect 1688 2517 1736 2523
rect 1896 2517 1928 2523
rect 2104 2517 2168 2523
rect 2216 2517 2312 2523
rect 2504 2517 2552 2523
rect 2776 2517 2872 2523
rect 2952 2517 3256 2523
rect 3288 2517 3496 2523
rect 3560 2517 3624 2523
rect 3912 2517 3992 2523
rect 4088 2517 4104 2523
rect 4312 2517 4424 2523
rect 4440 2517 4568 2523
rect 4648 2517 4744 2523
rect 4888 2517 4920 2523
rect 4984 2517 5128 2523
rect 5240 2517 5304 2523
rect 5320 2517 5416 2523
rect 5544 2517 5656 2523
rect 5752 2517 5768 2523
rect 6008 2517 6040 2523
rect 6056 2517 6312 2523
rect 6408 2517 6520 2523
rect 6536 2517 6744 2523
rect 7032 2517 7192 2523
rect 7416 2517 7480 2523
rect 7592 2517 7640 2523
rect 7656 2517 7864 2523
rect 7960 2517 8024 2523
rect 88 2497 312 2503
rect 808 2497 840 2503
rect 920 2497 968 2503
rect 1048 2497 1256 2503
rect 1576 2497 1624 2503
rect 2072 2497 2184 2503
rect 3528 2497 3912 2503
rect 4104 2497 4136 2503
rect 4760 2497 4792 2503
rect 4920 2497 4984 2503
rect 5256 2497 5720 2503
rect 5736 2497 6024 2503
rect 6328 2497 6712 2503
rect 6728 2497 6776 2503
rect 7000 2497 7032 2503
rect 7608 2497 7688 2503
rect 152 2477 360 2483
rect 776 2477 1016 2483
rect 1096 2477 1528 2483
rect 1624 2477 1688 2483
rect 2328 2477 2632 2483
rect 2808 2477 3048 2483
rect 3608 2477 4056 2483
rect 4264 2477 4776 2483
rect 5096 2477 5352 2483
rect 5368 2477 5544 2483
rect 5656 2477 5688 2483
rect 5704 2477 5832 2483
rect 5864 2477 6008 2483
rect 6024 2477 6344 2483
rect 6440 2477 6792 2483
rect 6808 2477 7160 2483
rect 7176 2477 7352 2483
rect 7368 2477 7416 2483
rect 7432 2477 7512 2483
rect 7528 2477 7736 2483
rect 1016 2457 1032 2463
rect 1064 2457 1400 2463
rect 1480 2457 1512 2463
rect 1528 2457 1752 2463
rect 1848 2457 2264 2463
rect 2680 2457 2744 2463
rect 2760 2457 4968 2463
rect 7000 2457 7096 2463
rect 7624 2457 7944 2463
rect 216 2437 328 2443
rect 1032 2437 1064 2443
rect 1208 2437 1288 2443
rect 1352 2437 1768 2443
rect 1896 2437 1992 2443
rect 2024 2437 2072 2443
rect 2280 2437 2392 2443
rect 2408 2437 2936 2443
rect 3864 2437 4072 2443
rect 4248 2437 5704 2443
rect 6744 2437 7048 2443
rect 7496 2437 7624 2443
rect 760 2397 792 2403
rect 984 2417 1256 2423
rect 1672 2417 2792 2423
rect 1128 2397 1304 2403
rect 2072 2397 2120 2403
rect 4072 2417 4328 2423
rect 3576 2397 3736 2403
rect 3752 2397 3864 2403
rect 5208 2417 6728 2423
rect 5928 2397 6200 2403
rect 7224 2417 7672 2423
rect 7720 2417 7784 2423
rect 7640 2397 7800 2403
rect 7816 2397 7848 2403
rect 7864 2397 7992 2403
rect 280 2377 408 2383
rect 424 2377 824 2383
rect 856 2377 1592 2383
rect 1624 2377 1736 2383
rect 1912 2377 3736 2383
rect 5896 2377 6136 2383
rect 6360 2377 6424 2383
rect 6584 2377 6595 2383
rect 6664 2377 7656 2383
rect -51 2357 712 2363
rect 872 2357 1048 2363
rect 1080 2357 1160 2363
rect 1176 2357 1576 2363
rect 1592 2357 1704 2363
rect 1768 2357 2712 2363
rect 3576 2357 4248 2363
rect 6184 2357 6744 2363
rect 6968 2357 7384 2363
rect 7560 2357 7656 2363
rect 376 2337 408 2343
rect 760 2337 808 2343
rect 824 2337 968 2343
rect 1000 2337 1187 2343
rect -51 2317 8 2323
rect 136 2317 296 2323
rect 328 2317 696 2323
rect 728 2317 984 2323
rect 1181 2323 1187 2337
rect 1208 2337 1224 2343
rect 1256 2337 1768 2343
rect 2168 2337 2248 2343
rect 2424 2337 3080 2343
rect 3416 2337 3496 2343
rect 3720 2337 3800 2343
rect 5464 2337 5480 2343
rect 5880 2337 5960 2343
rect 6344 2337 6840 2343
rect 7576 2337 7848 2343
rect 1181 2317 1240 2323
rect 1336 2317 1640 2323
rect 1752 2317 1800 2323
rect 1992 2317 2040 2323
rect 2296 2317 2344 2323
rect 2360 2317 3032 2323
rect 3160 2317 3480 2323
rect 3496 2317 3544 2323
rect 3560 2317 3768 2323
rect 3848 2317 4056 2323
rect 4312 2317 4360 2323
rect 4856 2317 4872 2323
rect 5480 2317 5512 2323
rect 5528 2317 5640 2323
rect 5656 2317 5704 2323
rect 5752 2317 5912 2323
rect 5928 2317 6312 2323
rect 6536 2317 6776 2323
rect 6808 2317 6904 2323
rect 7416 2317 7464 2323
rect 168 2297 200 2303
rect 216 2297 264 2303
rect 376 2297 408 2303
rect 728 2297 1064 2303
rect 1080 2297 1128 2303
rect 1832 2297 1880 2303
rect 1912 2297 1923 2303
rect 2120 2297 2296 2303
rect 2328 2297 2472 2303
rect 3064 2297 3144 2303
rect 3368 2297 3640 2303
rect 3800 2297 3880 2303
rect 4360 2297 4408 2303
rect 4888 2297 5240 2303
rect 5368 2297 5464 2303
rect 5672 2297 5816 2303
rect 5880 2297 6248 2303
rect 6296 2297 6307 2303
rect 6680 2297 6712 2303
rect 6776 2297 6824 2303
rect 6872 2297 6920 2303
rect 7160 2297 7272 2303
rect 7624 2297 7816 2303
rect 6253 2288 6259 2292
rect 184 2277 392 2283
rect 408 2277 568 2283
rect 584 2277 616 2283
rect 680 2277 1032 2283
rect 1272 2277 1336 2283
rect 1384 2277 1432 2283
rect 1768 2277 1864 2283
rect 2392 2277 2552 2283
rect 2888 2277 2984 2283
rect 3128 2277 3256 2283
rect 3336 2277 3432 2283
rect 3656 2277 3848 2283
rect 4376 2277 4840 2283
rect 4856 2277 4984 2283
rect 5016 2277 5624 2283
rect 5640 2277 5960 2283
rect 6280 2277 6392 2283
rect 6424 2277 6632 2283
rect 7208 2277 7352 2283
rect 7512 2277 7544 2283
rect 7560 2277 7720 2283
rect 1160 2257 1320 2263
rect 1480 2257 1832 2263
rect 1848 2257 2056 2263
rect 2440 2257 3768 2263
rect 4472 2257 4520 2263
rect 4840 2257 4936 2263
rect 5400 2257 5496 2263
rect 5512 2257 6024 2263
rect 6232 2257 6280 2263
rect 6408 2257 6472 2263
rect 6504 2257 6584 2263
rect 6600 2257 6984 2263
rect 7112 2257 7256 2263
rect 7272 2257 7320 2263
rect 7368 2257 7416 2263
rect 616 2237 952 2243
rect 968 2237 984 2243
rect 1000 2237 1288 2243
rect 1512 2237 1544 2243
rect 1576 2237 1608 2243
rect 1624 2237 2424 2243
rect 2568 2237 3192 2243
rect 3224 2237 4184 2243
rect 4296 2237 4344 2243
rect 4360 2237 4568 2243
rect 5112 2237 5528 2243
rect 5544 2237 5672 2243
rect 6024 2237 6072 2243
rect 6504 2237 6696 2243
rect 6712 2237 6888 2243
rect 6904 2237 6984 2243
rect 7176 2237 7400 2243
rect 1192 2217 1560 2223
rect 1624 2217 1688 2223
rect 648 2197 808 2203
rect 824 2197 872 2203
rect 888 2197 1368 2203
rect 2648 2217 3064 2223
rect 2072 2197 2296 2203
rect 2728 2197 2776 2203
rect 5848 2217 5896 2223
rect 4152 2197 4296 2203
rect 5304 2197 5544 2203
rect 5704 2197 5928 2203
rect 6264 2217 6504 2223
rect 7256 2217 7480 2223
rect 6200 2197 6664 2203
rect 6936 2197 7128 2203
rect 7144 2197 7288 2203
rect 7320 2197 7368 2203
rect 7592 2197 7704 2203
rect 792 2177 936 2183
rect 984 2177 1112 2183
rect 1464 2177 1592 2183
rect 2200 2177 3208 2183
rect 3224 2177 5064 2183
rect 5192 2177 5592 2183
rect 5640 2177 5784 2183
rect 5800 2177 6296 2183
rect 6312 2177 6440 2183
rect 6856 2177 7000 2183
rect 7416 2177 7976 2183
rect 552 2157 1096 2163
rect 1112 2157 2216 2163
rect 2232 2157 2264 2163
rect 2328 2157 3032 2163
rect 3160 2157 3208 2163
rect 3224 2157 3544 2163
rect 4280 2157 4312 2163
rect 4744 2157 4808 2163
rect 4936 2157 5176 2163
rect 5320 2157 5576 2163
rect 5592 2157 5752 2163
rect 7592 2157 7640 2163
rect 328 2137 456 2143
rect 840 2137 1032 2143
rect 1048 2137 1288 2143
rect 1368 2137 1416 2143
rect 1480 2137 1528 2143
rect 1928 2137 2168 2143
rect 2216 2137 2376 2143
rect 2392 2137 2456 2143
rect 2776 2137 2872 2143
rect 2904 2137 3096 2143
rect 3112 2137 3144 2143
rect 3576 2137 3592 2143
rect 3880 2137 3960 2143
rect 3992 2137 4136 2143
rect 4589 2137 4616 2143
rect 1677 2128 1683 2132
rect 104 2117 168 2123
rect 472 2117 552 2123
rect 792 2117 888 2123
rect 1208 2117 1416 2123
rect 1432 2117 1512 2123
rect 1576 2117 1608 2123
rect 1896 2117 2008 2123
rect 2232 2117 2328 2123
rect 2504 2117 2536 2123
rect 2696 2117 2787 2123
rect 696 2097 760 2103
rect 856 2097 1080 2103
rect 1224 2097 1544 2103
rect 1704 2097 1976 2103
rect 2040 2097 2328 2103
rect 2360 2097 2408 2103
rect 2456 2097 2488 2103
rect 2568 2097 2680 2103
rect 2781 2103 2787 2117
rect 2808 2117 2824 2123
rect 3064 2117 3128 2123
rect 3144 2117 3256 2123
rect 3432 2117 3512 2123
rect 3800 2117 3912 2123
rect 4104 2117 4168 2123
rect 4589 2123 4595 2137
rect 4680 2137 4760 2143
rect 4776 2137 5096 2143
rect 5192 2137 5352 2143
rect 5373 2137 5400 2143
rect 4504 2117 4595 2123
rect 4616 2117 4648 2123
rect 4728 2117 4792 2123
rect 5080 2117 5128 2123
rect 5373 2123 5379 2137
rect 5464 2137 5592 2143
rect 5672 2137 5784 2143
rect 6120 2137 6152 2143
rect 6792 2137 6920 2143
rect 7672 2137 7752 2143
rect 7768 2137 7880 2143
rect 5288 2117 5379 2123
rect 5400 2117 5432 2123
rect 5592 2117 5704 2123
rect 6024 2117 6264 2123
rect 6520 2117 6680 2123
rect 6856 2117 6952 2123
rect 7416 2117 7432 2123
rect 7528 2117 7560 2123
rect 7608 2117 7672 2123
rect 7704 2117 7880 2123
rect 2781 2097 2808 2103
rect 3000 2097 3032 2103
rect 3048 2097 3704 2103
rect 3912 2097 4104 2103
rect 4536 2097 4680 2103
rect 5768 2097 5848 2103
rect 5960 2097 5976 2103
rect 5992 2097 6072 2103
rect 6168 2097 6216 2103
rect 6408 2097 6472 2103
rect 6968 2097 7000 2103
rect 7032 2097 7656 2103
rect 7896 2097 7912 2103
rect 152 2077 504 2083
rect 552 2077 600 2083
rect 616 2077 648 2083
rect 1272 2077 1848 2083
rect 2696 2077 3112 2083
rect 3256 2077 3352 2083
rect 3912 2077 4008 2083
rect 4888 2077 4936 2083
rect 7416 2077 7464 2083
rect 7496 2077 7592 2083
rect 7640 2077 7768 2083
rect 7800 2077 7928 2083
rect 1736 2057 3208 2063
rect 3336 2057 3576 2063
rect 4360 2057 5848 2063
rect 888 2037 952 2043
rect 984 2037 1656 2043
rect 1672 2037 2888 2043
rect 2904 2037 3112 2043
rect 3592 2037 3624 2043
rect 3768 2037 4760 2043
rect 4776 2037 4888 2043
rect 7864 2037 7992 2043
rect 1784 2017 2568 2023
rect 1592 1997 1784 2003
rect 2328 1997 2344 2003
rect 3192 2017 3960 2023
rect 3976 2017 4040 2023
rect 4200 2017 4296 2023
rect 4312 2017 4840 2023
rect 3005 1997 3672 2003
rect 456 1977 984 1983
rect 1528 1977 2184 1983
rect 2872 1977 2936 1983
rect 3005 1983 3011 1997
rect 3688 1997 4824 2003
rect 2952 1977 3011 1983
rect 3208 1977 3912 1983
rect 3928 1977 4056 1983
rect 4152 1977 4264 1983
rect 4888 1977 5288 1983
rect 5880 1977 6456 1983
rect 88 1957 968 1963
rect 1112 1957 1128 1963
rect 1144 1957 1992 1963
rect 2952 1957 2968 1963
rect 3112 1957 3176 1963
rect 3320 1957 3368 1963
rect 3496 1957 4984 1963
rect 5000 1957 5224 1963
rect 5240 1957 5272 1963
rect 5944 1957 6184 1963
rect 6712 1957 6760 1963
rect 7640 1957 7688 1963
rect 7704 1957 7832 1963
rect 248 1937 280 1943
rect 344 1937 552 1943
rect 568 1937 824 1943
rect 1544 1937 1560 1943
rect 2504 1937 3416 1943
rect 3464 1937 3608 1943
rect 3880 1937 3992 1943
rect 4008 1937 4200 1943
rect 5112 1937 5256 1943
rect 5304 1937 5320 1943
rect 5880 1937 5944 1943
rect 5976 1937 5992 1943
rect 6344 1937 6568 1943
rect 6584 1937 6616 1943
rect 6680 1937 6696 1943
rect 6744 1937 7192 1943
rect 7736 1937 7944 1943
rect 568 1917 664 1923
rect 808 1917 888 1923
rect 1576 1917 1688 1923
rect 1768 1917 1864 1923
rect 3080 1917 3192 1923
rect 3480 1917 3528 1923
rect 4024 1917 4200 1923
rect 4216 1917 4328 1923
rect 4344 1917 4392 1923
rect 4568 1917 4728 1923
rect 4840 1917 5400 1923
rect 5416 1917 6280 1923
rect 6616 1917 6632 1923
rect 6680 1917 6728 1923
rect 6856 1917 6920 1923
rect 6936 1917 7032 1923
rect 7352 1917 7496 1923
rect 7832 1917 7928 1923
rect 3757 1908 3763 1912
rect 6493 1908 6499 1912
rect 56 1897 168 1903
rect 1288 1897 1320 1903
rect 1400 1897 1560 1903
rect 1688 1897 1768 1903
rect 1800 1897 2104 1903
rect 3064 1897 3091 1903
rect 269 1888 275 1892
rect 104 1877 184 1883
rect 504 1877 616 1883
rect 632 1877 664 1883
rect 680 1877 1272 1883
rect 1752 1877 2040 1883
rect 2056 1877 2088 1883
rect 2104 1877 2360 1883
rect 2440 1877 2472 1883
rect 2488 1877 2776 1883
rect 2792 1877 2840 1883
rect 2968 1877 3064 1883
rect 3085 1883 3091 1897
rect 3176 1897 3352 1903
rect 3400 1897 3432 1903
rect 3448 1897 3496 1903
rect 4168 1897 4216 1903
rect 4584 1897 4776 1903
rect 4872 1897 5432 1903
rect 5656 1897 5816 1903
rect 5848 1897 5960 1903
rect 6024 1897 6088 1903
rect 6696 1897 6707 1903
rect 6728 1897 6792 1903
rect 6920 1897 6936 1903
rect 6968 1897 7000 1903
rect 7016 1897 7064 1903
rect 7080 1897 7400 1903
rect 7528 1897 7656 1903
rect 7672 1897 7784 1903
rect 3085 1877 3480 1883
rect 3960 1877 4024 1883
rect 4712 1877 4744 1883
rect 4760 1877 4904 1883
rect 5000 1877 5192 1883
rect 5832 1877 5928 1883
rect 5960 1877 5976 1883
rect 6056 1877 6232 1883
rect 6696 1877 6808 1883
rect 6989 1877 7000 1883
rect 7048 1877 7160 1883
rect 7464 1877 7592 1883
rect 7021 1868 7027 1872
rect 136 1857 536 1863
rect 552 1857 584 1863
rect 616 1857 696 1863
rect 712 1857 1192 1863
rect 1256 1857 1480 1863
rect 1688 1857 1832 1863
rect 2904 1857 2984 1863
rect 3368 1857 4040 1863
rect 4056 1857 4232 1863
rect 4776 1857 5304 1863
rect 5320 1857 5944 1863
rect 6040 1857 6632 1863
rect 6680 1857 6776 1863
rect 7544 1857 7640 1863
rect 7656 1857 7768 1863
rect 472 1837 632 1843
rect 744 1837 792 1843
rect 1128 1837 1288 1843
rect 1400 1837 1416 1843
rect 2936 1837 3048 1843
rect 3272 1837 3416 1843
rect 3464 1837 5624 1843
rect 5912 1837 6104 1843
rect 6120 1837 6312 1843
rect 6328 1837 6616 1843
rect 376 1817 744 1823
rect 1240 1817 1352 1823
rect 1400 1817 1528 1823
rect 1720 1817 1832 1823
rect 56 1797 152 1803
rect 168 1797 536 1803
rect 792 1797 1784 1803
rect 3384 1817 3496 1823
rect 3288 1797 3368 1803
rect 3384 1797 3752 1803
rect 3768 1797 3896 1803
rect 4136 1817 4232 1823
rect 5496 1817 6024 1823
rect 4088 1797 4184 1803
rect 4237 1797 4280 1803
rect 56 1777 104 1783
rect 120 1777 184 1783
rect 200 1777 456 1783
rect 1208 1777 1400 1783
rect 1448 1777 1608 1783
rect 2024 1777 2056 1783
rect 2136 1777 2248 1783
rect 2568 1777 3336 1783
rect 3416 1777 3976 1783
rect 4237 1783 4243 1797
rect 4792 1797 4808 1803
rect 6104 1817 6280 1823
rect 6296 1817 6328 1823
rect 7272 1817 7464 1823
rect 7352 1797 7464 1803
rect 7480 1797 7752 1803
rect 3992 1777 4243 1783
rect 4264 1777 4968 1783
rect 5608 1777 6264 1783
rect 6280 1777 7240 1783
rect 584 1757 648 1763
rect 664 1757 840 1763
rect 1240 1757 1336 1763
rect 1464 1757 1512 1763
rect 1608 1757 1656 1763
rect 1944 1757 2264 1763
rect 3096 1757 3464 1763
rect 3544 1757 4424 1763
rect 4456 1757 4520 1763
rect 4680 1757 4744 1763
rect 4920 1757 5000 1763
rect 5592 1757 5640 1763
rect 5656 1757 5704 1763
rect 5768 1757 5976 1763
rect 6968 1757 7032 1763
rect 7112 1757 7224 1763
rect 7448 1757 7512 1763
rect -51 1737 8 1743
rect 392 1737 424 1743
rect 488 1737 872 1743
rect 888 1737 1032 1743
rect 1101 1737 1112 1743
rect 1336 1737 1352 1743
rect 1480 1737 1496 1743
rect 1528 1737 2136 1743
rect 2152 1737 2440 1743
rect 2456 1737 2856 1743
rect 3032 1737 3208 1743
rect 3640 1737 3656 1743
rect 3976 1737 4168 1743
rect 4200 1737 4296 1743
rect 4520 1737 4552 1743
rect 4813 1743 4819 1752
rect 4808 1737 4819 1743
rect 4920 1737 4952 1743
rect 5208 1737 5368 1743
rect 5672 1737 5688 1743
rect 5784 1737 5800 1743
rect 5992 1737 6168 1743
rect 6189 1737 6200 1743
rect 24 1717 104 1723
rect 136 1717 168 1723
rect 184 1717 216 1723
rect 264 1717 296 1723
rect 360 1717 456 1723
rect 696 1717 744 1723
rect 1432 1717 1544 1723
rect 1576 1717 1624 1723
rect 1704 1717 1715 1723
rect 1848 1717 1928 1723
rect 2088 1717 2168 1723
rect 2552 1717 2728 1723
rect 2904 1717 3032 1723
rect 3720 1717 3832 1723
rect 4072 1717 4104 1723
rect 4120 1717 4360 1723
rect 4408 1717 4488 1723
rect 4504 1717 4600 1723
rect 4808 1717 4952 1723
rect 4968 1717 5032 1723
rect 5544 1717 5560 1723
rect 5624 1717 6008 1723
rect 6189 1723 6195 1737
rect 6312 1737 6424 1743
rect 6760 1737 6808 1743
rect 7016 1737 7160 1743
rect 7256 1737 7368 1743
rect 7464 1737 7528 1743
rect 6088 1717 6195 1723
rect 6216 1717 6248 1723
rect 6264 1717 6344 1723
rect 6440 1717 6456 1723
rect 6488 1717 6520 1723
rect 6568 1717 6696 1723
rect 6712 1717 6760 1723
rect 6824 1717 7288 1723
rect 7560 1717 7768 1723
rect 7784 1717 7896 1723
rect -51 1697 200 1703
rect 216 1697 328 1703
rect 392 1697 408 1703
rect 440 1697 568 1703
rect 600 1697 616 1703
rect 728 1697 1240 1703
rect 1288 1697 1464 1703
rect 1496 1697 1656 1703
rect 1912 1697 1976 1703
rect 2360 1697 2504 1703
rect 2520 1697 2552 1703
rect 2568 1697 2632 1703
rect 2888 1697 3000 1703
rect 3624 1697 3704 1703
rect 3848 1697 3896 1703
rect 3917 1697 3992 1703
rect 184 1677 280 1683
rect 312 1677 952 1683
rect 984 1677 1032 1683
rect 1560 1677 1816 1683
rect 1832 1677 1880 1683
rect 1960 1677 3480 1683
rect 3512 1677 3800 1683
rect 3917 1683 3923 1697
rect 4104 1697 4216 1703
rect 4248 1697 4296 1703
rect 4349 1697 4360 1703
rect 4424 1697 4456 1703
rect 4488 1697 4616 1703
rect 4840 1697 5016 1703
rect 5037 1697 5048 1703
rect 5144 1697 5256 1703
rect 5976 1697 6536 1703
rect 6760 1697 6824 1703
rect 6920 1697 7032 1703
rect 7336 1697 7400 1703
rect 7512 1697 7688 1703
rect 3816 1677 3923 1683
rect 3944 1677 4120 1683
rect 4136 1677 4184 1683
rect 4872 1677 5144 1683
rect 5176 1677 5224 1683
rect 5864 1677 7080 1683
rect 7096 1677 7240 1683
rect 7528 1677 7544 1683
rect 1165 1668 1171 1672
rect 328 1657 392 1663
rect 424 1657 472 1663
rect 600 1657 1016 1663
rect 1496 1657 3416 1663
rect 3752 1657 3944 1663
rect 4008 1657 4136 1663
rect 4440 1657 5496 1663
rect 5704 1657 5720 1663
rect 5736 1657 5912 1663
rect 5928 1657 6136 1663
rect 6152 1657 6504 1663
rect 6552 1657 7336 1663
rect 7352 1657 7496 1663
rect 424 1637 536 1643
rect 648 1637 1624 1643
rect 1656 1637 1816 1643
rect 1848 1637 2376 1643
rect 4040 1637 4072 1643
rect 4168 1637 4200 1643
rect 4296 1637 4440 1643
rect 4792 1637 5240 1643
rect 6584 1637 7512 1643
rect 7528 1637 7960 1643
rect 3437 1628 3443 1632
rect 184 1597 568 1603
rect 1160 1617 1288 1623
rect 1592 1617 2184 1623
rect 1032 1597 2072 1603
rect 3672 1617 4168 1623
rect 4184 1617 4504 1623
rect 3144 1597 3320 1603
rect 3336 1597 4824 1603
rect 5560 1617 6136 1623
rect 6152 1617 6248 1623
rect 6264 1617 6296 1623
rect 5608 1597 5928 1603
rect 6520 1597 6664 1603
rect 120 1577 344 1583
rect 360 1577 680 1583
rect 1288 1577 1944 1583
rect 2120 1577 2792 1583
rect 3384 1577 3544 1583
rect 3608 1577 4088 1583
rect 4216 1577 5592 1583
rect 6808 1577 7064 1583
rect 24 1557 584 1563
rect 1144 1557 1160 1563
rect 1640 1557 1992 1563
rect 2248 1557 2312 1563
rect 2408 1557 2504 1563
rect 2680 1557 3736 1563
rect 3752 1557 3816 1563
rect 4104 1557 4200 1563
rect 4216 1557 4456 1563
rect 4888 1557 5128 1563
rect 5192 1557 5272 1563
rect 568 1537 600 1543
rect 1016 1537 1624 1543
rect 1656 1537 1736 1543
rect 1960 1537 2120 1543
rect 2152 1537 2424 1543
rect 2824 1537 2872 1543
rect 2904 1537 2936 1543
rect 3560 1537 3672 1543
rect 3688 1537 4488 1543
rect 4616 1537 4872 1543
rect 5096 1537 5320 1543
rect 5400 1537 5704 1543
rect 5720 1537 5752 1543
rect 5768 1537 5816 1543
rect 5896 1537 6280 1543
rect 6616 1537 6776 1543
rect 7720 1537 7768 1543
rect 477 1528 483 1532
rect 1789 1528 1795 1532
rect -51 1517 8 1523
rect 392 1517 440 1523
rect 1336 1517 1352 1523
rect 1480 1517 1704 1523
rect 1736 1517 1784 1523
rect 1800 1517 1848 1523
rect 1896 1517 2056 1523
rect 2104 1517 2152 1523
rect 2168 1517 2424 1523
rect 2824 1517 2888 1523
rect 2936 1517 3224 1523
rect 3640 1517 3896 1523
rect 3912 1517 3944 1523
rect 3960 1517 3976 1523
rect 3992 1517 4184 1523
rect 4296 1517 4392 1523
rect 4776 1517 4840 1523
rect 4904 1517 5208 1523
rect 5224 1517 5432 1523
rect 5848 1517 5880 1523
rect 6072 1517 6232 1523
rect 6328 1517 6360 1523
rect 6600 1517 6664 1523
rect 6776 1517 6888 1523
rect 6904 1517 6952 1523
rect 6968 1517 6984 1523
rect 7192 1517 7224 1523
rect 7256 1517 7512 1523
rect 7592 1517 7608 1523
rect 7752 1517 7864 1523
rect 461 1508 467 1512
rect 2781 1508 2787 1512
rect 4765 1508 4771 1512
rect 168 1497 216 1503
rect 232 1497 312 1503
rect 392 1497 408 1503
rect 584 1497 712 1503
rect 968 1497 1016 1503
rect 1160 1497 1336 1503
rect 1528 1497 2104 1503
rect 2296 1497 2312 1503
rect 2488 1497 2536 1503
rect 2744 1497 2760 1503
rect 2936 1497 3144 1503
rect 3592 1497 3624 1503
rect 5176 1497 5256 1503
rect 5272 1497 5352 1503
rect 5368 1497 5416 1503
rect 5576 1497 5736 1503
rect 5912 1497 6168 1503
rect 6216 1497 6248 1503
rect 6344 1497 6408 1503
rect 6504 1497 6568 1503
rect 6680 1497 6792 1503
rect 6808 1497 7048 1503
rect 7064 1497 7096 1503
rect 7480 1497 7592 1503
rect 7624 1497 7688 1503
rect 7704 1497 7992 1503
rect 8008 1497 8024 1503
rect 2733 1488 2739 1492
rect 408 1477 552 1483
rect 1432 1477 1624 1483
rect 1832 1477 1880 1483
rect 2200 1477 2344 1483
rect 2552 1477 2648 1483
rect 2744 1477 3128 1483
rect 3512 1477 3576 1483
rect 3592 1477 3832 1483
rect 3896 1477 4008 1483
rect 4424 1477 5544 1483
rect 5784 1477 5848 1483
rect 5944 1477 6216 1483
rect 6232 1477 6344 1483
rect 6637 1483 6643 1492
rect 6632 1477 6643 1483
rect 7064 1477 7080 1483
rect 7096 1477 7176 1483
rect 7261 1483 7267 1492
rect 7256 1477 7267 1483
rect 7304 1477 7384 1483
rect 7400 1477 7464 1483
rect 7560 1477 7848 1483
rect 6941 1468 6947 1472
rect 264 1457 392 1463
rect 1192 1457 1336 1463
rect 1352 1457 1672 1463
rect 1912 1457 2200 1463
rect 2296 1457 2392 1463
rect 2456 1457 3416 1463
rect 3432 1457 3448 1463
rect 3464 1457 4360 1463
rect 4712 1457 4792 1463
rect 5960 1457 6264 1463
rect 6280 1457 6344 1463
rect 6376 1457 6387 1463
rect 6424 1457 6552 1463
rect 6600 1457 6680 1463
rect 6696 1457 6872 1463
rect 6888 1457 6904 1463
rect 6984 1457 7032 1463
rect 7080 1457 7128 1463
rect 7272 1457 7384 1463
rect 7528 1457 7704 1463
rect 7720 1457 7736 1463
rect 248 1437 616 1443
rect 632 1437 680 1443
rect 696 1437 1528 1443
rect 1544 1437 1736 1443
rect 1752 1437 1800 1443
rect 1848 1437 1992 1443
rect 2136 1437 2248 1443
rect 2328 1437 3768 1443
rect 3928 1437 4168 1443
rect 4488 1437 6104 1443
rect 6120 1437 6584 1443
rect 6744 1437 7576 1443
rect 7640 1437 7704 1443
rect 1112 1417 1656 1423
rect 168 1397 536 1403
rect 1272 1397 1288 1403
rect 2024 1417 3768 1423
rect 3960 1417 3976 1423
rect 2088 1397 3320 1403
rect 3336 1397 3368 1403
rect 3384 1397 3512 1403
rect 4232 1417 4584 1423
rect 4152 1397 4216 1403
rect 4392 1397 4520 1403
rect 4536 1397 4664 1403
rect 4680 1397 4952 1403
rect 4968 1397 4984 1403
rect 6264 1417 6520 1423
rect 6584 1417 6744 1423
rect 6408 1397 7128 1403
rect 4237 1388 4243 1392
rect 280 1377 360 1383
rect 376 1377 552 1383
rect 1080 1377 1256 1383
rect 1512 1377 1560 1383
rect 1688 1377 2168 1383
rect 3336 1377 3400 1383
rect 3416 1377 3448 1383
rect 3512 1377 3656 1383
rect 3672 1377 4216 1383
rect 5880 1377 6168 1383
rect 6392 1377 6403 1383
rect 7384 1377 7656 1383
rect 56 1357 136 1363
rect 152 1357 531 1363
rect -51 1337 184 1343
rect 200 1337 248 1343
rect 525 1343 531 1357
rect 552 1357 856 1363
rect 1128 1357 1224 1363
rect 1240 1357 1576 1363
rect 1688 1357 1928 1363
rect 2280 1357 2376 1363
rect 3400 1357 3432 1363
rect 3448 1357 3496 1363
rect 3560 1357 3784 1363
rect 3864 1357 4008 1363
rect 4056 1357 4312 1363
rect 4344 1357 4376 1363
rect 4472 1357 4616 1363
rect 4776 1357 4872 1363
rect 5816 1357 6024 1363
rect 6360 1357 6488 1363
rect 6936 1357 6968 1363
rect 6984 1357 7304 1363
rect 7752 1357 7800 1363
rect 525 1337 584 1343
rect 616 1337 664 1343
rect 680 1337 872 1343
rect 984 1337 1096 1343
rect 1144 1337 1160 1343
rect 1192 1337 1656 1343
rect 1672 1337 1784 1343
rect 2248 1337 2360 1343
rect 2600 1337 2744 1343
rect 2808 1337 2856 1343
rect 2920 1337 2968 1343
rect 2984 1337 3176 1343
rect 3624 1337 3640 1343
rect 3656 1337 3736 1343
rect 3960 1337 4152 1343
rect 4184 1337 4632 1343
rect 4696 1337 4952 1343
rect 5128 1337 5224 1343
rect 5400 1337 5512 1343
rect 5528 1337 5624 1343
rect 5704 1337 5720 1343
rect 6248 1337 6296 1343
rect 6328 1337 6392 1343
rect 6536 1337 6680 1343
rect 6824 1337 6936 1343
rect 7240 1337 7464 1343
rect 7512 1337 7816 1343
rect 7880 1337 7944 1343
rect 413 1328 419 1332
rect 24 1317 104 1323
rect 184 1317 216 1323
rect 248 1317 328 1323
rect 424 1317 472 1323
rect 488 1317 536 1323
rect 600 1317 728 1323
rect 744 1317 808 1323
rect 840 1317 936 1323
rect 952 1317 1032 1323
rect 1112 1317 1192 1323
rect 1256 1317 1267 1323
rect 1288 1317 1464 1323
rect 1560 1317 1592 1323
rect 1608 1317 1720 1323
rect 1736 1317 1832 1323
rect 1848 1317 1880 1323
rect 1944 1317 2200 1323
rect 2216 1317 2280 1323
rect 2328 1317 2488 1323
rect 2744 1317 2872 1323
rect 2888 1317 2936 1323
rect 3576 1317 3672 1323
rect 3768 1317 4152 1323
rect 4440 1317 4456 1323
rect 4488 1317 4520 1323
rect 4536 1317 4776 1323
rect 4808 1317 4840 1323
rect 5000 1317 5176 1323
rect 5320 1317 5432 1323
rect 5528 1317 5539 1323
rect 5576 1317 5688 1323
rect 5704 1317 5736 1323
rect 6024 1317 6312 1323
rect 6424 1317 6520 1323
rect 6552 1317 6616 1323
rect 6872 1317 6920 1323
rect 6989 1323 6995 1332
rect 6984 1317 6995 1323
rect 7032 1317 7576 1323
rect 7608 1317 7688 1323
rect 7768 1317 7832 1323
rect 7864 1317 7960 1323
rect 2701 1308 2707 1312
rect 4797 1308 4803 1312
rect 5885 1308 5891 1312
rect -51 1297 8 1303
rect 184 1297 296 1303
rect 344 1297 456 1303
rect 520 1297 531 1303
rect 552 1297 648 1303
rect 664 1297 712 1303
rect 840 1297 888 1303
rect 1032 1297 1128 1303
rect 1336 1297 1576 1303
rect 1624 1297 1864 1303
rect 1928 1297 2264 1303
rect 2344 1297 2504 1303
rect 2520 1297 2568 1303
rect 2904 1297 3080 1303
rect 3576 1297 3608 1303
rect 3928 1297 3960 1303
rect 4008 1297 4056 1303
rect 4312 1297 4600 1303
rect 4616 1297 4760 1303
rect 4840 1297 4968 1303
rect 5240 1297 5400 1303
rect 5432 1297 5480 1303
rect 5997 1303 6003 1312
rect 6797 1308 6803 1312
rect 5992 1297 6003 1303
rect 7528 1297 7608 1303
rect 7704 1297 7768 1303
rect 6893 1288 6899 1292
rect 248 1277 280 1283
rect 328 1277 360 1283
rect 504 1277 760 1283
rect 776 1277 792 1283
rect 904 1277 1064 1283
rect 1288 1277 1640 1283
rect 1960 1277 2040 1283
rect 2584 1277 2664 1283
rect 3496 1277 3592 1283
rect 3608 1277 3704 1283
rect 3736 1277 3832 1283
rect 3848 1277 4184 1283
rect 4200 1277 4280 1283
rect 4648 1277 4824 1283
rect 5480 1277 5528 1283
rect 6216 1277 6808 1283
rect 7240 1277 7880 1283
rect 232 1257 616 1263
rect 648 1257 840 1263
rect 1480 1257 1816 1263
rect 1848 1257 1928 1263
rect 2504 1257 2616 1263
rect 3704 1257 3720 1263
rect 3741 1257 3896 1263
rect 376 1237 456 1243
rect 488 1237 1160 1243
rect 1176 1237 1352 1243
rect 1368 1237 1784 1243
rect 1800 1237 1928 1243
rect 3741 1243 3747 1257
rect 4088 1257 4168 1263
rect 4472 1257 4520 1263
rect 4552 1257 4632 1263
rect 5912 1257 6536 1263
rect 7496 1257 7576 1263
rect 2024 1237 3747 1243
rect 4312 1237 4344 1243
rect 4616 1237 4664 1243
rect 6680 1237 7848 1243
rect 3885 1228 3891 1232
rect 456 1217 504 1223
rect 760 1217 872 1223
rect 184 1197 536 1203
rect 568 1197 728 1203
rect 1320 1217 1528 1223
rect 1544 1217 1928 1223
rect 1944 1217 2088 1223
rect 1432 1197 1512 1203
rect 1528 1197 1672 1203
rect 1752 1197 1848 1203
rect 2056 1197 2696 1203
rect 3016 1197 4104 1203
rect 6120 1217 6776 1223
rect 6296 1197 6904 1203
rect 7352 1217 7512 1223
rect 136 1177 1048 1183
rect 1192 1177 1384 1183
rect 1400 1177 1464 1183
rect 1544 1177 1720 1183
rect 1800 1177 2152 1183
rect 2712 1177 4248 1183
rect 4408 1177 4616 1183
rect 5304 1177 5480 1183
rect 5496 1177 5528 1183
rect 6840 1177 6872 1183
rect 7064 1177 7272 1183
rect 7688 1177 7864 1183
rect 56 1157 72 1163
rect 104 1157 152 1163
rect 312 1157 472 1163
rect 584 1157 776 1163
rect 1064 1157 1560 1163
rect 1576 1157 2344 1163
rect 2360 1157 2600 1163
rect 2616 1157 2712 1163
rect 3688 1157 3752 1163
rect 3784 1157 4248 1163
rect 4376 1157 4504 1163
rect 4520 1157 4728 1163
rect 5896 1157 7080 1163
rect 7096 1157 7224 1163
rect 7256 1157 7352 1163
rect 7368 1157 7416 1163
rect 7432 1157 7480 1163
rect 7752 1157 7784 1163
rect 40 1137 200 1143
rect 248 1137 264 1143
rect 312 1137 424 1143
rect 504 1137 536 1143
rect 696 1137 984 1143
rect 1096 1137 1176 1143
rect 1256 1137 1496 1143
rect 1512 1137 2232 1143
rect 2632 1137 2808 1143
rect 3064 1137 3400 1143
rect 3448 1137 3560 1143
rect 3720 1137 3960 1143
rect 4456 1137 4568 1143
rect 4648 1137 4760 1143
rect 5640 1137 6152 1143
rect 6904 1137 7096 1143
rect 7320 1137 7448 1143
rect 7656 1137 7768 1143
rect 7800 1137 7896 1143
rect 3981 1128 3987 1132
rect -51 1117 120 1123
rect 136 1117 200 1123
rect 264 1117 360 1123
rect 520 1117 584 1123
rect 632 1117 664 1123
rect 856 1117 1576 1123
rect 2280 1117 2392 1123
rect 2408 1117 2456 1123
rect 2472 1117 2664 1123
rect 2744 1117 2760 1123
rect 2824 1117 2840 1123
rect 2888 1117 3144 1123
rect 3176 1117 3192 1123
rect 3208 1117 3336 1123
rect 3485 1117 3592 1123
rect 797 1108 803 1112
rect 56 1097 104 1103
rect 232 1097 408 1103
rect 440 1097 520 1103
rect 552 1097 776 1103
rect 824 1097 904 1103
rect 1160 1097 1171 1103
rect 1208 1097 1288 1103
rect 1592 1097 1624 1103
rect 1640 1097 1768 1103
rect 1821 1103 1827 1112
rect 1816 1097 1827 1103
rect 1912 1097 2296 1103
rect 2328 1097 2360 1103
rect 2744 1097 2792 1103
rect 3485 1103 3491 1117
rect 3608 1117 3688 1123
rect 3848 1117 3864 1123
rect 3896 1117 3944 1123
rect 4104 1117 4216 1123
rect 4328 1117 4536 1123
rect 4920 1117 4952 1123
rect 4984 1117 5096 1123
rect 5160 1117 5192 1123
rect 5208 1117 5400 1123
rect 6536 1117 6616 1123
rect 6968 1117 7016 1123
rect 7160 1117 7880 1123
rect 6013 1108 6019 1112
rect 2856 1097 3491 1103
rect 3512 1097 3544 1103
rect 3592 1097 3832 1103
rect 3880 1097 4056 1103
rect 4280 1097 4312 1103
rect 4584 1097 4616 1103
rect 4808 1097 4872 1103
rect 5128 1097 5208 1103
rect 5528 1097 5656 1103
rect 5832 1097 5864 1103
rect 6248 1097 6360 1103
rect 6376 1097 6408 1103
rect 6584 1097 6728 1103
rect 7000 1097 7827 1103
rect 200 1077 232 1083
rect 296 1077 488 1083
rect 504 1077 584 1083
rect 632 1077 664 1083
rect 696 1077 760 1083
rect 984 1077 1032 1083
rect 1224 1077 1256 1083
rect 1464 1077 1683 1083
rect 104 1057 168 1063
rect 408 1057 664 1063
rect 680 1057 712 1063
rect 744 1057 824 1063
rect 1480 1057 1512 1063
rect 1677 1063 1683 1077
rect 1704 1077 1800 1083
rect 1816 1077 1848 1083
rect 2376 1077 2424 1083
rect 2792 1077 2872 1083
rect 2888 1077 3160 1083
rect 3176 1077 3240 1083
rect 3384 1077 3416 1083
rect 3432 1077 3656 1083
rect 3784 1077 3816 1083
rect 3832 1077 4024 1083
rect 4104 1077 4296 1083
rect 4616 1077 4792 1083
rect 4856 1077 4984 1083
rect 5192 1077 5320 1083
rect 5464 1077 5576 1083
rect 5752 1077 5880 1083
rect 6104 1077 6152 1083
rect 6280 1077 6328 1083
rect 6664 1077 6744 1083
rect 6760 1077 6792 1083
rect 6936 1077 6984 1083
rect 7128 1077 7144 1083
rect 7224 1077 7288 1083
rect 7304 1077 7384 1083
rect 7560 1077 7704 1083
rect 7821 1083 7827 1097
rect 7848 1097 7912 1103
rect 7928 1097 7992 1103
rect 7821 1077 8024 1083
rect 1677 1057 1720 1063
rect 2152 1057 2296 1063
rect 2840 1057 2888 1063
rect 3320 1057 3352 1063
rect 3368 1057 3464 1063
rect 3800 1057 3880 1063
rect 3992 1057 4184 1063
rect 4200 1057 4344 1063
rect 4408 1057 4440 1063
rect 4568 1057 4856 1063
rect 4872 1057 4968 1063
rect 5224 1057 5304 1063
rect 5320 1057 5640 1063
rect 5960 1057 5976 1063
rect 6040 1057 6168 1063
rect 6456 1057 6584 1063
rect 6760 1057 6872 1063
rect 6904 1057 6936 1063
rect 7928 1057 7992 1063
rect 3757 1048 3763 1052
rect 6189 1048 6195 1052
rect 392 1037 424 1043
rect 1181 1037 1192 1043
rect 3288 1037 3512 1043
rect 4344 1037 4504 1043
rect 5496 1037 5784 1043
rect 6029 1037 6088 1043
rect 488 1017 1448 1023
rect 920 997 1672 1003
rect 2312 1017 2536 1023
rect 2552 1017 2968 1023
rect 2248 997 2440 1003
rect 3496 997 3512 1003
rect 3816 997 3960 1003
rect 6029 1023 6035 1037
rect 6408 1037 6632 1043
rect 6824 1037 6936 1043
rect 7848 1037 7864 1043
rect 7880 1037 7944 1043
rect 4296 1017 6035 1023
rect 5624 997 5832 1003
rect 6184 1017 6232 1023
rect 6552 1017 7480 1023
rect 6168 997 6392 1003
rect 6520 997 7112 1003
rect 7352 997 7544 1003
rect 7560 997 7608 1003
rect 1165 977 1176 983
rect 2184 977 2360 983
rect 2392 977 3576 983
rect 3720 977 3832 983
rect 4264 977 4344 983
rect 4440 977 4760 983
rect 4776 977 4952 983
rect 6008 977 6184 983
rect 6232 977 6488 983
rect 6520 977 6536 983
rect 6872 977 6883 983
rect 5629 968 5635 972
rect 72 957 264 963
rect 424 957 1144 963
rect 1240 957 1256 963
rect 1352 957 1400 963
rect 1896 957 2408 963
rect 3176 957 3384 963
rect 3400 957 3528 963
rect 3672 957 3992 963
rect 4088 957 4120 963
rect 4280 957 4408 963
rect 4440 957 4664 963
rect 4845 957 5240 963
rect 168 937 312 943
rect 408 937 536 943
rect 1208 937 1272 943
rect 1304 937 1320 943
rect 1336 937 1352 943
rect 1368 937 1784 943
rect 2408 937 2520 943
rect 2552 937 2664 943
rect 3176 937 3416 943
rect 3432 937 3464 943
rect 3560 937 3640 943
rect 3656 937 3736 943
rect 3800 937 3880 943
rect 4136 937 4168 943
rect 4845 943 4851 957
rect 5352 957 5480 963
rect 6056 957 6104 963
rect 6232 957 6248 963
rect 6280 957 6520 963
rect 6664 957 6728 963
rect 6776 957 6888 963
rect 7624 957 8008 963
rect 4184 937 4851 943
rect 4872 937 5176 943
rect 5288 937 5352 943
rect 5368 937 5432 943
rect 5944 937 6088 943
rect 6104 937 6264 943
rect 6424 937 6648 943
rect 6712 937 6824 943
rect 6888 937 7064 943
rect 7736 937 7832 943
rect 3485 928 3491 932
rect 5837 928 5843 932
rect 7517 928 7523 932
rect 136 917 232 923
rect 296 917 312 923
rect 328 917 376 923
rect 440 917 488 923
rect 504 917 552 923
rect 888 917 984 923
rect 1000 917 1064 923
rect 1256 917 1432 923
rect 1704 917 1816 923
rect 2200 917 2280 923
rect 2360 917 2456 923
rect 3080 917 3432 923
rect 3608 917 3640 923
rect 3784 917 3816 923
rect 3960 917 4120 923
rect 4168 917 4264 923
rect 4312 917 4344 923
rect 4360 917 4392 923
rect 4424 917 4456 923
rect 4520 917 4712 923
rect 4744 917 4920 923
rect 5160 917 5272 923
rect 6024 917 6472 923
rect 6504 917 6536 923
rect 6568 917 6600 923
rect 6792 917 6803 923
rect 6856 917 6904 923
rect 6920 917 6952 923
rect 7048 917 7272 923
rect 7864 917 7896 923
rect 232 897 408 903
rect 1000 897 1208 903
rect 1320 897 1416 903
rect 1512 897 2008 903
rect 2456 897 2696 903
rect 3624 897 3656 903
rect 3688 897 3800 903
rect 4104 897 4344 903
rect 4968 897 5128 903
rect 5256 897 5336 903
rect 5992 897 6136 903
rect 6152 897 6312 903
rect 6328 897 6568 903
rect 6616 897 6627 903
rect 6952 897 7000 903
rect 7112 897 7176 903
rect 7192 897 7240 903
rect 264 877 312 883
rect 1080 877 1336 883
rect 1576 877 2328 883
rect 2344 877 2376 883
rect 2392 877 2776 883
rect 2792 877 3288 883
rect 3528 877 3752 883
rect 3976 877 4120 883
rect 4168 877 4296 883
rect 4312 877 4376 883
rect 4808 877 4904 883
rect 5784 877 6504 883
rect 6728 877 6760 883
rect 6776 877 7704 883
rect 3496 857 3528 863
rect 3544 857 3688 863
rect 4136 857 4184 863
rect 4216 857 4392 863
rect 4424 857 4520 863
rect 4536 857 5912 863
rect 6136 857 6152 863
rect 6312 857 6856 863
rect 7224 857 7640 863
rect 2584 837 2632 843
rect 2648 837 5688 843
rect 6040 837 6168 843
rect 6344 837 6680 843
rect 6696 837 6760 843
rect 7000 837 7768 843
rect 392 817 696 823
rect 1160 817 1384 823
rect 1400 817 2088 823
rect 2440 817 2584 823
rect 4040 817 4168 823
rect 4200 817 4360 823
rect 4376 817 4632 823
rect 4104 797 4264 803
rect 4296 797 4344 803
rect 6680 797 6904 803
rect 7160 817 7512 823
rect 440 777 1240 783
rect 3784 777 4312 783
rect 5832 777 6152 783
rect 6168 777 6696 783
rect 6712 777 7320 783
rect 936 757 1000 763
rect 3512 757 3656 763
rect 4072 757 4120 763
rect 4184 757 6264 763
rect 6600 757 6760 763
rect 984 737 1048 743
rect 1080 737 1160 743
rect 1336 737 1608 743
rect 3096 737 3352 743
rect 3640 737 3832 743
rect 3928 737 4136 743
rect 4184 737 4456 743
rect 4936 737 5480 743
rect 5496 737 5528 743
rect 5544 737 5592 743
rect 6008 737 6216 743
rect 6248 737 6392 743
rect 7208 737 7336 743
rect 7480 737 7848 743
rect 344 717 392 723
rect 424 717 600 723
rect 1080 717 1256 723
rect 1384 717 1400 723
rect 1784 717 1864 723
rect 2008 717 2200 723
rect 3160 717 3256 723
rect 3560 717 3592 723
rect 3656 717 3688 723
rect 3944 717 4040 723
rect 4056 717 4104 723
rect 4136 717 4216 723
rect 4312 717 4392 723
rect 4472 717 4536 723
rect 4552 717 4760 723
rect 4952 717 5000 723
rect 5192 717 5416 723
rect 5464 717 5576 723
rect 5864 717 6760 723
rect 6776 717 7016 723
rect 7176 717 7240 723
rect 7496 717 7672 723
rect 7688 717 7832 723
rect 1069 708 1075 712
rect 264 697 312 703
rect 328 697 392 703
rect 408 697 424 703
rect 440 697 504 703
rect 1016 697 1032 703
rect 1144 697 1192 703
rect 1208 697 1443 703
rect 104 677 248 683
rect 728 677 760 683
rect 776 677 808 683
rect 824 677 888 683
rect 968 677 1016 683
rect 1032 677 1080 683
rect 1437 683 1443 697
rect 1496 697 1560 703
rect 1864 697 1992 703
rect 2136 697 2216 703
rect 2376 697 2632 703
rect 2904 697 2936 703
rect 2952 697 3000 703
rect 3032 697 3096 703
rect 3128 697 3160 703
rect 3592 697 3704 703
rect 3725 697 3736 703
rect 3752 697 3784 703
rect 3928 697 3960 703
rect 4008 697 4216 703
rect 4632 697 5368 703
rect 5432 697 5784 703
rect 5880 697 6072 703
rect 6152 697 6232 703
rect 6280 697 6312 703
rect 6328 697 6360 703
rect 6488 697 6824 703
rect 7048 697 7112 703
rect 7128 697 7208 703
rect 7224 697 7256 703
rect 7672 697 7688 703
rect 7752 697 7784 703
rect 7800 697 7976 703
rect 1437 677 1592 683
rect 1608 677 1832 683
rect 1928 677 2184 683
rect 2536 677 2600 683
rect 2616 677 2792 683
rect 2888 677 2920 683
rect 2936 677 3032 683
rect 3048 677 3448 683
rect 3464 677 3496 683
rect 3608 677 3768 683
rect 3880 677 4008 683
rect 4152 677 4200 683
rect 4392 677 4808 683
rect 4984 677 5176 683
rect 5320 677 5448 683
rect 5528 677 5656 683
rect 5752 677 5816 683
rect 5944 677 6280 683
rect 6360 677 6488 683
rect 6632 677 6728 683
rect 6808 677 7160 683
rect 7240 677 7480 683
rect 7496 677 7624 683
rect 7784 677 8008 683
rect 376 657 824 663
rect 1048 657 1304 663
rect 1816 657 2152 663
rect 2168 657 2328 663
rect 2600 657 3000 663
rect 3016 657 3128 663
rect 3693 657 3704 663
rect 3736 657 3880 663
rect 3912 657 4232 663
rect 4840 657 5288 663
rect 6392 657 6648 663
rect 6664 657 7016 663
rect 7928 657 7976 663
rect 808 637 920 643
rect 1176 637 1240 643
rect 1272 637 1768 643
rect 2504 637 2680 643
rect 2920 637 3160 643
rect 3528 637 4152 643
rect 4360 637 4648 643
rect 4680 637 4776 643
rect 5032 637 5384 643
rect 5400 637 5784 643
rect 5896 637 6184 643
rect 6200 637 6584 643
rect 6904 637 6915 643
rect 664 617 744 623
rect 760 617 840 623
rect 856 617 1064 623
rect 1080 617 1448 623
rect 1224 597 1736 603
rect 1816 597 1864 603
rect 2008 617 2488 623
rect 3064 617 3080 623
rect 2760 597 2808 603
rect 2904 597 3368 603
rect 4088 617 6024 623
rect 4344 597 4424 603
rect 4440 597 4712 603
rect 4728 597 4840 603
rect 4856 597 4888 603
rect 4920 597 5640 603
rect 6296 617 6808 623
rect 6232 597 6296 603
rect 6616 597 6632 603
rect 6696 597 7064 603
rect 216 577 360 583
rect 376 577 472 583
rect 1112 577 1448 583
rect 1645 577 1656 583
rect 1896 577 1944 583
rect 2648 577 3192 583
rect 3688 577 3811 583
rect 568 557 600 563
rect 616 557 664 563
rect 1384 557 1400 563
rect 1432 557 1928 563
rect 2792 557 3016 563
rect 3053 557 3064 563
rect 3720 557 3752 563
rect 3768 557 3784 563
rect 3805 563 3811 577
rect 3848 577 4104 583
rect 4280 577 4744 583
rect 4776 577 4840 583
rect 4856 577 5096 583
rect 5656 577 5880 583
rect 7784 577 7800 583
rect 3805 557 4040 563
rect 4200 557 4280 563
rect 4296 557 4408 563
rect 4840 557 4920 563
rect 4936 557 5224 563
rect 5240 557 5320 563
rect 5336 557 5432 563
rect 5464 557 5560 563
rect 5576 557 5672 563
rect 5704 557 6904 563
rect 7560 557 7848 563
rect 3037 548 3043 552
rect 104 537 328 543
rect 360 537 440 543
rect 472 537 504 543
rect 584 537 1480 543
rect 1688 537 1816 543
rect 2072 537 2120 543
rect 2280 537 2728 543
rect 3240 537 3299 543
rect 296 517 408 523
rect 424 517 488 523
rect 600 517 680 523
rect 744 517 792 523
rect 872 517 1032 523
rect 1352 517 1400 523
rect 1432 517 1448 523
rect 1912 517 2104 523
rect 2152 517 2163 523
rect 2157 508 2163 517
rect 2312 517 2376 523
rect 2568 517 2600 523
rect 2632 517 2760 523
rect 3224 517 3272 523
rect 3293 523 3299 537
rect 3512 537 3576 543
rect 4360 537 4488 543
rect 4616 537 4728 543
rect 4984 537 5144 543
rect 5368 537 5528 543
rect 5560 537 5864 543
rect 6328 537 6376 543
rect 6520 537 6712 543
rect 7032 537 7208 543
rect 7384 537 7448 543
rect 3293 517 3304 523
rect 3672 517 3752 523
rect 3768 517 4312 523
rect 4328 517 4360 523
rect 4904 517 5352 523
rect 5624 517 5688 523
rect 5752 517 5816 523
rect 5992 517 6168 523
rect 6296 517 6456 523
rect 7000 517 7032 523
rect 7816 517 7880 523
rect 376 497 552 503
rect 712 497 1160 503
rect 1517 497 1688 503
rect 264 477 312 483
rect 328 477 632 483
rect 1517 483 1523 497
rect 1864 497 1912 503
rect 2632 497 2904 503
rect 2920 497 3464 503
rect 3752 497 3880 503
rect 3912 497 4040 503
rect 4264 497 4280 503
rect 4808 497 5128 503
rect 5144 497 5176 503
rect 5192 497 5256 503
rect 5272 497 5304 503
rect 5352 497 5368 503
rect 5400 497 5512 503
rect 5672 497 5736 503
rect 6216 497 6264 503
rect 6360 497 6744 503
rect 7016 497 7368 503
rect 1789 488 1795 492
rect 1160 477 1523 483
rect 2205 477 2216 483
rect 3160 477 3224 483
rect 3256 477 4104 483
rect 4136 477 4216 483
rect 4408 477 5080 483
rect 5096 477 5224 483
rect 7032 477 7336 483
rect 7352 477 7544 483
rect 328 457 424 463
rect 456 457 488 463
rect 520 457 696 463
rect 1533 463 1539 472
rect 1528 457 1539 463
rect 1560 457 2040 463
rect 3256 457 3864 463
rect 3880 457 3976 463
rect 4344 457 4936 463
rect 6200 457 6344 463
rect 6568 457 6904 463
rect 40 437 344 443
rect 472 437 1240 443
rect 1272 437 1288 443
rect 1736 437 2136 443
rect 3400 437 3560 443
rect 3688 437 3864 443
rect 4216 437 5528 443
rect 6872 437 7432 443
rect 120 417 536 423
rect 792 417 840 423
rect 184 397 808 403
rect 840 397 888 403
rect 1464 417 1880 423
rect 2040 417 2504 423
rect 1448 397 2360 403
rect 3720 417 4616 423
rect 3560 397 3640 403
rect 4024 397 4568 403
rect 5512 417 5560 423
rect 264 377 344 383
rect 504 377 600 383
rect 632 377 1048 383
rect 1176 377 1571 383
rect 200 357 232 363
rect 312 357 328 363
rect 520 357 680 363
rect 1064 357 1544 363
rect 1565 363 1571 377
rect 1592 377 3096 383
rect 3112 377 3608 383
rect 3656 377 5464 383
rect 5480 377 7656 383
rect 1565 357 2424 363
rect 3128 357 3384 363
rect 3448 357 4248 363
rect 4264 357 4376 363
rect 4392 357 4568 363
rect 5928 357 6584 363
rect 6600 357 6632 363
rect 6648 357 6728 363
rect 29 348 35 352
rect 429 348 435 352
rect 56 337 152 343
rect 248 337 264 343
rect 312 337 424 343
rect 456 337 472 343
rect 552 337 968 343
rect 984 337 1032 343
rect 1080 337 1096 343
rect 1112 337 1304 343
rect 1336 337 1416 343
rect 1688 337 1864 343
rect 1880 337 1928 343
rect 1944 337 2120 343
rect 2136 337 2232 343
rect 2648 337 2776 343
rect 3096 337 3304 343
rect 4696 337 4856 343
rect 5128 337 5240 343
rect 6408 337 6728 343
rect 6744 337 6840 343
rect 6904 337 6984 343
rect 7000 337 7576 343
rect -51 303 -45 323
rect 56 317 104 323
rect 120 317 360 323
rect 376 317 552 323
rect 568 317 616 323
rect 1048 317 1176 323
rect 1192 317 1224 323
rect 1240 317 1384 323
rect 1400 317 1496 323
rect 2008 317 2056 323
rect 2568 317 2696 323
rect 2712 317 2744 323
rect 2760 317 2968 323
rect 2984 317 3160 323
rect 3288 317 3336 323
rect 3368 317 3880 323
rect 3896 317 3992 323
rect 4568 317 4616 323
rect 4824 317 4888 323
rect 4904 317 4936 323
rect 5176 317 5224 323
rect 5240 317 5288 323
rect 5304 317 5656 323
rect 5896 317 6392 323
rect 6536 317 6648 323
rect 6696 317 7016 323
rect 7144 317 7656 323
rect 7672 317 7704 323
rect 7800 317 7880 323
rect 4397 308 4403 312
rect -51 297 120 303
rect 136 297 200 303
rect 232 297 280 303
rect 344 297 360 303
rect 424 297 600 303
rect 696 297 712 303
rect 1016 297 1048 303
rect 1064 297 1352 303
rect 1368 297 1432 303
rect 1512 297 1560 303
rect 1736 297 1880 303
rect 2008 297 2024 303
rect 2104 297 2280 303
rect 2744 297 2840 303
rect 3208 297 3272 303
rect 3469 297 3480 303
rect 3896 297 3960 303
rect 4280 297 4328 303
rect 4776 297 4904 303
rect 5208 297 5320 303
rect 5416 297 5480 303
rect 5512 297 5720 303
rect 5752 297 6488 303
rect 6504 297 6616 303
rect 6968 297 7032 303
rect 7064 297 7128 303
rect 7160 297 7272 303
rect 7480 297 7512 303
rect 7560 297 7592 303
rect 7784 297 7864 303
rect 120 277 168 283
rect 344 277 664 283
rect 968 277 1512 283
rect 1656 277 1816 283
rect 2520 277 2728 283
rect 2776 277 3000 283
rect 3192 277 3320 283
rect 3336 277 3400 283
rect 3496 277 3640 283
rect 3704 277 3848 283
rect 4392 277 4472 283
rect 4600 277 5400 283
rect 5448 277 5464 283
rect 5480 277 5608 283
rect 6616 277 6696 283
rect 6952 277 7160 283
rect 7624 277 7720 283
rect 776 257 872 263
rect 888 257 1064 263
rect 1560 257 1848 263
rect 2072 257 2104 263
rect 2120 257 2616 263
rect 3032 257 3048 263
rect 4536 257 4744 263
rect 4824 257 4920 263
rect 5016 257 5208 263
rect 5224 257 5480 263
rect 5528 257 5944 263
rect 6040 257 6312 263
rect 6792 257 7224 263
rect 7432 257 7624 263
rect 7640 257 7752 263
rect 936 237 968 243
rect 1480 237 1736 243
rect 1944 237 2216 243
rect 2696 237 2840 243
rect 4632 237 4840 243
rect 6024 237 6104 243
rect 7576 237 7640 243
rect 7688 237 7864 243
rect 680 217 1576 223
rect 152 197 504 203
rect 1400 197 1928 203
rect 2040 217 2648 223
rect 2680 217 3496 223
rect 2344 197 2504 203
rect 4984 217 5880 223
rect 5896 217 5992 223
rect 4216 197 4392 203
rect 4552 197 4728 203
rect 5736 197 6008 203
rect 6120 217 6456 223
rect 6472 217 6616 223
rect 6632 217 6968 223
rect 6216 197 6360 203
rect 6392 197 6616 203
rect 1128 177 2792 183
rect 2808 177 3464 183
rect 3512 177 3528 183
rect 3992 177 4504 183
rect 5848 177 6184 183
rect 6200 177 6216 183
rect 6232 177 6440 183
rect 6968 177 7320 183
rect 7528 177 7544 183
rect 72 157 248 163
rect 392 157 600 163
rect 872 157 1000 163
rect 1016 157 1320 163
rect 1352 157 1592 163
rect 1784 157 1896 163
rect 1912 157 2184 163
rect 2200 157 2328 163
rect 2376 157 2600 163
rect 2872 157 3736 163
rect 3960 157 4168 163
rect 4200 157 4264 163
rect 4376 157 4472 163
rect 4488 157 4616 163
rect 5400 157 5528 163
rect 5640 157 5736 163
rect 5976 157 5992 163
rect 6008 157 6072 163
rect 6328 157 6504 163
rect 6632 157 6760 163
rect 6840 157 6888 163
rect 6904 157 6968 163
rect 7240 157 7464 163
rect 232 137 280 143
rect 296 137 312 143
rect 328 137 440 143
rect 488 137 888 143
rect 904 137 1080 143
rect 1272 137 1496 143
rect 1720 137 1992 143
rect 2344 137 2472 143
rect 2605 137 2632 143
rect 168 117 248 123
rect 440 117 536 123
rect 728 117 744 123
rect 968 117 1032 123
rect 1624 117 1672 123
rect 2248 117 2280 123
rect 2605 123 2611 137
rect 2920 137 3112 143
rect 3512 137 3576 143
rect 3592 137 3720 143
rect 4136 137 4216 143
rect 5080 137 5176 143
rect 5480 137 5560 143
rect 5672 137 5704 143
rect 5976 137 6040 143
rect 6344 137 6408 143
rect 6584 137 6712 143
rect 6936 137 7096 143
rect 7192 137 7288 143
rect 7736 137 7832 143
rect 2552 117 2611 123
rect 2632 117 2680 123
rect 2984 117 3048 123
rect 3080 117 3320 123
rect 3576 117 3608 123
rect 3752 117 4968 123
rect 5224 117 5272 123
rect 5512 117 5592 123
rect 5704 117 5832 123
rect 5976 117 6328 123
rect 6344 117 6376 123
rect 6536 117 6584 123
rect 6600 117 6856 123
rect 6872 117 6936 123
rect 7272 117 7304 123
rect 1528 97 1624 103
rect 2168 97 2248 103
rect 2488 97 2712 103
rect 2728 97 2936 103
rect 3048 97 3144 103
rect 3336 97 3464 103
rect 4312 97 4552 103
rect 5608 97 5960 103
rect 6040 97 6200 103
rect 7304 97 7416 103
rect 3464 17 3480 23
<< m4contact >>
rect 926 5602 954 5618
rect 2264 5612 2280 5628
rect 2958 5602 2986 5618
rect 3176 5612 3192 5628
rect 5022 5602 5050 5618
rect 7054 5602 7082 5618
rect 72 5492 88 5508
rect 2808 5492 2824 5508
rect 4216 5492 4232 5508
rect 2072 5472 2088 5488
rect 3176 5472 3192 5488
rect 7688 5472 7704 5488
rect 1080 5452 1096 5468
rect 7800 5452 7816 5468
rect 7720 5432 7736 5448
rect 1950 5402 1978 5418
rect 328 5372 344 5388
rect 3688 5392 3704 5408
rect 3998 5402 4026 5418
rect 6046 5402 6074 5418
rect 520 5352 536 5368
rect 1096 5352 1112 5368
rect 1576 5332 1592 5348
rect 1784 5332 1800 5348
rect 2264 5332 2280 5348
rect 7784 5312 7800 5328
rect 4408 5292 4424 5308
rect 6616 5292 6632 5308
rect 6024 5272 6040 5288
rect 7768 5272 7784 5288
rect 72 5252 88 5268
rect 1272 5252 1288 5268
rect 3480 5252 3496 5268
rect 6920 5252 6936 5268
rect 72 5232 88 5248
rect 3848 5232 3864 5248
rect 926 5202 954 5218
rect 2616 5212 2632 5228
rect 2958 5202 2986 5218
rect 5022 5202 5050 5218
rect 7054 5202 7082 5218
rect 7704 5172 7720 5188
rect 1416 5152 1432 5168
rect 4056 5152 4072 5168
rect 2264 5112 2280 5128
rect 2856 5112 2872 5128
rect 5656 5132 5672 5148
rect 3640 5112 3656 5128
rect 3848 5112 3864 5128
rect 4872 5112 4888 5128
rect 5976 5112 5992 5128
rect 7800 5112 7816 5128
rect 1016 5072 1032 5088
rect 2904 5072 2920 5088
rect 3752 5072 3768 5088
rect 7832 5072 7848 5088
rect 4888 5052 4904 5068
rect 5656 5052 5672 5068
rect 6488 5052 6504 5068
rect 7912 5052 7928 5068
rect 1950 5002 1978 5018
rect 3998 5002 4026 5018
rect 7928 5032 7944 5048
rect 6046 5002 6074 5018
rect 7816 4992 7832 5008
rect 1256 4972 1272 4988
rect 328 4952 344 4968
rect 472 4912 488 4928
rect 728 4912 744 4928
rect 6440 4932 6456 4948
rect 6680 4932 6696 4948
rect 7864 4932 7880 4948
rect 7896 4932 7912 4948
rect 3160 4912 3176 4928
rect 4088 4912 4104 4928
rect 4568 4912 4584 4928
rect 6344 4912 6360 4928
rect 6776 4912 6792 4928
rect 7848 4912 7864 4928
rect 328 4892 344 4908
rect 1080 4892 1096 4908
rect 2360 4892 2376 4908
rect 3720 4892 3736 4908
rect 4344 4892 4360 4908
rect 5944 4892 5960 4908
rect 6312 4892 6328 4908
rect 6392 4892 6408 4908
rect 1528 4872 1544 4888
rect 6024 4872 6040 4888
rect 6392 4852 6408 4868
rect 1368 4832 1384 4848
rect 2776 4832 2792 4848
rect 3656 4832 3672 4848
rect 3896 4832 3912 4848
rect 3928 4832 3944 4848
rect 632 4812 648 4828
rect 926 4802 954 4818
rect 2936 4812 2952 4828
rect 968 4792 984 4808
rect 2920 4792 2936 4808
rect 2958 4802 2986 4818
rect 3688 4792 3704 4808
rect 5022 4802 5050 4818
rect 6424 4792 6440 4808
rect 7054 4802 7082 4818
rect 7800 4812 7816 4828
rect 968 4752 984 4768
rect 2360 4752 2376 4768
rect 3384 4752 3400 4768
rect 3896 4752 3912 4768
rect 4408 4752 4424 4768
rect 888 4732 904 4748
rect 968 4732 984 4748
rect 1432 4732 1448 4748
rect 3176 4732 3192 4748
rect 3528 4732 3544 4748
rect 3896 4732 3912 4748
rect 3912 4732 3928 4748
rect 5080 4732 5096 4748
rect 5528 4732 5544 4748
rect 5688 4732 5704 4748
rect 6216 4732 6232 4748
rect 6632 4732 6648 4748
rect 952 4712 968 4728
rect 1320 4712 1336 4728
rect 3944 4712 3960 4728
rect 40 4692 56 4708
rect 424 4692 440 4708
rect 856 4692 872 4708
rect 1032 4692 1048 4708
rect 1512 4692 1528 4708
rect 2264 4692 2280 4708
rect 2840 4692 2856 4708
rect 4184 4692 4200 4708
rect 4280 4712 4312 4728
rect 4328 4712 4344 4728
rect 4408 4712 4424 4728
rect 4936 4712 4952 4728
rect 5416 4712 5432 4728
rect 5448 4712 5464 4728
rect 6952 4712 6968 4728
rect 7016 4712 7032 4728
rect 7384 4712 7400 4728
rect 4440 4692 4456 4708
rect 5112 4692 5128 4708
rect 7416 4692 7432 4708
rect 7704 4692 7720 4708
rect 1432 4672 1448 4688
rect 2808 4672 2824 4688
rect 3448 4672 3464 4688
rect 3480 4672 3496 4688
rect 3784 4672 3800 4688
rect 4280 4672 4296 4688
rect 4312 4672 4328 4688
rect 4968 4672 4984 4688
rect 6536 4672 6552 4688
rect 6584 4672 6600 4688
rect 6664 4672 6680 4688
rect 7128 4672 7144 4688
rect 3816 4652 3832 4668
rect 4152 4652 4168 4668
rect 5208 4652 5224 4668
rect 6248 4652 6264 4668
rect 6648 4652 6664 4668
rect 6728 4652 6744 4668
rect 344 4632 360 4648
rect 1512 4632 1528 4648
rect 1624 4632 1640 4648
rect 2264 4632 2280 4648
rect 4856 4632 4872 4648
rect 5320 4632 5336 4648
rect 6472 4632 6488 4648
rect 7400 4632 7416 4648
rect 904 4612 920 4628
rect 1928 4612 1944 4628
rect 1048 4592 1064 4608
rect 1950 4602 1978 4618
rect 2872 4592 2888 4608
rect 3998 4602 4026 4618
rect 4056 4612 4072 4628
rect 5752 4612 5768 4628
rect 5848 4612 5864 4628
rect 6046 4602 6074 4618
rect 6088 4592 6104 4608
rect 6232 4592 6248 4608
rect 6408 4592 6424 4608
rect 872 4572 888 4588
rect 1016 4572 1032 4588
rect 1208 4572 1224 4588
rect 1720 4572 1736 4588
rect 1832 4572 1848 4588
rect 1880 4572 1896 4588
rect 2760 4572 2776 4588
rect 4616 4572 4632 4588
rect 6712 4572 6728 4588
rect 6760 4572 6776 4588
rect 1128 4552 1144 4568
rect 4872 4552 4888 4568
rect 6408 4552 6424 4568
rect 6632 4552 6648 4568
rect 6680 4552 6696 4568
rect 7832 4552 7848 4568
rect 40 4532 56 4548
rect 312 4532 328 4548
rect 872 4532 888 4548
rect 1016 4532 1032 4548
rect 1096 4532 1112 4548
rect 1816 4532 1848 4548
rect 3784 4532 3800 4548
rect 5528 4532 5544 4548
rect 6648 4532 6664 4548
rect 312 4512 328 4528
rect 376 4512 392 4528
rect 1400 4512 1416 4528
rect 1480 4512 1496 4528
rect 1896 4512 1912 4528
rect 2056 4512 2072 4528
rect 3912 4512 3928 4528
rect 4824 4512 4840 4528
rect 5176 4512 5192 4528
rect 5192 4512 5208 4528
rect 6664 4512 6680 4528
rect 6984 4512 7000 4528
rect 520 4492 536 4508
rect 2072 4492 2088 4508
rect 4008 4492 4024 4508
rect 5912 4492 5928 4508
rect 5992 4492 6008 4508
rect 6088 4492 6104 4508
rect 3304 4472 3336 4488
rect 3816 4472 3832 4488
rect 3928 4472 3944 4488
rect 4200 4472 4216 4488
rect 328 4452 344 4468
rect 424 4452 440 4468
rect 3896 4452 3912 4468
rect 7480 4452 7496 4468
rect 488 4432 504 4448
rect 824 4432 840 4448
rect 2584 4432 2600 4448
rect 6424 4432 6440 4448
rect 6456 4432 6472 4448
rect 926 4402 954 4418
rect 2958 4402 2986 4418
rect 3992 4412 4008 4428
rect 3224 4392 3240 4408
rect 5022 4402 5050 4418
rect 6904 4392 6920 4408
rect 7054 4402 7082 4418
rect 1928 4372 1944 4388
rect 2856 4372 2872 4388
rect 2920 4372 2936 4388
rect 3160 4372 3176 4388
rect 3624 4372 3640 4388
rect 968 4352 984 4368
rect 3288 4352 3304 4368
rect 3672 4352 3688 4368
rect 4568 4352 4584 4368
rect 6168 4352 6184 4368
rect 632 4332 648 4348
rect 1528 4332 1544 4348
rect 2024 4332 2056 4348
rect 3976 4332 3992 4348
rect 6616 4332 6632 4348
rect 6664 4332 6680 4348
rect 344 4312 360 4328
rect 1272 4312 1288 4328
rect 3192 4312 3208 4328
rect 3224 4312 3240 4328
rect 3720 4312 3736 4328
rect 3912 4312 3928 4328
rect 6120 4312 6136 4328
rect 8 4292 24 4308
rect 1768 4292 1784 4308
rect 2008 4292 2024 4308
rect 3656 4292 3672 4308
rect 3848 4292 3864 4308
rect 5656 4292 5672 4308
rect 5976 4292 5992 4308
rect 6312 4292 6328 4308
rect 376 4272 392 4288
rect 3736 4272 3768 4288
rect 3896 4272 3912 4288
rect 3944 4272 3960 4288
rect 7016 4272 7032 4288
rect 3896 4252 3912 4268
rect 1368 4232 1384 4248
rect 1576 4192 1592 4208
rect 1950 4202 1978 4218
rect 3336 4212 3352 4228
rect 3998 4202 4026 4218
rect 5912 4212 5928 4228
rect 6046 4202 6074 4218
rect 6728 4212 6744 4228
rect 8 4172 24 4188
rect 2040 4172 2056 4188
rect 2920 4172 2936 4188
rect 3352 4172 3368 4188
rect 3544 4172 3560 4188
rect 3880 4172 3896 4188
rect 7160 4172 7176 4188
rect 2936 4152 2952 4168
rect 3672 4152 3688 4168
rect 4856 4152 4872 4168
rect 6456 4152 6472 4168
rect 2600 4132 2616 4148
rect 2824 4132 2840 4148
rect 3944 4132 3960 4148
rect 6488 4132 6504 4148
rect 6920 4132 6936 4148
rect 344 4112 360 4128
rect 776 4112 792 4128
rect 1096 4112 1112 4128
rect 888 4092 904 4108
rect 1672 4112 1688 4128
rect 1736 4112 1752 4128
rect 1816 4112 1832 4128
rect 2264 4112 2280 4128
rect 2792 4112 2808 4128
rect 2856 4112 2872 4128
rect 4344 4112 4360 4128
rect 5928 4112 5944 4128
rect 1848 4092 1864 4108
rect 3128 4092 3144 4108
rect 3224 4092 3240 4108
rect 3272 4092 3288 4108
rect 3416 4092 3432 4108
rect 3720 4092 3736 4108
rect 3800 4092 3816 4108
rect 4216 4092 4232 4108
rect 5640 4092 5656 4108
rect 1528 4072 1544 4088
rect 3320 4072 3336 4088
rect 3832 4072 3848 4088
rect 1848 4052 1864 4068
rect 6840 4052 6856 4068
rect 3976 4032 3992 4048
rect 926 4002 954 4018
rect 2024 3992 2040 4008
rect 2088 3992 2104 4008
rect 2958 4002 2986 4018
rect 5022 4002 5050 4018
rect 6440 4012 6456 4028
rect 6024 3992 6040 4008
rect 7054 4002 7082 4018
rect 2872 3972 2888 3988
rect 6008 3972 6024 3988
rect 312 3952 328 3968
rect 3416 3952 3432 3968
rect 3928 3952 3944 3968
rect 1400 3932 1416 3948
rect 1448 3932 1464 3948
rect 2104 3932 2120 3948
rect 2360 3932 2376 3948
rect 3528 3932 3544 3948
rect 360 3912 376 3928
rect 1048 3912 1064 3928
rect 1416 3912 1432 3928
rect 3912 3912 3928 3928
rect 4184 3912 4200 3928
rect 7752 3912 7768 3928
rect 200 3892 216 3908
rect 728 3892 744 3908
rect 824 3892 840 3908
rect 1400 3892 1416 3908
rect 1608 3892 1624 3908
rect 728 3872 744 3888
rect 1240 3872 1256 3888
rect 1496 3872 1512 3888
rect 1800 3872 1816 3888
rect 3688 3892 3704 3908
rect 3720 3892 3736 3908
rect 4680 3892 4696 3908
rect 4712 3892 4728 3908
rect 2536 3872 2552 3888
rect 3448 3872 3464 3888
rect 5912 3892 5928 3908
rect 5912 3872 5928 3888
rect 5992 3892 6008 3908
rect 6248 3872 6264 3888
rect 6760 3872 6776 3888
rect 6952 3872 6968 3888
rect 7512 3872 7528 3888
rect 1000 3852 1016 3868
rect 1416 3852 1432 3868
rect 4856 3852 4872 3868
rect 6632 3852 6648 3868
rect 6968 3852 6984 3868
rect 392 3832 408 3848
rect 1240 3832 1256 3848
rect 1272 3832 1288 3848
rect 3944 3832 3960 3848
rect 5960 3832 5976 3848
rect 6136 3832 6152 3848
rect 6232 3832 6248 3848
rect 1800 3812 1816 3828
rect 8 3792 24 3808
rect 1950 3802 1978 3818
rect 2776 3792 2792 3808
rect 3928 3792 3944 3808
rect 3998 3802 4026 3818
rect 5864 3812 5880 3828
rect 4760 3792 4776 3808
rect 5064 3792 5080 3808
rect 6046 3802 6074 3818
rect 6408 3812 6424 3828
rect 6984 3812 7000 3828
rect 2760 3772 2776 3788
rect 2952 3772 2968 3788
rect 3176 3772 3208 3788
rect 3592 3772 3608 3788
rect 1016 3752 1032 3768
rect 2824 3752 2840 3768
rect 4040 3772 4056 3788
rect 4184 3772 4200 3788
rect 4888 3772 4904 3788
rect 5720 3772 5736 3788
rect 6296 3772 6312 3788
rect 6840 3772 6856 3788
rect 6904 3772 6920 3788
rect 5912 3752 5928 3768
rect 6168 3752 6184 3768
rect 312 3732 328 3748
rect 1592 3732 1608 3748
rect 1736 3732 1768 3748
rect 1800 3732 1816 3748
rect 2104 3732 2136 3748
rect 2760 3732 2776 3748
rect 2776 3732 2792 3748
rect 3096 3732 3112 3748
rect 4024 3732 4040 3748
rect 8 3712 24 3728
rect 1272 3712 1288 3728
rect 1624 3712 1640 3728
rect 1688 3712 1704 3728
rect 1784 3712 1800 3728
rect 2584 3712 2600 3728
rect 2680 3712 2696 3728
rect 2808 3712 2824 3728
rect 2872 3712 2888 3728
rect 2952 3712 2968 3728
rect 3880 3712 3896 3728
rect 4824 3712 4840 3728
rect 5720 3712 5736 3728
rect 6536 3712 6552 3728
rect 2440 3692 2456 3708
rect 4088 3692 4104 3708
rect 5992 3692 6008 3708
rect 344 3672 360 3688
rect 1320 3672 1336 3688
rect 2584 3672 2600 3688
rect 3448 3672 3464 3688
rect 2008 3652 2024 3668
rect 5864 3652 5880 3668
rect 6088 3652 6104 3668
rect 7176 3652 7192 3668
rect 1576 3632 1592 3648
rect 5192 3632 5208 3648
rect 926 3602 954 3618
rect 2088 3612 2104 3628
rect 2392 3592 2408 3608
rect 2958 3602 2986 3618
rect 5022 3602 5050 3618
rect 7054 3602 7082 3618
rect 776 3572 792 3588
rect 2600 3572 2616 3588
rect 3272 3572 3288 3588
rect 3336 3572 3352 3588
rect 3928 3572 3944 3588
rect 7160 3572 7176 3588
rect 1128 3552 1144 3568
rect 1704 3532 1720 3548
rect 1784 3552 1800 3568
rect 4760 3552 4776 3568
rect 3224 3532 3240 3548
rect 3320 3532 3336 3548
rect 3848 3532 3864 3548
rect 3896 3532 3912 3548
rect 4712 3532 4728 3548
rect 424 3512 440 3528
rect 1528 3512 1544 3528
rect 2504 3512 2520 3528
rect 3128 3512 3144 3528
rect 3720 3512 3736 3528
rect 4536 3512 4552 3528
rect 5336 3512 5352 3528
rect 6696 3512 6712 3528
rect 6968 3512 6984 3528
rect 168 3492 184 3508
rect 968 3492 984 3508
rect 1016 3492 1032 3508
rect 2552 3492 2568 3508
rect 3432 3492 3448 3508
rect 3800 3492 3816 3508
rect 4856 3492 4872 3508
rect 5192 3492 5208 3508
rect 264 3472 280 3488
rect 1096 3472 1112 3488
rect 1688 3472 1704 3488
rect 2920 3472 2936 3488
rect 5640 3472 5656 3488
rect 6632 3472 6648 3488
rect 6952 3472 6968 3488
rect 1400 3452 1416 3468
rect 2024 3452 2040 3468
rect 2120 3452 2136 3468
rect 2616 3452 2632 3468
rect 3128 3452 3144 3468
rect 4888 3452 4920 3468
rect 5368 3452 5384 3468
rect 5432 3452 5448 3468
rect 6936 3452 6952 3468
rect 6968 3452 6984 3468
rect 248 3432 264 3448
rect 1560 3432 1576 3448
rect 2744 3432 2760 3448
rect 472 3392 488 3408
rect 648 3392 664 3408
rect 984 3392 1000 3408
rect 1768 3392 1784 3408
rect 1928 3392 1944 3408
rect 1950 3402 1978 3418
rect 3416 3432 3432 3448
rect 3064 3392 3080 3408
rect 3998 3402 4026 3418
rect 4888 3392 4904 3408
rect 6046 3402 6074 3418
rect 6216 3412 6232 3428
rect 6344 3412 6360 3428
rect 1176 3372 1192 3388
rect 1208 3352 1224 3368
rect 1368 3352 1384 3368
rect 1704 3352 1720 3368
rect 2776 3352 2792 3368
rect 1576 3332 1592 3348
rect 3176 3332 3192 3348
rect 4296 3332 4312 3348
rect 4760 3332 4776 3348
rect 152 3312 168 3328
rect 376 3312 392 3328
rect 392 3312 408 3328
rect 904 3312 920 3328
rect 1256 3312 1272 3328
rect 1560 3312 1576 3328
rect 3816 3312 3832 3328
rect 8 3292 24 3308
rect 1384 3292 1400 3308
rect 1800 3292 1816 3308
rect 2792 3292 2808 3308
rect 3096 3292 3112 3308
rect 3656 3292 3672 3308
rect 6024 3292 6040 3308
rect 7176 3292 7192 3308
rect 1208 3272 1224 3288
rect 1464 3272 1480 3288
rect 6984 3272 7000 3288
rect 7288 3272 7304 3288
rect 312 3252 328 3268
rect 360 3252 376 3268
rect 2280 3252 2296 3268
rect 2936 3232 2952 3248
rect 3368 3232 3384 3248
rect 5432 3232 5448 3248
rect 7752 3232 7768 3248
rect 926 3202 954 3218
rect 968 3212 984 3228
rect 2344 3212 2360 3228
rect 2936 3192 2952 3208
rect 2958 3202 2986 3218
rect 3064 3212 3080 3228
rect 4200 3212 4216 3228
rect 3640 3192 3656 3208
rect 5022 3202 5050 3218
rect 5064 3212 5080 3228
rect 5288 3212 5304 3228
rect 7054 3202 7082 3218
rect 728 3172 744 3188
rect 2264 3172 2280 3188
rect 6664 3172 6680 3188
rect 6728 3172 6744 3188
rect 6920 3172 6936 3188
rect 632 3152 648 3168
rect 1928 3152 1944 3168
rect 5064 3152 5080 3168
rect 440 3132 456 3148
rect 1368 3132 1384 3148
rect 2552 3132 2568 3148
rect 6456 3132 6472 3148
rect 7288 3132 7304 3148
rect 8056 3132 8072 3148
rect 2120 3112 2136 3128
rect 2392 3112 2408 3128
rect 2648 3112 2664 3128
rect 4760 3112 4776 3128
rect 360 3092 376 3108
rect 520 3092 536 3108
rect 872 3092 888 3108
rect 1256 3092 1272 3108
rect 2744 3092 2760 3108
rect 4072 3092 4088 3108
rect 5096 3092 5112 3108
rect 6120 3092 6136 3108
rect 6520 3092 6536 3108
rect 7816 3112 7832 3128
rect 8056 3092 8072 3108
rect 104 3072 120 3088
rect 968 3072 984 3088
rect 1992 3072 2008 3088
rect 2392 3072 2408 3088
rect 2888 3072 2904 3088
rect 2936 3072 2952 3088
rect 3016 3072 3032 3088
rect 3080 3072 3096 3088
rect 872 3052 888 3068
rect 2440 3052 2456 3068
rect 2824 3052 2840 3068
rect 904 3032 920 3048
rect 3224 3032 3240 3048
rect 1432 3012 1448 3028
rect 1950 3002 1978 3018
rect 5992 3032 6008 3048
rect 168 2972 184 2988
rect 424 2972 440 2988
rect 3998 3002 4026 3018
rect 6136 3032 6152 3048
rect 5320 2992 5336 3008
rect 5848 2992 5864 3008
rect 6046 3002 6074 3018
rect 7832 3012 7848 3028
rect 6952 2992 6968 3008
rect 648 2952 664 2968
rect 1336 2952 1352 2968
rect 1400 2952 1432 2968
rect 1912 2952 1928 2968
rect 2776 2972 2792 2988
rect 2904 2972 2920 2988
rect 3832 2952 3848 2968
rect 5304 2952 5320 2968
rect 440 2932 456 2948
rect 1560 2932 1592 2948
rect 2712 2932 2728 2948
rect 2872 2932 2888 2948
rect 248 2912 264 2928
rect 1624 2912 1640 2928
rect 1656 2912 1672 2928
rect 3544 2912 3560 2928
rect 6664 2912 6680 2928
rect 7448 2912 7464 2928
rect 424 2892 440 2908
rect 1720 2892 1736 2908
rect 3000 2892 3016 2908
rect 5080 2892 5096 2908
rect 5320 2892 5336 2908
rect 5912 2892 5928 2908
rect 2792 2852 2824 2868
rect 3032 2832 3048 2848
rect 3768 2832 3784 2848
rect 824 2792 840 2808
rect 926 2802 954 2818
rect 2056 2812 2072 2828
rect 2696 2812 2712 2828
rect 2808 2812 2824 2828
rect 2958 2802 2986 2818
rect 3592 2812 3608 2828
rect 4824 2812 4840 2828
rect 2024 2772 2040 2788
rect 5022 2802 5050 2818
rect 5832 2812 5848 2828
rect 6552 2812 6568 2828
rect 7054 2802 7082 2818
rect 6344 2772 6360 2788
rect 152 2752 168 2768
rect 1688 2752 1704 2768
rect 2648 2752 2664 2768
rect 3816 2752 3832 2768
rect 2488 2732 2504 2748
rect 600 2692 616 2708
rect 1176 2692 1192 2708
rect 1688 2692 1704 2708
rect 2024 2692 2040 2708
rect 2472 2692 2488 2708
rect 3080 2692 3096 2708
rect 6392 2712 6408 2728
rect 6008 2692 6024 2708
rect 7448 2692 7464 2708
rect 6104 2672 6120 2688
rect 6232 2672 6248 2688
rect 6488 2672 6504 2688
rect 5864 2652 5880 2668
rect 6824 2652 6840 2668
rect 1000 2632 1016 2648
rect 600 2612 616 2628
rect 808 2612 824 2628
rect 1464 2612 1480 2628
rect 264 2592 280 2608
rect 984 2592 1000 2608
rect 1736 2592 1752 2608
rect 1950 2602 1978 2618
rect 3998 2602 4026 2618
rect 5704 2612 5720 2628
rect 6046 2602 6074 2618
rect 6264 2612 6280 2628
rect 6312 2592 6328 2608
rect 7624 2592 7640 2608
rect 376 2572 392 2588
rect 904 2572 920 2588
rect 328 2552 344 2568
rect 2312 2572 2328 2588
rect 1448 2532 1464 2548
rect 2280 2532 2296 2548
rect 2744 2532 2760 2548
rect 7640 2532 7656 2548
rect 3544 2512 3560 2528
rect 6520 2512 6536 2528
rect 968 2492 984 2508
rect 1464 2492 1480 2508
rect 3032 2492 3048 2508
rect 5064 2492 5080 2508
rect 6776 2492 6792 2508
rect 376 2472 392 2488
rect 1016 2472 1032 2488
rect 1704 2472 1720 2488
rect 5848 2472 5864 2488
rect 7160 2472 7176 2488
rect 2264 2452 2280 2468
rect 1992 2432 2008 2448
rect 4200 2432 4216 2448
rect 5704 2432 5720 2448
rect 792 2392 808 2408
rect 926 2402 954 2418
rect 2958 2402 2986 2418
rect 3560 2392 3576 2408
rect 5022 2402 5050 2418
rect 7054 2402 7082 2418
rect 7800 2392 7816 2408
rect 7848 2392 7864 2408
rect 264 2372 280 2388
rect 1736 2372 1752 2388
rect 3736 2372 3768 2388
rect 6344 2372 6360 2388
rect 6568 2372 6584 2388
rect 1048 2352 1080 2368
rect 360 2332 376 2348
rect 296 2312 312 2328
rect 1192 2332 1208 2348
rect 1768 2332 1800 2348
rect 2024 2332 2040 2348
rect 2248 2332 2264 2348
rect 1736 2312 1752 2328
rect 2344 2312 2360 2328
rect 7624 2312 7640 2328
rect 408 2292 424 2308
rect 1896 2292 1912 2308
rect 2296 2292 2312 2308
rect 4680 2292 4696 2308
rect 5864 2292 5880 2308
rect 6248 2292 6264 2308
rect 6280 2292 6296 2308
rect 616 2272 632 2288
rect 4984 2272 5000 2288
rect 1464 2252 1480 2268
rect 3768 2252 3784 2268
rect 6216 2252 6232 2268
rect 6488 2252 6504 2268
rect 7416 2252 7432 2268
rect 1560 2232 1576 2248
rect 1608 2232 1624 2248
rect 3208 2232 3224 2248
rect 6984 2232 7000 2248
rect 1560 2212 1576 2228
rect 1950 2202 1978 2218
rect 3998 2202 4026 2218
rect 5832 2212 5848 2228
rect 4680 2192 4696 2208
rect 6046 2202 6074 2218
rect 6920 2192 6936 2208
rect 5592 2172 5608 2188
rect 6296 2172 6312 2188
rect 6824 2172 6840 2188
rect 2312 2152 2328 2168
rect 5576 2152 5592 2168
rect 7640 2152 7656 2168
rect 2376 2132 2392 2148
rect 3368 2132 3384 2148
rect 1672 2112 1688 2128
rect 840 2092 856 2108
rect 2440 2092 2456 2108
rect 4792 2112 4808 2128
rect 7160 2132 7176 2148
rect 6008 2112 6024 2128
rect 7688 2112 7704 2128
rect 7896 2112 7912 2128
rect 3032 2092 3048 2108
rect 3896 2092 3912 2108
rect 5848 2092 5864 2108
rect 5976 2092 5992 2108
rect 6392 2092 6408 2108
rect 536 2072 552 2088
rect 2264 2072 2280 2088
rect 3208 2052 3224 2068
rect 968 2032 984 2048
rect 2888 2032 2904 2048
rect 3752 2032 3768 2048
rect 926 2002 954 2018
rect 2958 2002 2986 2018
rect 3960 2012 3976 2028
rect 424 1972 440 1988
rect 2936 1972 2952 1988
rect 4824 1992 4840 2008
rect 5022 2002 5050 2018
rect 7054 2002 7082 2018
rect 5288 1972 5304 1988
rect 968 1952 984 1968
rect 1096 1952 1112 1968
rect 3096 1952 3112 1968
rect 232 1932 248 1948
rect 824 1932 840 1948
rect 2488 1932 2504 1948
rect 5288 1932 5304 1948
rect 4200 1912 4216 1928
rect 4760 1912 4776 1928
rect 4824 1912 4840 1928
rect 1016 1892 1032 1908
rect 1560 1892 1576 1908
rect 264 1872 280 1888
rect 3752 1892 3768 1908
rect 4856 1892 4872 1908
rect 5816 1892 5832 1908
rect 5960 1892 5976 1908
rect 6488 1892 6504 1908
rect 6680 1892 6696 1908
rect 7000 1872 7016 1888
rect 7016 1872 7048 1888
rect 6024 1852 6040 1868
rect 392 1832 408 1848
rect 1384 1832 1400 1848
rect 1950 1802 1978 1818
rect 3496 1812 3512 1828
rect 3944 1812 3960 1828
rect 3896 1792 3912 1808
rect 3998 1802 4026 1818
rect 6024 1812 6040 1828
rect 4184 1792 4200 1808
rect 2120 1772 2136 1788
rect 2552 1772 2568 1788
rect 6046 1802 6074 1818
rect 6280 1812 6296 1828
rect 6488 1792 6504 1808
rect 5592 1772 5608 1788
rect 7736 1772 7752 1788
rect 1448 1752 1464 1768
rect 2376 1752 2392 1768
rect 4424 1752 4440 1768
rect 4808 1752 4824 1768
rect 8 1732 24 1748
rect 1112 1732 1128 1748
rect 1352 1732 1368 1748
rect 1512 1732 1528 1748
rect 3656 1732 3672 1748
rect 4168 1732 4184 1748
rect 4184 1732 4200 1748
rect 120 1712 136 1728
rect 456 1712 472 1728
rect 792 1712 808 1728
rect 1336 1712 1352 1728
rect 1688 1712 1704 1728
rect 3688 1712 3704 1728
rect 6008 1712 6024 1728
rect 6808 1732 6824 1748
rect 6456 1712 6472 1728
rect 6552 1712 6568 1728
rect 6760 1712 6776 1728
rect 7480 1712 7496 1728
rect 7768 1712 7784 1728
rect 568 1692 584 1708
rect 712 1692 728 1708
rect 2136 1692 2152 1708
rect 2312 1692 2328 1708
rect 952 1672 968 1688
rect 1064 1672 1080 1688
rect 1160 1672 1176 1688
rect 1928 1672 1960 1688
rect 3496 1672 3512 1688
rect 4232 1692 4248 1708
rect 4360 1692 4376 1708
rect 5048 1692 5064 1708
rect 7400 1672 7416 1688
rect 4424 1652 4440 1668
rect 536 1632 552 1648
rect 1624 1632 1640 1648
rect 1816 1632 1832 1648
rect 3432 1632 3448 1648
rect 3512 1632 3528 1648
rect 840 1612 856 1628
rect 168 1592 184 1608
rect 926 1602 954 1618
rect 1016 1592 1032 1608
rect 2958 1602 2986 1618
rect 3128 1592 3144 1608
rect 4824 1592 4840 1608
rect 5022 1602 5050 1618
rect 6248 1612 6264 1628
rect 7054 1602 7082 1618
rect 1944 1572 1960 1588
rect 3352 1572 3368 1588
rect 8 1552 24 1568
rect 1624 1552 1640 1568
rect 3912 1552 3928 1568
rect 472 1532 488 1548
rect 1624 1532 1640 1548
rect 3544 1532 3560 1548
rect 3672 1532 3688 1548
rect 6520 1532 6536 1548
rect 6792 1532 6808 1548
rect 8 1512 24 1528
rect 1784 1512 1800 1528
rect 2920 1512 2936 1528
rect 3592 1512 3608 1528
rect 3944 1512 3960 1528
rect 3976 1512 3992 1528
rect 5576 1512 5592 1528
rect 5816 1512 5832 1528
rect 6568 1512 6584 1528
rect 7512 1512 7528 1528
rect 152 1492 168 1508
rect 456 1492 472 1508
rect 808 1492 824 1508
rect 2280 1492 2296 1508
rect 2776 1492 2792 1508
rect 4696 1492 4712 1508
rect 4760 1492 4776 1508
rect 7400 1492 7416 1508
rect 328 1472 344 1488
rect 1000 1472 1016 1488
rect 1816 1472 1832 1488
rect 2728 1472 2744 1488
rect 6616 1472 6632 1488
rect 6872 1472 6888 1488
rect 6936 1472 6952 1488
rect 7176 1472 7192 1488
rect 7240 1472 7256 1488
rect 1832 1452 1848 1468
rect 4696 1452 4712 1468
rect 6344 1452 6360 1468
rect 6360 1452 6376 1468
rect 6552 1452 6568 1468
rect 7384 1452 7400 1468
rect 7512 1452 7528 1468
rect 7736 1452 7752 1468
rect 6104 1432 6120 1448
rect 280 1412 296 1428
rect 1288 1392 1304 1408
rect 1950 1402 1978 1418
rect 3768 1412 3784 1428
rect 3320 1392 3336 1408
rect 3960 1392 3976 1408
rect 3998 1402 4026 1418
rect 5096 1412 5112 1428
rect 6024 1412 6040 1428
rect 4216 1392 4232 1408
rect 6046 1402 6074 1418
rect 264 1372 280 1388
rect 1672 1372 1688 1388
rect 3448 1372 3464 1388
rect 4232 1372 4248 1388
rect 6376 1372 6392 1388
rect 6888 1372 6904 1388
rect 248 1332 264 1348
rect 536 1352 552 1368
rect 2120 1352 2136 1368
rect 3496 1352 3512 1368
rect 4328 1352 4344 1368
rect 6344 1352 6360 1368
rect 7512 1352 7528 1368
rect 1128 1332 1144 1348
rect 1176 1332 1192 1348
rect 1656 1332 1672 1348
rect 3800 1332 3816 1348
rect 3880 1332 3896 1348
rect 4152 1332 4168 1348
rect 5688 1332 5704 1348
rect 6296 1332 6312 1348
rect 6520 1332 6536 1348
rect 6680 1332 6696 1348
rect 6808 1332 6824 1348
rect 232 1312 248 1328
rect 328 1312 344 1328
rect 408 1312 424 1328
rect 584 1312 600 1328
rect 824 1312 840 1328
rect 1240 1312 1256 1328
rect 1272 1312 1288 1328
rect 2696 1312 2712 1328
rect 4456 1312 4472 1328
rect 4776 1312 4792 1328
rect 4984 1312 5000 1328
rect 5512 1312 5528 1328
rect 5880 1312 5896 1328
rect 5992 1312 6024 1328
rect 6520 1312 6536 1328
rect 6792 1312 6808 1328
rect 6968 1312 6984 1328
rect 7016 1312 7032 1328
rect 7848 1312 7864 1328
rect 8 1292 24 1308
rect 504 1292 520 1308
rect 536 1292 552 1308
rect 3832 1292 3848 1308
rect 3864 1292 3880 1308
rect 4760 1292 4776 1308
rect 4792 1292 4808 1308
rect 6888 1292 6904 1308
rect 7928 1292 7944 1308
rect 312 1272 328 1288
rect 424 1272 440 1288
rect 472 1272 488 1288
rect 1928 1272 1944 1288
rect 3832 1272 3848 1288
rect 7224 1272 7240 1288
rect 7896 1272 7912 1288
rect 1432 1252 1448 1268
rect 1816 1252 1832 1268
rect 456 1232 472 1248
rect 1160 1232 1176 1248
rect 1784 1232 1800 1248
rect 1928 1232 1944 1248
rect 2008 1232 2024 1248
rect 4456 1252 4472 1268
rect 3816 1232 3832 1248
rect 3880 1232 3896 1248
rect 6664 1232 6680 1248
rect 536 1192 552 1208
rect 926 1202 954 1218
rect 1304 1212 1320 1228
rect 1288 1192 1304 1208
rect 1416 1192 1432 1208
rect 2958 1202 2986 1218
rect 3000 1192 3016 1208
rect 5022 1202 5050 1218
rect 7054 1202 7082 1218
rect 7848 1212 7864 1228
rect 72 1152 88 1168
rect 184 1152 200 1168
rect 472 1152 488 1168
rect 2728 1152 2744 1168
rect 3768 1152 3784 1168
rect 7224 1152 7240 1168
rect 7832 1152 7848 1168
rect 24 1132 40 1148
rect 264 1132 280 1148
rect 424 1132 440 1148
rect 1176 1132 1192 1148
rect 2856 1132 2872 1148
rect 3560 1132 3576 1148
rect 5624 1132 5640 1148
rect 840 1112 856 1128
rect 3144 1112 3160 1128
rect 120 1092 136 1108
rect 408 1092 424 1108
rect 776 1092 808 1108
rect 1144 1092 1160 1108
rect 1288 1092 1320 1108
rect 1400 1092 1416 1108
rect 1800 1092 1816 1108
rect 3688 1112 3704 1128
rect 3720 1112 3736 1128
rect 3784 1112 3800 1128
rect 3976 1112 3992 1128
rect 4968 1112 4984 1128
rect 3560 1092 3592 1108
rect 3848 1092 3864 1108
rect 6008 1092 6024 1108
rect 584 1072 600 1088
rect 664 1072 680 1088
rect 712 1052 728 1068
rect 2136 1072 2152 1088
rect 3768 1072 3784 1088
rect 4328 1072 4344 1088
rect 6744 1072 6760 1088
rect 7832 1092 7848 1108
rect 3752 1052 3768 1068
rect 4344 1052 4360 1068
rect 6168 1052 6200 1068
rect 6696 1052 6712 1068
rect 7720 1052 7736 1068
rect 7816 1052 7832 1068
rect 7912 1052 7928 1068
rect 1192 1032 1208 1048
rect 1432 1032 1448 1048
rect 1896 1032 1912 1048
rect 4248 1032 4264 1048
rect 472 1012 488 1028
rect 1672 992 1688 1008
rect 1950 1002 1978 1018
rect 3800 992 3816 1008
rect 3998 1002 4026 1018
rect 6264 1032 6280 1048
rect 6808 1032 6824 1048
rect 7864 1032 7880 1048
rect 6046 1002 6074 1018
rect 6168 1012 6184 1028
rect 7480 1012 7496 1028
rect 1176 972 1192 988
rect 2376 972 2392 988
rect 3832 972 3848 988
rect 6184 972 6200 988
rect 6488 972 6504 988
rect 6856 972 6872 988
rect 1880 952 1896 968
rect 4136 952 4152 968
rect 392 932 408 948
rect 1800 932 1816 948
rect 3480 932 3496 948
rect 3784 932 3800 948
rect 5624 952 5640 968
rect 6216 952 6232 968
rect 4856 932 4872 948
rect 6296 932 6312 948
rect 6392 932 6408 948
rect 120 912 136 928
rect 280 912 296 928
rect 616 912 632 928
rect 1064 912 1080 928
rect 1896 912 1912 928
rect 4120 912 4136 928
rect 4392 912 4408 928
rect 4712 912 4728 928
rect 5832 912 5848 928
rect 6536 912 6552 928
rect 6776 912 6792 928
rect 7512 912 7528 928
rect 7848 912 7864 928
rect 2008 892 2024 908
rect 2696 892 2712 908
rect 3656 892 3672 908
rect 6600 892 6616 908
rect 6808 892 6824 908
rect 312 872 328 888
rect 4200 852 4216 868
rect 4408 852 4424 868
rect 6296 852 6312 868
rect 6024 832 6040 848
rect 376 812 392 828
rect 926 802 954 818
rect 2958 802 2986 818
rect 3592 812 3608 828
rect 5022 802 5050 818
rect 6280 792 6296 808
rect 7054 802 7082 818
rect 424 772 440 788
rect 6696 772 6712 788
rect 6264 752 6280 768
rect 3912 732 3928 748
rect 4168 732 4184 748
rect 5976 732 5992 748
rect 6744 732 6760 748
rect 3032 712 3048 728
rect 3784 712 3800 728
rect 4120 712 4136 728
rect 6760 712 6776 728
rect 7832 712 7848 728
rect 968 692 984 708
rect 1064 692 1096 708
rect 1416 672 1432 688
rect 3096 692 3112 708
rect 3576 692 3592 708
rect 3736 692 3752 708
rect 3816 692 3832 708
rect 3976 692 3992 708
rect 7784 692 7800 708
rect 3032 672 3048 688
rect 3768 672 3784 688
rect 3832 672 3848 688
rect 4376 672 4392 688
rect 5464 672 5480 688
rect 6728 672 6744 688
rect 7480 672 7496 688
rect 3000 652 3016 668
rect 3592 652 3608 668
rect 3704 652 3720 668
rect 3880 652 3912 668
rect 7016 652 7032 668
rect 4344 632 4360 648
rect 6888 632 6904 648
rect 1800 592 1816 608
rect 1950 602 1978 618
rect 1992 612 2008 628
rect 3512 612 3528 628
rect 3998 602 4026 618
rect 6024 612 6040 628
rect 4888 592 4904 608
rect 6046 602 6074 618
rect 1656 572 1672 588
rect 1256 552 1272 568
rect 1400 552 1416 568
rect 3016 552 3032 568
rect 3064 552 3080 568
rect 3752 552 3768 568
rect 4744 572 4760 588
rect 5448 552 5464 568
rect 344 532 360 548
rect 3032 532 3048 548
rect 408 512 424 528
rect 1416 512 1432 528
rect 1624 512 1640 528
rect 2136 512 2152 528
rect 2616 512 2632 528
rect 3768 532 3784 548
rect 4888 512 4904 528
rect 312 472 328 488
rect 2600 492 2616 508
rect 3896 492 3912 508
rect 4248 492 4264 508
rect 4792 492 4808 508
rect 1784 472 1800 488
rect 2216 472 2232 488
rect 3240 472 3256 488
rect 4120 472 4136 488
rect 488 452 504 468
rect 1512 452 1528 468
rect 1544 452 1560 468
rect 6184 452 6200 468
rect 24 432 40 448
rect 3864 432 3880 448
rect 616 412 632 428
rect 808 392 824 408
rect 926 402 954 418
rect 2536 392 2552 408
rect 2958 402 2986 418
rect 5022 402 5050 418
rect 7054 402 7082 418
rect 344 372 360 388
rect 1544 352 1560 368
rect 24 332 40 348
rect 264 332 280 348
rect 424 332 440 348
rect 1064 332 1080 348
rect 2120 332 2136 348
rect 2776 332 2792 348
rect 2856 332 2872 348
rect 3432 332 3448 348
rect 6728 332 6744 348
rect 616 312 632 328
rect 1384 312 1400 328
rect 6680 312 6696 328
rect 7880 312 7896 328
rect 328 292 344 308
rect 3480 292 3496 308
rect 4392 292 4408 308
rect 5736 292 5752 308
rect 5464 272 5480 288
rect 1950 202 1978 218
rect 3000 192 3016 208
rect 3998 202 4026 218
rect 5880 212 5896 228
rect 6046 202 6074 218
rect 3464 172 3480 188
rect 3496 172 3512 188
rect 3736 152 3752 168
rect 280 132 296 148
rect 3672 112 3688 128
rect 3736 112 3752 128
rect 5960 112 5976 128
rect 4136 92 4152 108
rect 926 2 954 18
rect 1832 12 1848 28
rect 2696 12 2712 28
rect 2958 2 2986 18
rect 3448 12 3464 28
rect 4328 12 4344 28
rect 5022 2 5050 18
rect 7054 2 7082 18
<< metal4 >>
rect 954 5606 960 5614
rect 77 5268 83 5492
rect 77 5248 83 5252
rect 333 4968 339 5372
rect 333 4908 339 4952
rect 45 4548 51 4692
rect 317 4528 323 4532
rect 332 4516 340 4524
rect 13 4188 19 4292
rect 317 3968 323 4512
rect 333 4468 339 4516
rect 349 4328 355 4632
rect 381 4288 387 4512
rect 429 4468 435 4692
rect 13 3728 19 3792
rect 92 3083 100 3084
rect 92 3077 104 3083
rect 92 3076 100 3077
rect 157 2768 163 3312
rect 173 2988 179 3492
rect 13 1528 19 1552
rect 13 1284 19 1292
rect 12 1276 20 1284
rect 29 448 35 1132
rect 125 1108 131 1712
rect 157 1508 163 2752
rect 173 1608 179 2972
rect 253 2928 259 3432
rect 269 2608 275 3472
rect 317 3268 323 3732
rect 349 3688 355 4112
rect 365 3268 371 3912
rect 397 3328 403 3832
rect 237 1328 243 1932
rect 269 1888 275 2372
rect 333 1488 339 2552
rect 365 2348 371 3092
rect 381 2588 387 3312
rect 429 2988 435 3512
rect 477 3408 483 4912
rect 525 4508 531 5352
rect 954 5206 960 5214
rect 637 4348 643 4812
rect 637 3168 643 4332
rect 733 3908 739 4912
rect 954 4806 960 4814
rect 973 4768 979 4792
rect 876 4756 884 4764
rect 877 4588 883 4756
rect 844 4443 852 4444
rect 840 4437 852 4443
rect 844 4436 852 4437
rect 652 3436 660 3444
rect 653 3408 659 3436
rect 733 3188 739 3872
rect 781 3588 787 4112
rect 893 4108 899 4732
rect 844 3903 852 3904
rect 840 3897 852 3903
rect 844 3896 852 3897
rect 909 3328 915 4612
rect 954 4406 960 4414
rect 973 4368 979 4732
rect 1021 4588 1027 5072
rect 1085 4908 1091 5452
rect 1978 5406 1984 5414
rect 1052 4703 1060 4704
rect 1048 4697 1060 4703
rect 1052 4696 1060 4697
rect 1021 4548 1027 4572
rect 954 4006 960 4014
rect 1053 3928 1059 4592
rect 1101 4548 1107 5352
rect 1244 4983 1252 4984
rect 1244 4977 1256 4983
rect 1244 4976 1252 4977
rect 1212 4696 1220 4704
rect 1213 4588 1219 4696
rect 954 3606 960 3614
rect 1021 3508 1027 3752
rect 973 3228 979 3492
rect 954 3206 960 3214
rect 445 2948 451 3132
rect 524 3116 532 3124
rect 525 3108 531 3116
rect 860 3103 868 3104
rect 860 3097 872 3103
rect 860 3096 868 3097
rect 653 2944 659 2952
rect 652 2936 660 2944
rect 412 2903 420 2904
rect 412 2897 424 2903
rect 412 2896 420 2897
rect 605 2628 611 2692
rect 253 1304 259 1332
rect 252 1296 260 1304
rect 172 1163 180 1164
rect 172 1157 184 1163
rect 172 1156 180 1157
rect 269 1148 275 1372
rect 125 928 131 1092
rect 29 348 35 432
rect 269 348 275 1132
rect 285 928 291 1412
rect 285 148 291 912
rect 317 888 323 1272
rect 317 488 323 872
rect 333 308 339 1312
rect 381 828 387 2472
rect 397 948 403 1832
rect 413 1328 419 2292
rect 413 1108 419 1312
rect 429 1288 435 1972
rect 461 1508 467 1712
rect 541 1648 547 2072
rect 460 1316 468 1324
rect 461 1248 467 1316
rect 477 1288 483 1532
rect 541 1368 547 1632
rect 524 1303 532 1304
rect 520 1297 532 1303
rect 524 1296 532 1297
rect 541 1284 547 1292
rect 540 1276 548 1284
rect 540 1256 548 1264
rect 541 1208 547 1256
rect 349 388 355 532
rect 413 528 419 1092
rect 429 788 435 1132
rect 477 1028 483 1152
rect 589 1088 595 1312
rect 621 964 627 2272
rect 797 1728 803 2392
rect 717 1068 723 1692
rect 797 1108 803 1712
rect 813 1524 819 2612
rect 829 1948 835 2792
rect 909 2588 915 3032
rect 954 2806 960 2814
rect 973 2508 979 3072
rect 989 2608 995 3392
rect 954 2406 960 2414
rect 812 1516 820 1524
rect 813 1508 819 1516
rect 829 1328 835 1932
rect 845 1628 851 2092
rect 954 2006 960 2014
rect 973 1968 979 2032
rect 956 1716 964 1724
rect 957 1688 963 1716
rect 845 1128 851 1612
rect 954 1606 960 1614
rect 1005 1488 1011 2632
rect 1021 2488 1027 3492
rect 1101 3488 1107 4112
rect 1133 3568 1139 4552
rect 1277 4328 1283 5252
rect 1340 4723 1348 4724
rect 1336 4717 1348 4723
rect 1340 4716 1348 4717
rect 1373 4248 1379 4832
rect 1405 3948 1411 4512
rect 1421 3928 1427 5152
rect 1437 4688 1443 4732
rect 1517 4648 1523 4692
rect 1500 4523 1508 4524
rect 1496 4517 1508 4523
rect 1500 4516 1508 4517
rect 1533 4348 1539 4872
rect 1533 4088 1539 4332
rect 1581 4208 1587 5332
rect 1724 4736 1732 4744
rect 1612 4643 1620 4644
rect 1612 4637 1624 4643
rect 1612 4636 1620 4637
rect 1725 4588 1731 4736
rect 1405 3884 1411 3892
rect 1404 3876 1412 3884
rect 1245 3848 1251 3872
rect 1436 3863 1444 3864
rect 1432 3857 1444 3863
rect 1436 3856 1444 3857
rect 1277 3728 1283 3832
rect 1324 3696 1332 3704
rect 1325 3688 1331 3696
rect 1021 1908 1027 2472
rect 1053 2344 1059 2352
rect 1052 2336 1060 2344
rect 1021 1608 1027 1892
rect 1069 1688 1075 2352
rect 1101 1968 1107 3472
rect 1181 2708 1187 3372
rect 1213 3288 1219 3352
rect 1261 3108 1267 3312
rect 1373 3148 1379 3352
rect 1405 2968 1411 3452
rect 1437 2984 1443 3012
rect 1436 2976 1444 2984
rect 1324 2963 1332 2964
rect 1324 2957 1336 2963
rect 1324 2956 1332 2957
rect 1453 2548 1459 3932
rect 1516 3883 1524 3884
rect 1512 3877 1524 3883
rect 1516 3876 1524 3877
rect 1533 3528 1539 4072
rect 1596 3756 1604 3764
rect 1597 3748 1603 3756
rect 1565 3328 1571 3432
rect 1581 3348 1587 3632
rect 1469 2628 1475 3272
rect 1565 2948 1571 3312
rect 1100 1743 1108 1744
rect 1100 1737 1112 1743
rect 1100 1736 1108 1737
rect 1341 1704 1347 1712
rect 1357 1704 1363 1732
rect 1340 1696 1348 1704
rect 1356 1696 1364 1704
rect 1148 1343 1156 1344
rect 1144 1337 1156 1343
rect 1148 1336 1156 1337
rect 1165 1248 1171 1672
rect 1276 1336 1284 1344
rect 954 1206 960 1214
rect 1181 1148 1187 1332
rect 1277 1328 1283 1336
rect 1260 1323 1268 1324
rect 1256 1317 1268 1323
rect 1260 1316 1268 1317
rect 1293 1208 1299 1392
rect 1309 1108 1315 1212
rect 1164 1103 1172 1104
rect 1160 1097 1172 1103
rect 1164 1096 1172 1097
rect 1180 1043 1188 1044
rect 1180 1037 1192 1043
rect 1180 1036 1188 1037
rect 1164 983 1172 984
rect 1164 977 1176 983
rect 1164 976 1172 977
rect 620 956 628 964
rect 621 928 627 956
rect 954 806 960 814
rect 429 348 435 772
rect 1069 708 1075 912
rect 988 703 996 704
rect 984 697 996 703
rect 988 696 996 697
rect 1100 703 1108 704
rect 1096 697 1108 703
rect 1100 696 1108 697
rect 812 516 820 524
rect 492 496 500 504
rect 493 468 499 496
rect 621 328 627 412
rect 813 408 819 516
rect 954 406 960 414
rect 1069 348 1075 692
rect 1261 544 1267 552
rect 1260 536 1268 544
rect 1389 328 1395 1832
rect 1453 1768 1459 2532
rect 1469 2268 1475 2492
rect 1613 2248 1619 3892
rect 1629 2928 1635 3712
rect 1565 2228 1571 2232
rect 1565 1908 1571 2212
rect 1629 1568 1635 1632
rect 1629 1504 1635 1532
rect 1628 1496 1636 1504
rect 1661 1348 1667 2912
rect 1677 2128 1683 4112
rect 1741 3748 1747 4112
rect 1773 3884 1779 4292
rect 1772 3876 1780 3884
rect 1693 3488 1699 3712
rect 1709 3524 1715 3532
rect 1708 3516 1716 3524
rect 1709 3104 1715 3352
rect 1708 3096 1716 3104
rect 1693 2708 1699 2752
rect 1709 2488 1715 3096
rect 1741 2608 1747 3732
rect 1773 3408 1779 3876
rect 1789 3728 1795 5332
rect 1978 5006 1984 5014
rect 1884 4656 1892 4664
rect 1885 4588 1891 4656
rect 1837 4548 1843 4572
rect 1900 4536 1908 4544
rect 1821 4128 1827 4532
rect 1901 4528 1907 4536
rect 1933 4388 1939 4612
rect 1978 4606 1984 4614
rect 1978 4206 1984 4214
rect 1853 4068 1859 4092
rect 1805 3828 1811 3872
rect 1805 3748 1811 3812
rect 1978 3806 1984 3814
rect 1741 2328 1747 2372
rect 1789 2348 1795 3552
rect 1805 3308 1811 3732
rect 2013 3668 2019 4292
rect 2029 4008 2035 4332
rect 2045 4188 2051 4332
rect 2029 3468 2035 3992
rect 1978 3406 1984 3414
rect 1933 3168 1939 3392
rect 1978 3006 1984 3014
rect 1900 2963 1908 2964
rect 1900 2957 1912 2963
rect 1900 2956 1908 2957
rect 2061 2828 2067 4512
rect 2077 4508 2083 5472
rect 2269 5348 2275 5612
rect 2986 5606 2992 5614
rect 2269 4708 2275 5112
rect 2365 4768 2371 4892
rect 2269 4128 2275 4632
rect 2093 3628 2099 3992
rect 2109 3748 2115 3932
rect 2125 3128 2131 3452
rect 2269 3188 2275 4112
rect 2365 3948 2371 4752
rect 2589 4384 2595 4432
rect 2588 4376 2596 4384
rect 2556 3883 2564 3884
rect 2552 3877 2564 3883
rect 2556 3876 2564 3877
rect 2589 3728 2595 4376
rect 2029 2708 2035 2772
rect 1978 2606 1984 2614
rect 2252 2496 2260 2504
rect 1773 2304 1779 2332
rect 1772 2296 1780 2304
rect 1677 1388 1683 2112
rect 1708 1723 1716 1724
rect 1704 1717 1716 1723
rect 1708 1716 1716 1717
rect 1789 1528 1795 2332
rect 1916 2303 1924 2304
rect 1912 2297 1924 2303
rect 1916 2296 1924 2297
rect 1978 2206 1984 2214
rect 1978 1806 1984 1814
rect 1821 1488 1827 1632
rect 1452 1263 1460 1264
rect 1448 1257 1460 1263
rect 1452 1256 1460 1257
rect 1405 1084 1411 1092
rect 1404 1076 1412 1084
rect 1421 688 1427 1192
rect 1437 944 1443 1032
rect 1677 1008 1683 1372
rect 1821 1268 1827 1472
rect 1436 936 1444 944
rect 1644 583 1652 584
rect 1644 577 1656 583
rect 1644 576 1652 577
rect 1416 557 1427 563
rect 1421 528 1427 557
rect 1629 504 1635 512
rect 1628 496 1636 504
rect 1789 488 1795 1232
rect 1820 1103 1828 1104
rect 1816 1097 1828 1103
rect 1820 1096 1828 1097
rect 1805 608 1811 932
rect 1532 463 1540 464
rect 1528 457 1540 463
rect 1532 456 1540 457
rect 1549 368 1555 452
rect 1837 28 1843 1452
rect 1933 1288 1939 1672
rect 1949 1588 1955 1672
rect 1978 1406 1984 1414
rect 1933 1248 1939 1272
rect 1901 928 1907 1032
rect 1978 1006 1984 1014
rect 1997 628 2003 2432
rect 2253 2348 2259 2496
rect 2269 2468 2275 3172
rect 2285 2548 2291 3252
rect 2029 2324 2035 2332
rect 2028 2316 2036 2324
rect 2269 2088 2275 2452
rect 2317 2168 2323 2572
rect 2349 2328 2355 3212
rect 2397 3128 2403 3592
rect 2445 3068 2451 3692
rect 2524 3523 2532 3524
rect 2520 3517 2532 3523
rect 2524 3516 2532 3517
rect 2557 3148 2563 3492
rect 2589 3444 2595 3672
rect 2605 3588 2611 4132
rect 2621 3468 2627 5212
rect 2765 3788 2771 4572
rect 2781 3808 2787 4832
rect 2813 4688 2819 5492
rect 3181 5488 3187 5612
rect 5050 5606 5056 5614
rect 7082 5606 7088 5614
rect 4026 5406 4032 5414
rect 2986 5206 2992 5214
rect 2844 4716 2852 4724
rect 2845 4708 2851 4716
rect 2588 3436 2596 3444
rect 2125 1368 2131 1772
rect 2317 1708 2323 2152
rect 2381 1768 2387 2132
rect 2445 2108 2451 3052
rect 2493 1948 2499 2732
rect 2557 1788 2563 3132
rect 2653 2768 2659 3112
rect 2749 3108 2755 3432
rect 2781 3368 2787 3732
rect 2813 3728 2819 4672
rect 2861 4388 2867 5112
rect 2829 3768 2835 4132
rect 2844 4123 2852 4124
rect 2844 4117 2856 4123
rect 2844 4116 2852 4117
rect 2877 3988 2883 4592
rect 2877 3704 2883 3712
rect 2876 3696 2884 3704
rect 2013 908 2019 1232
rect 1978 606 1984 614
rect 2125 348 2131 1352
rect 2141 1088 2147 1692
rect 2300 1503 2308 1504
rect 2296 1497 2308 1503
rect 2300 1496 2308 1497
rect 2701 1328 2707 2812
rect 2749 2548 2755 3092
rect 2781 1508 2787 2972
rect 2797 2868 2803 3292
rect 2829 2964 2835 3052
rect 2828 2956 2836 2964
rect 2813 2828 2819 2852
rect 2893 2048 2899 3072
rect 2909 2988 2915 5072
rect 2925 4388 2931 4792
rect 2925 4164 2931 4172
rect 2941 4168 2947 4812
rect 2986 4806 2992 4814
rect 2986 4406 2992 4414
rect 3165 4388 3171 4912
rect 2924 4156 2932 4164
rect 2986 4006 2992 4014
rect 2940 3783 2948 3784
rect 2940 3777 2952 3783
rect 2940 3776 2948 3777
rect 2956 3736 2964 3744
rect 2957 3728 2963 3736
rect 2986 3606 2992 3614
rect 2925 1528 2931 3472
rect 2941 3208 2947 3232
rect 3069 3228 3075 3392
rect 3101 3308 3107 3732
rect 3133 3528 3139 4092
rect 3181 3788 3187 4732
rect 3485 4688 3491 5252
rect 3308 4576 3316 4584
rect 3292 4536 3300 4544
rect 3229 4328 3235 4392
rect 3293 4368 3299 4536
rect 3309 4488 3315 4576
rect 3229 4108 3235 4312
rect 3229 3548 3235 4092
rect 3277 3588 3283 4092
rect 3325 4088 3331 4472
rect 3341 3588 3347 4212
rect 3357 4164 3363 4172
rect 3356 4156 3364 4164
rect 3421 3968 3427 4092
rect 3356 3696 3364 3704
rect 2986 3206 2992 3214
rect 3036 3083 3044 3084
rect 3032 3077 3044 3083
rect 3036 3076 3044 3077
rect 2941 1988 2947 3072
rect 3085 3064 3091 3072
rect 3084 3056 3092 3064
rect 2988 2903 2996 2904
rect 2988 2897 3000 2903
rect 2988 2896 2996 2897
rect 2986 2806 2992 2814
rect 3037 2508 3043 2832
rect 2986 2406 2992 2414
rect 2986 2006 2992 2014
rect 2986 1606 2992 1614
rect 2733 1168 2739 1472
rect 2380 1036 2388 1044
rect 2381 988 2387 1036
rect 2156 523 2164 524
rect 2152 517 2164 523
rect 2156 516 2164 517
rect 2621 503 2627 512
rect 2616 497 2627 503
rect 2204 483 2212 484
rect 2204 477 2216 483
rect 2204 476 2212 477
rect 2540 436 2548 444
rect 2541 408 2547 436
rect 1978 206 1984 214
rect 2701 28 2707 892
rect 2781 348 2787 1492
rect 2986 1206 2992 1214
rect 2861 348 2867 1132
rect 3005 984 3011 1192
rect 3004 976 3012 984
rect 2986 806 2992 814
rect 3037 728 3043 2092
rect 3101 1968 3107 3292
rect 3133 1608 3139 3452
rect 3229 2904 3235 3032
rect 3228 2896 3236 2904
rect 3213 2068 3219 2232
rect 3325 1408 3331 3532
rect 3357 1588 3363 3696
rect 3421 3448 3427 3952
rect 3533 3904 3539 3932
rect 3532 3896 3540 3904
rect 3453 3688 3459 3872
rect 3437 3464 3443 3492
rect 3436 3456 3444 3464
rect 3373 2148 3379 3232
rect 3549 2928 3555 4172
rect 3549 2528 3555 2912
rect 3597 2828 3603 3772
rect 3645 3208 3651 5112
rect 3661 4308 3667 4832
rect 3693 4808 3699 5392
rect 3853 5128 3859 5232
rect 3677 4168 3683 4352
rect 3725 4328 3731 4892
rect 3757 4288 3763 5072
rect 4026 5006 4032 5014
rect 3916 4976 3924 4984
rect 3901 4768 3907 4832
rect 3917 4748 3923 4976
rect 3933 4744 3939 4832
rect 3932 4736 3940 4744
rect 3789 4548 3795 4672
rect 3821 4488 3827 4652
rect 3901 4468 3907 4732
rect 3949 4704 3955 4712
rect 3948 4696 3956 4704
rect 4061 4628 4067 5152
rect 4026 4606 4032 4614
rect 4012 4516 4020 4524
rect 4013 4508 4019 4516
rect 3724 4283 3732 4284
rect 3724 4277 3736 4283
rect 3724 4276 3732 4277
rect 3788 4103 3796 4104
rect 3788 4097 3800 4103
rect 3788 4096 3796 4097
rect 3725 3908 3731 4092
rect 3501 1688 3507 1812
rect 3149 1084 3155 1112
rect 3148 1076 3156 1084
rect 2986 406 2992 414
rect 3005 208 3011 652
rect 3037 548 3043 672
rect 3052 563 3060 564
rect 3052 557 3064 563
rect 3052 556 3060 557
rect 3245 464 3251 472
rect 3244 456 3252 464
rect 3437 348 3443 1632
rect 3453 28 3459 1372
rect 3485 564 3491 932
rect 3484 556 3492 564
rect 3468 303 3476 304
rect 3468 297 3480 303
rect 3468 296 3476 297
rect 3469 188 3475 296
rect 3501 188 3507 1352
rect 3517 628 3523 1632
rect 3549 1548 3555 2512
rect 3565 1148 3571 2392
rect 3661 1748 3667 3292
rect 3693 1728 3699 3892
rect 3725 3528 3731 3892
rect 3757 2048 3763 2372
rect 3773 2268 3779 2832
rect 3821 2768 3827 3312
rect 3837 2968 3843 4072
rect 3853 3548 3859 4292
rect 3901 4288 3907 4452
rect 3885 3728 3891 4172
rect 3901 3548 3907 4252
rect 3917 3928 3923 4312
rect 3933 3968 3939 4472
rect 3996 4436 4004 4444
rect 3997 4428 4003 4436
rect 3949 4104 3955 4132
rect 3948 4096 3956 4104
rect 3981 4048 3987 4332
rect 4026 4206 4032 4214
rect 4026 3806 4032 3814
rect 4044 3796 4052 3804
rect 3933 3588 3939 3792
rect 4045 3788 4051 3796
rect 4028 3776 4036 3784
rect 4029 3748 4035 3776
rect 4093 3708 4099 4912
rect 4189 3788 4195 3912
rect 4026 3406 4032 3414
rect 4205 3228 4211 4472
rect 4221 4108 4227 5492
rect 6074 5406 6080 5414
rect 4300 4736 4308 4744
rect 4316 4736 4324 4744
rect 4301 4728 4307 4736
rect 4285 4688 4291 4712
rect 4317 4688 4323 4736
rect 4333 4644 4339 4712
rect 4332 4636 4340 4644
rect 4349 4128 4355 4892
rect 4413 4768 4419 5292
rect 5050 5206 5056 5214
rect 4412 4736 4420 4744
rect 4444 4736 4452 4744
rect 4413 4728 4419 4736
rect 4445 4708 4451 4736
rect 4573 4368 4579 4912
rect 4621 4564 4627 4572
rect 4620 4556 4628 4564
rect 4700 3903 4708 3904
rect 4696 3897 4708 3903
rect 4700 3896 4708 3897
rect 4717 3548 4723 3892
rect 4765 3568 4771 3792
rect 4829 3728 4835 4512
rect 4861 4168 4867 4632
rect 4877 4568 4883 5112
rect 5661 5068 5667 5132
rect 4524 3523 4532 3524
rect 4524 3517 4536 3523
rect 4524 3516 4532 3517
rect 4765 3348 4771 3552
rect 4861 3508 4867 3852
rect 4893 3804 4899 5052
rect 5050 4806 5056 4814
rect 5116 4736 5124 4744
rect 5085 4724 5091 4732
rect 5084 4716 5092 4724
rect 4941 4684 4947 4712
rect 5117 4708 5123 4736
rect 4940 4676 4948 4684
rect 4988 4683 4996 4684
rect 4984 4677 4996 4683
rect 4988 4676 4996 4677
rect 5421 4644 5427 4712
rect 5453 4704 5459 4712
rect 5452 4696 5460 4704
rect 5420 4636 5428 4644
rect 5325 4624 5331 4632
rect 5324 4616 5332 4624
rect 5533 4548 5539 4732
rect 5181 4504 5187 4512
rect 5180 4496 5188 4504
rect 5050 4406 5056 4414
rect 5050 4006 5056 4014
rect 4892 3796 4900 3804
rect 4893 3788 4899 3796
rect 5050 3606 5056 3614
rect 4908 3516 4916 3524
rect 4909 3468 4915 3516
rect 4893 3408 4899 3452
rect 4316 3343 4324 3344
rect 4312 3337 4324 3343
rect 4316 3336 4324 3337
rect 5069 3228 5075 3792
rect 5197 3648 5203 4512
rect 5661 4308 5667 5052
rect 5932 4903 5940 4904
rect 5932 4897 5944 4903
rect 5932 4896 5940 4897
rect 5693 4684 5699 4732
rect 5692 4676 5700 4684
rect 5772 4623 5780 4624
rect 5768 4617 5780 4623
rect 5772 4616 5780 4617
rect 5196 3516 5204 3524
rect 5197 3508 5203 3516
rect 5341 3504 5347 3512
rect 5340 3496 5348 3504
rect 5645 3488 5651 4092
rect 5725 3728 5731 3772
rect 5388 3463 5396 3464
rect 5384 3457 5396 3463
rect 5388 3456 5396 3457
rect 5437 3248 5443 3452
rect 5050 3206 5056 3214
rect 5069 3168 5075 3212
rect 4077 3084 4083 3092
rect 4076 3076 4084 3084
rect 4026 3006 4032 3014
rect 4026 2606 4032 2614
rect 4026 2206 4032 2214
rect 3757 1908 3763 2032
rect 3901 1808 3907 2092
rect 3612 1523 3620 1524
rect 3608 1517 3620 1523
rect 3612 1516 3620 1517
rect 3565 1108 3571 1132
rect 3581 708 3587 1092
rect 3597 668 3603 812
rect 3677 128 3683 1532
rect 3773 1168 3779 1412
rect 3868 1343 3876 1344
rect 3868 1337 3880 1343
rect 3868 1336 3876 1337
rect 3708 1123 3716 1124
rect 3708 1117 3720 1123
rect 3708 1116 3716 1117
rect 3693 1104 3699 1112
rect 3789 1104 3795 1112
rect 3692 1096 3700 1104
rect 3788 1096 3796 1104
rect 3724 703 3732 704
rect 3724 697 3736 703
rect 3724 696 3732 697
rect 3692 663 3700 664
rect 3692 657 3704 663
rect 3692 656 3700 657
rect 3757 568 3763 1052
rect 3773 688 3779 1072
rect 3805 1008 3811 1332
rect 3821 708 3827 1232
rect 3837 988 3843 1272
rect 3853 1084 3859 1092
rect 3852 1076 3860 1084
rect 3836 696 3844 704
rect 3837 688 3843 696
rect 3772 556 3780 564
rect 3773 548 3779 556
rect 3869 448 3875 1292
rect 3885 668 3891 1232
rect 3917 748 3923 1552
rect 3949 1528 3955 1812
rect 3965 1408 3971 2012
rect 4205 1928 4211 2432
rect 4685 2208 4691 2292
rect 4026 1806 4032 1814
rect 4189 1748 4195 1792
rect 4348 1703 4356 1704
rect 4348 1697 4360 1703
rect 4348 1696 4356 1697
rect 4429 1668 4435 1752
rect 4765 1524 4771 1912
rect 4764 1516 4772 1524
rect 3981 1128 3987 1512
rect 4765 1508 4771 1516
rect 4701 1468 4707 1492
rect 4220 1456 4228 1464
rect 4026 1406 4032 1414
rect 4221 1408 4227 1456
rect 4236 1436 4244 1444
rect 4237 1388 4243 1436
rect 4156 1376 4164 1384
rect 4157 1348 4163 1376
rect 4333 1344 4339 1352
rect 4332 1336 4340 1344
rect 4764 1336 4772 1344
rect 4461 1268 4467 1312
rect 4765 1308 4771 1336
rect 4797 1308 4803 2112
rect 4829 2008 4835 2812
rect 5050 2806 5056 2814
rect 5084 2503 5092 2504
rect 5080 2497 5092 2503
rect 5084 2496 5092 2497
rect 5050 2406 5056 2414
rect 4813 1744 4819 1752
rect 4812 1736 4820 1744
rect 4829 1608 4835 1912
rect 4026 1006 4032 1014
rect 4125 704 4131 712
rect 4124 696 4132 704
rect 3981 684 3987 692
rect 3980 676 3988 684
rect 4026 606 4032 614
rect 3900 536 3908 544
rect 3901 508 3907 536
rect 4026 206 4032 214
rect 3741 128 3747 152
rect 4141 108 4147 952
rect 4173 584 4179 732
rect 4205 724 4211 852
rect 4204 716 4212 724
rect 4172 576 4180 584
rect 4253 508 4259 1032
rect 4333 28 4339 1072
rect 4349 648 4355 1052
rect 4716 956 4724 964
rect 4717 928 4723 956
rect 4397 308 4403 912
rect 4413 444 4419 852
rect 4748 636 4756 644
rect 4749 588 4755 636
rect 4797 508 4803 1292
rect 4861 948 4867 1892
rect 4989 1328 4995 2272
rect 5050 2006 5056 2014
rect 5036 1703 5044 1704
rect 5036 1697 5048 1703
rect 5036 1696 5044 1697
rect 5050 1606 5056 1614
rect 5101 1428 5107 3092
rect 5293 1988 5299 3212
rect 5324 3036 5332 3044
rect 5325 3008 5331 3036
rect 5853 3008 5859 4612
rect 5932 4503 5940 4504
rect 5928 4497 5940 4503
rect 5932 4496 5940 4497
rect 5917 3908 5923 4212
rect 5933 4128 5939 4496
rect 5981 4308 5987 5112
rect 6029 4888 6035 5272
rect 6074 5006 6080 5014
rect 6236 4743 6244 4744
rect 6232 4737 6244 4743
rect 6236 4736 6244 4737
rect 6092 4636 6100 4644
rect 6074 4606 6080 4614
rect 6093 4608 6099 4636
rect 6093 4508 6099 4592
rect 6237 4584 6243 4592
rect 6236 4576 6244 4584
rect 5997 3908 6003 4492
rect 6074 4206 6080 4214
rect 5869 3668 5875 3812
rect 5917 3768 5923 3872
rect 5965 3764 5971 3832
rect 5964 3756 5972 3764
rect 5308 2976 5316 2984
rect 5309 2968 5315 2976
rect 5340 2903 5348 2904
rect 5336 2897 5348 2903
rect 5340 2896 5348 2897
rect 5709 2448 5715 2612
rect 5837 2228 5843 2812
rect 5869 2668 5875 3652
rect 5917 2908 5923 3752
rect 5997 3708 6003 3892
rect 5997 3048 6003 3692
rect 6013 2708 6019 3972
rect 6029 3308 6035 3992
rect 6074 3806 6080 3814
rect 6093 3668 6099 4492
rect 6140 4323 6148 4324
rect 6136 4317 6148 4323
rect 6140 4316 6148 4317
rect 6156 3843 6164 3844
rect 6152 3837 6164 3843
rect 6156 3836 6164 3837
rect 6173 3768 6179 4352
rect 6253 3888 6259 4652
rect 6317 4308 6323 4892
rect 6074 3406 6080 3414
rect 6074 3006 6080 3014
rect 5293 1948 5299 1972
rect 5581 1528 5587 2152
rect 5597 1788 5603 2172
rect 5708 1343 5716 1344
rect 5704 1337 5716 1343
rect 5708 1336 5716 1337
rect 5532 1323 5540 1324
rect 5528 1317 5540 1323
rect 5532 1316 5540 1317
rect 5050 1206 5056 1214
rect 5629 968 5635 1132
rect 5837 928 5843 2212
rect 5853 2108 5859 2472
rect 5869 2308 5875 2652
rect 6013 2128 6019 2692
rect 6074 2606 6080 2614
rect 6074 2206 6080 2214
rect 5050 806 5056 814
rect 4893 528 4899 592
rect 4412 436 4420 444
rect 5050 406 5056 414
rect 5469 288 5475 672
rect 5885 228 5891 1312
rect 5965 128 5971 1892
rect 5981 748 5987 2092
rect 6013 1728 6019 2112
rect 6029 1828 6035 1852
rect 6074 1806 6080 1814
rect 6013 1328 6019 1712
rect 6028 1476 6036 1484
rect 6029 1428 6035 1476
rect 6109 1448 6115 2672
rect 6221 2268 6227 3412
rect 6237 2688 6243 3832
rect 6316 3783 6324 3784
rect 6312 3777 6324 3783
rect 6316 3776 6324 3777
rect 6349 3428 6355 4912
rect 6397 4868 6403 4892
rect 6413 4568 6419 4592
rect 6413 3828 6419 4552
rect 6429 4448 6435 4792
rect 6445 4028 6451 4932
rect 6476 4656 6484 4664
rect 6477 4648 6483 4656
rect 6476 4443 6484 4444
rect 6472 4437 6484 4443
rect 6476 4436 6484 4437
rect 6461 3148 6467 4152
rect 6493 4148 6499 5052
rect 6604 4683 6612 4684
rect 6600 4677 6612 4683
rect 6604 4676 6612 4677
rect 6541 4664 6547 4672
rect 6540 4656 6548 4664
rect 6621 4348 6627 5292
rect 6637 4568 6643 4732
rect 6653 4548 6659 4652
rect 6669 4528 6675 4672
rect 6685 4568 6691 4932
rect 6781 4904 6787 4912
rect 6780 4896 6788 4904
rect 6748 4663 6756 4664
rect 6744 4657 6756 4663
rect 6748 4656 6756 4657
rect 6717 4564 6723 4572
rect 6716 4556 6724 4564
rect 6765 4544 6771 4572
rect 6764 4536 6772 4544
rect 6556 3723 6564 3724
rect 6552 3717 6564 3723
rect 6556 3716 6564 3717
rect 6637 3488 6643 3852
rect 6669 3188 6675 4332
rect 6733 3188 6739 4212
rect 6269 2604 6275 2612
rect 6268 2596 6276 2604
rect 6349 2388 6355 2772
rect 6300 2303 6308 2304
rect 6296 2297 6308 2303
rect 6300 2296 6308 2297
rect 6253 1628 6259 2292
rect 6074 1406 6080 1414
rect 5997 1304 6003 1312
rect 5996 1296 6004 1304
rect 6013 1108 6019 1312
rect 6173 1028 6179 1052
rect 6074 1006 6080 1014
rect 6189 988 6195 1052
rect 6029 628 6035 832
rect 6074 606 6080 614
rect 6189 468 6195 972
rect 6236 963 6244 964
rect 6232 957 6244 963
rect 6236 956 6244 957
rect 6269 768 6275 1032
rect 6285 808 6291 1812
rect 6301 1348 6307 2172
rect 6397 2108 6403 2712
rect 6461 1728 6467 3132
rect 6540 3103 6548 3104
rect 6536 3097 6548 3103
rect 6540 3096 6548 3097
rect 6493 2268 6499 2672
rect 6493 1808 6499 1892
rect 6525 1548 6531 2512
rect 6557 1728 6563 2812
rect 6588 2383 6596 2384
rect 6584 2377 6596 2383
rect 6588 2376 6596 2377
rect 6380 1463 6388 1464
rect 6376 1457 6388 1463
rect 6380 1456 6388 1457
rect 6349 1368 6355 1452
rect 6396 1383 6404 1384
rect 6392 1377 6404 1383
rect 6396 1376 6404 1377
rect 6525 1348 6531 1532
rect 6573 1444 6579 1512
rect 6636 1483 6644 1484
rect 6632 1477 6644 1483
rect 6636 1476 6644 1477
rect 6572 1436 6580 1444
rect 6669 1248 6675 2912
rect 6781 2508 6787 4896
rect 6845 3788 6851 4052
rect 6909 3788 6915 4392
rect 6925 4148 6931 5252
rect 7082 5206 7088 5214
rect 7082 4806 7088 4814
rect 6940 4723 6948 4724
rect 6940 4717 6952 4723
rect 6940 4716 6948 4717
rect 6957 3488 6963 3872
rect 6973 3528 6979 3852
rect 6989 3828 6995 4512
rect 7021 4288 7027 4712
rect 7082 4406 7088 4414
rect 7082 4006 7088 4014
rect 7082 3606 7088 3614
rect 7165 3588 7171 4172
rect 6829 2188 6835 2652
rect 6925 2208 6931 3172
rect 6957 3008 6963 3472
rect 6988 3463 6996 3464
rect 6984 3457 6996 3463
rect 6988 3456 6996 3457
rect 7181 3308 7187 3652
rect 6989 2248 6995 3272
rect 7082 3206 7088 3214
rect 7293 3148 7299 3272
rect 7082 2806 7088 2814
rect 7082 2406 7088 2414
rect 7165 2148 7171 2472
rect 7082 2006 7088 2014
rect 6700 1903 6708 1904
rect 6696 1897 6708 1903
rect 6700 1896 6708 1897
rect 6988 1883 6996 1884
rect 6988 1877 7000 1883
rect 6988 1876 6996 1877
rect 6301 868 6307 932
rect 6397 924 6403 932
rect 6396 916 6404 924
rect 6620 903 6628 904
rect 6616 897 6628 903
rect 6620 896 6628 897
rect 6685 328 6691 1332
rect 6701 788 6707 1052
rect 6749 748 6755 1072
rect 6765 728 6771 1712
rect 6797 1328 6803 1532
rect 6813 1348 6819 1732
rect 6941 1464 6947 1472
rect 6940 1456 6948 1464
rect 6893 1308 6899 1372
rect 7021 1328 7027 1872
rect 7082 1606 7088 1614
rect 7180 1496 7188 1504
rect 7181 1488 7187 1496
rect 7260 1483 7268 1484
rect 7256 1477 7268 1483
rect 7260 1476 7268 1477
rect 7389 1468 7395 4712
rect 7405 1688 7411 4632
rect 7421 2268 7427 4692
rect 7453 2708 7459 2912
rect 7485 1728 7491 4452
rect 7532 3883 7540 3884
rect 7528 3877 7540 3883
rect 7532 3876 7540 3877
rect 7629 2328 7635 2592
rect 7645 2168 7651 2532
rect 7693 2128 7699 5472
rect 7709 4708 7715 5172
rect 7420 1503 7428 1504
rect 7416 1497 7428 1503
rect 7420 1496 7428 1497
rect 6988 1323 6996 1324
rect 6984 1317 6996 1323
rect 6988 1316 6996 1317
rect 6796 923 6804 924
rect 6792 917 6804 923
rect 6796 916 6804 917
rect 6813 908 6819 1032
rect 6876 983 6884 984
rect 6872 977 6884 983
rect 6876 976 6884 977
rect 6733 348 6739 672
rect 7021 668 7027 1312
rect 7082 1206 7088 1214
rect 7229 1168 7235 1272
rect 7485 1028 7491 1712
rect 7517 1468 7523 1512
rect 7082 806 7088 814
rect 7485 688 7491 1012
rect 7517 928 7523 1352
rect 7725 1068 7731 5432
rect 7757 3248 7763 3912
rect 7741 1468 7747 1772
rect 7773 1728 7779 5272
rect 7789 708 7795 5312
rect 7805 5128 7811 5452
rect 7805 4828 7811 5112
rect 7805 2408 7811 4812
rect 7821 3144 7827 4992
rect 7837 4568 7843 5072
rect 7852 4936 7860 4944
rect 7853 4928 7859 4936
rect 7884 4943 7892 4944
rect 7884 4937 7896 4943
rect 7884 4936 7892 4937
rect 7820 3136 7828 3144
rect 7821 1068 7827 3112
rect 7837 1168 7843 3012
rect 7853 1328 7859 2392
rect 7837 728 7843 1092
rect 7853 928 7859 1212
rect 7869 1048 7875 4932
rect 7884 3136 7892 3144
rect 6908 643 6916 644
rect 6904 637 6916 643
rect 6908 636 6916 637
rect 7082 406 7088 414
rect 7885 328 7891 3136
rect 7901 1288 7907 2112
rect 7917 1068 7923 5052
rect 7933 1308 7939 5032
rect 8061 3108 8067 3132
rect 6074 206 6080 214
rect 954 6 960 14
rect 2986 6 2992 14
rect 5050 6 5056 14
rect 7082 6 7088 14
use FILL  FILL_BUFX4_315
timestamp 1515882711
transform -1 0 24 0 1 5410
box 0 0 16 200
use BUFX4  BUFX4_315
timestamp 1515882711
transform -1 0 88 0 1 5410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_251
timestamp 1515882711
transform -1 0 104 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_251
timestamp 1515882711
transform -1 0 296 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_263
timestamp 1515882711
transform 1 0 296 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_263
timestamp 1515882711
transform 1 0 312 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_197
timestamp 1515882711
transform -1 0 520 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_197
timestamp 1515882711
transform -1 0 712 0 1 5410
box 0 0 192 200
use FILL  FILL_AOI21X1_30
timestamp 1515882711
transform 1 0 712 0 1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_30
timestamp 1515882711
transform 1 0 728 0 1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_106
timestamp 1515882711
transform 1 0 792 0 1 5410
box 0 0 48 200
use NOR2X1  NOR2X1_124
timestamp 1515882711
transform -1 0 888 0 1 5410
box 0 0 48 200
use FILL  FILL_AOI21X1_48
timestamp 1515882711
transform -1 0 904 0 1 5410
box 0 0 16 200
use FILL  FILL_27_0_0
timestamp 1515882711
transform -1 0 920 0 1 5410
box 0 0 16 200
use FILL  FILL_27_0_1
timestamp 1515882711
transform -1 0 936 0 1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_48
timestamp 1515882711
transform -1 0 1000 0 1 5410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_215
timestamp 1515882711
transform 1 0 1000 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_215
timestamp 1515882711
transform 1 0 1016 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_184
timestamp 1515882711
transform 1 0 1208 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_184
timestamp 1515882711
transform 1 0 1224 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_228
timestamp 1515882711
transform -1 0 1432 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_228
timestamp 1515882711
transform -1 0 1624 0 1 5410
box 0 0 192 200
use FILL  FILL_NAND2X1_152
timestamp 1515882711
transform -1 0 1640 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_152
timestamp 1515882711
transform -1 0 1688 0 1 5410
box 0 0 48 200
use FILL  FILL_INVX2_3
timestamp 1515882711
transform 1 0 1688 0 1 5410
box 0 0 16 200
use INVX2  INVX2_3
timestamp 1515882711
transform 1 0 1704 0 1 5410
box 0 0 32 200
use FILL  FILL_BUFX4_278
timestamp 1515882711
transform -1 0 1752 0 1 5410
box 0 0 16 200
use BUFX4  BUFX4_278
timestamp 1515882711
transform -1 0 1816 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_154
timestamp 1515882711
transform 1 0 1816 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_154
timestamp 1515882711
transform 1 0 1832 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_3
timestamp 1515882711
transform -1 0 1896 0 1 5410
box 0 0 16 200
use FILL  FILL_27_1_0
timestamp 1515882711
transform -1 0 1912 0 1 5410
box 0 0 16 200
use FILL  FILL_27_1_1
timestamp 1515882711
transform -1 0 1928 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1515882711
transform -1 0 2120 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_448
timestamp 1515882711
transform -1 0 2184 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_381
timestamp 1515882711
transform 1 0 2184 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_381
timestamp 1515882711
transform 1 0 2200 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_7
timestamp 1515882711
transform 1 0 2248 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1515882711
transform 1 0 2264 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_449
timestamp 1515882711
transform -1 0 2520 0 1 5410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_4
timestamp 1515882711
transform 1 0 2520 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1515882711
transform 1 0 2536 0 1 5410
box 0 0 192 200
use FILL  FILL_INVX1_22
timestamp 1515882711
transform 1 0 2728 0 1 5410
box 0 0 16 200
use INVX1  INVX1_22
timestamp 1515882711
transform 1 0 2744 0 1 5410
box 0 0 32 200
use FILL  FILL_BUFX2_31
timestamp 1515882711
transform 1 0 2776 0 1 5410
box 0 0 16 200
use BUFX2  BUFX2_31
timestamp 1515882711
transform 1 0 2792 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_40
timestamp 1515882711
transform 1 0 2840 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_39
timestamp 1515882711
transform 1 0 2888 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_56
timestamp 1515882711
transform 1 0 2936 0 1 5410
box 0 0 48 200
use FILL  FILL_27_2_0
timestamp 1515882711
transform 1 0 2984 0 1 5410
box 0 0 16 200
use FILL  FILL_27_2_1
timestamp 1515882711
transform 1 0 3000 0 1 5410
box 0 0 16 200
use BUFX2  BUFX2_58
timestamp 1515882711
transform 1 0 3016 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_55
timestamp 1515882711
transform 1 0 3064 0 1 5410
box 0 0 48 200
use FILL  FILL_BUFX2_16
timestamp 1515882711
transform -1 0 3128 0 1 5410
box 0 0 16 200
use BUFX2  BUFX2_16
timestamp 1515882711
transform -1 0 3176 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_60
timestamp 1515882711
transform 1 0 3176 0 1 5410
box 0 0 48 200
use FILL  FILL_BUFX2_28
timestamp 1515882711
transform 1 0 3224 0 1 5410
box 0 0 16 200
use BUFX2  BUFX2_28
timestamp 1515882711
transform 1 0 3240 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_37
timestamp 1515882711
transform 1 0 3288 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_337
timestamp 1515882711
transform -1 0 3352 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_337
timestamp 1515882711
transform -1 0 3544 0 1 5410
box 0 0 192 200
use FILL  FILL_NAND2X1_363
timestamp 1515882711
transform 1 0 3544 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_363
timestamp 1515882711
transform 1 0 3560 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_430
timestamp 1515882711
transform -1 0 3672 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_429
timestamp 1515882711
transform 1 0 3672 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_362
timestamp 1515882711
transform -1 0 3752 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_362
timestamp 1515882711
transform -1 0 3800 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_336
timestamp 1515882711
transform -1 0 3816 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_336
timestamp 1515882711
transform -1 0 4008 0 1 5410
box 0 0 192 200
use FILL  FILL_27_3_0
timestamp 1515882711
transform 1 0 4008 0 1 5410
box 0 0 16 200
use FILL  FILL_27_3_1
timestamp 1515882711
transform 1 0 4024 0 1 5410
box 0 0 16 200
use FILL  FILL_BUFX2_7
timestamp 1515882711
transform 1 0 4040 0 1 5410
box 0 0 16 200
use BUFX2  BUFX2_7
timestamp 1515882711
transform 1 0 4056 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_47
timestamp 1515882711
transform 1 0 4104 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_36
timestamp 1515882711
transform 1 0 4152 0 1 5410
box 0 0 48 200
use BUFX2  BUFX2_61
timestamp 1515882711
transform 1 0 4200 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_39
timestamp 1515882711
transform -1 0 4264 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_39
timestamp 1515882711
transform -1 0 4456 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_109
timestamp 1515882711
transform 1 0 4456 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_109
timestamp 1515882711
transform 1 0 4472 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_109
timestamp 1515882711
transform 1 0 4664 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_93
timestamp 1515882711
transform 1 0 4728 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_93
timestamp 1515882711
transform 1 0 4744 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_331
timestamp 1515882711
transform 1 0 4792 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_331
timestamp 1515882711
transform 1 0 4808 0 1 5410
box 0 0 192 200
use FILL  FILL_27_4_0
timestamp 1515882711
transform 1 0 5000 0 1 5410
box 0 0 16 200
use FILL  FILL_27_4_1
timestamp 1515882711
transform 1 0 5016 0 1 5410
box 0 0 16 200
use OAI21X1  OAI21X1_335
timestamp 1515882711
transform 1 0 5032 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_390
timestamp 1515882711
transform -1 0 5112 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_390
timestamp 1515882711
transform -1 0 5160 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_357
timestamp 1515882711
transform 1 0 5160 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_395
timestamp 1515882711
transform -1 0 5240 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_395
timestamp 1515882711
transform -1 0 5288 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_2
timestamp 1515882711
transform 1 0 5288 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1515882711
transform 1 0 5304 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_97
timestamp 1515882711
transform -1 0 5512 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_97
timestamp 1515882711
transform -1 0 5704 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_108
timestamp 1515882711
transform -1 0 5720 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_108
timestamp 1515882711
transform -1 0 5912 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_108
timestamp 1515882711
transform -1 0 5976 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_91
timestamp 1515882711
transform 1 0 5976 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_73
timestamp 1515882711
transform -1 0 6056 0 1 5410
box 0 0 16 200
use FILL  FILL_27_5_0
timestamp 1515882711
transform -1 0 6072 0 1 5410
box 0 0 16 200
use FILL  FILL_27_5_1
timestamp 1515882711
transform -1 0 6088 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_73
timestamp 1515882711
transform -1 0 6136 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_91
timestamp 1515882711
transform -1 0 6152 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_91
timestamp 1515882711
transform -1 0 6344 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_287
timestamp 1515882711
transform -1 0 6360 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_287
timestamp 1515882711
transform -1 0 6552 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_103
timestamp 1515882711
transform 1 0 6552 0 1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_85
timestamp 1515882711
transform -1 0 6632 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_85
timestamp 1515882711
transform -1 0 6680 0 1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_103
timestamp 1515882711
transform 1 0 6680 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_103
timestamp 1515882711
transform 1 0 6696 0 1 5410
box 0 0 192 200
use FILL  FILL_NAND2X1_104
timestamp 1515882711
transform 1 0 6888 0 1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_104
timestamp 1515882711
transform 1 0 6904 0 1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_121
timestamp 1515882711
transform -1 0 7016 0 1 5410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_121
timestamp 1515882711
transform -1 0 7032 0 1 5410
box 0 0 16 200
use FILL  FILL_27_6_0
timestamp 1515882711
transform -1 0 7048 0 1 5410
box 0 0 16 200
use FILL  FILL_27_6_1
timestamp 1515882711
transform -1 0 7064 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_121
timestamp 1515882711
transform -1 0 7256 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_325
timestamp 1515882711
transform 1 0 7256 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_325
timestamp 1515882711
transform 1 0 7272 0 1 5410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_322
timestamp 1515882711
transform -1 0 7480 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_322
timestamp 1515882711
transform -1 0 7672 0 1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_150
timestamp 1515882711
transform 1 0 7672 0 1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_130
timestamp 1515882711
transform -1 0 7800 0 1 5410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_130
timestamp 1515882711
transform 1 0 7800 0 1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_130
timestamp 1515882711
transform 1 0 7816 0 1 5410
box 0 0 192 200
use FILL  FILL_28_1
timestamp 1515882711
transform 1 0 8008 0 1 5410
box 0 0 16 200
use FILL  FILL_28_2
timestamp 1515882711
transform 1 0 8024 0 1 5410
box 0 0 16 200
use FILL  FILL_28_3
timestamp 1515882711
transform 1 0 8040 0 1 5410
box 0 0 16 200
use FILL  FILL_DFFPOSX1_255
timestamp 1515882711
transform -1 0 24 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_255
timestamp 1515882711
transform -1 0 216 0 -1 5410
box 0 0 192 200
use NOR2X1  NOR2X1_75
timestamp 1515882711
transform 1 0 216 0 -1 5410
box 0 0 48 200
use FILL  FILL_AOI21X1_63
timestamp 1515882711
transform -1 0 280 0 -1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_63
timestamp 1515882711
transform -1 0 344 0 -1 5410
box 0 0 64 200
use FILL  FILL_AOI21X1_34
timestamp 1515882711
transform 1 0 344 0 -1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_34
timestamp 1515882711
transform 1 0 360 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_35
timestamp 1515882711
transform 1 0 424 0 -1 5410
box 0 0 48 200
use FILL  FILL_AOI21X1_7
timestamp 1515882711
transform 1 0 472 0 -1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_7
timestamp 1515882711
transform 1 0 488 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_83
timestamp 1515882711
transform -1 0 600 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_219
timestamp 1515882711
transform 1 0 600 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_219
timestamp 1515882711
transform 1 0 616 0 -1 5410
box 0 0 192 200
use FILL  FILL_AOI21X1_52
timestamp 1515882711
transform 1 0 808 0 -1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_52
timestamp 1515882711
transform 1 0 824 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_128
timestamp 1515882711
transform 1 0 888 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_0_0
timestamp 1515882711
transform -1 0 952 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_0_1
timestamp 1515882711
transform -1 0 968 0 -1 5410
box 0 0 16 200
use FILL  FILL_INVX2_30
timestamp 1515882711
transform -1 0 984 0 -1 5410
box 0 0 16 200
use INVX2  INVX2_30
timestamp 1515882711
transform -1 0 1016 0 -1 5410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_181
timestamp 1515882711
transform -1 0 1032 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_181
timestamp 1515882711
transform -1 0 1224 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_164
timestamp 1515882711
transform 1 0 1224 0 -1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_149
timestamp 1515882711
transform -1 0 1304 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_149
timestamp 1515882711
transform -1 0 1352 0 -1 5410
box 0 0 48 200
use FILL  FILL_INVX2_33
timestamp 1515882711
transform 1 0 1352 0 -1 5410
box 0 0 16 200
use INVX2  INVX2_33
timestamp 1515882711
transform 1 0 1368 0 -1 5410
box 0 0 32 200
use FILL  FILL_BUFX4_308
timestamp 1515882711
transform -1 0 1416 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_308
timestamp 1515882711
transform -1 0 1480 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_167
timestamp 1515882711
transform 1 0 1480 0 -1 5410
box 0 0 64 200
use FILL  FILL_AOI21X1_60
timestamp 1515882711
transform 1 0 1544 0 -1 5410
box 0 0 16 200
use AOI21X1  AOI21X1_60
timestamp 1515882711
transform 1 0 1560 0 -1 5410
box 0 0 64 200
use NOR2X1  NOR2X1_136
timestamp 1515882711
transform -1 0 1672 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_186
timestamp 1515882711
transform -1 0 1688 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_186
timestamp 1515882711
transform -1 0 1880 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_170
timestamp 1515882711
transform -1 0 1944 0 -1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_148
timestamp 1515882711
transform -1 0 1960 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_1_0
timestamp 1515882711
transform -1 0 1976 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_1_1
timestamp 1515882711
transform -1 0 1992 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_148
timestamp 1515882711
transform -1 0 2040 0 -1 5410
box 0 0 48 200
use FILL  FILL_BUFX4_294
timestamp 1515882711
transform 1 0 2040 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_294
timestamp 1515882711
transform 1 0 2056 0 -1 5410
box 0 0 64 200
use FILL  FILL_INVX1_17
timestamp 1515882711
transform 1 0 2120 0 -1 5410
box 0 0 16 200
use INVX1  INVX1_17
timestamp 1515882711
transform 1 0 2136 0 -1 5410
box 0 0 32 200
use FILL  FILL_NAND2X1_380
timestamp 1515882711
transform -1 0 2184 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_380
timestamp 1515882711
transform -1 0 2232 0 -1 5410
box 0 0 48 200
use FILL  FILL_NAND2X1_384
timestamp 1515882711
transform 1 0 2232 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_384
timestamp 1515882711
transform 1 0 2248 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_452
timestamp 1515882711
transform -1 0 2360 0 -1 5410
box 0 0 64 200
use FILL  FILL_INVX1_39
timestamp 1515882711
transform -1 0 2376 0 -1 5410
box 0 0 16 200
use INVX1  INVX1_39
timestamp 1515882711
transform -1 0 2408 0 -1 5410
box 0 0 32 200
use FILL  FILL_BUFX4_231
timestamp 1515882711
transform -1 0 2424 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_231
timestamp 1515882711
transform -1 0 2488 0 -1 5410
box 0 0 64 200
use FILL  FILL_INVX8_13
timestamp 1515882711
transform 1 0 2488 0 -1 5410
box 0 0 16 200
use INVX8  INVX8_13
timestamp 1515882711
transform 1 0 2504 0 -1 5410
box 0 0 80 200
use FILL  FILL_BUFX4_224
timestamp 1515882711
transform 1 0 2584 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_224
timestamp 1515882711
transform 1 0 2600 0 -1 5410
box 0 0 64 200
use FILL  FILL_INVX8_7
timestamp 1515882711
transform 1 0 2664 0 -1 5410
box 0 0 16 200
use INVX8  INVX8_7
timestamp 1515882711
transform 1 0 2680 0 -1 5410
box 0 0 80 200
use FILL  FILL_NAND2X1_245
timestamp 1515882711
transform -1 0 2776 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_245
timestamp 1515882711
transform -1 0 2824 0 -1 5410
box 0 0 48 200
use FILL  FILL_BUFX2_30
timestamp 1515882711
transform 1 0 2824 0 -1 5410
box 0 0 16 200
use BUFX2  BUFX2_30
timestamp 1515882711
transform 1 0 2840 0 -1 5410
box 0 0 48 200
use FILL  FILL_BUFX2_19
timestamp 1515882711
transform 1 0 2888 0 -1 5410
box 0 0 16 200
use BUFX2  BUFX2_19
timestamp 1515882711
transform 1 0 2904 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_343
timestamp 1515882711
transform 1 0 2952 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_2_0
timestamp 1515882711
transform 1 0 2968 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_2_1
timestamp 1515882711
transform 1 0 2984 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_343
timestamp 1515882711
transform 1 0 3000 0 -1 5410
box 0 0 192 200
use FILL  FILL_BUFX2_21
timestamp 1515882711
transform -1 0 3208 0 -1 5410
box 0 0 16 200
use BUFX2  BUFX2_21
timestamp 1515882711
transform -1 0 3256 0 -1 5410
box 0 0 48 200
use FILL  FILL_NAND2X1_222
timestamp 1515882711
transform 1 0 3256 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_222
timestamp 1515882711
transform 1 0 3272 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_241
timestamp 1515882711
transform -1 0 3384 0 -1 5410
box 0 0 64 200
use FILL  FILL_INVX1_24
timestamp 1515882711
transform -1 0 3400 0 -1 5410
box 0 0 16 200
use INVX1  INVX1_24
timestamp 1515882711
transform -1 0 3432 0 -1 5410
box 0 0 32 200
use OAI21X1  OAI21X1_436
timestamp 1515882711
transform -1 0 3496 0 -1 5410
box 0 0 64 200
use FILL  FILL_INVX1_51
timestamp 1515882711
transform -1 0 3512 0 -1 5410
box 0 0 16 200
use INVX1  INVX1_51
timestamp 1515882711
transform -1 0 3544 0 -1 5410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_38
timestamp 1515882711
transform -1 0 3560 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_38
timestamp 1515882711
transform -1 0 3752 0 -1 5410
box 0 0 192 200
use FILL  FILL_NAND2X1_215
timestamp 1515882711
transform 1 0 3752 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_215
timestamp 1515882711
transform 1 0 3768 0 -1 5410
box 0 0 48 200
use FILL  FILL_BUFX2_13
timestamp 1515882711
transform 1 0 3816 0 -1 5410
box 0 0 16 200
use BUFX2  BUFX2_13
timestamp 1515882711
transform 1 0 3832 0 -1 5410
box 0 0 48 200
use BUFX2  BUFX2_52
timestamp 1515882711
transform 1 0 3880 0 -1 5410
box 0 0 48 200
use FILL  FILL_NAND2X1_23
timestamp 1515882711
transform 1 0 3928 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_23
timestamp 1515882711
transform 1 0 3944 0 -1 5410
box 0 0 48 200
use FILL  FILL_26_3_0
timestamp 1515882711
transform -1 0 4008 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_3_1
timestamp 1515882711
transform -1 0 4024 0 -1 5410
box 0 0 16 200
use OAI21X1  OAI21X1_44
timestamp 1515882711
transform -1 0 4088 0 -1 5410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_44
timestamp 1515882711
transform -1 0 4104 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_44
timestamp 1515882711
transform -1 0 4296 0 -1 5410
box 0 0 192 200
use FILL  FILL_NAND2X1_18
timestamp 1515882711
transform 1 0 4296 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_18
timestamp 1515882711
transform 1 0 4312 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_39
timestamp 1515882711
transform -1 0 4424 0 -1 5410
box 0 0 64 200
use FILL  FILL_BUFX2_27
timestamp 1515882711
transform -1 0 4440 0 -1 5410
box 0 0 16 200
use BUFX2  BUFX2_27
timestamp 1515882711
transform -1 0 4488 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_319
timestamp 1515882711
transform -1 0 4504 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_319
timestamp 1515882711
transform -1 0 4696 0 -1 5410
box 0 0 192 200
use FILL  FILL_MUX2X1_5
timestamp 1515882711
transform 1 0 4696 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_5
timestamp 1515882711
transform 1 0 4712 0 -1 5410
box 0 0 96 200
use NAND2X1  NAND2X1_408
timestamp 1515882711
transform 1 0 4808 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_95
timestamp 1515882711
transform 1 0 4856 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_95
timestamp 1515882711
transform 1 0 4872 0 -1 5410
box 0 0 192 200
use FILL  FILL_26_4_0
timestamp 1515882711
transform -1 0 5080 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_4_1
timestamp 1515882711
transform -1 0 5096 0 -1 5410
box 0 0 16 200
use FILL  FILL_MUX2X1_16
timestamp 1515882711
transform -1 0 5112 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_16
timestamp 1515882711
transform -1 0 5208 0 -1 5410
box 0 0 96 200
use FILL  FILL_NAND2X1_77
timestamp 1515882711
transform 1 0 5208 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_77
timestamp 1515882711
transform 1 0 5224 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_95
timestamp 1515882711
transform -1 0 5336 0 -1 5410
box 0 0 64 200
use FILL  FILL_MUX2X1_22
timestamp 1515882711
transform -1 0 5352 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_22
timestamp 1515882711
transform -1 0 5448 0 -1 5410
box 0 0 96 200
use FILL  FILL_NAND2X1_80
timestamp 1515882711
transform 1 0 5448 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_80
timestamp 1515882711
transform 1 0 5464 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_97
timestamp 1515882711
transform -1 0 5576 0 -1 5410
box 0 0 64 200
use FILL  FILL_BUFX4_321
timestamp 1515882711
transform -1 0 5592 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_321
timestamp 1515882711
transform -1 0 5656 0 -1 5410
box 0 0 64 200
use FILL  FILL_BUFX4_279
timestamp 1515882711
transform 1 0 5656 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_279
timestamp 1515882711
transform 1 0 5672 0 -1 5410
box 0 0 64 200
use FILL  FILL_BUFX4_282
timestamp 1515882711
transform -1 0 5752 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_282
timestamp 1515882711
transform -1 0 5816 0 -1 5410
box 0 0 64 200
use FILL  FILL_BUFX4_235
timestamp 1515882711
transform -1 0 5832 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_235
timestamp 1515882711
transform -1 0 5896 0 -1 5410
box 0 0 64 200
use FILL  FILL_NAND2X1_92
timestamp 1515882711
transform -1 0 5912 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_92
timestamp 1515882711
transform -1 0 5960 0 -1 5410
box 0 0 48 200
use FILL  FILL_BUFX4_318
timestamp 1515882711
transform -1 0 5976 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_318
timestamp 1515882711
transform -1 0 6040 0 -1 5410
box 0 0 64 200
use FILL  FILL_MUX2X1_3
timestamp 1515882711
transform 1 0 6040 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_5_0
timestamp 1515882711
transform 1 0 6056 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_5_1
timestamp 1515882711
transform 1 0 6072 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_3
timestamp 1515882711
transform 1 0 6088 0 -1 5410
box 0 0 96 200
use FILL  FILL_NAND2X1_346
timestamp 1515882711
transform 1 0 6184 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_346
timestamp 1515882711
transform 1 0 6200 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_290
timestamp 1515882711
transform -1 0 6312 0 -1 5410
box 0 0 64 200
use FILL  FILL_BUFX4_81
timestamp 1515882711
transform 1 0 6312 0 -1 5410
box 0 0 16 200
use BUFX4  BUFX4_81
timestamp 1515882711
transform 1 0 6328 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_412
timestamp 1515882711
transform 1 0 6392 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_401
timestamp 1515882711
transform -1 0 6504 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_57
timestamp 1515882711
transform 1 0 6504 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_57
timestamp 1515882711
transform 1 0 6520 0 -1 5410
box 0 0 192 200
use FILL  FILL_MUX2X1_39
timestamp 1515882711
transform -1 0 6728 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_39
timestamp 1515882711
transform -1 0 6824 0 -1 5410
box 0 0 96 200
use FILL  FILL_MUX2X1_38
timestamp 1515882711
transform -1 0 6840 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_38
timestamp 1515882711
transform -1 0 6936 0 -1 5410
box 0 0 96 200
use OAI21X1  OAI21X1_474
timestamp 1515882711
transform 1 0 6936 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_419
timestamp 1515882711
transform -1 0 7048 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_330
timestamp 1515882711
transform -1 0 7064 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_6_0
timestamp 1515882711
transform -1 0 7080 0 -1 5410
box 0 0 16 200
use FILL  FILL_26_6_1
timestamp 1515882711
transform -1 0 7096 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_330
timestamp 1515882711
transform -1 0 7288 0 -1 5410
box 0 0 192 200
use OAI21X1  OAI21X1_468
timestamp 1515882711
transform 1 0 7288 0 -1 5410
box 0 0 64 200
use OAI21X1  OAI21X1_465
timestamp 1515882711
transform 1 0 7352 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_411
timestamp 1515882711
transform -1 0 7464 0 -1 5410
box 0 0 48 200
use FILL  FILL_MUX2X1_14
timestamp 1515882711
transform 1 0 7464 0 -1 5410
box 0 0 16 200
use MUX2X1  MUX2X1_14
timestamp 1515882711
transform 1 0 7480 0 -1 5410
box 0 0 96 200
use FILL  FILL_NAND2X1_115
timestamp 1515882711
transform 1 0 7576 0 -1 5410
box 0 0 16 200
use NAND2X1  NAND2X1_115
timestamp 1515882711
transform 1 0 7592 0 -1 5410
box 0 0 48 200
use OAI21X1  OAI21X1_483
timestamp 1515882711
transform 1 0 7640 0 -1 5410
box 0 0 64 200
use NAND2X1  NAND2X1_430
timestamp 1515882711
transform -1 0 7752 0 -1 5410
box 0 0 48 200
use NAND2X1  NAND2X1_433
timestamp 1515882711
transform 1 0 7752 0 -1 5410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_304
timestamp 1515882711
transform -1 0 7816 0 -1 5410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_304
timestamp 1515882711
transform -1 0 8008 0 -1 5410
box 0 0 192 200
use FILL  FILL_27_1
timestamp 1515882711
transform -1 0 8024 0 -1 5410
box 0 0 16 200
use FILL  FILL_27_2
timestamp 1515882711
transform -1 0 8040 0 -1 5410
box 0 0 16 200
use FILL  FILL_27_3
timestamp 1515882711
transform -1 0 8056 0 -1 5410
box 0 0 16 200
use FILL  FILL_DFFPOSX1_162
timestamp 1515882711
transform 1 0 8 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_162
timestamp 1515882711
transform 1 0 24 0 1 5010
box 0 0 192 200
use NOR2X1  NOR2X1_88
timestamp 1515882711
transform -1 0 264 0 1 5010
box 0 0 48 200
use FILL  FILL_AOI21X1_13
timestamp 1515882711
transform -1 0 280 0 1 5010
box 0 0 16 200
use AOI21X1  AOI21X1_13
timestamp 1515882711
transform -1 0 344 0 1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_174
timestamp 1515882711
transform 1 0 344 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_174
timestamp 1515882711
transform 1 0 360 0 1 5010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_234
timestamp 1515882711
transform 1 0 552 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_234
timestamp 1515882711
transform 1 0 568 0 1 5010
box 0 0 192 200
use FILL  FILL_INVX2_15
timestamp 1515882711
transform 1 0 760 0 1 5010
box 0 0 16 200
use INVX2  INVX2_15
timestamp 1515882711
transform 1 0 776 0 1 5010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_209
timestamp 1515882711
transform -1 0 824 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_209
timestamp 1515882711
transform -1 0 1016 0 1 5010
box 0 0 192 200
use FILL  FILL_25_0_0
timestamp 1515882711
transform 1 0 1016 0 1 5010
box 0 0 16 200
use FILL  FILL_25_0_1
timestamp 1515882711
transform 1 0 1032 0 1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_182
timestamp 1515882711
transform 1 0 1048 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_166
timestamp 1515882711
transform -1 0 1128 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_166
timestamp 1515882711
transform -1 0 1176 0 1 5010
box 0 0 48 200
use FILL  FILL_INVX2_14
timestamp 1515882711
transform -1 0 1192 0 1 5010
box 0 0 16 200
use INVX2  INVX2_14
timestamp 1515882711
transform -1 0 1224 0 1 5010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_233
timestamp 1515882711
transform -1 0 1240 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_233
timestamp 1515882711
transform -1 0 1432 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_181
timestamp 1515882711
transform 1 0 1432 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_165
timestamp 1515882711
transform -1 0 1512 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_165
timestamp 1515882711
transform -1 0 1560 0 1 5010
box 0 0 48 200
use FILL  FILL_INVX2_29
timestamp 1515882711
transform -1 0 1576 0 1 5010
box 0 0 16 200
use INVX2  INVX2_29
timestamp 1515882711
transform -1 0 1608 0 1 5010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_180
timestamp 1515882711
transform -1 0 1624 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_180
timestamp 1515882711
transform -1 0 1816 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_163
timestamp 1515882711
transform 1 0 1816 0 1 5010
box 0 0 64 200
use FILL  FILL_INVX8_14
timestamp 1515882711
transform -1 0 1896 0 1 5010
box 0 0 16 200
use INVX8  INVX8_14
timestamp 1515882711
transform -1 0 1976 0 1 5010
box 0 0 80 200
use FILL  FILL_25_1_0
timestamp 1515882711
transform 1 0 1976 0 1 5010
box 0 0 16 200
use FILL  FILL_25_1_1
timestamp 1515882711
transform 1 0 1992 0 1 5010
box 0 0 16 200
use FILL  FILL_NAND2X1_170
timestamp 1515882711
transform 1 0 2008 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_170
timestamp 1515882711
transform 1 0 2024 0 1 5010
box 0 0 48 200
use FILL  FILL_BUFX4_312
timestamp 1515882711
transform 1 0 2072 0 1 5010
box 0 0 16 200
use BUFX4  BUFX4_312
timestamp 1515882711
transform 1 0 2088 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_177
timestamp 1515882711
transform -1 0 2168 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_177
timestamp 1515882711
transform -1 0 2216 0 1 5010
box 0 0 48 200
use FILL  FILL_NAND2X1_160
timestamp 1515882711
transform 1 0 2216 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_160
timestamp 1515882711
transform 1 0 2232 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_25
timestamp 1515882711
transform 1 0 2280 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_3
timestamp 1515882711
transform -1 0 2360 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_3
timestamp 1515882711
transform -1 0 2408 0 1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_273
timestamp 1515882711
transform 1 0 2408 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_273
timestamp 1515882711
transform 1 0 2424 0 1 5010
box 0 0 192 200
use FILL  FILL_NAND2X1_392
timestamp 1515882711
transform 1 0 2616 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_392
timestamp 1515882711
transform 1 0 2632 0 1 5010
box 0 0 48 200
use FILL  FILL_BUFX4_78
timestamp 1515882711
transform -1 0 2696 0 1 5010
box 0 0 16 200
use BUFX4  BUFX4_78
timestamp 1515882711
transform -1 0 2760 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_270
timestamp 1515882711
transform -1 0 2824 0 1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_230
timestamp 1515882711
transform 1 0 2824 0 1 5010
box 0 0 16 200
use BUFX4  BUFX4_230
timestamp 1515882711
transform 1 0 2840 0 1 5010
box 0 0 64 200
use FILL  FILL_BUFX2_17
timestamp 1515882711
transform 1 0 2904 0 1 5010
box 0 0 16 200
use BUFX2  BUFX2_17
timestamp 1515882711
transform 1 0 2920 0 1 5010
box 0 0 48 200
use FILL  FILL_NAND2X1_221
timestamp 1515882711
transform -1 0 2984 0 1 5010
box 0 0 16 200
use FILL  FILL_25_2_0
timestamp 1515882711
transform -1 0 3000 0 1 5010
box 0 0 16 200
use FILL  FILL_25_2_1
timestamp 1515882711
transform -1 0 3016 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_221
timestamp 1515882711
transform -1 0 3064 0 1 5010
box 0 0 48 200
use FILL  FILL_NAND2X1_214
timestamp 1515882711
transform -1 0 3080 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_214
timestamp 1515882711
transform -1 0 3128 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_42
timestamp 1515882711
transform 1 0 3128 0 1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_270
timestamp 1515882711
transform 1 0 3176 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_270
timestamp 1515882711
transform 1 0 3192 0 1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_450
timestamp 1515882711
transform 1 0 3384 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_21
timestamp 1515882711
transform -1 0 3496 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_240
timestamp 1515882711
transform -1 0 3560 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_262
timestamp 1515882711
transform 1 0 3560 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_262
timestamp 1515882711
transform 1 0 3576 0 1 5010
box 0 0 48 200
use FILL  FILL_NAND2X1_369
timestamp 1515882711
transform -1 0 3640 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_369
timestamp 1515882711
transform -1 0 3688 0 1 5010
box 0 0 48 200
use FILL  FILL_BUFX2_14
timestamp 1515882711
transform 1 0 3688 0 1 5010
box 0 0 16 200
use BUFX2  BUFX2_14
timestamp 1515882711
transform 1 0 3704 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_53
timestamp 1515882711
transform 1 0 3752 0 1 5010
box 0 0 48 200
use BUFX2  BUFX2_63
timestamp 1515882711
transform 1 0 3800 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_231
timestamp 1515882711
transform -1 0 3912 0 1 5010
box 0 0 64 200
use FILL  FILL_INVX1_18
timestamp 1515882711
transform -1 0 3928 0 1 5010
box 0 0 16 200
use INVX1  INVX1_18
timestamp 1515882711
transform -1 0 3960 0 1 5010
box 0 0 32 200
use FILL  FILL_NAND2X1_17
timestamp 1515882711
transform 1 0 3960 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_17
timestamp 1515882711
transform 1 0 3976 0 1 5010
box 0 0 48 200
use FILL  FILL_25_3_0
timestamp 1515882711
transform -1 0 4040 0 1 5010
box 0 0 16 200
use FILL  FILL_25_3_1
timestamp 1515882711
transform -1 0 4056 0 1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_38
timestamp 1515882711
transform -1 0 4120 0 1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_73
timestamp 1515882711
transform -1 0 4136 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_73
timestamp 1515882711
transform -1 0 4328 0 1 5010
box 0 0 192 200
use FILL  FILL_NAND2X1_54
timestamp 1515882711
transform 1 0 4328 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_54
timestamp 1515882711
transform 1 0 4344 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_73
timestamp 1515882711
transform -1 0 4456 0 1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_246
timestamp 1515882711
transform 1 0 4456 0 1 5010
box 0 0 16 200
use BUFX4  BUFX4_246
timestamp 1515882711
transform 1 0 4472 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_80
timestamp 1515882711
transform 1 0 4536 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_61
timestamp 1515882711
transform -1 0 4616 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_61
timestamp 1515882711
transform -1 0 4664 0 1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_80
timestamp 1515882711
transform -1 0 4680 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_80
timestamp 1515882711
transform -1 0 4872 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_463
timestamp 1515882711
transform -1 0 4936 0 1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_114
timestamp 1515882711
transform -1 0 5000 0 1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_114
timestamp 1515882711
transform -1 0 5016 0 1 5010
box 0 0 16 200
use FILL  FILL_25_4_0
timestamp 1515882711
transform -1 0 5032 0 1 5010
box 0 0 16 200
use FILL  FILL_25_4_1
timestamp 1515882711
transform -1 0 5048 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_114
timestamp 1515882711
transform -1 0 5240 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_92
timestamp 1515882711
transform -1 0 5304 0 1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_92
timestamp 1515882711
transform 1 0 5304 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_92
timestamp 1515882711
transform 1 0 5320 0 1 5010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_128
timestamp 1515882711
transform -1 0 5528 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_128
timestamp 1515882711
transform -1 0 5720 0 1 5010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_318
timestamp 1515882711
transform 1 0 5720 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_318
timestamp 1515882711
transform 1 0 5736 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_462
timestamp 1515882711
transform 1 0 5928 0 1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_407
timestamp 1515882711
transform -1 0 6040 0 1 5010
box 0 0 48 200
use FILL  FILL_MUX2X1_2
timestamp 1515882711
transform 1 0 6040 0 1 5010
box 0 0 16 200
use FILL  FILL_25_5_0
timestamp 1515882711
transform 1 0 6056 0 1 5010
box 0 0 16 200
use FILL  FILL_25_5_1
timestamp 1515882711
transform 1 0 6072 0 1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_2
timestamp 1515882711
transform 1 0 6088 0 1 5010
box 0 0 96 200
use FILL  FILL_DFFPOSX1_302
timestamp 1515882711
transform 1 0 6184 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_302
timestamp 1515882711
transform 1 0 6200 0 1 5010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_94
timestamp 1515882711
transform 1 0 6392 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_94
timestamp 1515882711
transform 1 0 6408 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_323
timestamp 1515882711
transform 1 0 6600 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_379
timestamp 1515882711
transform -1 0 6680 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_379
timestamp 1515882711
transform -1 0 6728 0 1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_320
timestamp 1515882711
transform -1 0 6744 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_320
timestamp 1515882711
transform -1 0 6936 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_139
timestamp 1515882711
transform -1 0 7000 0 1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_139
timestamp 1515882711
transform -1 0 7016 0 1 5010
box 0 0 16 200
use FILL  FILL_25_6_0
timestamp 1515882711
transform -1 0 7032 0 1 5010
box 0 0 16 200
use FILL  FILL_25_6_1
timestamp 1515882711
transform -1 0 7048 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_139
timestamp 1515882711
transform -1 0 7240 0 1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_116
timestamp 1515882711
transform 1 0 7240 0 1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_98
timestamp 1515882711
transform -1 0 7320 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_98
timestamp 1515882711
transform -1 0 7368 0 1 5010
box 0 0 48 200
use NAND2X1  NAND2X1_414
timestamp 1515882711
transform -1 0 7416 0 1 5010
box 0 0 48 200
use FILL  FILL_MUX2X1_11
timestamp 1515882711
transform -1 0 7432 0 1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_11
timestamp 1515882711
transform -1 0 7528 0 1 5010
box 0 0 96 200
use FILL  FILL_NAND2X1_95
timestamp 1515882711
transform -1 0 7544 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_95
timestamp 1515882711
transform -1 0 7592 0 1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_111
timestamp 1515882711
transform -1 0 7656 0 1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_111
timestamp 1515882711
transform -1 0 7672 0 1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_111
timestamp 1515882711
transform -1 0 7864 0 1 5010
box 0 0 192 200
use FILL  FILL_NAND2X1_128
timestamp 1515882711
transform -1 0 7880 0 1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_128
timestamp 1515882711
transform -1 0 7928 0 1 5010
box 0 0 48 200
use FILL  FILL_BUFX4_297
timestamp 1515882711
transform 1 0 7928 0 1 5010
box 0 0 16 200
use BUFX4  BUFX4_297
timestamp 1515882711
transform 1 0 7944 0 1 5010
box 0 0 64 200
use FILL  FILL_26_1
timestamp 1515882711
transform 1 0 8008 0 1 5010
box 0 0 16 200
use FILL  FILL_26_2
timestamp 1515882711
transform 1 0 8024 0 1 5010
box 0 0 16 200
use FILL  FILL_26_3
timestamp 1515882711
transform 1 0 8040 0 1 5010
box 0 0 16 200
use FILL  FILL_BUFX4_10
timestamp 1515882711
transform -1 0 24 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_10
timestamp 1515882711
transform -1 0 88 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_296
timestamp 1515882711
transform -1 0 152 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_252
timestamp 1515882711
transform 1 0 152 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_153
timestamp 1515882711
transform -1 0 280 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_108
timestamp 1515882711
transform -1 0 344 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_109
timestamp 1515882711
transform -1 0 408 0 -1 5010
box 0 0 64 200
use FILL  FILL_AOI21X1_25
timestamp 1515882711
transform 1 0 408 0 -1 5010
box 0 0 16 200
use AOI21X1  AOI21X1_25
timestamp 1515882711
transform 1 0 424 0 -1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_101
timestamp 1515882711
transform -1 0 536 0 -1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_202
timestamp 1515882711
transform 1 0 536 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_202
timestamp 1515882711
transform 1 0 552 0 -1 5010
box 0 0 192 200
use FILL  FILL_AOI21X1_35
timestamp 1515882711
transform 1 0 744 0 -1 5010
box 0 0 16 200
use AOI21X1  AOI21X1_35
timestamp 1515882711
transform 1 0 760 0 -1 5010
box 0 0 64 200
use NOR2X1  NOR2X1_110
timestamp 1515882711
transform 1 0 824 0 -1 5010
box 0 0 48 200
use NOR2X1  NOR2X1_118
timestamp 1515882711
transform 1 0 872 0 -1 5010
box 0 0 48 200
use FILL  FILL_AOI21X1_42
timestamp 1515882711
transform -1 0 936 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_0_0
timestamp 1515882711
transform -1 0 952 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_0_1
timestamp 1515882711
transform -1 0 968 0 -1 5010
box 0 0 16 200
use AOI21X1  AOI21X1_42
timestamp 1515882711
transform -1 0 1032 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_105
timestamp 1515882711
transform -1 0 1096 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_370
timestamp 1515882711
transform -1 0 1160 0 -1 5010
box 0 0 64 200
use NOR3X1  NOR3X1_30
timestamp 1515882711
transform -1 0 1288 0 -1 5010
box 0 0 128 200
use NAND3X1  NAND3X1_249
timestamp 1515882711
transform 1 0 1288 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_246
timestamp 1515882711
transform -1 0 1416 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_104
timestamp 1515882711
transform 1 0 1416 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_369
timestamp 1515882711
transform -1 0 1544 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_50
timestamp 1515882711
transform -1 0 1608 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_228
timestamp 1515882711
transform -1 0 1672 0 -1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_245
timestamp 1515882711
transform 1 0 1672 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_245
timestamp 1515882711
transform 1 0 1688 0 -1 5010
box 0 0 192 200
use FILL  FILL_INVX2_26
timestamp 1515882711
transform 1 0 1880 0 -1 5010
box 0 0 16 200
use INVX2  INVX2_26
timestamp 1515882711
transform 1 0 1896 0 -1 5010
box 0 0 32 200
use FILL  FILL_24_1_0
timestamp 1515882711
transform 1 0 1928 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_1_1
timestamp 1515882711
transform 1 0 1944 0 -1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_193
timestamp 1515882711
transform 1 0 1960 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_291
timestamp 1515882711
transform 1 0 2024 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_291
timestamp 1515882711
transform 1 0 2040 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_29
timestamp 1515882711
transform -1 0 2120 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_29
timestamp 1515882711
transform -1 0 2184 0 -1 5010
box 0 0 64 200
use FILL  FILL_INVX8_17
timestamp 1515882711
transform 1 0 2184 0 -1 5010
box 0 0 16 200
use INVX8  INVX8_17
timestamp 1515882711
transform 1 0 2200 0 -1 5010
box 0 0 80 200
use OAI21X1  OAI21X1_32
timestamp 1515882711
transform 1 0 2280 0 -1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_10
timestamp 1515882711
transform -1 0 2360 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_10
timestamp 1515882711
transform -1 0 2408 0 -1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_281
timestamp 1515882711
transform 1 0 2408 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_281
timestamp 1515882711
transform 1 0 2424 0 -1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_460
timestamp 1515882711
transform -1 0 2680 0 -1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_15
timestamp 1515882711
transform 1 0 2680 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1515882711
transform 1 0 2696 0 -1 5010
box 0 0 192 200
use FILL  FILL_INVX1_77
timestamp 1515882711
transform 1 0 2888 0 -1 5010
box 0 0 16 200
use INVX1  INVX1_77
timestamp 1515882711
transform 1 0 2904 0 -1 5010
box 0 0 32 200
use FILL  FILL_NAND2X1_299
timestamp 1515882711
transform -1 0 2952 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_299
timestamp 1515882711
transform -1 0 3000 0 -1 5010
box 0 0 48 200
use FILL  FILL_24_2_0
timestamp 1515882711
transform -1 0 3016 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_2_1
timestamp 1515882711
transform -1 0 3032 0 -1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_340
timestamp 1515882711
transform -1 0 3096 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX2_2
timestamp 1515882711
transform 1 0 3096 0 -1 5010
box 0 0 16 200
use BUFX2  BUFX2_2
timestamp 1515882711
transform 1 0 3112 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_230
timestamp 1515882711
transform -1 0 3224 0 -1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_269
timestamp 1515882711
transform -1 0 3240 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_269
timestamp 1515882711
transform -1 0 3432 0 -1 5010
box 0 0 192 200
use NAND2X1  NAND2X1_449
timestamp 1515882711
transform 1 0 3432 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_20
timestamp 1515882711
transform -1 0 3544 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_291
timestamp 1515882711
transform 1 0 3544 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_265
timestamp 1515882711
transform -1 0 3672 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_122
timestamp 1515882711
transform -1 0 3736 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX2_25
timestamp 1515882711
transform 1 0 3736 0 -1 5010
box 0 0 16 200
use BUFX2  BUFX2_25
timestamp 1515882711
transform 1 0 3752 0 -1 5010
box 0 0 48 200
use NAND3X1  NAND3X1_110
timestamp 1515882711
transform -1 0 3864 0 -1 5010
box 0 0 64 200
use NAND3X1  NAND3X1_254
timestamp 1515882711
transform 1 0 3864 0 -1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_216
timestamp 1515882711
transform 1 0 3928 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_216
timestamp 1515882711
transform 1 0 3944 0 -1 5010
box 0 0 48 200
use FILL  FILL_24_3_0
timestamp 1515882711
transform -1 0 4008 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_3_1
timestamp 1515882711
transform -1 0 4024 0 -1 5010
box 0 0 16 200
use OAI21X1  OAI21X1_233
timestamp 1515882711
transform -1 0 4088 0 -1 5010
box 0 0 64 200
use FILL  FILL_INVX1_19
timestamp 1515882711
transform -1 0 4104 0 -1 5010
box 0 0 16 200
use INVX1  INVX1_19
timestamp 1515882711
transform -1 0 4136 0 -1 5010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_113
timestamp 1515882711
transform 1 0 4136 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_113
timestamp 1515882711
transform 1 0 4152 0 -1 5010
box 0 0 192 200
use FILL  FILL_NAND2X1_146
timestamp 1515882711
transform 1 0 4344 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_146
timestamp 1515882711
transform 1 0 4360 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_113
timestamp 1515882711
transform -1 0 4472 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_52
timestamp 1515882711
transform 1 0 4472 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_52
timestamp 1515882711
transform 1 0 4488 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_31
timestamp 1515882711
transform 1 0 4552 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_31
timestamp 1515882711
transform 1 0 4568 0 -1 5010
box 0 0 64 200
use FILL  FILL_INVX1_52
timestamp 1515882711
transform 1 0 4632 0 -1 5010
box 0 0 16 200
use INVX1  INVX1_52
timestamp 1515882711
transform 1 0 4648 0 -1 5010
box 0 0 32 200
use FILL  FILL_NAND2X1_96
timestamp 1515882711
transform -1 0 4696 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_96
timestamp 1515882711
transform -1 0 4744 0 -1 5010
box 0 0 48 200
use FILL  FILL_MUX2X1_15
timestamp 1515882711
transform 1 0 4744 0 -1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_15
timestamp 1515882711
transform 1 0 4760 0 -1 5010
box 0 0 96 200
use OAI21X1  OAI21X1_466
timestamp 1515882711
transform 1 0 4856 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_412
timestamp 1515882711
transform -1 0 4968 0 -1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_323
timestamp 1515882711
transform -1 0 4984 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_4_0
timestamp 1515882711
transform -1 0 5000 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_4_1
timestamp 1515882711
transform -1 0 5016 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_323
timestamp 1515882711
transform -1 0 5208 0 -1 5010
box 0 0 192 200
use FILL  FILL_NAND2X1_74
timestamp 1515882711
transform 1 0 5208 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_74
timestamp 1515882711
transform 1 0 5224 0 -1 5010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_298
timestamp 1515882711
transform 1 0 5272 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_298
timestamp 1515882711
transform 1 0 5288 0 -1 5010
box 0 0 192 200
use FILL  FILL_MUX2X1_7
timestamp 1515882711
transform 1 0 5480 0 -1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_7
timestamp 1515882711
transform 1 0 5496 0 -1 5010
box 0 0 96 200
use OAI21X1  OAI21X1_301
timestamp 1515882711
transform 1 0 5592 0 -1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_111
timestamp 1515882711
transform 1 0 5656 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_111
timestamp 1515882711
transform 1 0 5672 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_128
timestamp 1515882711
transform -1 0 5784 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_87
timestamp 1515882711
transform -1 0 5800 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_87
timestamp 1515882711
transform -1 0 5864 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_121
timestamp 1515882711
transform -1 0 5880 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_121
timestamp 1515882711
transform -1 0 5944 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_131
timestamp 1515882711
transform 1 0 5944 0 -1 5010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_131
timestamp 1515882711
transform -1 0 6024 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_5_0
timestamp 1515882711
transform -1 0 6040 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_5_1
timestamp 1515882711
transform -1 0 6056 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_131
timestamp 1515882711
transform -1 0 6248 0 -1 5010
box 0 0 192 200
use OAI21X1  OAI21X1_480
timestamp 1515882711
transform 1 0 6248 0 -1 5010
box 0 0 64 200
use NAND2X1  NAND2X1_428
timestamp 1515882711
transform -1 0 6360 0 -1 5010
box 0 0 48 200
use FILL  FILL_BUFX4_267
timestamp 1515882711
transform 1 0 6360 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_267
timestamp 1515882711
transform 1 0 6376 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_94
timestamp 1515882711
transform 1 0 6440 0 -1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_76
timestamp 1515882711
transform -1 0 6520 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_76
timestamp 1515882711
transform -1 0 6568 0 -1 5010
box 0 0 48 200
use FILL  FILL_BUFX4_114
timestamp 1515882711
transform 1 0 6568 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_114
timestamp 1515882711
transform 1 0 6584 0 -1 5010
box 0 0 64 200
use FILL  FILL_MUX2X1_13
timestamp 1515882711
transform 1 0 6648 0 -1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_13
timestamp 1515882711
transform 1 0 6664 0 -1 5010
box 0 0 96 200
use FILL  FILL_BUFX4_122
timestamp 1515882711
transform 1 0 6760 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_122
timestamp 1515882711
transform 1 0 6776 0 -1 5010
box 0 0 64 200
use FILL  FILL_BUFX4_247
timestamp 1515882711
transform 1 0 6840 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_247
timestamp 1515882711
transform 1 0 6856 0 -1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_123
timestamp 1515882711
transform -1 0 6936 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_123
timestamp 1515882711
transform -1 0 6984 0 -1 5010
box 0 0 48 200
use FILL  FILL_BUFX4_249
timestamp 1515882711
transform 1 0 6984 0 -1 5010
box 0 0 16 200
use BUFX4  BUFX4_249
timestamp 1515882711
transform 1 0 7000 0 -1 5010
box 0 0 64 200
use FILL  FILL_MUX2X1_40
timestamp 1515882711
transform 1 0 7064 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_6_0
timestamp 1515882711
transform 1 0 7080 0 -1 5010
box 0 0 16 200
use FILL  FILL_24_6_1
timestamp 1515882711
transform 1 0 7096 0 -1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_40
timestamp 1515882711
transform 1 0 7112 0 -1 5010
box 0 0 96 200
use FILL  FILL_DFFPOSX1_116
timestamp 1515882711
transform 1 0 7208 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_116
timestamp 1515882711
transform 1 0 7224 0 -1 5010
box 0 0 192 200
use FILL  FILL_MUX2X1_21
timestamp 1515882711
transform -1 0 7432 0 -1 5010
box 0 0 16 200
use MUX2X1  MUX2X1_21
timestamp 1515882711
transform -1 0 7528 0 -1 5010
box 0 0 96 200
use FILL  FILL_INVX1_32
timestamp 1515882711
transform -1 0 7544 0 -1 5010
box 0 0 16 200
use INVX1  INVX1_32
timestamp 1515882711
transform -1 0 7576 0 -1 5010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_148
timestamp 1515882711
transform -1 0 7592 0 -1 5010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_148
timestamp 1515882711
transform -1 0 7784 0 -1 5010
box 0 0 192 200
use FILL  FILL_NAND2X1_136
timestamp 1515882711
transform -1 0 7800 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_136
timestamp 1515882711
transform -1 0 7848 0 -1 5010
box 0 0 48 200
use OAI21X1  OAI21X1_148
timestamp 1515882711
transform 1 0 7848 0 -1 5010
box 0 0 64 200
use OAI21X1  OAI21X1_149
timestamp 1515882711
transform 1 0 7912 0 -1 5010
box 0 0 64 200
use FILL  FILL_NAND2X1_133
timestamp 1515882711
transform 1 0 7976 0 -1 5010
box 0 0 16 200
use NAND2X1  NAND2X1_133
timestamp 1515882711
transform 1 0 7992 0 -1 5010
box 0 0 48 200
use FILL  FILL_25_1
timestamp 1515882711
transform -1 0 8056 0 -1 5010
box 0 0 16 200
use FILL  FILL_AOI21X1_17
timestamp 1515882711
transform 1 0 8 0 1 4610
box 0 0 16 200
use AOI21X1  AOI21X1_17
timestamp 1515882711
transform 1 0 24 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_93
timestamp 1515882711
transform -1 0 136 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_295
timestamp 1515882711
transform 1 0 136 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_152
timestamp 1515882711
transform 1 0 200 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_154
timestamp 1515882711
transform -1 0 328 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_107
timestamp 1515882711
transform -1 0 392 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_106
timestamp 1515882711
transform 1 0 392 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_253
timestamp 1515882711
transform 1 0 456 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_251
timestamp 1515882711
transform 1 0 520 0 1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_242
timestamp 1515882711
transform 1 0 584 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_242
timestamp 1515882711
transform 1 0 600 0 1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_292
timestamp 1515882711
transform -1 0 856 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_149
timestamp 1515882711
transform 1 0 856 0 1 4610
box 0 0 64 200
use FILL  FILL_23_0_0
timestamp 1515882711
transform -1 0 936 0 1 4610
box 0 0 16 200
use FILL  FILL_23_0_1
timestamp 1515882711
transform -1 0 952 0 1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_150
timestamp 1515882711
transform -1 0 1016 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_189
timestamp 1515882711
transform 1 0 1016 0 1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_174
timestamp 1515882711
transform -1 0 1096 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_174
timestamp 1515882711
transform -1 0 1144 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_387
timestamp 1515882711
transform -1 0 1208 0 1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_35
timestamp 1515882711
transform -1 0 1336 0 1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_386
timestamp 1515882711
transform -1 0 1400 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_227
timestamp 1515882711
transform -1 0 1464 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_265
timestamp 1515882711
transform -1 0 1528 0 1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_46
timestamp 1515882711
transform -1 0 1656 0 1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_226
timestamp 1515882711
transform -1 0 1720 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_49
timestamp 1515882711
transform 1 0 1720 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_336
timestamp 1515882711
transform -1 0 1848 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_337
timestamp 1515882711
transform -1 0 1912 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_418
timestamp 1515882711
transform -1 0 1976 0 1 4610
box 0 0 64 200
use FILL  FILL_23_1_0
timestamp 1515882711
transform 1 0 1976 0 1 4610
box 0 0 16 200
use FILL  FILL_23_1_1
timestamp 1515882711
transform 1 0 1992 0 1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_185
timestamp 1515882711
transform 1 0 2008 0 1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_238
timestamp 1515882711
transform 1 0 2072 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_238
timestamp 1515882711
transform 1 0 2088 0 1 4610
box 0 0 192 200
use FILL  FILL_NAND2X1_151
timestamp 1515882711
transform -1 0 2296 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_151
timestamp 1515882711
transform -1 0 2344 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_175
timestamp 1515882711
transform -1 0 2408 0 1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_212
timestamp 1515882711
transform -1 0 2424 0 1 4610
box 0 0 16 200
use BUFX4  BUFX4_212
timestamp 1515882711
transform -1 0 2488 0 1 4610
box 0 0 64 200
use FILL  FILL_INVX2_8
timestamp 1515882711
transform -1 0 2504 0 1 4610
box 0 0 16 200
use INVX2  INVX2_8
timestamp 1515882711
transform -1 0 2536 0 1 4610
box 0 0 32 200
use FILL  FILL_DFFPOSX1_192
timestamp 1515882711
transform -1 0 2552 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_192
timestamp 1515882711
transform -1 0 2744 0 1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_159
timestamp 1515882711
transform -1 0 2808 0 1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_388
timestamp 1515882711
transform 1 0 2808 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_388
timestamp 1515882711
transform 1 0 2824 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_302
timestamp 1515882711
transform -1 0 2936 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_456
timestamp 1515882711
transform -1 0 3000 0 1 4610
box 0 0 64 200
use FILL  FILL_23_2_0
timestamp 1515882711
transform 1 0 3000 0 1 4610
box 0 0 16 200
use FILL  FILL_23_2_1
timestamp 1515882711
transform 1 0 3016 0 1 4610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_11
timestamp 1515882711
transform 1 0 3032 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1515882711
transform 1 0 3048 0 1 4610
box 0 0 192 200
use FILL  FILL_INVX1_61
timestamp 1515882711
transform 1 0 3240 0 1 4610
box 0 0 16 200
use INVX1  INVX1_61
timestamp 1515882711
transform 1 0 3256 0 1 4610
box 0 0 32 200
use FILL  FILL_NAND2X1_276
timestamp 1515882711
transform -1 0 3304 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_276
timestamp 1515882711
transform -1 0 3352 0 1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_5
timestamp 1515882711
transform -1 0 3368 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_5
timestamp 1515882711
transform -1 0 3416 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_27
timestamp 1515882711
transform -1 0 3480 0 1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_275
timestamp 1515882711
transform 1 0 3480 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_275
timestamp 1515882711
transform 1 0 3496 0 1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_126
timestamp 1515882711
transform -1 0 3752 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_50
timestamp 1515882711
transform 1 0 3752 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_376
timestamp 1515882711
transform -1 0 3864 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_59
timestamp 1515882711
transform -1 0 3928 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_242
timestamp 1515882711
transform -1 0 3992 0 1 4610
box 0 0 64 200
use FILL  FILL_23_3_0
timestamp 1515882711
transform 1 0 3992 0 1 4610
box 0 0 16 200
use FILL  FILL_23_3_1
timestamp 1515882711
transform 1 0 4008 0 1 4610
box 0 0 16 200
use NOR2X1  NOR2X1_160
timestamp 1515882711
transform 1 0 4024 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_269
timestamp 1515882711
transform -1 0 4136 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_372
timestamp 1515882711
transform 1 0 4136 0 1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_237
timestamp 1515882711
transform -1 0 4264 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_232
timestamp 1515882711
transform 1 0 4264 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_157
timestamp 1515882711
transform -1 0 4376 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_258
timestamp 1515882711
transform -1 0 4440 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_48
timestamp 1515882711
transform -1 0 4488 0 1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_115
timestamp 1515882711
transform -1 0 4552 0 1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_53
timestamp 1515882711
transform 1 0 4552 0 1 4610
box 0 0 16 200
use BUFX4  BUFX4_53
timestamp 1515882711
transform 1 0 4568 0 1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_82
timestamp 1515882711
transform 1 0 4632 0 1 4610
box 0 0 16 200
use BUFX4  BUFX4_82
timestamp 1515882711
transform 1 0 4648 0 1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_20
timestamp 1515882711
transform -1 0 4728 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_20
timestamp 1515882711
transform -1 0 4920 0 1 4610
box 0 0 192 200
use NOR3X1  NOR3X1_8
timestamp 1515882711
transform -1 0 5048 0 1 4610
box 0 0 128 200
use FILL  FILL_23_4_0
timestamp 1515882711
transform -1 0 5064 0 1 4610
box 0 0 16 200
use FILL  FILL_23_4_1
timestamp 1515882711
transform -1 0 5080 0 1 4610
box 0 0 16 200
use NOR2X1  NOR2X1_4
timestamp 1515882711
transform -1 0 5128 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_5
timestamp 1515882711
transform -1 0 5176 0 1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_15
timestamp 1515882711
transform 1 0 5176 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_55
timestamp 1515882711
transform -1 0 5304 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_159
timestamp 1515882711
transform -1 0 5352 0 1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_12
timestamp 1515882711
transform -1 0 5432 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_49
timestamp 1515882711
transform -1 0 5480 0 1 4610
box 0 0 48 200
use FILL  FILL_MUX2X1_6
timestamp 1515882711
transform 1 0 5480 0 1 4610
box 0 0 16 200
use MUX2X1  MUX2X1_6
timestamp 1515882711
transform 1 0 5496 0 1 4610
box 0 0 96 200
use FILL  FILL_NAND2X1_357
timestamp 1515882711
transform 1 0 5592 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_357
timestamp 1515882711
transform 1 0 5608 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_269
timestamp 1515882711
transform 1 0 5656 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_388
timestamp 1515882711
transform 1 0 5720 0 1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_109
timestamp 1515882711
transform -1 0 5800 0 1 4610
box 0 0 16 200
use BUFX4  BUFX4_109
timestamp 1515882711
transform -1 0 5864 0 1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_80
timestamp 1515882711
transform 1 0 5864 0 1 4610
box 0 0 16 200
use BUFX4  BUFX4_80
timestamp 1515882711
transform 1 0 5880 0 1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_116
timestamp 1515882711
transform -1 0 5960 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_116
timestamp 1515882711
transform -1 0 6008 0 1 4610
box 0 0 48 200
use FILL  FILL_MUX2X1_17
timestamp 1515882711
transform 1 0 6008 0 1 4610
box 0 0 16 200
use FILL  FILL_23_5_0
timestamp 1515882711
transform 1 0 6024 0 1 4610
box 0 0 16 200
use FILL  FILL_23_5_1
timestamp 1515882711
transform 1 0 6040 0 1 4610
box 0 0 16 200
use MUX2X1  MUX2X1_17
timestamp 1515882711
transform 1 0 6056 0 1 4610
box 0 0 96 200
use OAI22X1  OAI22X1_11
timestamp 1515882711
transform 1 0 6152 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_47
timestamp 1515882711
transform -1 0 6280 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_154
timestamp 1515882711
transform 1 0 6280 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_371
timestamp 1515882711
transform -1 0 6392 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_156
timestamp 1515882711
transform 1 0 6392 0 1 4610
box 0 0 48 200
use NOR3X1  NOR3X1_47
timestamp 1515882711
transform 1 0 6440 0 1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_229
timestamp 1515882711
transform -1 0 6632 0 1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_165
timestamp 1515882711
transform -1 0 6680 0 1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_14
timestamp 1515882711
transform 1 0 6680 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_53
timestamp 1515882711
transform -1 0 6808 0 1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_27
timestamp 1515882711
transform -1 0 6856 0 1 4610
box 0 0 48 200
use OAI22X1  OAI22X1_7
timestamp 1515882711
transform -1 0 6936 0 1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_71
timestamp 1515882711
transform -1 0 6984 0 1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_384
timestamp 1515882711
transform 1 0 6984 0 1 4610
box 0 0 64 200
use FILL  FILL_23_6_0
timestamp 1515882711
transform -1 0 7064 0 1 4610
box 0 0 16 200
use FILL  FILL_23_6_1
timestamp 1515882711
transform -1 0 7080 0 1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_491
timestamp 1515882711
transform -1 0 7144 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_439
timestamp 1515882711
transform -1 0 7192 0 1 4610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_313
timestamp 1515882711
transform -1 0 7208 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_313
timestamp 1515882711
transform -1 0 7400 0 1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_125
timestamp 1515882711
transform -1 0 7464 0 1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_110
timestamp 1515882711
transform 1 0 7464 0 1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_110
timestamp 1515882711
transform 1 0 7480 0 1 4610
box 0 0 48 200
use FILL  FILL_MUX2X1_4
timestamp 1515882711
transform 1 0 7528 0 1 4610
box 0 0 16 200
use MUX2X1  MUX2X1_4
timestamp 1515882711
transform 1 0 7544 0 1 4610
box 0 0 96 200
use FILL  FILL_BUFX4_296
timestamp 1515882711
transform 1 0 7640 0 1 4610
box 0 0 16 200
use BUFX4  BUFX4_296
timestamp 1515882711
transform 1 0 7656 0 1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_479
timestamp 1515882711
transform 1 0 7720 0 1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_427
timestamp 1515882711
transform -1 0 7832 0 1 4610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_301
timestamp 1515882711
transform 1 0 7832 0 1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_301
timestamp 1515882711
transform 1 0 7848 0 1 4610
box 0 0 192 200
use FILL  FILL_24_1
timestamp 1515882711
transform 1 0 8040 0 1 4610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_166
timestamp 1515882711
transform 1 0 8 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_166
timestamp 1515882711
transform 1 0 24 0 -1 4610
box 0 0 192 200
use NAND3X1  NAND3X1_297
timestamp 1515882711
transform -1 0 280 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_294
timestamp 1515882711
transform 1 0 280 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_151
timestamp 1515882711
transform 1 0 344 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_250
timestamp 1515882711
transform 1 0 408 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_231
timestamp 1515882711
transform -1 0 536 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_232
timestamp 1515882711
transform -1 0 600 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_229
timestamp 1515882711
transform 1 0 600 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_51
timestamp 1515882711
transform 1 0 664 0 -1 4610
box 0 0 64 200
use FILL  FILL_INVX2_22
timestamp 1515882711
transform 1 0 728 0 -1 4610
box 0 0 16 200
use INVX2  INVX2_22
timestamp 1515882711
transform 1 0 744 0 -1 4610
box 0 0 32 200
use NOR3X1  NOR3X1_31
timestamp 1515882711
transform -1 0 904 0 -1 4610
box 0 0 128 200
use FILL  FILL_22_0_0
timestamp 1515882711
transform 1 0 904 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_0_1
timestamp 1515882711
transform 1 0 920 0 -1 4610
box 0 0 16 200
use OAI21X1  OAI21X1_374
timestamp 1515882711
transform 1 0 936 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_237
timestamp 1515882711
transform 1 0 1000 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_373
timestamp 1515882711
transform 1 0 1064 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_48
timestamp 1515882711
transform -1 0 1256 0 -1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_236
timestamp 1515882711
transform -1 0 1320 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_293
timestamp 1515882711
transform 1 0 1320 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_266
timestamp 1515882711
transform -1 0 1448 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_7
timestamp 1515882711
transform 1 0 1448 0 -1 4610
box 0 0 128 200
use NAND3X1  NAND3X1_227
timestamp 1515882711
transform -1 0 1640 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_22
timestamp 1515882711
transform -1 0 1768 0 -1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_417
timestamp 1515882711
transform -1 0 1832 0 -1 4610
box 0 0 64 200
use NOR3X1  NOR3X1_42
timestamp 1515882711
transform -1 0 1960 0 -1 4610
box 0 0 128 200
use FILL  FILL_22_1_0
timestamp 1515882711
transform -1 0 1976 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_1_1
timestamp 1515882711
transform -1 0 1992 0 -1 4610
box 0 0 16 200
use FILL  FILL_BUFX4_144
timestamp 1515882711
transform -1 0 2008 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_144
timestamp 1515882711
transform -1 0 2072 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_141
timestamp 1515882711
transform 1 0 2072 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_141
timestamp 1515882711
transform 1 0 2088 0 -1 4610
box 0 0 64 200
use FILL  FILL_INVX2_18
timestamp 1515882711
transform -1 0 2168 0 -1 4610
box 0 0 16 200
use INVX2  INVX2_18
timestamp 1515882711
transform -1 0 2200 0 -1 4610
box 0 0 32 200
use FILL  FILL_INVX2_32
timestamp 1515882711
transform -1 0 2216 0 -1 4610
box 0 0 16 200
use INVX2  INVX2_32
timestamp 1515882711
transform -1 0 2248 0 -1 4610
box 0 0 32 200
use OAI21X1  OAI21X1_166
timestamp 1515882711
transform 1 0 2248 0 -1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_183
timestamp 1515882711
transform -1 0 2328 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_183
timestamp 1515882711
transform -1 0 2520 0 -1 4610
box 0 0 192 200
use FILL  FILL_INVX8_2
timestamp 1515882711
transform 1 0 2520 0 -1 4610
box 0 0 16 200
use INVX8  INVX8_2
timestamp 1515882711
transform 1 0 2536 0 -1 4610
box 0 0 80 200
use FILL  FILL_NAND2X1_386
timestamp 1515882711
transform 1 0 2616 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_386
timestamp 1515882711
transform 1 0 2632 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_454
timestamp 1515882711
transform -1 0 2744 0 -1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_9
timestamp 1515882711
transform 1 0 2744 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1515882711
transform 1 0 2760 0 -1 4610
box 0 0 192 200
use FILL  FILL_INVX1_50
timestamp 1515882711
transform 1 0 2952 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_0
timestamp 1515882711
transform 1 0 2968 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_2_1
timestamp 1515882711
transform 1 0 2984 0 -1 4610
box 0 0 16 200
use INVX1  INVX1_50
timestamp 1515882711
transform 1 0 3000 0 -1 4610
box 0 0 32 200
use FILL  FILL_NAND2X1_261
timestamp 1515882711
transform -1 0 3048 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_261
timestamp 1515882711
transform -1 0 3096 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_289
timestamp 1515882711
transform -1 0 3160 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_292
timestamp 1515882711
transform 1 0 3160 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_398
timestamp 1515882711
transform 1 0 3224 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_177
timestamp 1515882711
transform 1 0 3288 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_320
timestamp 1515882711
transform 1 0 3352 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_321
timestamp 1515882711
transform 1 0 3416 0 -1 4610
box 0 0 64 200
use NAND3X1  NAND3X1_178
timestamp 1515882711
transform -1 0 3544 0 -1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_331
timestamp 1515882711
transform 1 0 3544 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_331
timestamp 1515882711
transform 1 0 3560 0 -1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_227
timestamp 1515882711
transform 1 0 3608 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_227
timestamp 1515882711
transform 1 0 3624 0 -1 4610
box 0 0 48 200
use FILL  FILL_BUFX4_217
timestamp 1515882711
transform -1 0 3688 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_217
timestamp 1515882711
transform -1 0 3752 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_342
timestamp 1515882711
transform 1 0 3752 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_420
timestamp 1515882711
transform 1 0 3816 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_29
timestamp 1515882711
transform -1 0 3928 0 -1 4610
box 0 0 48 200
use NAND3X1  NAND3X1_255
timestamp 1515882711
transform 1 0 3928 0 -1 4610
box 0 0 64 200
use FILL  FILL_22_3_0
timestamp 1515882711
transform 1 0 3992 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_3_1
timestamp 1515882711
transform 1 0 4008 0 -1 4610
box 0 0 16 200
use NAND3X1  NAND3X1_111
timestamp 1515882711
transform 1 0 4024 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_72
timestamp 1515882711
transform -1 0 4136 0 -1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_329
timestamp 1515882711
transform 1 0 4136 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_329
timestamp 1515882711
transform 1 0 4152 0 -1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_218
timestamp 1515882711
transform 1 0 4200 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_218
timestamp 1515882711
transform 1 0 4216 0 -1 4610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_76
timestamp 1515882711
transform -1 0 4280 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_76
timestamp 1515882711
transform -1 0 4472 0 -1 4610
box 0 0 192 200
use FILL  FILL_NAND2X1_58
timestamp 1515882711
transform 1 0 4472 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_58
timestamp 1515882711
transform 1 0 4488 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_76
timestamp 1515882711
transform -1 0 4600 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_50
timestamp 1515882711
transform -1 0 4616 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_50
timestamp 1515882711
transform -1 0 4680 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_293
timestamp 1515882711
transform 1 0 4680 0 -1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_217
timestamp 1515882711
transform -1 0 4760 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_217
timestamp 1515882711
transform -1 0 4808 0 -1 4610
box 0 0 48 200
use NAND2X1  NAND2X1_409
timestamp 1515882711
transform 1 0 4808 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_334
timestamp 1515882711
transform -1 0 4920 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_195
timestamp 1515882711
transform 1 0 4920 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_195
timestamp 1515882711
transform 1 0 4936 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_216
timestamp 1515882711
transform -1 0 5016 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_4_0
timestamp 1515882711
transform -1 0 5032 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_4_1
timestamp 1515882711
transform -1 0 5048 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_216
timestamp 1515882711
transform -1 0 5112 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_203
timestamp 1515882711
transform -1 0 5128 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_203
timestamp 1515882711
transform -1 0 5192 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_158
timestamp 1515882711
transform -1 0 5240 0 -1 4610
box 0 0 48 200
use NOR3X1  NOR3X1_2
timestamp 1515882711
transform 1 0 5240 0 -1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_239
timestamp 1515882711
transform 1 0 5368 0 -1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_220
timestamp 1515882711
transform -1 0 5448 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_220
timestamp 1515882711
transform -1 0 5496 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_375
timestamp 1515882711
transform -1 0 5560 0 -1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_330
timestamp 1515882711
transform -1 0 5576 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_330
timestamp 1515882711
transform -1 0 5624 0 -1 4610
box 0 0 48 200
use FILL  FILL_BUFX4_248
timestamp 1515882711
transform 1 0 5624 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_248
timestamp 1515882711
transform 1 0 5640 0 -1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_244
timestamp 1515882711
transform -1 0 5720 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_244
timestamp 1515882711
transform -1 0 5768 0 -1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_338
timestamp 1515882711
transform -1 0 5784 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_338
timestamp 1515882711
transform -1 0 5832 0 -1 4610
box 0 0 48 200
use FILL  FILL_BUFX4_84
timestamp 1515882711
transform -1 0 5848 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_84
timestamp 1515882711
transform -1 0 5912 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_200
timestamp 1515882711
transform 1 0 5912 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_200
timestamp 1515882711
transform 1 0 5928 0 -1 4610
box 0 0 64 200
use NOR2X1  NOR2X1_11
timestamp 1515882711
transform 1 0 5992 0 -1 4610
box 0 0 48 200
use FILL  FILL_22_5_0
timestamp 1515882711
transform 1 0 6040 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_5_1
timestamp 1515882711
transform 1 0 6056 0 -1 4610
box 0 0 16 200
use OAI22X1  OAI22X1_2
timestamp 1515882711
transform 1 0 6072 0 -1 4610
box 0 0 80 200
use NOR2X1  NOR2X1_10
timestamp 1515882711
transform -1 0 6200 0 -1 4610
box 0 0 48 200
use NOR3X1  NOR3X1_13
timestamp 1515882711
transform 1 0 6200 0 -1 4610
box 0 0 128 200
use FILL  FILL_NAND2X1_328
timestamp 1515882711
transform -1 0 6344 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_328
timestamp 1515882711
transform -1 0 6392 0 -1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_213
timestamp 1515882711
transform 1 0 6392 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_213
timestamp 1515882711
transform 1 0 6408 0 -1 4610
box 0 0 48 200
use NOR3X1  NOR3X1_6
timestamp 1515882711
transform -1 0 6584 0 -1 4610
box 0 0 128 200
use NOR2X1  NOR2X1_164
timestamp 1515882711
transform -1 0 6632 0 -1 4610
box 0 0 48 200
use NOR2X1  NOR2X1_28
timestamp 1515882711
transform -1 0 6680 0 -1 4610
box 0 0 48 200
use NOR3X1  NOR3X1_24
timestamp 1515882711
transform 1 0 6680 0 -1 4610
box 0 0 128 200
use OAI21X1  OAI21X1_339
timestamp 1515882711
transform 1 0 6808 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_259
timestamp 1515882711
transform 1 0 6872 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_419
timestamp 1515882711
transform -1 0 7000 0 -1 4610
box 0 0 64 200
use FILL  FILL_NAND2X1_237
timestamp 1515882711
transform -1 0 7016 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_237
timestamp 1515882711
transform -1 0 7064 0 -1 4610
box 0 0 48 200
use FILL  FILL_NAND2X1_336
timestamp 1515882711
transform -1 0 7080 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_6_0
timestamp 1515882711
transform -1 0 7096 0 -1 4610
box 0 0 16 200
use FILL  FILL_22_6_1
timestamp 1515882711
transform -1 0 7112 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_336
timestamp 1515882711
transform -1 0 7160 0 -1 4610
box 0 0 48 200
use OAI21X1  OAI21X1_258
timestamp 1515882711
transform -1 0 7224 0 -1 4610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_127
timestamp 1515882711
transform 1 0 7224 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_127
timestamp 1515882711
transform 1 0 7240 0 -1 4610
box 0 0 192 200
use OAI21X1  OAI21X1_127
timestamp 1515882711
transform -1 0 7496 0 -1 4610
box 0 0 64 200
use FILL  FILL_BUFX4_273
timestamp 1515882711
transform 1 0 7496 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_273
timestamp 1515882711
transform 1 0 7512 0 -1 4610
box 0 0 64 200
use OAI21X1  OAI21X1_484
timestamp 1515882711
transform 1 0 7576 0 -1 4610
box 0 0 64 200
use NAND2X1  NAND2X1_432
timestamp 1515882711
transform -1 0 7688 0 -1 4610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_305
timestamp 1515882711
transform -1 0 7704 0 -1 4610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_305
timestamp 1515882711
transform -1 0 7896 0 -1 4610
box 0 0 192 200
use FILL  FILL_NAND2X1_132
timestamp 1515882711
transform -1 0 7912 0 -1 4610
box 0 0 16 200
use NAND2X1  NAND2X1_132
timestamp 1515882711
transform -1 0 7960 0 -1 4610
box 0 0 48 200
use FILL  FILL_BUFX4_287
timestamp 1515882711
transform 1 0 7960 0 -1 4610
box 0 0 16 200
use BUFX4  BUFX4_287
timestamp 1515882711
transform 1 0 7976 0 -1 4610
box 0 0 64 200
use FILL  FILL_23_1
timestamp 1515882711
transform -1 0 8056 0 -1 4610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_252
timestamp 1515882711
transform -1 0 24 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_252
timestamp 1515882711
transform -1 0 216 0 1 4210
box 0 0 192 200
use NAND3X1  NAND3X1_262
timestamp 1515882711
transform -1 0 280 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_119
timestamp 1515882711
transform 1 0 280 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_121
timestamp 1515882711
transform 1 0 344 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_120
timestamp 1515882711
transform 1 0 408 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_230
timestamp 1515882711
transform -1 0 536 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_264
timestamp 1515882711
transform 1 0 536 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_263
timestamp 1515882711
transform 1 0 600 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_53
timestamp 1515882711
transform 1 0 664 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_52
timestamp 1515882711
transform 1 0 728 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_54
timestamp 1515882711
transform 1 0 792 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_315
timestamp 1515882711
transform 1 0 856 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_315
timestamp 1515882711
transform 1 0 872 0 1 4210
box 0 0 48 200
use FILL  FILL_21_0_0
timestamp 1515882711
transform -1 0 936 0 1 4210
box 0 0 16 200
use FILL  FILL_21_0_1
timestamp 1515882711
transform -1 0 952 0 1 4210
box 0 0 16 200
use NAND3X1  NAND3X1_117
timestamp 1515882711
transform -1 0 1016 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_260
timestamp 1515882711
transform 1 0 1016 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_116
timestamp 1515882711
transform 1 0 1080 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_259
timestamp 1515882711
transform 1 0 1144 0 1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_301
timestamp 1515882711
transform -1 0 1224 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_301
timestamp 1515882711
transform -1 0 1288 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_150
timestamp 1515882711
transform -1 0 1304 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_150
timestamp 1515882711
transform -1 0 1352 0 1 4210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_216
timestamp 1515882711
transform -1 0 1368 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_216
timestamp 1515882711
transform -1 0 1560 0 1 4210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_218
timestamp 1515882711
transform 1 0 1560 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_218
timestamp 1515882711
transform 1 0 1576 0 1 4210
box 0 0 192 200
use FILL  FILL_AOI21X1_51
timestamp 1515882711
transform 1 0 1768 0 1 4210
box 0 0 16 200
use AOI21X1  AOI21X1_51
timestamp 1515882711
transform 1 0 1784 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_127
timestamp 1515882711
transform -1 0 1896 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_139
timestamp 1515882711
transform -1 0 1960 0 1 4210
box 0 0 64 200
use FILL  FILL_21_1_0
timestamp 1515882711
transform 1 0 1960 0 1 4210
box 0 0 16 200
use FILL  FILL_21_1_1
timestamp 1515882711
transform 1 0 1976 0 1 4210
box 0 0 16 200
use NAND3X1  NAND3X1_282
timestamp 1515882711
transform 1 0 1992 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_256
timestamp 1515882711
transform -1 0 2120 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_383
timestamp 1515882711
transform -1 0 2184 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_172
timestamp 1515882711
transform -1 0 2200 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_172
timestamp 1515882711
transform -1 0 2248 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_184
timestamp 1515882711
transform 1 0 2248 0 1 4210
box 0 0 64 200
use FILL  FILL_INVX2_17
timestamp 1515882711
transform -1 0 2328 0 1 4210
box 0 0 16 200
use INVX2  INVX2_17
timestamp 1515882711
transform -1 0 2360 0 1 4210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_237
timestamp 1515882711
transform -1 0 2376 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_237
timestamp 1515882711
transform -1 0 2568 0 1 4210
box 0 0 192 200
use FILL  FILL_INVX1_33
timestamp 1515882711
transform -1 0 2584 0 1 4210
box 0 0 16 200
use INVX1  INVX1_33
timestamp 1515882711
transform -1 0 2616 0 1 4210
box 0 0 32 200
use FILL  FILL_NAND2X1_238
timestamp 1515882711
transform -1 0 2632 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_238
timestamp 1515882711
transform -1 0 2680 0 1 4210
box 0 0 48 200
use FILL  FILL_BUFX4_244
timestamp 1515882711
transform -1 0 2696 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_244
timestamp 1515882711
transform -1 0 2760 0 1 4210
box 0 0 64 200
use FILL  FILL_INVX8_16
timestamp 1515882711
transform 1 0 2760 0 1 4210
box 0 0 16 200
use INVX8  INVX8_16
timestamp 1515882711
transform 1 0 2776 0 1 4210
box 0 0 80 200
use NAND3X1  NAND3X1_148
timestamp 1515882711
transform -1 0 2920 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_4
timestamp 1515882711
transform -1 0 2984 0 1 4210
box 0 0 64 200
use FILL  FILL_21_2_0
timestamp 1515882711
transform -1 0 3000 0 1 4210
box 0 0 16 200
use FILL  FILL_21_2_1
timestamp 1515882711
transform -1 0 3016 0 1 4210
box 0 0 16 200
use NOR2X1  NOR2X1_12
timestamp 1515882711
transform -1 0 3064 0 1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_181
timestamp 1515882711
transform -1 0 3128 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_291
timestamp 1515882711
transform -1 0 3192 0 1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_61
timestamp 1515882711
transform -1 0 3240 0 1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_343
timestamp 1515882711
transform -1 0 3256 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_343
timestamp 1515882711
transform -1 0 3304 0 1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_265
timestamp 1515882711
transform -1 0 3320 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_265
timestamp 1515882711
transform -1 0 3368 0 1 4210
box 0 0 48 200
use FILL  FILL_BUFX4_196
timestamp 1515882711
transform -1 0 3384 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_196
timestamp 1515882711
transform -1 0 3448 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_266
timestamp 1515882711
transform -1 0 3512 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_123
timestamp 1515882711
transform -1 0 3576 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_125
timestamp 1515882711
transform 1 0 3576 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_268
timestamp 1515882711
transform 1 0 3640 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_74
timestamp 1515882711
transform -1 0 3768 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_55
timestamp 1515882711
transform -1 0 3832 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_233
timestamp 1515882711
transform 1 0 3832 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_257
timestamp 1515882711
transform -1 0 3960 0 1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_114
timestamp 1515882711
transform 1 0 3960 0 1 4210
box 0 0 64 200
use FILL  FILL_21_3_0
timestamp 1515882711
transform -1 0 4040 0 1 4210
box 0 0 16 200
use FILL  FILL_21_3_1
timestamp 1515882711
transform -1 0 4056 0 1 4210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_74
timestamp 1515882711
transform -1 0 4072 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_74
timestamp 1515882711
transform -1 0 4264 0 1 4210
box 0 0 192 200
use FILL  FILL_INVX1_36
timestamp 1515882711
transform -1 0 4280 0 1 4210
box 0 0 16 200
use INVX1  INVX1_36
timestamp 1515882711
transform -1 0 4312 0 1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_234
timestamp 1515882711
transform -1 0 4376 0 1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_146
timestamp 1515882711
transform -1 0 4392 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_146
timestamp 1515882711
transform -1 0 4584 0 1 4210
box 0 0 192 200
use FILL  FILL_BUFX4_245
timestamp 1515882711
transform -1 0 4600 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_245
timestamp 1515882711
transform -1 0 4664 0 1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_30
timestamp 1515882711
transform 1 0 4664 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_30
timestamp 1515882711
transform 1 0 4680 0 1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_45
timestamp 1515882711
transform -1 0 4760 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_45
timestamp 1515882711
transform -1 0 4824 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_263
timestamp 1515882711
transform 1 0 4824 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_263
timestamp 1515882711
transform 1 0 4840 0 1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_212
timestamp 1515882711
transform 1 0 4888 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_212
timestamp 1515882711
transform 1 0 4904 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_179
timestamp 1515882711
transform -1 0 5016 0 1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_179
timestamp 1515882711
transform -1 0 5032 0 1 4210
box 0 0 16 200
use FILL  FILL_21_4_0
timestamp 1515882711
transform -1 0 5048 0 1 4210
box 0 0 16 200
use FILL  FILL_21_4_1
timestamp 1515882711
transform -1 0 5064 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_179
timestamp 1515882711
transform -1 0 5256 0 1 4210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_309
timestamp 1515882711
transform 1 0 5256 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_309
timestamp 1515882711
transform 1 0 5272 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_312
timestamp 1515882711
transform -1 0 5528 0 1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_321
timestamp 1515882711
transform 1 0 5528 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_321
timestamp 1515882711
transform 1 0 5544 0 1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_464
timestamp 1515882711
transform 1 0 5736 0 1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_410
timestamp 1515882711
transform 1 0 5800 0 1 4210
box 0 0 48 200
use FILL  FILL_MUX2X1_8
timestamp 1515882711
transform -1 0 5864 0 1 4210
box 0 0 16 200
use MUX2X1  MUX2X1_8
timestamp 1515882711
transform -1 0 5960 0 1 4210
box 0 0 96 200
use OAI21X1  OAI21X1_129
timestamp 1515882711
transform 1 0 5960 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_114
timestamp 1515882711
transform -1 0 6040 0 1 4210
box 0 0 16 200
use FILL  FILL_21_5_0
timestamp 1515882711
transform -1 0 6056 0 1 4210
box 0 0 16 200
use FILL  FILL_21_5_1
timestamp 1515882711
transform -1 0 6072 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_114
timestamp 1515882711
transform -1 0 6120 0 1 4210
box 0 0 48 200
use NOR2X1  NOR2X1_60
timestamp 1515882711
transform -1 0 6168 0 1 4210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_129
timestamp 1515882711
transform 1 0 6168 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_129
timestamp 1515882711
transform 1 0 6184 0 1 4210
box 0 0 192 200
use NAND2X1  NAND2X1_429
timestamp 1515882711
transform 1 0 6376 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_482
timestamp 1515882711
transform -1 0 6488 0 1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_67
timestamp 1515882711
transform 1 0 6488 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_67
timestamp 1515882711
transform 1 0 6504 0 1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_269
timestamp 1515882711
transform -1 0 6584 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_269
timestamp 1515882711
transform -1 0 6648 0 1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_191
timestamp 1515882711
transform -1 0 6664 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_191
timestamp 1515882711
transform -1 0 6728 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_120
timestamp 1515882711
transform 1 0 6728 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_120
timestamp 1515882711
transform 1 0 6744 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_136
timestamp 1515882711
transform -1 0 6856 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_298
timestamp 1515882711
transform -1 0 6872 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_298
timestamp 1515882711
transform -1 0 6920 0 1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_353
timestamp 1515882711
transform 1 0 6920 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_353
timestamp 1515882711
transform 1 0 6936 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_488
timestamp 1515882711
transform -1 0 7048 0 1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_310
timestamp 1515882711
transform -1 0 7064 0 1 4210
box 0 0 16 200
use FILL  FILL_21_6_0
timestamp 1515882711
transform -1 0 7080 0 1 4210
box 0 0 16 200
use FILL  FILL_21_6_1
timestamp 1515882711
transform -1 0 7096 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_310
timestamp 1515882711
transform -1 0 7288 0 1 4210
box 0 0 192 200
use FILL  FILL_BUFX4_189
timestamp 1515882711
transform 1 0 7288 0 1 4210
box 0 0 16 200
use BUFX4  BUFX4_189
timestamp 1515882711
transform 1 0 7304 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_228
timestamp 1515882711
transform 1 0 7368 0 1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_211
timestamp 1515882711
transform 1 0 7432 0 1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_211
timestamp 1515882711
transform 1 0 7448 0 1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_501
timestamp 1515882711
transform 1 0 7496 0 1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_500
timestamp 1515882711
transform -1 0 7624 0 1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_283
timestamp 1515882711
transform -1 0 7640 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_283
timestamp 1515882711
transform -1 0 7832 0 1 4210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_149
timestamp 1515882711
transform 1 0 7832 0 1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_149
timestamp 1515882711
transform 1 0 7848 0 1 4210
box 0 0 192 200
use FILL  FILL_22_1
timestamp 1515882711
transform 1 0 8040 0 1 4210
box 0 0 16 200
use NAND3X1  NAND3X1_273
timestamp 1515882711
transform -1 0 72 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_46
timestamp 1515882711
transform 1 0 72 0 -1 4210
box 0 0 48 200
use FILL  FILL_AOI21X1_45
timestamp 1515882711
transform -1 0 136 0 -1 4210
box 0 0 16 200
use AOI21X1  AOI21X1_45
timestamp 1515882711
transform -1 0 200 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_130
timestamp 1515882711
transform 1 0 200 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_132
timestamp 1515882711
transform -1 0 328 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_118
timestamp 1515882711
transform -1 0 392 0 -1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_163
timestamp 1515882711
transform -1 0 408 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_163
timestamp 1515882711
transform -1 0 600 0 -1 4210
box 0 0 192 200
use FILL  FILL_BUFX4_22
timestamp 1515882711
transform -1 0 616 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_22
timestamp 1515882711
transform -1 0 680 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_182
timestamp 1515882711
transform 1 0 680 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_182
timestamp 1515882711
transform 1 0 696 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_270
timestamp 1515882711
transform -1 0 808 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_127
timestamp 1515882711
transform 1 0 808 0 -1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_97
timestamp 1515882711
transform -1 0 888 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_97
timestamp 1515882711
transform -1 0 952 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_0_0
timestamp 1515882711
transform -1 0 968 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_0_1
timestamp 1515882711
transform -1 0 984 0 -1 4210
box 0 0 16 200
use FILL  FILL_INVX2_31
timestamp 1515882711
transform -1 0 1000 0 -1 4210
box 0 0 16 200
use INVX2  INVX2_31
timestamp 1515882711
transform -1 0 1032 0 -1 4210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_182
timestamp 1515882711
transform -1 0 1048 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_182
timestamp 1515882711
transform -1 0 1240 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_165
timestamp 1515882711
transform 1 0 1240 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_125
timestamp 1515882711
transform 1 0 1304 0 -1 4210
box 0 0 48 200
use FILL  FILL_AOI21X1_49
timestamp 1515882711
transform -1 0 1368 0 -1 4210
box 0 0 16 200
use AOI21X1  AOI21X1_49
timestamp 1515882711
transform -1 0 1432 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_271
timestamp 1515882711
transform -1 0 1496 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_128
timestamp 1515882711
transform 1 0 1496 0 -1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_124
timestamp 1515882711
transform 1 0 1560 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_124
timestamp 1515882711
transform 1 0 1576 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_138
timestamp 1515882711
transform -1 0 1704 0 -1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_93
timestamp 1515882711
transform 1 0 1704 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_93
timestamp 1515882711
transform 1 0 1720 0 -1 4210
box 0 0 64 200
use NOR3X1  NOR3X1_5
timestamp 1515882711
transform -1 0 1912 0 -1 4210
box 0 0 128 200
use OAI21X1  OAI21X1_255
timestamp 1515882711
transform -1 0 1976 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_1_0
timestamp 1515882711
transform -1 0 1992 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_1_1
timestamp 1515882711
transform -1 0 2008 0 -1 4210
box 0 0 16 200
use OAI21X1  OAI21X1_382
timestamp 1515882711
transform -1 0 2072 0 -1 4210
box 0 0 64 200
use NOR3X1  NOR3X1_33
timestamp 1515882711
transform 1 0 2072 0 -1 4210
box 0 0 128 200
use FILL  FILL_BUFX4_179
timestamp 1515882711
transform -1 0 2216 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_179
timestamp 1515882711
transform -1 0 2280 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_169
timestamp 1515882711
transform -1 0 2296 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_169
timestamp 1515882711
transform -1 0 2344 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_383
timestamp 1515882711
transform 1 0 2344 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_383
timestamp 1515882711
transform 1 0 2360 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_451
timestamp 1515882711
transform -1 0 2472 0 -1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_6
timestamp 1515882711
transform 1 0 2472 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1515882711
transform 1 0 2488 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_260
timestamp 1515882711
transform -1 0 2744 0 -1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_238
timestamp 1515882711
transform -1 0 2760 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_238
timestamp 1515882711
transform -1 0 2824 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_385
timestamp 1515882711
transform 1 0 2824 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_54
timestamp 1515882711
transform -1 0 2936 0 -1 4210
box 0 0 48 200
use FILL  FILL_BUFX4_234
timestamp 1515882711
transform 1 0 2936 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_0
timestamp 1515882711
transform 1 0 2952 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_2_1
timestamp 1515882711
transform 1 0 2968 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_234
timestamp 1515882711
transform 1 0 2984 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_262
timestamp 1515882711
transform 1 0 3048 0 -1 4210
box 0 0 64 200
use NOR2X1  NOR2X1_3
timestamp 1515882711
transform -1 0 3160 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_287
timestamp 1515882711
transform 1 0 3160 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_144
timestamp 1515882711
transform 1 0 3224 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_242
timestamp 1515882711
transform 1 0 3288 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_242
timestamp 1515882711
transform 1 0 3304 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_337
timestamp 1515882711
transform -1 0 3368 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_337
timestamp 1515882711
transform -1 0 3416 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_288
timestamp 1515882711
transform 1 0 3416 0 -1 4210
box 0 0 64 200
use NAND3X1  NAND3X1_145
timestamp 1515882711
transform -1 0 3544 0 -1 4210
box 0 0 64 200
use FILL  FILL_BUFX4_32
timestamp 1515882711
transform 1 0 3544 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_32
timestamp 1515882711
transform 1 0 3560 0 -1 4210
box 0 0 64 200
use FILL  FILL_INVX1_25
timestamp 1515882711
transform -1 0 3640 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_25
timestamp 1515882711
transform -1 0 3672 0 -1 4210
box 0 0 32 200
use FILL  FILL_NAND2X1_55
timestamp 1515882711
transform 1 0 3672 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_55
timestamp 1515882711
transform 1 0 3688 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_243
timestamp 1515882711
transform 1 0 3736 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_354
timestamp 1515882711
transform 1 0 3800 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_354
timestamp 1515882711
transform 1 0 3816 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_304
timestamp 1515882711
transform 1 0 3864 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_304
timestamp 1515882711
transform 1 0 3880 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_263
timestamp 1515882711
transform -1 0 3992 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_240
timestamp 1515882711
transform 1 0 3992 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_3_0
timestamp 1515882711
transform 1 0 4008 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_3_1
timestamp 1515882711
transform 1 0 4024 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_240
timestamp 1515882711
transform 1 0 4040 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_179
timestamp 1515882711
transform 1 0 4088 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_179
timestamp 1515882711
transform 1 0 4104 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_146
timestamp 1515882711
transform -1 0 4216 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_225
timestamp 1515882711
transform 1 0 4216 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_225
timestamp 1515882711
transform 1 0 4232 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_157
timestamp 1515882711
transform 1 0 4280 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_157
timestamp 1515882711
transform 1 0 4296 0 -1 4210
box 0 0 48 200
use FILL  FILL_INVX1_20
timestamp 1515882711
transform -1 0 4360 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_20
timestamp 1515882711
transform -1 0 4392 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_481
timestamp 1515882711
transform 1 0 4392 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_442
timestamp 1515882711
transform -1 0 4504 0 -1 4210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_23
timestamp 1515882711
transform -1 0 4520 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_23
timestamp 1515882711
transform -1 0 4712 0 -1 4210
box 0 0 192 200
use FILL  FILL_NAND2X1_241
timestamp 1515882711
transform -1 0 4728 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_241
timestamp 1515882711
transform -1 0 4776 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_36
timestamp 1515882711
transform 1 0 4776 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_36
timestamp 1515882711
transform 1 0 4792 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_55
timestamp 1515882711
transform -1 0 4904 0 -1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_55
timestamp 1515882711
transform -1 0 4920 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_55
timestamp 1515882711
transform -1 0 5112 0 -1 4210
box 0 0 192 200
use FILL  FILL_20_4_0
timestamp 1515882711
transform 1 0 5112 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_4_1
timestamp 1515882711
transform 1 0 5128 0 -1 4210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_93
timestamp 1515882711
transform 1 0 5144 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_93
timestamp 1515882711
transform 1 0 5160 0 -1 4210
box 0 0 192 200
use FILL  FILL_MUX2X1_9
timestamp 1515882711
transform 1 0 5352 0 -1 4210
box 0 0 16 200
use MUX2X1  MUX2X1_9
timestamp 1515882711
transform 1 0 5368 0 -1 4210
box 0 0 96 200
use FILL  FILL_NAND2X1_368
timestamp 1515882711
transform 1 0 5464 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_368
timestamp 1515882711
transform 1 0 5480 0 -1 4210
box 0 0 48 200
use FILL  FILL_NAND2X1_75
timestamp 1515882711
transform 1 0 5528 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_75
timestamp 1515882711
transform 1 0 5544 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_93
timestamp 1515882711
transform -1 0 5656 0 -1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_110
timestamp 1515882711
transform 1 0 5656 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_110
timestamp 1515882711
transform 1 0 5672 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_110
timestamp 1515882711
transform 1 0 5864 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_94
timestamp 1515882711
transform 1 0 5928 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_94
timestamp 1515882711
transform 1 0 5944 0 -1 4210
box 0 0 48 200
use FILL  FILL_BUFX4_69
timestamp 1515882711
transform -1 0 6008 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_69
timestamp 1515882711
transform -1 0 6072 0 -1 4210
box 0 0 64 200
use FILL  FILL_20_5_0
timestamp 1515882711
transform 1 0 6072 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_5_1
timestamp 1515882711
transform 1 0 6088 0 -1 4210
box 0 0 16 200
use FILL  FILL_BUFX4_199
timestamp 1515882711
transform 1 0 6104 0 -1 4210
box 0 0 16 200
use BUFX4  BUFX4_199
timestamp 1515882711
transform 1 0 6120 0 -1 4210
box 0 0 64 200
use FILL  FILL_MUX2X1_10
timestamp 1515882711
transform 1 0 6184 0 -1 4210
box 0 0 16 200
use MUX2X1  MUX2X1_10
timestamp 1515882711
transform 1 0 6200 0 -1 4210
box 0 0 96 200
use FILL  FILL_DFFPOSX1_303
timestamp 1515882711
transform -1 0 6312 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_303
timestamp 1515882711
transform -1 0 6504 0 -1 4210
box 0 0 192 200
use FILL  FILL_MUX2X1_30
timestamp 1515882711
transform 1 0 6504 0 -1 4210
box 0 0 16 200
use MUX2X1  MUX2X1_30
timestamp 1515882711
transform 1 0 6520 0 -1 4210
box 0 0 96 200
use FILL  FILL_DFFPOSX1_136
timestamp 1515882711
transform -1 0 6632 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_136
timestamp 1515882711
transform -1 0 6824 0 -1 4210
box 0 0 192 200
use FILL  FILL_NAND2X1_236
timestamp 1515882711
transform 1 0 6824 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_236
timestamp 1515882711
transform 1 0 6840 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_486
timestamp 1515882711
transform -1 0 6952 0 -1 4210
box 0 0 64 200
use NAND2X1  NAND2X1_436
timestamp 1515882711
transform 1 0 6952 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_144
timestamp 1515882711
transform 1 0 7000 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_130
timestamp 1515882711
transform -1 0 7080 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_6_0
timestamp 1515882711
transform -1 0 7096 0 -1 4210
box 0 0 16 200
use FILL  FILL_20_6_1
timestamp 1515882711
transform -1 0 7112 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_130
timestamp 1515882711
transform -1 0 7160 0 -1 4210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_144
timestamp 1515882711
transform 1 0 7160 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_144
timestamp 1515882711
transform 1 0 7176 0 -1 4210
box 0 0 192 200
use FILL  FILL_INVX1_16
timestamp 1515882711
transform 1 0 7368 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_16
timestamp 1515882711
transform 1 0 7384 0 -1 4210
box 0 0 32 200
use OAI21X1  OAI21X1_267
timestamp 1515882711
transform -1 0 7480 0 -1 4210
box 0 0 64 200
use FILL  FILL_INVX1_38
timestamp 1515882711
transform -1 0 7496 0 -1 4210
box 0 0 16 200
use INVX1  INVX1_38
timestamp 1515882711
transform -1 0 7528 0 -1 4210
box 0 0 32 200
use FILL  FILL_NAND2X1_243
timestamp 1515882711
transform 1 0 7528 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_243
timestamp 1515882711
transform 1 0 7544 0 -1 4210
box 0 0 48 200
use OAI21X1  OAI21X1_509
timestamp 1515882711
transform 1 0 7592 0 -1 4210
box 0 0 64 200
use OAI21X1  OAI21X1_510
timestamp 1515882711
transform -1 0 7720 0 -1 4210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_288
timestamp 1515882711
transform -1 0 7736 0 -1 4210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_288
timestamp 1515882711
transform -1 0 7928 0 -1 4210
box 0 0 192 200
use OAI21X1  OAI21X1_147
timestamp 1515882711
transform 1 0 7928 0 -1 4210
box 0 0 64 200
use FILL  FILL_NAND2X1_134
timestamp 1515882711
transform -1 0 8008 0 -1 4210
box 0 0 16 200
use NAND2X1  NAND2X1_134
timestamp 1515882711
transform -1 0 8056 0 -1 4210
box 0 0 48 200
use NAND3X1  NAND3X1_274
timestamp 1515882711
transform -1 0 72 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_275
timestamp 1515882711
transform -1 0 136 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_272
timestamp 1515882711
transform -1 0 200 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_131
timestamp 1515882711
transform 1 0 200 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_129
timestamp 1515882711
transform 1 0 264 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_261
timestamp 1515882711
transform -1 0 392 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_91
timestamp 1515882711
transform 1 0 392 0 1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_90
timestamp 1515882711
transform 1 0 440 0 1 3810
box 0 0 48 200
use FILL  FILL_AOI21X1_14
timestamp 1515882711
transform -1 0 504 0 1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_14
timestamp 1515882711
transform -1 0 568 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_180
timestamp 1515882711
transform -1 0 584 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_180
timestamp 1515882711
transform -1 0 648 0 1 3810
box 0 0 64 200
use FILL  FILL_AOI21X1_32
timestamp 1515882711
transform 1 0 648 0 1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_32
timestamp 1515882711
transform 1 0 664 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_108
timestamp 1515882711
transform -1 0 776 0 1 3810
box 0 0 48 200
use NOR3X1  NOR3X1_3
timestamp 1515882711
transform -1 0 904 0 1 3810
box 0 0 128 200
use FILL  FILL_19_0_0
timestamp 1515882711
transform -1 0 920 0 1 3810
box 0 0 16 200
use FILL  FILL_19_0_1
timestamp 1515882711
transform -1 0 936 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_245
timestamp 1515882711
transform -1 0 1000 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_377
timestamp 1515882711
transform -1 0 1064 0 1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_107
timestamp 1515882711
transform -1 0 1112 0 1 3810
box 0 0 48 200
use FILL  FILL_AOI21X1_31
timestamp 1515882711
transform -1 0 1128 0 1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_31
timestamp 1515882711
transform -1 0 1192 0 1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_32
timestamp 1515882711
transform -1 0 1320 0 1 3810
box 0 0 128 200
use FILL  FILL_BUFX4_54
timestamp 1515882711
transform -1 0 1336 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_54
timestamp 1515882711
transform -1 0 1400 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_247
timestamp 1515882711
transform 1 0 1400 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_378
timestamp 1515882711
transform 1 0 1464 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_113
timestamp 1515882711
transform -1 0 1544 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_113
timestamp 1515882711
transform -1 0 1608 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_281
timestamp 1515882711
transform -1 0 1672 0 1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_240
timestamp 1515882711
transform 1 0 1672 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_240
timestamp 1515882711
transform 1 0 1688 0 1 3810
box 0 0 192 200
use FILL  FILL_INVX2_20
timestamp 1515882711
transform 1 0 1880 0 1 3810
box 0 0 16 200
use INVX2  INVX2_20
timestamp 1515882711
transform 1 0 1896 0 1 3810
box 0 0 32 200
use FILL  FILL_19_1_0
timestamp 1515882711
transform 1 0 1928 0 1 3810
box 0 0 16 200
use FILL  FILL_19_1_1
timestamp 1515882711
transform 1 0 1944 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_187
timestamp 1515882711
transform 1 0 1960 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_183
timestamp 1515882711
transform 1 0 2024 0 1 3810
box 0 0 64 200
use FILL  FILL_INVX2_16
timestamp 1515882711
transform -1 0 2104 0 1 3810
box 0 0 16 200
use INVX2  INVX2_16
timestamp 1515882711
transform -1 0 2136 0 1 3810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_236
timestamp 1515882711
transform 1 0 2136 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_236
timestamp 1515882711
transform 1 0 2152 0 1 3810
box 0 0 192 200
use FILL  FILL_DFFPOSX1_5
timestamp 1515882711
transform 1 0 2344 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1515882711
transform 1 0 2360 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_23
timestamp 1515882711
transform 1 0 2552 0 1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_272
timestamp 1515882711
transform 1 0 2616 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_272
timestamp 1515882711
transform 1 0 2632 0 1 3810
box 0 0 192 200
use NOR2X1  NOR2X1_6
timestamp 1515882711
transform 1 0 2824 0 1 3810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_277
timestamp 1515882711
transform 1 0 2872 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_0
timestamp 1515882711
transform 1 0 2888 0 1 3810
box 0 0 16 200
use FILL  FILL_19_2_1
timestamp 1515882711
transform 1 0 2904 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_277
timestamp 1515882711
transform 1 0 2920 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_309
timestamp 1515882711
transform 1 0 3112 0 1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_7
timestamp 1515882711
transform 1 0 3176 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_7
timestamp 1515882711
transform 1 0 3192 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_29
timestamp 1515882711
transform -1 0 3304 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_254
timestamp 1515882711
transform -1 0 3320 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_254
timestamp 1515882711
transform -1 0 3384 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_38
timestamp 1515882711
transform -1 0 3400 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_38
timestamp 1515882711
transform -1 0 3464 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_290
timestamp 1515882711
transform 1 0 3464 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_147
timestamp 1515882711
transform 1 0 3528 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_257
timestamp 1515882711
transform 1 0 3592 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_257
timestamp 1515882711
transform 1 0 3608 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_40
timestamp 1515882711
transform 1 0 3672 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_40
timestamp 1515882711
transform 1 0 3688 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_234
timestamp 1515882711
transform 1 0 3752 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_56
timestamp 1515882711
transform -1 0 3880 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_58
timestamp 1515882711
transform -1 0 3944 0 1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_236
timestamp 1515882711
transform 1 0 3944 0 1 3810
box 0 0 64 200
use FILL  FILL_19_3_0
timestamp 1515882711
transform 1 0 4008 0 1 3810
box 0 0 16 200
use FILL  FILL_19_3_1
timestamp 1515882711
transform 1 0 4024 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_244
timestamp 1515882711
transform 1 0 4040 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_51
timestamp 1515882711
transform 1 0 4104 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_51
timestamp 1515882711
transform 1 0 4120 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_343
timestamp 1515882711
transform -1 0 4248 0 1 3810
box 0 0 64 200
use FILL  FILL_INVX1_80
timestamp 1515882711
transform -1 0 4264 0 1 3810
box 0 0 16 200
use INVX1  INVX1_80
timestamp 1515882711
transform -1 0 4296 0 1 3810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_85
timestamp 1515882711
transform -1 0 4312 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_85
timestamp 1515882711
transform -1 0 4504 0 1 3810
box 0 0 192 200
use FILL  FILL_NAND2X1_66
timestamp 1515882711
transform 1 0 4504 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_66
timestamp 1515882711
transform 1 0 4520 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_85
timestamp 1515882711
transform -1 0 4632 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_124
timestamp 1515882711
transform -1 0 4696 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_264
timestamp 1515882711
transform -1 0 4760 0 1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_124
timestamp 1515882711
transform -1 0 4776 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_124
timestamp 1515882711
transform -1 0 4968 0 1 3810
box 0 0 192 200
use NAND2X1  NAND2X1_431
timestamp 1515882711
transform 1 0 4968 0 1 3810
box 0 0 48 200
use FILL  FILL_19_4_0
timestamp 1515882711
transform -1 0 5032 0 1 3810
box 0 0 16 200
use FILL  FILL_19_4_1
timestamp 1515882711
transform -1 0 5048 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_470
timestamp 1515882711
transform -1 0 5112 0 1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_22
timestamp 1515882711
transform -1 0 5128 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_22
timestamp 1515882711
transform -1 0 5320 0 1 3810
box 0 0 192 200
use FILL  FILL_INVX1_37
timestamp 1515882711
transform -1 0 5336 0 1 3810
box 0 0 16 200
use INVX1  INVX1_37
timestamp 1515882711
transform -1 0 5368 0 1 3810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_59
timestamp 1515882711
transform -1 0 5384 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_59
timestamp 1515882711
transform -1 0 5576 0 1 3810
box 0 0 192 200
use FILL  FILL_NAND2X1_39
timestamp 1515882711
transform 1 0 5576 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_39
timestamp 1515882711
transform 1 0 5592 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_59
timestamp 1515882711
transform -1 0 5704 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_118
timestamp 1515882711
transform -1 0 5720 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_118
timestamp 1515882711
transform -1 0 5784 0 1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_117
timestamp 1515882711
transform 1 0 5784 0 1 3810
box 0 0 16 200
use BUFX4  BUFX4_117
timestamp 1515882711
transform 1 0 5800 0 1 3810
box 0 0 64 200
use OAI22X1  OAI22X1_13
timestamp 1515882711
transform 1 0 5864 0 1 3810
box 0 0 80 200
use NOR2X1  NOR2X1_51
timestamp 1515882711
transform -1 0 5992 0 1 3810
box 0 0 48 200
use NOR2X1  NOR2X1_162
timestamp 1515882711
transform 1 0 5992 0 1 3810
box 0 0 48 200
use FILL  FILL_19_5_0
timestamp 1515882711
transform 1 0 6040 0 1 3810
box 0 0 16 200
use FILL  FILL_19_5_1
timestamp 1515882711
transform 1 0 6056 0 1 3810
box 0 0 16 200
use NOR2X1  NOR2X1_161
timestamp 1515882711
transform 1 0 6072 0 1 3810
box 0 0 48 200
use NOR3X1  NOR3X1_4
timestamp 1515882711
transform 1 0 6120 0 1 3810
box 0 0 128 200
use OAI21X1  OAI21X1_249
timestamp 1515882711
transform 1 0 6248 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_380
timestamp 1515882711
transform 1 0 6312 0 1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_332
timestamp 1515882711
transform -1 0 6392 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_332
timestamp 1515882711
transform -1 0 6440 0 1 3810
box 0 0 48 200
use FILL  FILL_NAND2X1_229
timestamp 1515882711
transform -1 0 6456 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_229
timestamp 1515882711
transform -1 0 6504 0 1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_406
timestamp 1515882711
transform 1 0 6504 0 1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_286
timestamp 1515882711
transform 1 0 6568 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_286
timestamp 1515882711
transform 1 0 6584 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_508
timestamp 1515882711
transform 1 0 6776 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_507
timestamp 1515882711
transform -1 0 6904 0 1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_434
timestamp 1515882711
transform -1 0 6952 0 1 3810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_307
timestamp 1515882711
transform 1 0 6952 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_307
timestamp 1515882711
transform 1 0 6968 0 1 3810
box 0 0 192 200
use FILL  FILL_19_6_0
timestamp 1515882711
transform 1 0 7160 0 1 3810
box 0 0 16 200
use FILL  FILL_19_6_1
timestamp 1515882711
transform 1 0 7176 0 1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_153
timestamp 1515882711
transform 1 0 7192 0 1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_139
timestamp 1515882711
transform -1 0 7272 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_139
timestamp 1515882711
transform -1 0 7320 0 1 3810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_153
timestamp 1515882711
transform 1 0 7320 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_153
timestamp 1515882711
transform 1 0 7336 0 1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_248
timestamp 1515882711
transform -1 0 7592 0 1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_228
timestamp 1515882711
transform 1 0 7592 0 1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_228
timestamp 1515882711
transform 1 0 7608 0 1 3810
box 0 0 48 200
use FILL  FILL_INVX1_27
timestamp 1515882711
transform -1 0 7672 0 1 3810
box 0 0 16 200
use INVX1  INVX1_27
timestamp 1515882711
transform -1 0 7704 0 1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_505
timestamp 1515882711
transform 1 0 7704 0 1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_506
timestamp 1515882711
transform -1 0 7832 0 1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_147
timestamp 1515882711
transform 1 0 7832 0 1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_147
timestamp 1515882711
transform 1 0 7848 0 1 3810
box 0 0 192 200
use FILL  FILL_20_1
timestamp 1515882711
transform 1 0 8040 0 1 3810
box 0 0 16 200
use FILL  FILL_DFFPOSX1_253
timestamp 1515882711
transform -1 0 24 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_253
timestamp 1515882711
transform -1 0 216 0 -1 3810
box 0 0 192 200
use NOR2X1  NOR2X1_57
timestamp 1515882711
transform 1 0 216 0 -1 3810
box 0 0 48 200
use FILL  FILL_AOI21X1_56
timestamp 1515882711
transform -1 0 280 0 -1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_56
timestamp 1515882711
transform -1 0 344 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_164
timestamp 1515882711
transform -1 0 360 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_164
timestamp 1515882711
transform -1 0 552 0 -1 3810
box 0 0 192 200
use FILL  FILL_AOI21X1_15
timestamp 1515882711
transform -1 0 568 0 -1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_15
timestamp 1515882711
transform -1 0 632 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_199
timestamp 1515882711
transform 1 0 632 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_199
timestamp 1515882711
transform 1 0 648 0 -1 3810
box 0 0 192 200
use BUFX2  BUFX2_44
timestamp 1515882711
transform -1 0 888 0 -1 3810
box 0 0 48 200
use FILL  FILL_BUFX4_166
timestamp 1515882711
transform 1 0 888 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_0
timestamp 1515882711
transform 1 0 904 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_0_1
timestamp 1515882711
transform 1 0 920 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_166
timestamp 1515882711
transform 1 0 936 0 -1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_132
timestamp 1515882711
transform -1 0 1016 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_132
timestamp 1515882711
transform -1 0 1080 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_198
timestamp 1515882711
transform -1 0 1096 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_198
timestamp 1515882711
transform -1 0 1288 0 -1 3810
box 0 0 192 200
use FILL  FILL_BUFX2_4
timestamp 1515882711
transform -1 0 1304 0 -1 3810
box 0 0 16 200
use BUFX2  BUFX2_4
timestamp 1515882711
transform -1 0 1352 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_280
timestamp 1515882711
transform -1 0 1416 0 -1 3810
box 0 0 64 200
use FILL  FILL_AOI21X1_50
timestamp 1515882711
transform 1 0 1416 0 -1 3810
box 0 0 16 200
use AOI21X1  AOI21X1_50
timestamp 1515882711
transform 1 0 1432 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_126
timestamp 1515882711
transform 1 0 1496 0 -1 3810
box 0 0 48 200
use NAND3X1  NAND3X1_137
timestamp 1515882711
transform -1 0 1608 0 -1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_133
timestamp 1515882711
transform 1 0 1608 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_133
timestamp 1515882711
transform 1 0 1624 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_395
timestamp 1515882711
transform -1 0 1752 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_285
timestamp 1515882711
transform -1 0 1816 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_396
timestamp 1515882711
transform -1 0 1880 0 -1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_37
timestamp 1515882711
transform 1 0 1880 0 -1 3810
box 0 0 128 200
use FILL  FILL_18_1_0
timestamp 1515882711
transform -1 0 2024 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_1_1
timestamp 1515882711
transform -1 0 2040 0 -1 3810
box 0 0 16 200
use FILL  FILL_NAND2X1_167
timestamp 1515882711
transform -1 0 2056 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_167
timestamp 1515882711
transform -1 0 2104 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_286
timestamp 1515882711
transform 1 0 2104 0 -1 3810
box 0 0 64 200
use NOR3X1  NOR3X1_11
timestamp 1515882711
transform 1 0 2168 0 -1 3810
box 0 0 128 200
use FILL  FILL_INVX8_15
timestamp 1515882711
transform -1 0 2312 0 -1 3810
box 0 0 16 200
use INVX8  INVX8_15
timestamp 1515882711
transform -1 0 2392 0 -1 3810
box 0 0 80 200
use FILL  FILL_NAND2X1_382
timestamp 1515882711
transform 1 0 2392 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_382
timestamp 1515882711
transform 1 0 2408 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_450
timestamp 1515882711
transform -1 0 2520 0 -1 3810
box 0 0 64 200
use FILL  FILL_INVX1_28
timestamp 1515882711
transform 1 0 2520 0 -1 3810
box 0 0 16 200
use INVX1  INVX1_28
timestamp 1515882711
transform 1 0 2536 0 -1 3810
box 0 0 32 200
use NAND3X1  NAND3X1_203
timestamp 1515882711
transform -1 0 2632 0 -1 3810
box 0 0 64 200
use NAND2X1  NAND2X1_452
timestamp 1515882711
transform -1 0 2680 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_389
timestamp 1515882711
transform 1 0 2680 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_56
timestamp 1515882711
transform -1 0 2792 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_272
timestamp 1515882711
transform 1 0 2792 0 -1 3810
box 0 0 64 200
use FILL  FILL_BUFX4_21
timestamp 1515882711
transform 1 0 2856 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_21
timestamp 1515882711
transform 1 0 2872 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_65
timestamp 1515882711
transform 1 0 2936 0 -1 3810
box 0 0 48 200
use FILL  FILL_18_2_0
timestamp 1515882711
transform 1 0 2984 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_2_1
timestamp 1515882711
transform 1 0 3000 0 -1 3810
box 0 0 16 200
use OAI21X1  OAI21X1_407
timestamp 1515882711
transform 1 0 3016 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_311
timestamp 1515882711
transform -1 0 3144 0 -1 3810
box 0 0 64 200
use NAND3X1  NAND3X1_26
timestamp 1515882711
transform -1 0 3208 0 -1 3810
box 0 0 64 200
use NOR2X1  NOR2X1_19
timestamp 1515882711
transform -1 0 3256 0 -1 3810
box 0 0 48 200
use FILL  FILL_BUFX4_184
timestamp 1515882711
transform -1 0 3272 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_184
timestamp 1515882711
transform -1 0 3336 0 -1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_281
timestamp 1515882711
transform -1 0 3352 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_281
timestamp 1515882711
transform -1 0 3400 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_261
timestamp 1515882711
transform -1 0 3464 0 -1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_239
timestamp 1515882711
transform 1 0 3464 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_239
timestamp 1515882711
transform 1 0 3480 0 -1 3810
box 0 0 48 200
use FILL  FILL_NAND2X1_348
timestamp 1515882711
transform -1 0 3544 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_348
timestamp 1515882711
transform -1 0 3592 0 -1 3810
box 0 0 48 200
use FILL  FILL_INVX1_35
timestamp 1515882711
transform -1 0 3608 0 -1 3810
box 0 0 16 200
use INVX1  INVX1_35
timestamp 1515882711
transform -1 0 3640 0 -1 3810
box 0 0 32 200
use FILL  FILL_NAND2X1_365
timestamp 1515882711
transform 1 0 3640 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_365
timestamp 1515882711
transform 1 0 3656 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_432
timestamp 1515882711
transform -1 0 3768 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_339
timestamp 1515882711
transform -1 0 3784 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_339
timestamp 1515882711
transform -1 0 3976 0 -1 3810
box 0 0 192 200
use FILL  FILL_BUFX4_207
timestamp 1515882711
transform -1 0 3992 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_0
timestamp 1515882711
transform -1 0 4008 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_3_1
timestamp 1515882711
transform -1 0 4024 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_207
timestamp 1515882711
transform -1 0 4088 0 -1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_20
timestamp 1515882711
transform 1 0 4088 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_20
timestamp 1515882711
transform 1 0 4104 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_41
timestamp 1515882711
transform -1 0 4216 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_41
timestamp 1515882711
transform -1 0 4232 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_41
timestamp 1515882711
transform -1 0 4424 0 -1 3810
box 0 0 192 200
use FILL  FILL_NAND2X1_302
timestamp 1515882711
transform 1 0 4424 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_302
timestamp 1515882711
transform 1 0 4440 0 -1 3810
box 0 0 48 200
use FILL  FILL_NAND2X1_226
timestamp 1515882711
transform 1 0 4488 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_226
timestamp 1515882711
transform 1 0 4504 0 -1 3810
box 0 0 48 200
use FILL  FILL_NAND2X1_268
timestamp 1515882711
transform 1 0 4552 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_268
timestamp 1515882711
transform 1 0 4568 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_235
timestamp 1515882711
transform -1 0 4680 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_344
timestamp 1515882711
transform 1 0 4680 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_235
timestamp 1515882711
transform -1 0 4760 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_235
timestamp 1515882711
transform -1 0 4952 0 -1 3810
box 0 0 192 200
use FILL  FILL_NAND2X1_303
timestamp 1515882711
transform -1 0 4968 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_303
timestamp 1515882711
transform -1 0 5016 0 -1 3810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_32
timestamp 1515882711
transform -1 0 5032 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_4_0
timestamp 1515882711
transform -1 0 5048 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_4_1
timestamp 1515882711
transform -1 0 5064 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_32
timestamp 1515882711
transform -1 0 5256 0 -1 3810
box 0 0 192 200
use FILL  FILL_NAND2X1_79
timestamp 1515882711
transform 1 0 5256 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_79
timestamp 1515882711
transform 1 0 5272 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_57
timestamp 1515882711
transform -1 0 5384 0 -1 3810
box 0 0 64 200
use FILL  FILL_INVX1_64
timestamp 1515882711
transform -1 0 5400 0 -1 3810
box 0 0 16 200
use INVX1  INVX1_64
timestamp 1515882711
transform -1 0 5432 0 -1 3810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_64
timestamp 1515882711
transform -1 0 5448 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_64
timestamp 1515882711
transform -1 0 5640 0 -1 3810
box 0 0 192 200
use FILL  FILL_NAND2X1_44
timestamp 1515882711
transform 1 0 5640 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_44
timestamp 1515882711
transform 1 0 5656 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_64
timestamp 1515882711
transform -1 0 5768 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_24
timestamp 1515882711
transform 1 0 5768 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_24
timestamp 1515882711
transform 1 0 5784 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_379
timestamp 1515882711
transform 1 0 5976 0 -1 3810
box 0 0 64 200
use FILL  FILL_18_5_0
timestamp 1515882711
transform -1 0 6056 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_5_1
timestamp 1515882711
transform -1 0 6072 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_397
timestamp 1515882711
transform -1 0 6120 0 -1 3810
box 0 0 48 200
use FILL  FILL_MUX2X1_29
timestamp 1515882711
transform -1 0 6136 0 -1 3810
box 0 0 16 200
use MUX2X1  MUX2X1_29
timestamp 1515882711
transform -1 0 6232 0 -1 3810
box 0 0 96 200
use NOR2X1  NOR2X1_18
timestamp 1515882711
transform -1 0 6280 0 -1 3810
box 0 0 48 200
use NOR3X1  NOR3X1_17
timestamp 1515882711
transform 1 0 6280 0 -1 3810
box 0 0 128 200
use NOR2X1  NOR2X1_17
timestamp 1515882711
transform -1 0 6456 0 -1 3810
box 0 0 48 200
use OAI22X1  OAI22X1_4
timestamp 1515882711
transform 1 0 6456 0 -1 3810
box 0 0 80 200
use NOR2X1  NOR2X1_64
timestamp 1515882711
transform -1 0 6584 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_308
timestamp 1515882711
transform 1 0 6584 0 -1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_347
timestamp 1515882711
transform -1 0 6664 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_347
timestamp 1515882711
transform -1 0 6712 0 -1 3810
box 0 0 48 200
use FILL  FILL_NAND2X1_275
timestamp 1515882711
transform -1 0 6728 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_275
timestamp 1515882711
transform -1 0 6776 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_397
timestamp 1515882711
transform 1 0 6776 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_288
timestamp 1515882711
transform 1 0 6840 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_238
timestamp 1515882711
transform -1 0 6968 0 -1 3810
box 0 0 64 200
use FILL  FILL_INVX1_21
timestamp 1515882711
transform -1 0 6984 0 -1 3810
box 0 0 16 200
use INVX1  INVX1_21
timestamp 1515882711
transform -1 0 7016 0 -1 3810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_145
timestamp 1515882711
transform -1 0 7032 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_6_0
timestamp 1515882711
transform -1 0 7048 0 -1 3810
box 0 0 16 200
use FILL  FILL_18_6_1
timestamp 1515882711
transform -1 0 7064 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_145
timestamp 1515882711
transform -1 0 7256 0 -1 3810
box 0 0 192 200
use OAI21X1  OAI21X1_145
timestamp 1515882711
transform 1 0 7256 0 -1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_131
timestamp 1515882711
transform 1 0 7320 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_131
timestamp 1515882711
transform 1 0 7336 0 -1 3810
box 0 0 48 200
use FILL  FILL_BUFX4_262
timestamp 1515882711
transform -1 0 7400 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_262
timestamp 1515882711
transform -1 0 7464 0 -1 3810
box 0 0 64 200
use FILL  FILL_INVX1_60
timestamp 1515882711
transform 1 0 7464 0 -1 3810
box 0 0 16 200
use INVX1  INVX1_60
timestamp 1515882711
transform 1 0 7480 0 -1 3810
box 0 0 32 200
use OAI21X1  OAI21X1_307
timestamp 1515882711
transform 1 0 7512 0 -1 3810
box 0 0 64 200
use FILL  FILL_NAND2X1_274
timestamp 1515882711
transform 1 0 7576 0 -1 3810
box 0 0 16 200
use NAND2X1  NAND2X1_274
timestamp 1515882711
transform 1 0 7592 0 -1 3810
box 0 0 48 200
use OAI21X1  OAI21X1_7
timestamp 1515882711
transform 1 0 7640 0 -1 3810
box 0 0 64 200
use OAI21X1  OAI21X1_6
timestamp 1515882711
transform -1 0 7768 0 -1 3810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_292
timestamp 1515882711
transform 1 0 7768 0 -1 3810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_292
timestamp 1515882711
transform 1 0 7784 0 -1 3810
box 0 0 192 200
use FILL  FILL_BUFX4_261
timestamp 1515882711
transform -1 0 7992 0 -1 3810
box 0 0 16 200
use BUFX4  BUFX4_261
timestamp 1515882711
transform -1 0 8056 0 -1 3810
box 0 0 64 200
use BUFX2  BUFX2_38
timestamp 1515882711
transform -1 0 56 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_221
timestamp 1515882711
transform -1 0 72 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_221
timestamp 1515882711
transform -1 0 136 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX2_29
timestamp 1515882711
transform -1 0 152 0 1 3410
box 0 0 16 200
use BUFX2  BUFX2_29
timestamp 1515882711
transform -1 0 200 0 1 3410
box 0 0 48 200
use BUFX2  BUFX2_54
timestamp 1515882711
transform -1 0 248 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_151
timestamp 1515882711
transform 1 0 248 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_151
timestamp 1515882711
transform 1 0 264 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX2_15
timestamp 1515882711
transform -1 0 344 0 1 3410
box 0 0 16 200
use BUFX2  BUFX2_15
timestamp 1515882711
transform -1 0 392 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_220
timestamp 1515882711
transform 1 0 392 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_220
timestamp 1515882711
transform 1 0 408 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_148
timestamp 1515882711
transform -1 0 488 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_148
timestamp 1515882711
transform -1 0 552 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_55
timestamp 1515882711
transform -1 0 568 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_55
timestamp 1515882711
transform -1 0 632 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_173
timestamp 1515882711
transform -1 0 648 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_173
timestamp 1515882711
transform -1 0 712 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_56
timestamp 1515882711
transform 1 0 712 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_56
timestamp 1515882711
transform 1 0 728 0 1 3410
box 0 0 64 200
use FILL  FILL_INVX2_5
timestamp 1515882711
transform 1 0 792 0 1 3410
box 0 0 16 200
use INVX2  INVX2_5
timestamp 1515882711
transform 1 0 808 0 1 3410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_188
timestamp 1515882711
transform -1 0 856 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_0
timestamp 1515882711
transform -1 0 872 0 1 3410
box 0 0 16 200
use FILL  FILL_17_0_1
timestamp 1515882711
transform -1 0 888 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_188
timestamp 1515882711
transform -1 0 1080 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_172
timestamp 1515882711
transform 1 0 1080 0 1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_156
timestamp 1515882711
transform -1 0 1160 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_156
timestamp 1515882711
transform -1 0 1208 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_17
timestamp 1515882711
transform 1 0 1208 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_17
timestamp 1515882711
transform 1 0 1224 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_182
timestamp 1515882711
transform 1 0 1288 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_182
timestamp 1515882711
transform 1 0 1304 0 1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_217
timestamp 1515882711
transform 1 0 1368 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_217
timestamp 1515882711
transform 1 0 1384 0 1 3410
box 0 0 192 200
use FILL  FILL_AOI21X1_33
timestamp 1515882711
transform -1 0 1592 0 1 3410
box 0 0 16 200
use AOI21X1  AOI21X1_33
timestamp 1515882711
transform -1 0 1656 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_171
timestamp 1515882711
transform -1 0 1720 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_314
timestamp 1515882711
transform 1 0 1720 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_172
timestamp 1515882711
transform -1 0 1848 0 1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_221
timestamp 1515882711
transform -1 0 1864 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_0
timestamp 1515882711
transform -1 0 1880 0 1 3410
box 0 0 16 200
use FILL  FILL_17_1_1
timestamp 1515882711
transform -1 0 1896 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_221
timestamp 1515882711
transform -1 0 2088 0 1 3410
box 0 0 192 200
use NAND3X1  NAND3X1_315
timestamp 1515882711
transform -1 0 2152 0 1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_130
timestamp 1515882711
transform 1 0 2152 0 1 3410
box 0 0 48 200
use FILL  FILL_AOI21X1_54
timestamp 1515882711
transform -1 0 2216 0 1 3410
box 0 0 16 200
use AOI21X1  AOI21X1_54
timestamp 1515882711
transform -1 0 2280 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_115
timestamp 1515882711
transform -1 0 2296 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_115
timestamp 1515882711
transform -1 0 2360 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_219
timestamp 1515882711
transform -1 0 2376 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_219
timestamp 1515882711
transform -1 0 2440 0 1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_230
timestamp 1515882711
transform 1 0 2440 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_230
timestamp 1515882711
transform 1 0 2456 0 1 3410
box 0 0 48 200
use NOR2X1  NOR2X1_163
timestamp 1515882711
transform -1 0 2552 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_7
timestamp 1515882711
transform -1 0 2568 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_7
timestamp 1515882711
transform -1 0 2632 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_256
timestamp 1515882711
transform -1 0 2648 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_256
timestamp 1515882711
transform -1 0 2712 0 1 3410
box 0 0 64 200
use FILL  FILL_INVX8_4
timestamp 1515882711
transform -1 0 2728 0 1 3410
box 0 0 16 200
use INVX8  INVX8_4
timestamp 1515882711
transform -1 0 2808 0 1 3410
box 0 0 80 200
use NAND3X1  NAND3X1_155
timestamp 1515882711
transform -1 0 2872 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_298
timestamp 1515882711
transform -1 0 2936 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_59
timestamp 1515882711
transform 1 0 2936 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_0
timestamp 1515882711
transform 1 0 2952 0 1 3410
box 0 0 16 200
use FILL  FILL_17_2_1
timestamp 1515882711
transform 1 0 2968 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_59
timestamp 1515882711
transform 1 0 2984 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_22
timestamp 1515882711
transform 1 0 3048 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_199
timestamp 1515882711
transform 1 0 3112 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_39
timestamp 1515882711
transform 1 0 3176 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_39
timestamp 1515882711
transform 1 0 3192 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_180
timestamp 1515882711
transform 1 0 3256 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_3
timestamp 1515882711
transform 1 0 3320 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_23
timestamp 1515882711
transform 1 0 3384 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_25
timestamp 1515882711
transform -1 0 3512 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_202
timestamp 1515882711
transform 1 0 3512 0 1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_200
timestamp 1515882711
transform 1 0 3576 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_176
timestamp 1515882711
transform 1 0 3640 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_176
timestamp 1515882711
transform 1 0 3656 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_116
timestamp 1515882711
transform 1 0 3720 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_116
timestamp 1515882711
transform 1 0 3736 0 1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_184
timestamp 1515882711
transform 1 0 3800 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_184
timestamp 1515882711
transform 1 0 3816 0 1 3410
box 0 0 48 200
use FILL  FILL_NAND2X1_186
timestamp 1515882711
transform 1 0 3864 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_186
timestamp 1515882711
transform 1 0 3880 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_156
timestamp 1515882711
transform 1 0 3928 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_156
timestamp 1515882711
transform 1 0 3944 0 1 3410
box 0 0 64 200
use FILL  FILL_17_3_0
timestamp 1515882711
transform -1 0 4024 0 1 3410
box 0 0 16 200
use FILL  FILL_17_3_1
timestamp 1515882711
transform -1 0 4040 0 1 3410
box 0 0 16 200
use FILL  FILL_INVX1_26
timestamp 1515882711
transform -1 0 4056 0 1 3410
box 0 0 16 200
use INVX1  INVX1_26
timestamp 1515882711
transform -1 0 4088 0 1 3410
box 0 0 32 200
use FILL  FILL_NAND2X1_29
timestamp 1515882711
transform -1 0 4104 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_29
timestamp 1515882711
transform -1 0 4152 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_50
timestamp 1515882711
transform -1 0 4216 0 1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_50
timestamp 1515882711
transform 1 0 4216 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_50
timestamp 1515882711
transform 1 0 4232 0 1 3410
box 0 0 192 200
use FILL  FILL_INVX1_79
timestamp 1515882711
transform 1 0 4424 0 1 3410
box 0 0 16 200
use INVX1  INVX1_79
timestamp 1515882711
transform 1 0 4440 0 1 3410
box 0 0 32 200
use OAI21X1  OAI21X1_341
timestamp 1515882711
transform 1 0 4472 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_264
timestamp 1515882711
transform -1 0 4552 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_264
timestamp 1515882711
transform -1 0 4616 0 1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_233
timestamp 1515882711
transform 1 0 4616 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_233
timestamp 1515882711
transform 1 0 4632 0 1 3410
box 0 0 48 200
use FILL  FILL_INVX1_81
timestamp 1515882711
transform -1 0 4696 0 1 3410
box 0 0 16 200
use INVX1  INVX1_81
timestamp 1515882711
transform -1 0 4728 0 1 3410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_21
timestamp 1515882711
transform -1 0 4744 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_21
timestamp 1515882711
transform -1 0 4936 0 1 3410
box 0 0 192 200
use NAND2X1  NAND2X1_420
timestamp 1515882711
transform 1 0 4936 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_445
timestamp 1515882711
transform -1 0 5048 0 1 3410
box 0 0 64 200
use FILL  FILL_17_4_0
timestamp 1515882711
transform 1 0 5048 0 1 3410
box 0 0 16 200
use FILL  FILL_17_4_1
timestamp 1515882711
transform 1 0 5064 0 1 3410
box 0 0 16 200
use FILL  FILL_BUFX4_13
timestamp 1515882711
transform 1 0 5080 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_13
timestamp 1515882711
transform 1 0 5096 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_295
timestamp 1515882711
transform -1 0 5176 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_295
timestamp 1515882711
transform -1 0 5240 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_218
timestamp 1515882711
transform 1 0 5240 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_218
timestamp 1515882711
transform 1 0 5256 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_314
timestamp 1515882711
transform -1 0 5384 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_294
timestamp 1515882711
transform -1 0 5448 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_263
timestamp 1515882711
transform 1 0 5448 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_263
timestamp 1515882711
transform 1 0 5464 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_305
timestamp 1515882711
transform 1 0 5528 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_305
timestamp 1515882711
transform 1 0 5544 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_320
timestamp 1515882711
transform 1 0 5608 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_320
timestamp 1515882711
transform 1 0 5624 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_83
timestamp 1515882711
transform -1 0 5704 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_83
timestamp 1515882711
transform -1 0 5768 0 1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_99
timestamp 1515882711
transform 1 0 5768 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_99
timestamp 1515882711
transform 1 0 5784 0 1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_99
timestamp 1515882711
transform 1 0 5976 0 1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_82
timestamp 1515882711
transform -1 0 6056 0 1 3410
box 0 0 16 200
use FILL  FILL_17_5_0
timestamp 1515882711
transform -1 0 6072 0 1 3410
box 0 0 16 200
use FILL  FILL_17_5_1
timestamp 1515882711
transform -1 0 6088 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_82
timestamp 1515882711
transform -1 0 6136 0 1 3410
box 0 0 48 200
use FILL  FILL_BUFX4_112
timestamp 1515882711
transform -1 0 6152 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_112
timestamp 1515882711
transform -1 0 6216 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_299
timestamp 1515882711
transform 1 0 6216 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_299
timestamp 1515882711
transform 1 0 6232 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_298
timestamp 1515882711
transform 1 0 6296 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_298
timestamp 1515882711
transform 1 0 6312 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_88
timestamp 1515882711
transform 1 0 6376 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_88
timestamp 1515882711
transform 1 0 6392 0 1 3410
box 0 0 64 200
use FILL  FILL_MUX2X1_28
timestamp 1515882711
transform 1 0 6456 0 1 3410
box 0 0 16 200
use MUX2X1  MUX2X1_28
timestamp 1515882711
transform 1 0 6472 0 1 3410
box 0 0 96 200
use NAND2X1  NAND2X1_416
timestamp 1515882711
transform 1 0 6568 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_471
timestamp 1515882711
transform -1 0 6680 0 1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_284
timestamp 1515882711
transform 1 0 6680 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_284
timestamp 1515882711
transform 1 0 6696 0 1 3410
box 0 0 192 200
use FILL  FILL_NAND2X1_219
timestamp 1515882711
transform -1 0 6904 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_219
timestamp 1515882711
transform -1 0 6952 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_504
timestamp 1515882711
transform 1 0 6952 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_502
timestamp 1515882711
transform -1 0 7080 0 1 3410
box 0 0 64 200
use FILL  FILL_17_6_0
timestamp 1515882711
transform -1 0 7096 0 1 3410
box 0 0 16 200
use FILL  FILL_17_6_1
timestamp 1515882711
transform -1 0 7112 0 1 3410
box 0 0 16 200
use FILL  FILL_MUX2X1_24
timestamp 1515882711
transform -1 0 7128 0 1 3410
box 0 0 16 200
use MUX2X1  MUX2X1_24
timestamp 1515882711
transform -1 0 7224 0 1 3410
box 0 0 96 200
use OAI21X1  OAI21X1_338
timestamp 1515882711
transform 1 0 7224 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_34
timestamp 1515882711
transform 1 0 7288 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_34
timestamp 1515882711
transform 1 0 7304 0 1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_297
timestamp 1515882711
transform 1 0 7368 0 1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_297
timestamp 1515882711
transform 1 0 7384 0 1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_12
timestamp 1515882711
transform 1 0 7432 0 1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_14
timestamp 1515882711
transform -1 0 7560 0 1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_295
timestamp 1515882711
transform -1 0 7576 0 1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_295
timestamp 1515882711
transform -1 0 7768 0 1 3410
box 0 0 192 200
use FILL  FILL_BUFX4_36
timestamp 1515882711
transform 1 0 7768 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_36
timestamp 1515882711
transform 1 0 7784 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_154
timestamp 1515882711
transform -1 0 7864 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_154
timestamp 1515882711
transform -1 0 7928 0 1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_155
timestamp 1515882711
transform 1 0 7928 0 1 3410
box 0 0 16 200
use BUFX4  BUFX4_155
timestamp 1515882711
transform 1 0 7944 0 1 3410
box 0 0 64 200
use FILL  FILL_18_1
timestamp 1515882711
transform 1 0 8008 0 1 3410
box 0 0 16 200
use FILL  FILL_18_2
timestamp 1515882711
transform 1 0 8024 0 1 3410
box 0 0 16 200
use FILL  FILL_18_3
timestamp 1515882711
transform 1 0 8040 0 1 3410
box 0 0 16 200
use FILL  FILL_BUFX4_57
timestamp 1515882711
transform -1 0 24 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_57
timestamp 1515882711
transform -1 0 88 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_136
timestamp 1515882711
transform -1 0 104 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_136
timestamp 1515882711
transform -1 0 168 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_19
timestamp 1515882711
transform -1 0 232 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_21
timestamp 1515882711
transform -1 0 296 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_18
timestamp 1515882711
transform 1 0 296 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_195
timestamp 1515882711
transform 1 0 360 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_196
timestamp 1515882711
transform 1 0 424 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_239
timestamp 1515882711
transform -1 0 504 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_239
timestamp 1515882711
transform -1 0 568 0 -1 3410
box 0 0 64 200
use NOR3X1  NOR3X1_16
timestamp 1515882711
transform -1 0 696 0 -1 3410
box 0 0 128 200
use OAI21X1  OAI21X1_306
timestamp 1515882711
transform -1 0 760 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_16
timestamp 1515882711
transform -1 0 824 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_305
timestamp 1515882711
transform -1 0 888 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_405
timestamp 1515882711
transform -1 0 952 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_0_0
timestamp 1515882711
transform -1 0 968 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_0_1
timestamp 1515882711
transform -1 0 984 0 -1 3410
box 0 0 16 200
use OAI21X1  OAI21X1_404
timestamp 1515882711
transform -1 0 1048 0 -1 3410
box 0 0 64 200
use NOR3X1  NOR3X1_39
timestamp 1515882711
transform 1 0 1048 0 -1 3410
box 0 0 128 200
use NAND3X1  NAND3X1_141
timestamp 1515882711
transform 1 0 1176 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_284
timestamp 1515882711
transform 1 0 1240 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_143
timestamp 1515882711
transform 1 0 1304 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_286
timestamp 1515882711
transform 1 0 1368 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_317
timestamp 1515882711
transform -1 0 1496 0 -1 3410
box 0 0 64 200
use NAND3X1  NAND3X1_174
timestamp 1515882711
transform 1 0 1496 0 -1 3410
box 0 0 64 200
use NOR2X1  NOR2X1_109
timestamp 1515882711
transform -1 0 1608 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_319
timestamp 1515882711
transform 1 0 1608 0 -1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_200
timestamp 1515882711
transform -1 0 1688 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_200
timestamp 1515882711
transform -1 0 1880 0 -1 3410
box 0 0 192 200
use FILL  FILL_BUFX4_317
timestamp 1515882711
transform -1 0 1896 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_317
timestamp 1515882711
transform -1 0 1960 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_1_0
timestamp 1515882711
transform -1 0 1976 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_1_1
timestamp 1515882711
transform -1 0 1992 0 -1 3410
box 0 0 16 200
use FILL  FILL_BUFX4_90
timestamp 1515882711
transform -1 0 2008 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_90
timestamp 1515882711
transform -1 0 2072 0 -1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_271
timestamp 1515882711
transform 1 0 2072 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_271
timestamp 1515882711
transform 1 0 2088 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_22
timestamp 1515882711
transform 1 0 2280 0 -1 3410
box 0 0 64 200
use NAND2X1  NAND2X1_451
timestamp 1515882711
transform -1 0 2392 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_250
timestamp 1515882711
transform 1 0 2392 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_252
timestamp 1515882711
transform 1 0 2456 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_255
timestamp 1515882711
transform -1 0 2536 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_255
timestamp 1515882711
transform -1 0 2600 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_234
timestamp 1515882711
transform -1 0 2616 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_234
timestamp 1515882711
transform -1 0 2664 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_299
timestamp 1515882711
transform -1 0 2728 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_250
timestamp 1515882711
transform 1 0 2728 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_250
timestamp 1515882711
transform 1 0 2744 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_156
timestamp 1515882711
transform 1 0 2792 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_339
timestamp 1515882711
transform 1 0 2856 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_339
timestamp 1515882711
transform 1 0 2872 0 -1 3410
box 0 0 48 200
use NAND3X1  NAND3X1_158
timestamp 1515882711
transform -1 0 2984 0 -1 3410
box 0 0 64 200
use FILL  FILL_16_2_0
timestamp 1515882711
transform 1 0 2984 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_2_1
timestamp 1515882711
transform 1 0 3000 0 -1 3410
box 0 0 16 200
use FILL  FILL_NAND2X1_277
timestamp 1515882711
transform 1 0 3016 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_277
timestamp 1515882711
transform 1 0 3032 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_310
timestamp 1515882711
transform -1 0 3144 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_101
timestamp 1515882711
transform 1 0 3144 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_101
timestamp 1515882711
transform 1 0 3160 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_241
timestamp 1515882711
transform -1 0 3240 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_241
timestamp 1515882711
transform -1 0 3304 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_371
timestamp 1515882711
transform 1 0 3304 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_371
timestamp 1515882711
transform 1 0 3320 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_438
timestamp 1515882711
transform -1 0 3432 0 -1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_345
timestamp 1515882711
transform -1 0 3448 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_345
timestamp 1515882711
transform -1 0 3640 0 -1 3410
box 0 0 192 200
use FILL  FILL_BUFX4_98
timestamp 1515882711
transform -1 0 3656 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_98
timestamp 1515882711
transform -1 0 3720 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_99
timestamp 1515882711
transform -1 0 3736 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_99
timestamp 1515882711
transform -1 0 3800 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_160
timestamp 1515882711
transform 1 0 3800 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_160
timestamp 1515882711
transform 1 0 3816 0 -1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_56
timestamp 1515882711
transform 1 0 3880 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_56
timestamp 1515882711
transform 1 0 3896 0 -1 3410
box 0 0 192 200
use FILL  FILL_16_3_0
timestamp 1515882711
transform 1 0 4088 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_3_1
timestamp 1515882711
transform 1 0 4104 0 -1 3410
box 0 0 16 200
use FILL  FILL_NAND2X1_37
timestamp 1515882711
transform 1 0 4120 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_37
timestamp 1515882711
transform 1 0 4136 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_56
timestamp 1515882711
transform -1 0 4248 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX2_22
timestamp 1515882711
transform -1 0 4264 0 -1 3410
box 0 0 16 200
use BUFX2  BUFX2_22
timestamp 1515882711
transform -1 0 4312 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_273
timestamp 1515882711
transform -1 0 4376 0 -1 3410
box 0 0 64 200
use FILL  FILL_INVX1_41
timestamp 1515882711
transform -1 0 4392 0 -1 3410
box 0 0 16 200
use INVX1  INVX1_41
timestamp 1515882711
transform -1 0 4424 0 -1 3410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_77
timestamp 1515882711
transform -1 0 4440 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_77
timestamp 1515882711
transform -1 0 4632 0 -1 3410
box 0 0 192 200
use FILL  FILL_NAND2X1_59
timestamp 1515882711
transform -1 0 4648 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_59
timestamp 1515882711
transform -1 0 4696 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_77
timestamp 1515882711
transform -1 0 4760 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_67
timestamp 1515882711
transform 1 0 4760 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_48
timestamp 1515882711
transform -1 0 4840 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_48
timestamp 1515882711
transform -1 0 4888 0 -1 3410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_67
timestamp 1515882711
transform -1 0 4904 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_67
timestamp 1515882711
transform -1 0 5096 0 -1 3410
box 0 0 192 200
use FILL  FILL_16_4_0
timestamp 1515882711
transform -1 0 5112 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_4_1
timestamp 1515882711
transform -1 0 5128 0 -1 3410
box 0 0 16 200
use FILL  FILL_BUFX4_9
timestamp 1515882711
transform -1 0 5144 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_9
timestamp 1515882711
transform -1 0 5208 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_300
timestamp 1515882711
transform 1 0 5208 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_300
timestamp 1515882711
transform 1 0 5224 0 -1 3410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_348
timestamp 1515882711
transform -1 0 5288 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_348
timestamp 1515882711
transform -1 0 5480 0 -1 3410
box 0 0 192 200
use FILL  FILL_NAND2X1_374
timestamp 1515882711
transform 1 0 5480 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_374
timestamp 1515882711
transform 1 0 5496 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_441
timestamp 1515882711
transform -1 0 5608 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_280
timestamp 1515882711
transform 1 0 5608 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_280
timestamp 1515882711
transform 1 0 5624 0 -1 3410
box 0 0 48 200
use FILL  FILL_NAND2X1_46
timestamp 1515882711
transform 1 0 5672 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_46
timestamp 1515882711
transform 1 0 5688 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_24
timestamp 1515882711
transform -1 0 5800 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_2
timestamp 1515882711
transform 1 0 5800 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_24
timestamp 1515882711
transform -1 0 5880 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_24
timestamp 1515882711
transform -1 0 5928 0 -1 3410
box 0 0 48 200
use FILL  FILL_NAND2X1_264
timestamp 1515882711
transform -1 0 5944 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_264
timestamp 1515882711
transform -1 0 5992 0 -1 3410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_27
timestamp 1515882711
transform -1 0 6008 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_5_0
timestamp 1515882711
transform -1 0 6024 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_5_1
timestamp 1515882711
transform -1 0 6040 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_27
timestamp 1515882711
transform -1 0 6232 0 -1 3410
box 0 0 192 200
use FILL  FILL_BUFX4_283
timestamp 1515882711
transform -1 0 6248 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_283
timestamp 1515882711
transform -1 0 6312 0 -1 3410
box 0 0 64 200
use FILL  FILL_BUFX4_91
timestamp 1515882711
transform 1 0 6312 0 -1 3410
box 0 0 16 200
use BUFX4  BUFX4_91
timestamp 1515882711
transform 1 0 6328 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_118
timestamp 1515882711
transform 1 0 6392 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_100
timestamp 1515882711
transform -1 0 6472 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_100
timestamp 1515882711
transform -1 0 6520 0 -1 3410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_118
timestamp 1515882711
transform -1 0 6536 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_118
timestamp 1515882711
transform -1 0 6728 0 -1 3410
box 0 0 192 200
use FILL  FILL_DFFPOSX1_327
timestamp 1515882711
transform -1 0 6744 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_327
timestamp 1515882711
transform -1 0 6936 0 -1 3410
box 0 0 192 200
use FILL  FILL_INVX1_23
timestamp 1515882711
transform 1 0 6936 0 -1 3410
box 0 0 16 200
use INVX1  INVX1_23
timestamp 1515882711
transform 1 0 6952 0 -1 3410
box 0 0 32 200
use FILL  FILL_NAND2X1_260
timestamp 1515882711
transform -1 0 7000 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_260
timestamp 1515882711
transform -1 0 7048 0 -1 3410
box 0 0 48 200
use FILL  FILL_NAND2X1_342
timestamp 1515882711
transform -1 0 7064 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_6_0
timestamp 1515882711
transform -1 0 7080 0 -1 3410
box 0 0 16 200
use FILL  FILL_16_6_1
timestamp 1515882711
transform -1 0 7096 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_342
timestamp 1515882711
transform -1 0 7144 0 -1 3410
box 0 0 48 200
use FILL  FILL_NAND2X1_118
timestamp 1515882711
transform 1 0 7144 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_118
timestamp 1515882711
transform 1 0 7160 0 -1 3410
box 0 0 48 200
use OAI21X1  OAI21X1_133
timestamp 1515882711
transform -1 0 7272 0 -1 3410
box 0 0 64 200
use OAI21X1  OAI21X1_156
timestamp 1515882711
transform -1 0 7336 0 -1 3410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_133
timestamp 1515882711
transform -1 0 7352 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_133
timestamp 1515882711
transform -1 0 7544 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_151
timestamp 1515882711
transform 1 0 7544 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_137
timestamp 1515882711
transform -1 0 7624 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_137
timestamp 1515882711
transform -1 0 7672 0 -1 3410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_151
timestamp 1515882711
transform 1 0 7672 0 -1 3410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_151
timestamp 1515882711
transform 1 0 7688 0 -1 3410
box 0 0 192 200
use OAI21X1  OAI21X1_287
timestamp 1515882711
transform 1 0 7880 0 -1 3410
box 0 0 64 200
use FILL  FILL_NAND2X1_259
timestamp 1515882711
transform -1 0 7960 0 -1 3410
box 0 0 16 200
use NAND2X1  NAND2X1_259
timestamp 1515882711
transform -1 0 8008 0 -1 3410
box 0 0 48 200
use FILL  FILL_17_1
timestamp 1515882711
transform -1 0 8024 0 -1 3410
box 0 0 16 200
use FILL  FILL_17_2
timestamp 1515882711
transform -1 0 8040 0 -1 3410
box 0 0 16 200
use FILL  FILL_17_3
timestamp 1515882711
transform -1 0 8056 0 -1 3410
box 0 0 16 200
use FILL  FILL_NAND2X1_181
timestamp 1515882711
transform 1 0 8 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_181
timestamp 1515882711
transform 1 0 24 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_139
timestamp 1515882711
transform -1 0 120 0 1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_20
timestamp 1515882711
transform -1 0 184 0 1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_260
timestamp 1515882711
transform 1 0 184 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_260
timestamp 1515882711
transform 1 0 200 0 1 3010
box 0 0 192 200
use NAND3X1  NAND3X1_198
timestamp 1515882711
transform 1 0 392 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_213
timestamp 1515882711
transform -1 0 472 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_213
timestamp 1515882711
transform -1 0 536 0 1 3010
box 0 0 64 200
use FILL  FILL_INVX8_9
timestamp 1515882711
transform 1 0 536 0 1 3010
box 0 0 16 200
use INVX8  INVX8_9
timestamp 1515882711
transform 1 0 552 0 1 3010
box 0 0 80 200
use NAND3X1  NAND3X1_17
timestamp 1515882711
transform -1 0 696 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_170
timestamp 1515882711
transform -1 0 712 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_170
timestamp 1515882711
transform -1 0 776 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_193
timestamp 1515882711
transform -1 0 840 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_194
timestamp 1515882711
transform 1 0 840 0 1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_165
timestamp 1515882711
transform 1 0 904 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_0
timestamp 1515882711
transform 1 0 920 0 1 3010
box 0 0 16 200
use FILL  FILL_15_0_1
timestamp 1515882711
transform 1 0 936 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_165
timestamp 1515882711
transform 1 0 952 0 1 3010
box 0 0 192 200
use FILL  FILL_AOI21X1_16
timestamp 1515882711
transform -1 0 1160 0 1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_16
timestamp 1515882711
transform -1 0 1224 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_283
timestamp 1515882711
transform -1 0 1288 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_140
timestamp 1515882711
transform 1 0 1288 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_142
timestamp 1515882711
transform -1 0 1416 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_285
timestamp 1515882711
transform 1 0 1416 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_173
timestamp 1515882711
transform -1 0 1544 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_176
timestamp 1515882711
transform 1 0 1544 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_316
timestamp 1515882711
transform 1 0 1608 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_318
timestamp 1515882711
transform 1 0 1672 0 1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_254
timestamp 1515882711
transform -1 0 1752 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_254
timestamp 1515882711
transform -1 0 1944 0 1 3010
box 0 0 192 200
use FILL  FILL_15_1_0
timestamp 1515882711
transform 1 0 1944 0 1 3010
box 0 0 16 200
use FILL  FILL_15_1_1
timestamp 1515882711
transform 1 0 1960 0 1 3010
box 0 0 16 200
use NOR2X1  NOR2X1_68
timestamp 1515882711
transform 1 0 1976 0 1 3010
box 0 0 48 200
use FILL  FILL_AOI21X1_62
timestamp 1515882711
transform -1 0 2040 0 1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_62
timestamp 1515882711
transform -1 0 2104 0 1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_180
timestamp 1515882711
transform -1 0 2120 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_180
timestamp 1515882711
transform -1 0 2168 0 1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_258
timestamp 1515882711
transform -1 0 2184 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_258
timestamp 1515882711
transform -1 0 2376 0 1 3010
box 0 0 192 200
use NOR2X1  NOR2X1_52
timestamp 1515882711
transform 1 0 2376 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_381
timestamp 1515882711
transform 1 0 2424 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_276
timestamp 1515882711
transform 1 0 2488 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_279
timestamp 1515882711
transform -1 0 2616 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_277
timestamp 1515882711
transform -1 0 2680 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_309
timestamp 1515882711
transform -1 0 2696 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_309
timestamp 1515882711
transform -1 0 2760 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_301
timestamp 1515882711
transform -1 0 2824 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_79
timestamp 1515882711
transform -1 0 2840 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_79
timestamp 1515882711
transform -1 0 2904 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_236
timestamp 1515882711
transform 1 0 2904 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_236
timestamp 1515882711
transform 1 0 2920 0 1 3010
box 0 0 64 200
use FILL  FILL_15_2_0
timestamp 1515882711
transform 1 0 2984 0 1 3010
box 0 0 16 200
use FILL  FILL_15_2_1
timestamp 1515882711
transform 1 0 3000 0 1 3010
box 0 0 16 200
use FILL  FILL_NAND2X1_189
timestamp 1515882711
transform 1 0 3016 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_189
timestamp 1515882711
transform 1 0 3032 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_146
timestamp 1515882711
transform 1 0 3080 0 1 3010
box 0 0 48 200
use FILL  FILL_INVX1_62
timestamp 1515882711
transform -1 0 3144 0 1 3010
box 0 0 16 200
use INVX1  INVX1_62
timestamp 1515882711
transform -1 0 3176 0 1 3010
box 0 0 32 200
use FILL  FILL_NAND2X1_231
timestamp 1515882711
transform 1 0 3176 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_231
timestamp 1515882711
transform 1 0 3192 0 1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_338
timestamp 1515882711
transform 1 0 3240 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_338
timestamp 1515882711
transform 1 0 3256 0 1 3010
box 0 0 192 200
use FILL  FILL_NAND2X1_364
timestamp 1515882711
transform 1 0 3448 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_364
timestamp 1515882711
transform 1 0 3464 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_431
timestamp 1515882711
transform -1 0 3576 0 1 3010
box 0 0 64 200
use FILL  FILL_INVX1_67
timestamp 1515882711
transform 1 0 3576 0 1 3010
box 0 0 16 200
use INVX1  INVX1_67
timestamp 1515882711
transform 1 0 3592 0 1 3010
box 0 0 32 200
use FILL  FILL_NAND2X1_232
timestamp 1515882711
transform 1 0 3624 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_232
timestamp 1515882711
transform 1 0 3640 0 1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_135
timestamp 1515882711
transform -1 0 3704 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_135
timestamp 1515882711
transform -1 0 3896 0 1 3010
box 0 0 192 200
use FILL  FILL_NAND2X1_168
timestamp 1515882711
transform 1 0 3896 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_168
timestamp 1515882711
transform 1 0 3912 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_135
timestamp 1515882711
transform -1 0 4024 0 1 3010
box 0 0 64 200
use FILL  FILL_15_3_0
timestamp 1515882711
transform 1 0 4024 0 1 3010
box 0 0 16 200
use FILL  FILL_15_3_1
timestamp 1515882711
transform 1 0 4040 0 1 3010
box 0 0 16 200
use FILL  FILL_NAND2X1_185
timestamp 1515882711
transform 1 0 4056 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_185
timestamp 1515882711
transform 1 0 4072 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_313
timestamp 1515882711
transform -1 0 4184 0 1 3010
box 0 0 64 200
use FILL  FILL_INVX1_63
timestamp 1515882711
transform 1 0 4184 0 1 3010
box 0 0 16 200
use INVX1  INVX1_63
timestamp 1515882711
transform 1 0 4200 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_58
timestamp 1515882711
transform 1 0 4232 0 1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_38
timestamp 1515882711
transform -1 0 4312 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_38
timestamp 1515882711
transform -1 0 4360 0 1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_58
timestamp 1515882711
transform 1 0 4360 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_58
timestamp 1515882711
transform 1 0 4376 0 1 3010
box 0 0 192 200
use FILL  FILL_INVX1_31
timestamp 1515882711
transform 1 0 4568 0 1 3010
box 0 0 16 200
use INVX1  INVX1_31
timestamp 1515882711
transform 1 0 4584 0 1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_254
timestamp 1515882711
transform 1 0 4616 0 1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_248
timestamp 1515882711
transform -1 0 4696 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_248
timestamp 1515882711
transform -1 0 4744 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_157
timestamp 1515882711
transform -1 0 4808 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_75
timestamp 1515882711
transform -1 0 4824 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_75
timestamp 1515882711
transform -1 0 4888 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_2
timestamp 1515882711
transform -1 0 4904 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_2
timestamp 1515882711
transform -1 0 4968 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_73
timestamp 1515882711
transform -1 0 4984 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_73
timestamp 1515882711
transform -1 0 5048 0 1 3010
box 0 0 64 200
use FILL  FILL_15_4_0
timestamp 1515882711
transform 1 0 5048 0 1 3010
box 0 0 16 200
use FILL  FILL_15_4_1
timestamp 1515882711
transform 1 0 5064 0 1 3010
box 0 0 16 200
use FILL  FILL_BUFX4_103
timestamp 1515882711
transform 1 0 5080 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_103
timestamp 1515882711
transform 1 0 5096 0 1 3010
box 0 0 64 200
use FILL  FILL_AND2X2_2
timestamp 1515882711
transform -1 0 5176 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_2
timestamp 1515882711
transform -1 0 5240 0 1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_101
timestamp 1515882711
transform -1 0 5256 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_101
timestamp 1515882711
transform -1 0 5304 0 1 3010
box 0 0 48 200
use FILL  FILL_NAND2X1_50
timestamp 1515882711
transform -1 0 5320 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_50
timestamp 1515882711
transform -1 0 5368 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_78
timestamp 1515882711
transform 1 0 5368 0 1 3010
box 0 0 48 200
use FILL  FILL_INVX1_53
timestamp 1515882711
transform -1 0 5432 0 1 3010
box 0 0 16 200
use INVX1  INVX1_53
timestamp 1515882711
transform -1 0 5464 0 1 3010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_62
timestamp 1515882711
transform -1 0 5480 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_62
timestamp 1515882711
transform -1 0 5672 0 1 3010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_29
timestamp 1515882711
transform -1 0 5688 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_29
timestamp 1515882711
transform -1 0 5880 0 1 3010
box 0 0 192 200
use FILL  FILL_AND2X2_5
timestamp 1515882711
transform -1 0 5896 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_5
timestamp 1515882711
transform -1 0 5960 0 1 3010
box 0 0 64 200
use FILL  FILL_INVX2_1
timestamp 1515882711
transform 1 0 5960 0 1 3010
box 0 0 16 200
use INVX2  INVX2_1
timestamp 1515882711
transform 1 0 5976 0 1 3010
box 0 0 32 200
use FILL  FILL_BUFX4_209
timestamp 1515882711
transform 1 0 6008 0 1 3010
box 0 0 16 200
use FILL  FILL_15_5_0
timestamp 1515882711
transform 1 0 6024 0 1 3010
box 0 0 16 200
use FILL  FILL_15_5_1
timestamp 1515882711
transform 1 0 6040 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_209
timestamp 1515882711
transform 1 0 6056 0 1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_1
timestamp 1515882711
transform -1 0 6136 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_1
timestamp 1515882711
transform -1 0 6184 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_444
timestamp 1515882711
transform -1 0 6232 0 1 3010
box 0 0 48 200
use FILL  FILL_INVX1_12
timestamp 1515882711
transform -1 0 6248 0 1 3010
box 0 0 16 200
use INVX1  INVX1_12
timestamp 1515882711
transform -1 0 6280 0 1 3010
box 0 0 32 200
use FILL  FILL_NAND2X1_290
timestamp 1515882711
transform -1 0 6296 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_290
timestamp 1515882711
transform -1 0 6344 0 1 3010
box 0 0 48 200
use FILL  FILL_INVX1_1
timestamp 1515882711
transform -1 0 6360 0 1 3010
box 0 0 16 200
use INVX1  INVX1_1
timestamp 1515882711
transform -1 0 6392 0 1 3010
box 0 0 32 200
use FILL  FILL_BUFX4_71
timestamp 1515882711
transform -1 0 6408 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_71
timestamp 1515882711
transform -1 0 6472 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_422
timestamp 1515882711
transform 1 0 6472 0 1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_111
timestamp 1515882711
transform -1 0 6568 0 1 3010
box 0 0 48 200
use FILL  FILL_AND2X2_6
timestamp 1515882711
transform -1 0 6584 0 1 3010
box 0 0 16 200
use AND2X2  AND2X2_6
timestamp 1515882711
transform -1 0 6648 0 1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_423
timestamp 1515882711
transform -1 0 6696 0 1 3010
box 0 0 48 200
use FILL  FILL_NAND2X1_106
timestamp 1515882711
transform 1 0 6696 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_106
timestamp 1515882711
transform 1 0 6712 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_441
timestamp 1515882711
transform 1 0 6760 0 1 3010
box 0 0 48 200
use FILL  FILL_INVX4_1
timestamp 1515882711
transform -1 0 6824 0 1 3010
box 0 0 16 200
use INVX4  INVX4_1
timestamp 1515882711
transform -1 0 6872 0 1 3010
box 0 0 48 200
use FILL  FILL_BUFX4_192
timestamp 1515882711
transform 1 0 6872 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_192
timestamp 1515882711
transform 1 0 6888 0 1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_126
timestamp 1515882711
transform -1 0 6968 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_126
timestamp 1515882711
transform -1 0 7016 0 1 3010
box 0 0 48 200
use FILL  FILL_INVX1_76
timestamp 1515882711
transform 1 0 7016 0 1 3010
box 0 0 16 200
use INVX1  INVX1_76
timestamp 1515882711
transform 1 0 7032 0 1 3010
box 0 0 32 200
use FILL  FILL_NAND2X1_142
timestamp 1515882711
transform 1 0 7064 0 1 3010
box 0 0 16 200
use FILL  FILL_15_6_0
timestamp 1515882711
transform 1 0 7080 0 1 3010
box 0 0 16 200
use FILL  FILL_15_6_1
timestamp 1515882711
transform 1 0 7096 0 1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_142
timestamp 1515882711
transform 1 0 7112 0 1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_156
timestamp 1515882711
transform -1 0 7176 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_156
timestamp 1515882711
transform -1 0 7368 0 1 3010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_290
timestamp 1515882711
transform 1 0 7368 0 1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_290
timestamp 1515882711
transform 1 0 7384 0 1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_3
timestamp 1515882711
transform 1 0 7576 0 1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_513
timestamp 1515882711
transform 1 0 7640 0 1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_122
timestamp 1515882711
transform 1 0 7704 0 1 3010
box 0 0 48 200
use NAND2X1  NAND2X1_443
timestamp 1515882711
transform -1 0 7800 0 1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_159
timestamp 1515882711
transform -1 0 7864 0 1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_1
timestamp 1515882711
transform 1 0 7864 0 1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_259
timestamp 1515882711
transform 1 0 7928 0 1 3010
box 0 0 16 200
use BUFX4  BUFX4_259
timestamp 1515882711
transform 1 0 7944 0 1 3010
box 0 0 64 200
use FILL  FILL_16_1
timestamp 1515882711
transform 1 0 8008 0 1 3010
box 0 0 16 200
use FILL  FILL_16_2
timestamp 1515882711
transform 1 0 8024 0 1 3010
box 0 0 16 200
use FILL  FILL_16_3
timestamp 1515882711
transform 1 0 8040 0 1 3010
box 0 0 16 200
use FILL  FILL_INVX1_56
timestamp 1515882711
transform 1 0 8 0 -1 3010
box 0 0 16 200
use INVX1  INVX1_56
timestamp 1515882711
transform 1 0 24 0 -1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_141
timestamp 1515882711
transform -1 0 104 0 -1 3010
box 0 0 48 200
use FILL  FILL_INVX1_45
timestamp 1515882711
transform 1 0 104 0 -1 3010
box 0 0 16 200
use INVX1  INVX1_45
timestamp 1515882711
transform 1 0 120 0 -1 3010
box 0 0 32 200
use NOR2X1  NOR2X1_140
timestamp 1515882711
transform -1 0 200 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_80
timestamp 1515882711
transform 1 0 200 0 -1 3010
box 0 0 48 200
use FILL  FILL_AOI21X1_4
timestamp 1515882711
transform -1 0 264 0 -1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_4
timestamp 1515882711
transform -1 0 328 0 -1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_211
timestamp 1515882711
transform -1 0 344 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_211
timestamp 1515882711
transform -1 0 408 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_142
timestamp 1515882711
transform -1 0 456 0 -1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_206
timestamp 1515882711
transform 1 0 456 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_206
timestamp 1515882711
transform 1 0 472 0 -1 3010
box 0 0 192 200
use FILL  FILL_AOI21X1_39
timestamp 1515882711
transform 1 0 664 0 -1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_39
timestamp 1515882711
transform 1 0 680 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_115
timestamp 1515882711
transform -1 0 792 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_95
timestamp 1515882711
transform -1 0 840 0 -1 3010
box 0 0 48 200
use FILL  FILL_AOI21X1_19
timestamp 1515882711
transform -1 0 856 0 -1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_19
timestamp 1515882711
transform -1 0 920 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_169
timestamp 1515882711
transform 1 0 920 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_0
timestamp 1515882711
transform 1 0 936 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_0_1
timestamp 1515882711
transform 1 0 952 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_169
timestamp 1515882711
transform 1 0 968 0 -1 3010
box 0 0 192 200
use NOR2X1  NOR2X1_92
timestamp 1515882711
transform -1 0 1208 0 -1 3010
box 0 0 48 200
use FILL  FILL_AOI21X1_37
timestamp 1515882711
transform 1 0 1208 0 -1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_37
timestamp 1515882711
transform 1 0 1224 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_113
timestamp 1515882711
transform -1 0 1336 0 -1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_204
timestamp 1515882711
transform 1 0 1336 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_204
timestamp 1515882711
transform 1 0 1352 0 -1 3010
box 0 0 192 200
use NAND3X1  NAND3X1_175
timestamp 1515882711
transform -1 0 1608 0 -1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_129
timestamp 1515882711
transform 1 0 1608 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_129
timestamp 1515882711
transform 1 0 1624 0 -1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_242
timestamp 1515882711
transform -1 0 1704 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_242
timestamp 1515882711
transform -1 0 1768 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_138
timestamp 1515882711
transform 1 0 1768 0 -1 3010
box 0 0 48 200
use FILL  FILL_INVX1_34
timestamp 1515882711
transform -1 0 1832 0 -1 3010
box 0 0 16 200
use INVX1  INVX1_34
timestamp 1515882711
transform -1 0 1864 0 -1 3010
box 0 0 32 200
use FILL  FILL_NAND2X1_183
timestamp 1515882711
transform -1 0 1880 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_183
timestamp 1515882711
transform -1 0 1928 0 -1 3010
box 0 0 48 200
use FILL  FILL_AND2X2_7
timestamp 1515882711
transform 1 0 1928 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_0
timestamp 1515882711
transform 1 0 1944 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_1_1
timestamp 1515882711
transform 1 0 1960 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_7
timestamp 1515882711
transform 1 0 1976 0 -1 3010
box 0 0 64 200
use NOR2X1  NOR2X1_77
timestamp 1515882711
transform -1 0 2088 0 -1 3010
box 0 0 48 200
use FILL  FILL_AOI21X1_2
timestamp 1515882711
transform -1 0 2104 0 -1 3010
box 0 0 16 200
use AOI21X1  AOI21X1_2
timestamp 1515882711
transform -1 0 2168 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_134
timestamp 1515882711
transform -1 0 2232 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_333
timestamp 1515882711
transform 1 0 2232 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_333
timestamp 1515882711
transform 1 0 2248 0 -1 3010
box 0 0 48 200
use NAND3X1  NAND3X1_136
timestamp 1515882711
transform 1 0 2296 0 -1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_232
timestamp 1515882711
transform -1 0 2376 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_232
timestamp 1515882711
transform -1 0 2440 0 -1 3010
box 0 0 64 200
use NAND3X1  NAND3X1_133
timestamp 1515882711
transform -1 0 2504 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_40
timestamp 1515882711
transform 1 0 2504 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_40
timestamp 1515882711
transform 1 0 2520 0 -1 3010
box 0 0 192 200
use FILL  FILL_INVX1_29
timestamp 1515882711
transform 1 0 2712 0 -1 3010
box 0 0 16 200
use INVX1  INVX1_29
timestamp 1515882711
transform 1 0 2728 0 -1 3010
box 0 0 32 200
use OAI21X1  OAI21X1_251
timestamp 1515882711
transform 1 0 2760 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_19
timestamp 1515882711
transform 1 0 2824 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_19
timestamp 1515882711
transform 1 0 2840 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_40
timestamp 1515882711
transform -1 0 2952 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_2_0
timestamp 1515882711
transform -1 0 2968 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_2_1
timestamp 1515882711
transform -1 0 2984 0 -1 3010
box 0 0 16 200
use OAI21X1  OAI21X1_253
timestamp 1515882711
transform -1 0 3048 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_26
timestamp 1515882711
transform -1 0 3064 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_26
timestamp 1515882711
transform -1 0 3112 0 -1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_47
timestamp 1515882711
transform -1 0 3128 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_47
timestamp 1515882711
transform -1 0 3320 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_47
timestamp 1515882711
transform -1 0 3384 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_75
timestamp 1515882711
transform -1 0 3448 0 -1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_89
timestamp 1515882711
transform -1 0 3464 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_89
timestamp 1515882711
transform -1 0 3528 0 -1 3010
box 0 0 64 200
use FILL  FILL_BUFX4_205
timestamp 1515882711
transform 1 0 3528 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_205
timestamp 1515882711
transform 1 0 3544 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_82
timestamp 1515882711
transform 1 0 3608 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_82
timestamp 1515882711
transform 1 0 3624 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_82
timestamp 1515882711
transform 1 0 3816 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_63
timestamp 1515882711
transform 1 0 3880 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_63
timestamp 1515882711
transform 1 0 3896 0 -1 3010
box 0 0 48 200
use FILL  FILL_BUFX4_47
timestamp 1515882711
transform -1 0 3960 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_47
timestamp 1515882711
transform -1 0 4024 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_3_0
timestamp 1515882711
transform 1 0 4024 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_3_1
timestamp 1515882711
transform 1 0 4040 0 -1 3010
box 0 0 16 200
use FILL  FILL_NAND2X1_278
timestamp 1515882711
transform 1 0 4056 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_278
timestamp 1515882711
transform 1 0 4072 0 -1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_201
timestamp 1515882711
transform -1 0 4136 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_201
timestamp 1515882711
transform -1 0 4328 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_201
timestamp 1515882711
transform 1 0 4328 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_235
timestamp 1515882711
transform 1 0 4392 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_235
timestamp 1515882711
transform 1 0 4408 0 -1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_157
timestamp 1515882711
transform 1 0 4456 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_157
timestamp 1515882711
transform 1 0 4472 0 -1 3010
box 0 0 192 200
use FILL  FILL_NAND2X1_190
timestamp 1515882711
transform 1 0 4664 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_190
timestamp 1515882711
transform 1 0 4680 0 -1 3010
box 0 0 48 200
use FILL  FILL_AND2X2_9
timestamp 1515882711
transform -1 0 4744 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_9
timestamp 1515882711
transform -1 0 4808 0 -1 3010
box 0 0 64 200
use NAND2X1  NAND2X1_445
timestamp 1515882711
transform -1 0 4856 0 -1 3010
box 0 0 48 200
use FILL  FILL_NAND2X1_12
timestamp 1515882711
transform 1 0 4856 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_12
timestamp 1515882711
transform 1 0 4872 0 -1 3010
box 0 0 48 200
use FILL  FILL_NAND2X1_358
timestamp 1515882711
transform 1 0 4920 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_358
timestamp 1515882711
transform 1 0 4936 0 -1 3010
box 0 0 48 200
use FILL  FILL_AND2X2_1
timestamp 1515882711
transform -1 0 5000 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_4_0
timestamp 1515882711
transform -1 0 5016 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_4_1
timestamp 1515882711
transform -1 0 5032 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_1
timestamp 1515882711
transform -1 0 5096 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_31
timestamp 1515882711
transform -1 0 5112 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_31
timestamp 1515882711
transform -1 0 5160 0 -1 3010
box 0 0 48 200
use FILL  FILL_NAND2X1_112
timestamp 1515882711
transform 1 0 5160 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_112
timestamp 1515882711
transform 1 0 5176 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_133
timestamp 1515882711
transform 1 0 5224 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_1
timestamp 1515882711
transform 1 0 5272 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_144
timestamp 1515882711
transform -1 0 5368 0 -1 3010
box 0 0 48 200
use FILL  FILL_AND2X2_3
timestamp 1515882711
transform -1 0 5384 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_3
timestamp 1515882711
transform -1 0 5448 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_42
timestamp 1515882711
transform 1 0 5448 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_42
timestamp 1515882711
transform 1 0 5464 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_62
timestamp 1515882711
transform -1 0 5576 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_100
timestamp 1515882711
transform 1 0 5576 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_100
timestamp 1515882711
transform 1 0 5592 0 -1 3010
box 0 0 192 200
use FILL  FILL_NAND2X1_69
timestamp 1515882711
transform -1 0 5800 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_69
timestamp 1515882711
transform -1 0 5848 0 -1 3010
box 0 0 48 200
use FILL  FILL_AND2X2_4
timestamp 1515882711
transform -1 0 5864 0 -1 3010
box 0 0 16 200
use AND2X2  AND2X2_4
timestamp 1515882711
transform -1 0 5928 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_301
timestamp 1515882711
transform -1 0 5944 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_301
timestamp 1515882711
transform -1 0 5992 0 -1 3010
box 0 0 48 200
use FILL  FILL_BUFX4_108
timestamp 1515882711
transform 1 0 5992 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_108
timestamp 1515882711
transform 1 0 6008 0 -1 3010
box 0 0 64 200
use FILL  FILL_14_5_0
timestamp 1515882711
transform 1 0 6072 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_5_1
timestamp 1515882711
transform 1 0 6088 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_403
timestamp 1515882711
transform 1 0 6104 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_89
timestamp 1515882711
transform 1 0 6152 0 -1 3010
box 0 0 48 200
use NOR2X1  NOR2X1_100
timestamp 1515882711
transform -1 0 6248 0 -1 3010
box 0 0 48 200
use FILL  FILL_NAND2X1_87
timestamp 1515882711
transform -1 0 6264 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_87
timestamp 1515882711
transform -1 0 6312 0 -1 3010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_328
timestamp 1515882711
transform -1 0 6328 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_328
timestamp 1515882711
transform -1 0 6520 0 -1 3010
box 0 0 192 200
use OR2X2  OR2X2_1
timestamp 1515882711
transform 1 0 6520 0 -1 3010
box 0 0 64 200
use FILL  FILL_NAND2X1_109
timestamp 1515882711
transform -1 0 6600 0 -1 3010
box 0 0 16 200
use NAND2X1  NAND2X1_109
timestamp 1515882711
transform -1 0 6648 0 -1 3010
box 0 0 48 200
use OAI21X1  OAI21X1_126
timestamp 1515882711
transform -1 0 6712 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_126
timestamp 1515882711
transform -1 0 6728 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_126
timestamp 1515882711
transform -1 0 6920 0 -1 3010
box 0 0 192 200
use FILL  FILL_BUFX4_272
timestamp 1515882711
transform 1 0 6920 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_272
timestamp 1515882711
transform 1 0 6936 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_499
timestamp 1515882711
transform 1 0 7000 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_279
timestamp 1515882711
transform 1 0 7064 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_6_0
timestamp 1515882711
transform 1 0 7080 0 -1 3010
box 0 0 16 200
use FILL  FILL_14_6_1
timestamp 1515882711
transform 1 0 7096 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_279
timestamp 1515882711
transform 1 0 7112 0 -1 3010
box 0 0 192 200
use OAI21X1  OAI21X1_498
timestamp 1515882711
transform -1 0 7368 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_293
timestamp 1515882711
transform -1 0 7384 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_293
timestamp 1515882711
transform -1 0 7576 0 -1 3010
box 0 0 192 200
use FILL  FILL_BUFX4_153
timestamp 1515882711
transform -1 0 7592 0 -1 3010
box 0 0 16 200
use BUFX4  BUFX4_153
timestamp 1515882711
transform -1 0 7656 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_494
timestamp 1515882711
transform 1 0 7656 0 -1 3010
box 0 0 64 200
use OAI21X1  OAI21X1_495
timestamp 1515882711
transform -1 0 7784 0 -1 3010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_257
timestamp 1515882711
transform -1 0 7800 0 -1 3010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_257
timestamp 1515882711
transform -1 0 7992 0 -1 3010
box 0 0 192 200
use FILL  FILL_INVX1_49
timestamp 1515882711
transform 1 0 7992 0 -1 3010
box 0 0 16 200
use INVX1  INVX1_49
timestamp 1515882711
transform 1 0 8008 0 -1 3010
box 0 0 32 200
use FILL  FILL_15_1
timestamp 1515882711
transform -1 0 8056 0 -1 3010
box 0 0 16 200
use FILL  FILL_DFFPOSX1_171
timestamp 1515882711
transform -1 0 24 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_171
timestamp 1515882711
transform -1 0 216 0 1 2610
box 0 0 192 200
use NOR2X1  NOR2X1_97
timestamp 1515882711
transform 1 0 216 0 1 2610
box 0 0 48 200
use FILL  FILL_BUFX4_134
timestamp 1515882711
transform -1 0 280 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_134
timestamp 1515882711
transform -1 0 344 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_175
timestamp 1515882711
transform -1 0 360 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_175
timestamp 1515882711
transform -1 0 552 0 1 2610
box 0 0 192 200
use FILL  FILL_DFFPOSX1_225
timestamp 1515882711
transform 1 0 552 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_225
timestamp 1515882711
transform 1 0 568 0 1 2610
box 0 0 192 200
use FILL  FILL_BUFX4_92
timestamp 1515882711
transform -1 0 776 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_92
timestamp 1515882711
transform -1 0 840 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_226
timestamp 1515882711
transform 1 0 840 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_226
timestamp 1515882711
transform 1 0 856 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_11
timestamp 1515882711
transform 1 0 920 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_0
timestamp 1515882711
transform 1 0 936 0 1 2610
box 0 0 16 200
use FILL  FILL_13_0_1
timestamp 1515882711
transform 1 0 952 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_11
timestamp 1515882711
transform 1 0 968 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_172
timestamp 1515882711
transform 1 0 1032 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_172
timestamp 1515882711
transform 1 0 1048 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_19
timestamp 1515882711
transform 1 0 1112 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_19
timestamp 1515882711
transform 1 0 1128 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_250
timestamp 1515882711
transform -1 0 1208 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_250
timestamp 1515882711
transform -1 0 1400 0 1 2610
box 0 0 192 200
use NOR2X1  NOR2X1_24
timestamp 1515882711
transform 1 0 1400 0 1 2610
box 0 0 48 200
use FILL  FILL_AOI21X1_23
timestamp 1515882711
transform -1 0 1464 0 1 2610
box 0 0 16 200
use AOI21X1  AOI21X1_23
timestamp 1515882711
transform -1 0 1528 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_214
timestamp 1515882711
transform -1 0 1544 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_214
timestamp 1515882711
transform -1 0 1736 0 1 2610
box 0 0 192 200
use FILL  FILL_BUFX4_137
timestamp 1515882711
transform -1 0 1752 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_137
timestamp 1515882711
transform -1 0 1816 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_62
timestamp 1515882711
transform 1 0 1816 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_62
timestamp 1515882711
transform 1 0 1832 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_142
timestamp 1515882711
transform -1 0 1912 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_142
timestamp 1515882711
transform -1 0 1976 0 1 2610
box 0 0 64 200
use FILL  FILL_13_1_0
timestamp 1515882711
transform 1 0 1976 0 1 2610
box 0 0 16 200
use FILL  FILL_13_1_1
timestamp 1515882711
transform 1 0 1992 0 1 2610
box 0 0 16 200
use FILL  FILL_BUFX4_250
timestamp 1515882711
transform 1 0 2008 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_250
timestamp 1515882711
transform 1 0 2024 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_212
timestamp 1515882711
transform 1 0 2088 0 1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_102
timestamp 1515882711
transform 1 0 2152 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_327
timestamp 1515882711
transform -1 0 2232 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_327
timestamp 1515882711
transform -1 0 2280 0 1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_100
timestamp 1515882711
transform 1 0 2280 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_37
timestamp 1515882711
transform -1 0 2360 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_37
timestamp 1515882711
transform -1 0 2552 0 1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_16
timestamp 1515882711
transform 1 0 2552 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_16
timestamp 1515882711
transform 1 0 2568 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_37
timestamp 1515882711
transform -1 0 2680 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_335
timestamp 1515882711
transform -1 0 2696 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_335
timestamp 1515882711
transform -1 0 2888 0 1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_361
timestamp 1515882711
transform 1 0 2888 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_361
timestamp 1515882711
transform 1 0 2904 0 1 2610
box 0 0 48 200
use FILL  FILL_13_2_0
timestamp 1515882711
transform -1 0 2968 0 1 2610
box 0 0 16 200
use FILL  FILL_13_2_1
timestamp 1515882711
transform -1 0 2984 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_428
timestamp 1515882711
transform -1 0 3048 0 1 2610
box 0 0 64 200
use FILL  FILL_INVX1_30
timestamp 1515882711
transform -1 0 3064 0 1 2610
box 0 0 16 200
use INVX1  INVX1_30
timestamp 1515882711
transform -1 0 3096 0 1 2610
box 0 0 32 200
use FILL  FILL_NAND2X1_192
timestamp 1515882711
transform 1 0 3096 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_192
timestamp 1515882711
transform 1 0 3112 0 1 2610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_75
timestamp 1515882711
transform -1 0 3176 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_75
timestamp 1515882711
transform -1 0 3368 0 1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_56
timestamp 1515882711
transform 1 0 3368 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_56
timestamp 1515882711
transform 1 0 3384 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_274
timestamp 1515882711
transform -1 0 3496 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_249
timestamp 1515882711
transform 1 0 3496 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_249
timestamp 1515882711
transform 1 0 3512 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_222
timestamp 1515882711
transform -1 0 3624 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_2
timestamp 1515882711
transform 1 0 3624 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_2
timestamp 1515882711
transform 1 0 3640 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_492
timestamp 1515882711
transform -1 0 3752 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_25
timestamp 1515882711
transform -1 0 3768 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_25
timestamp 1515882711
transform -1 0 3960 0 1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_208
timestamp 1515882711
transform 1 0 3960 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_208
timestamp 1515882711
transform 1 0 3976 0 1 2610
box 0 0 48 200
use FILL  FILL_13_3_0
timestamp 1515882711
transform 1 0 4024 0 1 2610
box 0 0 16 200
use FILL  FILL_13_3_1
timestamp 1515882711
transform 1 0 4040 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_223
timestamp 1515882711
transform 1 0 4056 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_19
timestamp 1515882711
transform -1 0 4136 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_19
timestamp 1515882711
transform -1 0 4328 0 1 2610
box 0 0 192 200
use FILL  FILL_BUFX4_265
timestamp 1515882711
transform -1 0 4344 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_265
timestamp 1515882711
transform -1 0 4408 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_333
timestamp 1515882711
transform -1 0 4424 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_333
timestamp 1515882711
transform -1 0 4616 0 1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_359
timestamp 1515882711
transform 1 0 4616 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_359
timestamp 1515882711
transform 1 0 4632 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_426
timestamp 1515882711
transform -1 0 4744 0 1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_74
timestamp 1515882711
transform -1 0 4760 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_74
timestamp 1515882711
transform -1 0 4824 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_135
timestamp 1515882711
transform 1 0 4824 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_135
timestamp 1515882711
transform 1 0 4840 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_101
timestamp 1515882711
transform -1 0 4952 0 1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_101
timestamp 1515882711
transform -1 0 4968 0 1 2610
box 0 0 16 200
use FILL  FILL_13_4_0
timestamp 1515882711
transform -1 0 4984 0 1 2610
box 0 0 16 200
use FILL  FILL_13_4_1
timestamp 1515882711
transform -1 0 5000 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_101
timestamp 1515882711
transform -1 0 5192 0 1 2610
box 0 0 192 200
use FILL  FILL_DFFPOSX1_87
timestamp 1515882711
transform -1 0 5208 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_87
timestamp 1515882711
transform -1 0 5400 0 1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_70
timestamp 1515882711
transform 1 0 5400 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_70
timestamp 1515882711
transform 1 0 5416 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_87
timestamp 1515882711
transform -1 0 5528 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_100
timestamp 1515882711
transform 1 0 5528 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_83
timestamp 1515882711
transform -1 0 5608 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_83
timestamp 1515882711
transform -1 0 5656 0 1 2610
box 0 0 48 200
use NOR3X1  NOR3X1_19
timestamp 1515882711
transform -1 0 5784 0 1 2610
box 0 0 128 200
use NOR2X1  NOR2X1_21
timestamp 1515882711
transform -1 0 5832 0 1 2610
box 0 0 48 200
use OAI22X1  OAI22X1_5
timestamp 1515882711
transform 1 0 5832 0 1 2610
box 0 0 80 200
use NOR2X1  NOR2X1_20
timestamp 1515882711
transform 1 0 5912 0 1 2610
box 0 0 48 200
use FILL  FILL_MUX2X1_31
timestamp 1515882711
transform -1 0 5976 0 1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_31
timestamp 1515882711
transform -1 0 6072 0 1 2610
box 0 0 96 200
use FILL  FILL_13_5_0
timestamp 1515882711
transform 1 0 6072 0 1 2610
box 0 0 16 200
use FILL  FILL_13_5_1
timestamp 1515882711
transform 1 0 6088 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_410
timestamp 1515882711
transform 1 0 6104 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_318
timestamp 1515882711
transform 1 0 6168 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_349
timestamp 1515882711
transform -1 0 6248 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_349
timestamp 1515882711
transform -1 0 6296 0 1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_417
timestamp 1515882711
transform 1 0 6296 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_472
timestamp 1515882711
transform -1 0 6408 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_137
timestamp 1515882711
transform 1 0 6408 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_121
timestamp 1515882711
transform -1 0 6488 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_121
timestamp 1515882711
transform -1 0 6536 0 1 2610
box 0 0 48 200
use FILL  FILL_MUX2X1_33
timestamp 1515882711
transform 1 0 6536 0 1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_33
timestamp 1515882711
transform 1 0 6552 0 1 2610
box 0 0 96 200
use FILL  FILL_DFFPOSX1_311
timestamp 1515882711
transform -1 0 6664 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_311
timestamp 1515882711
transform -1 0 6856 0 1 2610
box 0 0 192 200
use NAND2X1  NAND2X1_437
timestamp 1515882711
transform 1 0 6856 0 1 2610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_143
timestamp 1515882711
transform 1 0 6904 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_143
timestamp 1515882711
transform 1 0 6920 0 1 2610
box 0 0 192 200
use FILL  FILL_13_6_0
timestamp 1515882711
transform 1 0 7112 0 1 2610
box 0 0 16 200
use FILL  FILL_13_6_1
timestamp 1515882711
transform 1 0 7128 0 1 2610
box 0 0 16 200
use OAI21X1  OAI21X1_143
timestamp 1515882711
transform 1 0 7144 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_129
timestamp 1515882711
transform -1 0 7224 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_129
timestamp 1515882711
transform -1 0 7272 0 1 2610
box 0 0 48 200
use FILL  FILL_BUFX4_37
timestamp 1515882711
transform 1 0 7272 0 1 2610
box 0 0 16 200
use BUFX4  BUFX4_37
timestamp 1515882711
transform 1 0 7288 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_282
timestamp 1515882711
transform 1 0 7352 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_282
timestamp 1515882711
transform 1 0 7368 0 1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_8
timestamp 1515882711
transform -1 0 7480 0 1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1515882711
transform -1 0 7544 0 1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_187
timestamp 1515882711
transform 1 0 7544 0 1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_187
timestamp 1515882711
transform 1 0 7560 0 1 2610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_141
timestamp 1515882711
transform -1 0 7624 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_141
timestamp 1515882711
transform -1 0 7816 0 1 2610
box 0 0 192 200
use FILL  FILL_DFFPOSX1_285
timestamp 1515882711
transform -1 0 7832 0 1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_285
timestamp 1515882711
transform -1 0 8024 0 1 2610
box 0 0 192 200
use FILL  FILL_14_1
timestamp 1515882711
transform 1 0 8024 0 1 2610
box 0 0 16 200
use FILL  FILL_14_2
timestamp 1515882711
transform 1 0 8040 0 1 2610
box 0 0 16 200
use FILL  FILL_BUFX4_227
timestamp 1515882711
transform -1 0 24 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_227
timestamp 1515882711
transform -1 0 88 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_147
timestamp 1515882711
transform -1 0 104 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_147
timestamp 1515882711
transform -1 0 168 0 -1 2610
box 0 0 64 200
use FILL  FILL_AOI21X1_21
timestamp 1515882711
transform 1 0 168 0 -1 2610
box 0 0 16 200
use AOI21X1  AOI21X1_21
timestamp 1515882711
transform 1 0 184 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_102
timestamp 1515882711
transform -1 0 296 0 -1 2610
box 0 0 48 200
use FILL  FILL_AOI21X1_26
timestamp 1515882711
transform -1 0 312 0 -1 2610
box 0 0 16 200
use AOI21X1  AOI21X1_26
timestamp 1515882711
transform -1 0 376 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_313
timestamp 1515882711
transform -1 0 392 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_313
timestamp 1515882711
transform -1 0 456 0 -1 2610
box 0 0 64 200
use FILL  FILL_AOI21X1_57
timestamp 1515882711
transform 1 0 456 0 -1 2610
box 0 0 16 200
use AOI21X1  AOI21X1_57
timestamp 1515882711
transform 1 0 472 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_132
timestamp 1515882711
transform -1 0 584 0 -1 2610
box 0 0 48 200
use FILL  FILL_BUFX4_210
timestamp 1515882711
transform 1 0 584 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_210
timestamp 1515882711
transform 1 0 600 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_169
timestamp 1515882711
transform -1 0 680 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_169
timestamp 1515882711
transform -1 0 744 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_178
timestamp 1515882711
transform 1 0 744 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_178
timestamp 1515882711
transform 1 0 760 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_97
timestamp 1515882711
transform -1 0 888 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_157
timestamp 1515882711
transform -1 0 952 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_0_0
timestamp 1515882711
transform 1 0 952 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_0_1
timestamp 1515882711
transform 1 0 968 0 -1 2610
box 0 0 16 200
use NAND3X1  NAND3X1_190
timestamp 1515882711
transform 1 0 984 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_179
timestamp 1515882711
transform 1 0 1048 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_135
timestamp 1515882711
transform -1 0 1128 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_135
timestamp 1515882711
transform -1 0 1192 0 -1 2610
box 0 0 64 200
use NOR3X1  NOR3X1_44
timestamp 1515882711
transform -1 0 1320 0 -1 2610
box 0 0 128 200
use OAI21X1  OAI21X1_215
timestamp 1515882711
transform 1 0 1320 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_135
timestamp 1515882711
transform -1 0 1448 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_216
timestamp 1515882711
transform 1 0 1448 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_146
timestamp 1515882711
transform -1 0 1576 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_94
timestamp 1515882711
transform -1 0 1640 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_123
timestamp 1515882711
transform 1 0 1640 0 -1 2610
box 0 0 48 200
use FILL  FILL_AOI21X1_47
timestamp 1515882711
transform -1 0 1704 0 -1 2610
box 0 0 16 200
use AOI21X1  AOI21X1_47
timestamp 1515882711
transform -1 0 1768 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_201
timestamp 1515882711
transform -1 0 1784 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_201
timestamp 1515882711
transform -1 0 1848 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_235
timestamp 1515882711
transform -1 0 1912 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_153
timestamp 1515882711
transform 1 0 1912 0 -1 2610
box 0 0 48 200
use FILL  FILL_12_1_0
timestamp 1515882711
transform -1 0 1976 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_1_1
timestamp 1515882711
transform -1 0 1992 0 -1 2610
box 0 0 16 200
use FILL  FILL_NAND2X1_210
timestamp 1515882711
transform -1 0 2008 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_210
timestamp 1515882711
transform -1 0 2056 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_224
timestamp 1515882711
transform 1 0 2056 0 -1 2610
box 0 0 64 200
use NOR2X1  NOR2X1_45
timestamp 1515882711
transform -1 0 2168 0 -1 2610
box 0 0 48 200
use NAND3X1  NAND3X1_201
timestamp 1515882711
transform -1 0 2232 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_221
timestamp 1515882711
transform -1 0 2296 0 -1 2610
box 0 0 64 200
use NAND3X1  NAND3X1_99
timestamp 1515882711
transform -1 0 2360 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_367
timestamp 1515882711
transform -1 0 2424 0 -1 2610
box 0 0 64 200
use FILL  FILL_INVX1_13
timestamp 1515882711
transform 1 0 2424 0 -1 2610
box 0 0 16 200
use INVX1  INVX1_13
timestamp 1515882711
transform 1 0 2440 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_220
timestamp 1515882711
transform 1 0 2472 0 -1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_207
timestamp 1515882711
transform 1 0 2536 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_207
timestamp 1515882711
transform 1 0 2552 0 -1 2610
box 0 0 48 200
use FILL  FILL_BUFX4_127
timestamp 1515882711
transform -1 0 2616 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_127
timestamp 1515882711
transform -1 0 2680 0 -1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_14
timestamp 1515882711
transform -1 0 2696 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_14
timestamp 1515882711
transform -1 0 2744 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_34
timestamp 1515882711
transform -1 0 2808 0 -1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_34
timestamp 1515882711
transform 1 0 2808 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_34
timestamp 1515882711
transform 1 0 2824 0 -1 2610
box 0 0 192 200
use FILL  FILL_12_2_0
timestamp 1515882711
transform 1 0 3016 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_2_1
timestamp 1515882711
transform 1 0 3032 0 -1 2610
box 0 0 16 200
use FILL  FILL_INVX1_2
timestamp 1515882711
transform 1 0 3048 0 -1 2610
box 0 0 16 200
use INVX1  INVX1_2
timestamp 1515882711
transform 1 0 3064 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_200
timestamp 1515882711
transform 1 0 3096 0 -1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_17
timestamp 1515882711
transform 1 0 3160 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_17
timestamp 1515882711
transform 1 0 3176 0 -1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_194
timestamp 1515882711
transform -1 0 3384 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_194
timestamp 1515882711
transform -1 0 3432 0 -1 2610
box 0 0 48 200
use FILL  FILL_NAND2X1_223
timestamp 1515882711
transform 1 0 3432 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_223
timestamp 1515882711
transform 1 0 3448 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_1
timestamp 1515882711
transform -1 0 3560 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_206
timestamp 1515882711
transform -1 0 3576 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_206
timestamp 1515882711
transform -1 0 3640 0 -1 2610
box 0 0 64 200
use FILL  FILL_INVX1_14
timestamp 1515882711
transform -1 0 3656 0 -1 2610
box 0 0 16 200
use INVX1  INVX1_14
timestamp 1515882711
transform -1 0 3688 0 -1 2610
box 0 0 32 200
use FILL  FILL_BUFX4_159
timestamp 1515882711
transform -1 0 3704 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_159
timestamp 1515882711
transform -1 0 3768 0 -1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_53
timestamp 1515882711
transform 1 0 3768 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_53
timestamp 1515882711
transform 1 0 3784 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_72
timestamp 1515882711
transform -1 0 3896 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_225
timestamp 1515882711
transform -1 0 3960 0 -1 2610
box 0 0 64 200
use FILL  FILL_INVX1_15
timestamp 1515882711
transform -1 0 3976 0 -1 2610
box 0 0 16 200
use INVX1  INVX1_15
timestamp 1515882711
transform -1 0 4008 0 -1 2610
box 0 0 32 200
use FILL  FILL_12_3_0
timestamp 1515882711
transform 1 0 4008 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_3_1
timestamp 1515882711
transform 1 0 4024 0 -1 2610
box 0 0 16 200
use FILL  FILL_NAND2X1_209
timestamp 1515882711
transform 1 0 4040 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_209
timestamp 1515882711
transform 1 0 4056 0 -1 2610
box 0 0 48 200
use NAND2X1  NAND2X1_398
timestamp 1515882711
transform -1 0 4152 0 -1 2610
box 0 0 48 200
use FILL  FILL_NAND2X1_34
timestamp 1515882711
transform 1 0 4152 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_34
timestamp 1515882711
transform 1 0 4168 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_54
timestamp 1515882711
transform -1 0 4280 0 -1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_54
timestamp 1515882711
transform -1 0 4296 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_54
timestamp 1515882711
transform -1 0 4488 0 -1 2610
box 0 0 192 200
use FILL  FILL_DFFPOSX1_346
timestamp 1515882711
transform -1 0 4504 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_346
timestamp 1515882711
transform -1 0 4696 0 -1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_372
timestamp 1515882711
transform 1 0 4696 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_372
timestamp 1515882711
transform 1 0 4712 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_439
timestamp 1515882711
transform -1 0 4824 0 -1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_246
timestamp 1515882711
transform 1 0 4824 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_246
timestamp 1515882711
transform 1 0 4840 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_212
timestamp 1515882711
transform -1 0 4952 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_128
timestamp 1515882711
transform 1 0 4952 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_128
timestamp 1515882711
transform 1 0 4968 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_4_0
timestamp 1515882711
transform 1 0 5032 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_4_1
timestamp 1515882711
transform 1 0 5048 0 -1 2610
box 0 0 16 200
use FILL  FILL_BUFX4_186
timestamp 1515882711
transform 1 0 5064 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_186
timestamp 1515882711
transform 1 0 5080 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_125
timestamp 1515882711
transform 1 0 5144 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_125
timestamp 1515882711
transform 1 0 5160 0 -1 2610
box 0 0 64 200
use FILL  FILL_MUX2X1_12
timestamp 1515882711
transform 1 0 5224 0 -1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_12
timestamp 1515882711
transform 1 0 5240 0 -1 2610
box 0 0 96 200
use FILL  FILL_BUFX4_188
timestamp 1515882711
transform 1 0 5336 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_188
timestamp 1515882711
transform 1 0 5352 0 -1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_35
timestamp 1515882711
transform 1 0 5416 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_35
timestamp 1515882711
transform 1 0 5432 0 -1 2610
box 0 0 192 200
use OAI21X1  OAI21X1_390
timestamp 1515882711
transform 1 0 5624 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_399
timestamp 1515882711
transform -1 0 5736 0 -1 2610
box 0 0 48 200
use FILL  FILL_MUX2X1_32
timestamp 1515882711
transform 1 0 5736 0 -1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_32
timestamp 1515882711
transform 1 0 5752 0 -1 2610
box 0 0 96 200
use NOR2X1  NOR2X1_66
timestamp 1515882711
transform -1 0 5896 0 -1 2610
box 0 0 48 200
use FILL  FILL_BUFX4_119
timestamp 1515882711
transform -1 0 5912 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_119
timestamp 1515882711
transform -1 0 5976 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_123
timestamp 1515882711
transform -1 0 5992 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_123
timestamp 1515882711
transform -1 0 6056 0 -1 2610
box 0 0 64 200
use FILL  FILL_12_5_0
timestamp 1515882711
transform -1 0 6072 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_5_1
timestamp 1515882711
transform -1 0 6088 0 -1 2610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_119
timestamp 1515882711
transform -1 0 6104 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_119
timestamp 1515882711
transform -1 0 6296 0 -1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_102
timestamp 1515882711
transform 1 0 6296 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_102
timestamp 1515882711
transform 1 0 6312 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_119
timestamp 1515882711
transform -1 0 6424 0 -1 2610
box 0 0 64 200
use FILL  FILL_NAND2X1_283
timestamp 1515882711
transform 1 0 6424 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_283
timestamp 1515882711
transform 1 0 6440 0 -1 2610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_137
timestamp 1515882711
transform 1 0 6488 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_137
timestamp 1515882711
transform 1 0 6504 0 -1 2610
box 0 0 192 200
use FILL  FILL_BUFX4_120
timestamp 1515882711
transform 1 0 6696 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_120
timestamp 1515882711
transform 1 0 6712 0 -1 2610
box 0 0 64 200
use FILL  FILL_MUX2X1_48
timestamp 1515882711
transform 1 0 6776 0 -1 2610
box 0 0 16 200
use MUX2X1  MUX2X1_48
timestamp 1515882711
transform 1 0 6792 0 -1 2610
box 0 0 96 200
use OAI21X1  OAI21X1_489
timestamp 1515882711
transform -1 0 6952 0 -1 2610
box 0 0 64 200
use NAND2X1  NAND2X1_426
timestamp 1515882711
transform 1 0 6952 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_478
timestamp 1515882711
transform -1 0 7064 0 -1 2610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_300
timestamp 1515882711
transform -1 0 7080 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_6_0
timestamp 1515882711
transform -1 0 7096 0 -1 2610
box 0 0 16 200
use FILL  FILL_12_6_1
timestamp 1515882711
transform -1 0 7112 0 -1 2610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_300
timestamp 1515882711
transform -1 0 7304 0 -1 2610
box 0 0 192 200
use FILL  FILL_NAND2X1_204
timestamp 1515882711
transform -1 0 7320 0 -1 2610
box 0 0 16 200
use NAND2X1  NAND2X1_204
timestamp 1515882711
transform -1 0 7368 0 -1 2610
box 0 0 48 200
use OAI21X1  OAI21X1_217
timestamp 1515882711
transform -1 0 7432 0 -1 2610
box 0 0 64 200
use FILL  FILL_INVX1_10
timestamp 1515882711
transform 1 0 7432 0 -1 2610
box 0 0 16 200
use INVX1  INVX1_10
timestamp 1515882711
transform 1 0 7448 0 -1 2610
box 0 0 32 200
use OAI21X1  OAI21X1_317
timestamp 1515882711
transform -1 0 7544 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_310
timestamp 1515882711
transform -1 0 7560 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_310
timestamp 1515882711
transform -1 0 7624 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_141
timestamp 1515882711
transform 1 0 7624 0 -1 2610
box 0 0 64 200
use OAI21X1  OAI21X1_197
timestamp 1515882711
transform -1 0 7752 0 -1 2610
box 0 0 64 200
use FILL  FILL_INVX1_78
timestamp 1515882711
transform -1 0 7768 0 -1 2610
box 0 0 16 200
use INVX1  INVX1_78
timestamp 1515882711
transform -1 0 7800 0 -1 2610
box 0 0 32 200
use FILL  FILL_BUFX4_33
timestamp 1515882711
transform 1 0 7800 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_33
timestamp 1515882711
transform 1 0 7816 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_260
timestamp 1515882711
transform -1 0 7896 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_260
timestamp 1515882711
transform -1 0 7960 0 -1 2610
box 0 0 64 200
use FILL  FILL_BUFX4_258
timestamp 1515882711
transform -1 0 7976 0 -1 2610
box 0 0 16 200
use BUFX4  BUFX4_258
timestamp 1515882711
transform -1 0 8040 0 -1 2610
box 0 0 64 200
use FILL  FILL_13_1
timestamp 1515882711
transform -1 0 8056 0 -1 2610
box 0 0 16 200
use BUFX2  BUFX2_35
timestamp 1515882711
transform -1 0 56 0 1 2210
box 0 0 48 200
use FILL  FILL_BUFX2_23
timestamp 1515882711
transform -1 0 72 0 1 2210
box 0 0 16 200
use BUFX2  BUFX2_23
timestamp 1515882711
transform -1 0 120 0 1 2210
box 0 0 48 200
use FILL  FILL_AOI21X1_8
timestamp 1515882711
transform 1 0 120 0 1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_8
timestamp 1515882711
transform 1 0 136 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_84
timestamp 1515882711
transform -1 0 248 0 1 2210
box 0 0 48 200
use FILL  FILL_BUFX4_225
timestamp 1515882711
transform -1 0 264 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_225
timestamp 1515882711
transform -1 0 328 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_145
timestamp 1515882711
transform -1 0 344 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_145
timestamp 1515882711
transform -1 0 408 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_197
timestamp 1515882711
transform 1 0 408 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_280
timestamp 1515882711
transform -1 0 488 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_280
timestamp 1515882711
transform -1 0 552 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_149
timestamp 1515882711
transform 1 0 552 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_149
timestamp 1515882711
transform 1 0 568 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_222
timestamp 1515882711
transform -1 0 648 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_222
timestamp 1515882711
transform -1 0 712 0 1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_170
timestamp 1515882711
transform -1 0 728 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_170
timestamp 1515882711
transform -1 0 920 0 1 2210
box 0 0 192 200
use FILL  FILL_11_0_0
timestamp 1515882711
transform -1 0 936 0 1 2210
box 0 0 16 200
use FILL  FILL_11_0_1
timestamp 1515882711
transform -1 0 952 0 1 2210
box 0 0 16 200
use NAND3X1  NAND3X1_96
timestamp 1515882711
transform -1 0 1016 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_168
timestamp 1515882711
transform 1 0 1016 0 1 2210
box 0 0 64 200
use FILL  FILL_AOI21X1_40
timestamp 1515882711
transform 1 0 1080 0 1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_40
timestamp 1515882711
transform 1 0 1096 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_116
timestamp 1515882711
transform 1 0 1160 0 1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_98
timestamp 1515882711
transform -1 0 1272 0 1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_95
timestamp 1515882711
transform 1 0 1272 0 1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_87
timestamp 1515882711
transform 1 0 1336 0 1 2210
box 0 0 48 200
use FILL  FILL_AOI21X1_11
timestamp 1515882711
transform -1 0 1400 0 1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_11
timestamp 1515882711
transform -1 0 1464 0 1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_196
timestamp 1515882711
transform 1 0 1464 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_196
timestamp 1515882711
transform 1 0 1480 0 1 2210
box 0 0 192 200
use NAND3X1  NAND3X1_93
timestamp 1515882711
transform 1 0 1672 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_364
timestamp 1515882711
transform -1 0 1800 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_365
timestamp 1515882711
transform -1 0 1864 0 1 2210
box 0 0 64 200
use NOR3X1  NOR3X1_29
timestamp 1515882711
transform 1 0 1864 0 1 2210
box 0 0 128 200
use FILL  FILL_11_1_0
timestamp 1515882711
transform -1 0 2008 0 1 2210
box 0 0 16 200
use FILL  FILL_11_1_1
timestamp 1515882711
transform -1 0 2024 0 1 2210
box 0 0 16 200
use NAND3X1  NAND3X1_103
timestamp 1515882711
transform -1 0 2088 0 1 2210
box 0 0 64 200
use FILL  FILL_INVX8_5
timestamp 1515882711
transform -1 0 2104 0 1 2210
box 0 0 16 200
use INVX8  INVX8_5
timestamp 1515882711
transform -1 0 2184 0 1 2210
box 0 0 80 200
use FILL  FILL_BUFX4_185
timestamp 1515882711
transform -1 0 2200 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_185
timestamp 1515882711
transform -1 0 2264 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_30
timestamp 1515882711
transform 1 0 2264 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_8
timestamp 1515882711
transform -1 0 2344 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_8
timestamp 1515882711
transform -1 0 2392 0 1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_278
timestamp 1515882711
transform 1 0 2392 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_278
timestamp 1515882711
transform 1 0 2408 0 1 2210
box 0 0 192 200
use FILL  FILL_BUFX4_44
timestamp 1515882711
transform -1 0 2616 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_44
timestamp 1515882711
transform -1 0 2680 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_126
timestamp 1515882711
transform -1 0 2696 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_126
timestamp 1515882711
transform -1 0 2760 0 1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_265
timestamp 1515882711
transform 1 0 2760 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_265
timestamp 1515882711
transform 1 0 2776 0 1 2210
box 0 0 192 200
use FILL  FILL_11_2_0
timestamp 1515882711
transform -1 0 2984 0 1 2210
box 0 0 16 200
use FILL  FILL_11_2_1
timestamp 1515882711
transform -1 0 3000 0 1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_17
timestamp 1515882711
transform -1 0 3064 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_5
timestamp 1515882711
transform 1 0 3064 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_5
timestamp 1515882711
transform 1 0 3080 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_276
timestamp 1515882711
transform -1 0 3160 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_276
timestamp 1515882711
transform -1 0 3224 0 1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_79
timestamp 1515882711
transform 1 0 3224 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_79
timestamp 1515882711
transform 1 0 3240 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_79
timestamp 1515882711
transform -1 0 3496 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_204
timestamp 1515882711
transform -1 0 3560 0 1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_70
timestamp 1515882711
transform -1 0 3576 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_70
timestamp 1515882711
transform -1 0 3768 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_70
timestamp 1515882711
transform 1 0 3768 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_51
timestamp 1515882711
transform 1 0 3832 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_51
timestamp 1515882711
transform 1 0 3848 0 1 2210
box 0 0 48 200
use FILL  FILL_INVX1_42
timestamp 1515882711
transform -1 0 3912 0 1 2210
box 0 0 16 200
use INVX1  INVX1_42
timestamp 1515882711
transform -1 0 3944 0 1 2210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_72
timestamp 1515882711
transform -1 0 3960 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_0
timestamp 1515882711
transform -1 0 3976 0 1 2210
box 0 0 16 200
use FILL  FILL_11_3_1
timestamp 1515882711
transform -1 0 3992 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_72
timestamp 1515882711
transform -1 0 4184 0 1 2210
box 0 0 192 200
use NAND3X1  NAND3X1_37
timestamp 1515882711
transform -1 0 4248 0 1 2210
box 0 0 64 200
use FILL  FILL_INVX1_4
timestamp 1515882711
transform -1 0 4264 0 1 2210
box 0 0 16 200
use INVX1  INVX1_4
timestamp 1515882711
transform -1 0 4296 0 1 2210
box 0 0 32 200
use OAI21X1  OAI21X1_320
timestamp 1515882711
transform -1 0 4360 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_285
timestamp 1515882711
transform 1 0 4360 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_285
timestamp 1515882711
transform 1 0 4376 0 1 2210
box 0 0 48 200
use FILL  FILL_INVX1_68
timestamp 1515882711
transform -1 0 4440 0 1 2210
box 0 0 16 200
use INVX1  INVX1_68
timestamp 1515882711
transform -1 0 4472 0 1 2210
box 0 0 32 200
use FILL  FILL_NAND2X1_27
timestamp 1515882711
transform -1 0 4488 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_27
timestamp 1515882711
transform -1 0 4536 0 1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_48
timestamp 1515882711
transform -1 0 4552 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_48
timestamp 1515882711
transform -1 0 4744 0 1 2210
box 0 0 192 200
use FILL  FILL_BUFX4_311
timestamp 1515882711
transform -1 0 4760 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_311
timestamp 1515882711
transform -1 0 4824 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_286
timestamp 1515882711
transform -1 0 4840 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_286
timestamp 1515882711
transform -1 0 4888 0 1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_212
timestamp 1515882711
transform -1 0 4904 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_212
timestamp 1515882711
transform -1 0 5096 0 1 2210
box 0 0 192 200
use FILL  FILL_11_4_0
timestamp 1515882711
transform 1 0 5096 0 1 2210
box 0 0 16 200
use FILL  FILL_11_4_1
timestamp 1515882711
transform 1 0 5112 0 1 2210
box 0 0 16 200
use FILL  FILL_BUFX4_274
timestamp 1515882711
transform 1 0 5128 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_274
timestamp 1515882711
transform 1 0 5144 0 1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_1
timestamp 1515882711
transform -1 0 5224 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1515882711
transform -1 0 5416 0 1 2210
box 0 0 192 200
use FILL  FILL_NAND2X1_312
timestamp 1515882711
transform 1 0 5416 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_312
timestamp 1515882711
transform 1 0 5432 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_257
timestamp 1515882711
transform -1 0 5544 0 1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_187
timestamp 1515882711
transform 1 0 5544 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_187
timestamp 1515882711
transform 1 0 5560 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_279
timestamp 1515882711
transform 1 0 5624 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_335
timestamp 1515882711
transform -1 0 5704 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_335
timestamp 1515882711
transform -1 0 5752 0 1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_223
timestamp 1515882711
transform 1 0 5752 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_223
timestamp 1515882711
transform 1 0 5768 0 1 2210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_107
timestamp 1515882711
transform 1 0 5960 0 1 2210
box 0 0 16 200
use FILL  FILL_11_5_0
timestamp 1515882711
transform 1 0 5976 0 1 2210
box 0 0 16 200
use FILL  FILL_11_5_1
timestamp 1515882711
transform 1 0 5992 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_107
timestamp 1515882711
transform 1 0 6008 0 1 2210
box 0 0 192 200
use OAI22X1  OAI22X1_10
timestamp 1515882711
transform -1 0 6280 0 1 2210
box 0 0 80 200
use NOR2X1  NOR2X1_44
timestamp 1515882711
transform -1 0 6328 0 1 2210
box 0 0 48 200
use FILL  FILL_MUX2X1_47
timestamp 1515882711
transform -1 0 6344 0 1 2210
box 0 0 16 200
use MUX2X1  MUX2X1_47
timestamp 1515882711
transform -1 0 6440 0 1 2210
box 0 0 96 200
use NOR2X1  NOR2X1_152
timestamp 1515882711
transform -1 0 6488 0 1 2210
box 0 0 48 200
use NOR3X1  NOR3X1_45
timestamp 1515882711
transform 1 0 6488 0 1 2210
box 0 0 128 200
use FILL  FILL_NAND2X1_72
timestamp 1515882711
transform 1 0 6616 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_72
timestamp 1515882711
transform 1 0 6632 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_89
timestamp 1515882711
transform -1 0 6744 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_218
timestamp 1515882711
transform 1 0 6744 0 1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_366
timestamp 1515882711
transform 1 0 6808 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_205
timestamp 1515882711
transform -1 0 6888 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_205
timestamp 1515882711
transform -1 0 6936 0 1 2210
box 0 0 48 200
use FILL  FILL_NAND2X1_326
timestamp 1515882711
transform 1 0 6936 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_326
timestamp 1515882711
transform 1 0 6952 0 1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_123
timestamp 1515882711
transform 1 0 7000 0 1 2210
box 0 0 16 200
use FILL  FILL_11_6_0
timestamp 1515882711
transform 1 0 7016 0 1 2210
box 0 0 16 200
use FILL  FILL_11_6_1
timestamp 1515882711
transform 1 0 7032 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_123
timestamp 1515882711
transform 1 0 7048 0 1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_123
timestamp 1515882711
transform 1 0 7240 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_107
timestamp 1515882711
transform -1 0 7320 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_107
timestamp 1515882711
transform -1 0 7368 0 1 2210
box 0 0 48 200
use NAND2X1  NAND2X1_424
timestamp 1515882711
transform 1 0 7368 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_476
timestamp 1515882711
transform -1 0 7480 0 1 2210
box 0 0 64 200
use FILL  FILL_INVX1_65
timestamp 1515882711
transform 1 0 7480 0 1 2210
box 0 0 16 200
use INVX1  INVX1_65
timestamp 1515882711
transform 1 0 7496 0 1 2210
box 0 0 32 200
use FILL  FILL_NAND2X1_140
timestamp 1515882711
transform 1 0 7528 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_140
timestamp 1515882711
transform 1 0 7544 0 1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_154
timestamp 1515882711
transform -1 0 7656 0 1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_127
timestamp 1515882711
transform -1 0 7672 0 1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_127
timestamp 1515882711
transform -1 0 7720 0 1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_154
timestamp 1515882711
transform -1 0 7736 0 1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_154
timestamp 1515882711
transform -1 0 7928 0 1 2210
box 0 0 192 200
use FILL  FILL_BUFX4_307
timestamp 1515882711
transform 1 0 7928 0 1 2210
box 0 0 16 200
use BUFX4  BUFX4_307
timestamp 1515882711
transform 1 0 7944 0 1 2210
box 0 0 64 200
use FILL  FILL_12_1
timestamp 1515882711
transform 1 0 8008 0 1 2210
box 0 0 16 200
use FILL  FILL_12_2
timestamp 1515882711
transform 1 0 8024 0 1 2210
box 0 0 16 200
use FILL  FILL_12_3
timestamp 1515882711
transform 1 0 8040 0 1 2210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_264
timestamp 1515882711
transform 1 0 8 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_264
timestamp 1515882711
transform 1 0 24 0 -1 2210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_172
timestamp 1515882711
transform 1 0 216 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_172
timestamp 1515882711
transform 1 0 232 0 -1 2210
box 0 0 192 200
use NOR2X1  NOR2X1_98
timestamp 1515882711
transform 1 0 424 0 -1 2210
box 0 0 48 200
use FILL  FILL_AOI21X1_22
timestamp 1515882711
transform -1 0 488 0 -1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_22
timestamp 1515882711
transform -1 0 552 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_240
timestamp 1515882711
transform 1 0 552 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_240
timestamp 1515882711
transform 1 0 568 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_7
timestamp 1515882711
transform -1 0 696 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_23
timestamp 1515882711
transform 1 0 696 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_23
timestamp 1515882711
transform 1 0 712 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_96
timestamp 1515882711
transform 1 0 776 0 -1 2210
box 0 0 48 200
use FILL  FILL_AOI21X1_20
timestamp 1515882711
transform -1 0 840 0 -1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_20
timestamp 1515882711
transform -1 0 904 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_0_0
timestamp 1515882711
transform 1 0 904 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1515882711
transform 1 0 920 0 -1 2210
box 0 0 16 200
use NAND3X1  NAND3X1_184
timestamp 1515882711
transform 1 0 936 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_207
timestamp 1515882711
transform 1 0 1000 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_207
timestamp 1515882711
transform 1 0 1016 0 -1 2210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_161
timestamp 1515882711
transform -1 0 1224 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_161
timestamp 1515882711
transform -1 0 1416 0 -1 2210
box 0 0 192 200
use NOR2X1  NOR2X1_105
timestamp 1515882711
transform -1 0 1464 0 -1 2210
box 0 0 48 200
use FILL  FILL_AOI21X1_29
timestamp 1515882711
transform -1 0 1480 0 -1 2210
box 0 0 16 200
use AOI21X1  AOI21X1_29
timestamp 1515882711
transform -1 0 1544 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_204
timestamp 1515882711
transform 1 0 1544 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_96
timestamp 1515882711
transform -1 0 1624 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_96
timestamp 1515882711
transform -1 0 1688 0 -1 2210
box 0 0 64 200
use FILL  FILL_INVX2_6
timestamp 1515882711
transform -1 0 1704 0 -1 2210
box 0 0 16 200
use INVX2  INVX2_6
timestamp 1515882711
transform -1 0 1736 0 -1 2210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_189
timestamp 1515882711
transform -1 0 1752 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_189
timestamp 1515882711
transform -1 0 1944 0 -1 2210
box 0 0 192 200
use FILL  FILL_10_1_0
timestamp 1515882711
transform 1 0 1944 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1515882711
transform 1 0 1960 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_173
timestamp 1515882711
transform 1 0 1976 0 -1 2210
box 0 0 64 200
use FILL  FILL_INVX2_13
timestamp 1515882711
transform -1 0 2056 0 -1 2210
box 0 0 16 200
use INVX2  INVX2_13
timestamp 1515882711
transform -1 0 2088 0 -1 2210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_232
timestamp 1515882711
transform -1 0 2104 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_232
timestamp 1515882711
transform -1 0 2296 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_180
timestamp 1515882711
transform 1 0 2296 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_146
timestamp 1515882711
transform -1 0 2376 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_146
timestamp 1515882711
transform -1 0 2440 0 -1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_389
timestamp 1515882711
transform 1 0 2440 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_389
timestamp 1515882711
transform 1 0 2456 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_458
timestamp 1515882711
transform -1 0 2568 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_267
timestamp 1515882711
transform 1 0 2568 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_267
timestamp 1515882711
transform 1 0 2584 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_19
timestamp 1515882711
transform 1 0 2776 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_448
timestamp 1515882711
transform -1 0 2888 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_219
timestamp 1515882711
transform 1 0 2888 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_446
timestamp 1515882711
transform 1 0 2952 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_2_0
timestamp 1515882711
transform 1 0 3000 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_2_1
timestamp 1515882711
transform 1 0 3016 0 -1 2210
box 0 0 16 200
use NAND3X1  NAND3X1_77
timestamp 1515882711
transform 1 0 3032 0 -1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_284
timestamp 1515882711
transform -1 0 3112 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_284
timestamp 1515882711
transform -1 0 3160 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_319
timestamp 1515882711
transform -1 0 3224 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_300
timestamp 1515882711
transform -1 0 3288 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_311
timestamp 1515882711
transform -1 0 3352 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_243
timestamp 1515882711
transform 1 0 3352 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_243
timestamp 1515882711
transform 1 0 3368 0 -1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_113
timestamp 1515882711
transform 1 0 3432 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_113
timestamp 1515882711
transform 1 0 3448 0 -1 2210
box 0 0 48 200
use FILL  FILL_NAND2X1_193
timestamp 1515882711
transform -1 0 3512 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_193
timestamp 1515882711
transform -1 0 3560 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_203
timestamp 1515882711
transform -1 0 3624 0 -1 2210
box 0 0 64 200
use FILL  FILL_INVX1_3
timestamp 1515882711
transform -1 0 3640 0 -1 2210
box 0 0 16 200
use INVX1  INVX1_3
timestamp 1515882711
transform -1 0 3672 0 -1 2210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_60
timestamp 1515882711
transform 1 0 3672 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_60
timestamp 1515882711
transform 1 0 3688 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_60
timestamp 1515882711
transform 1 0 3880 0 -1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_40
timestamp 1515882711
transform 1 0 3944 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_40
timestamp 1515882711
transform 1 0 3960 0 -1 2210
box 0 0 48 200
use FILL  FILL_10_3_0
timestamp 1515882711
transform 1 0 4008 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_3_1
timestamp 1515882711
transform 1 0 4024 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_321
timestamp 1515882711
transform 1 0 4040 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_33
timestamp 1515882711
transform 1 0 4104 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_22
timestamp 1515882711
transform -1 0 4216 0 -1 2210
box 0 0 48 200
use FILL  FILL_NAND2X1_288
timestamp 1515882711
transform -1 0 4232 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_288
timestamp 1515882711
transform -1 0 4280 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_34
timestamp 1515882711
transform 1 0 4280 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_52
timestamp 1515882711
transform -1 0 4360 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_52
timestamp 1515882711
transform -1 0 4552 0 -1 2210
box 0 0 192 200
use FILL  FILL_NAND2X1_32
timestamp 1515882711
transform 1 0 4552 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_32
timestamp 1515882711
transform 1 0 4568 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_52
timestamp 1515882711
transform -1 0 4680 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_48
timestamp 1515882711
transform -1 0 4744 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_158
timestamp 1515882711
transform 1 0 4744 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_158
timestamp 1515882711
transform 1 0 4760 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_322
timestamp 1515882711
transform -1 0 4888 0 -1 2210
box 0 0 64 200
use FILL  FILL_INVX1_69
timestamp 1515882711
transform -1 0 4904 0 -1 2210
box 0 0 16 200
use INVX1  INVX1_69
timestamp 1515882711
transform -1 0 4936 0 -1 2210
box 0 0 32 200
use FILL  FILL_BUFX4_76
timestamp 1515882711
transform 1 0 4936 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_76
timestamp 1515882711
transform 1 0 4952 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_275
timestamp 1515882711
transform 1 0 5016 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_4_0
timestamp 1515882711
transform 1 0 5032 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_4_1
timestamp 1515882711
transform 1 0 5048 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_275
timestamp 1515882711
transform 1 0 5064 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_83
timestamp 1515882711
transform -1 0 5144 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_83
timestamp 1515882711
transform -1 0 5336 0 -1 2210
box 0 0 192 200
use FILL  FILL_NAND2X1_64
timestamp 1515882711
transform 1 0 5336 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_64
timestamp 1515882711
transform 1 0 5352 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_83
timestamp 1515882711
transform -1 0 5464 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_105
timestamp 1515882711
transform 1 0 5464 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_105
timestamp 1515882711
transform 1 0 5480 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_105
timestamp 1515882711
transform 1 0 5672 0 -1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_88
timestamp 1515882711
transform -1 0 5752 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_88
timestamp 1515882711
transform -1 0 5800 0 -1 2210
box 0 0 48 200
use FILL  FILL_BUFX4_110
timestamp 1515882711
transform -1 0 5816 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_110
timestamp 1515882711
transform -1 0 5880 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_86
timestamp 1515882711
transform 1 0 5880 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_86
timestamp 1515882711
transform 1 0 5896 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_107
timestamp 1515882711
transform 1 0 5960 0 -1 2210
box 0 0 64 200
use FILL  FILL_NAND2X1_91
timestamp 1515882711
transform -1 0 6040 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_5_0
timestamp 1515882711
transform -1 0 6056 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_5_1
timestamp 1515882711
transform -1 0 6072 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_91
timestamp 1515882711
transform -1 0 6120 0 -1 2210
box 0 0 48 200
use FILL  FILL_MUX2X1_46
timestamp 1515882711
transform 1 0 6120 0 -1 2210
box 0 0 16 200
use MUX2X1  MUX2X1_46
timestamp 1515882711
transform 1 0 6136 0 -1 2210
box 0 0 96 200
use NOR2X1  NOR2X1_151
timestamp 1515882711
transform 1 0 6232 0 -1 2210
box 0 0 48 200
use FILL  FILL_BUFX4_1
timestamp 1515882711
transform 1 0 6280 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_1
timestamp 1515882711
transform 1 0 6296 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_89
timestamp 1515882711
transform -1 0 6376 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_89
timestamp 1515882711
transform -1 0 6568 0 -1 2210
box 0 0 192 200
use FILL  FILL_NAND2X1_320
timestamp 1515882711
transform -1 0 6584 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_320
timestamp 1515882711
transform -1 0 6632 0 -1 2210
box 0 0 48 200
use FILL  FILL_NAND2X1_188
timestamp 1515882711
transform 1 0 6632 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_188
timestamp 1515882711
transform 1 0 6648 0 -1 2210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_138
timestamp 1515882711
transform -1 0 6712 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_138
timestamp 1515882711
transform -1 0 6904 0 -1 2210
box 0 0 192 200
use FILL  FILL_NAND2X1_122
timestamp 1515882711
transform 1 0 6904 0 -1 2210
box 0 0 16 200
use NAND2X1  NAND2X1_122
timestamp 1515882711
transform 1 0 6920 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_138
timestamp 1515882711
transform -1 0 7032 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_193
timestamp 1515882711
transform -1 0 7048 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_6_0
timestamp 1515882711
transform -1 0 7064 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_6_1
timestamp 1515882711
transform -1 0 7080 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_193
timestamp 1515882711
transform -1 0 7144 0 -1 2210
box 0 0 64 200
use FILL  FILL_MUX2X1_23
timestamp 1515882711
transform 1 0 7144 0 -1 2210
box 0 0 16 200
use MUX2X1  MUX2X1_23
timestamp 1515882711
transform 1 0 7160 0 -1 2210
box 0 0 96 200
use FILL  FILL_DFFPOSX1_297
timestamp 1515882711
transform -1 0 7272 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_297
timestamp 1515882711
transform -1 0 7464 0 -1 2210
box 0 0 192 200
use FILL  FILL_BUFX4_152
timestamp 1515882711
transform -1 0 7480 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_152
timestamp 1515882711
transform -1 0 7544 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_10
timestamp 1515882711
transform 1 0 7544 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_11
timestamp 1515882711
transform -1 0 7672 0 -1 2210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_294
timestamp 1515882711
transform -1 0 7688 0 -1 2210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_294
timestamp 1515882711
transform -1 0 7880 0 -1 2210
box 0 0 192 200
use OAI21X1  OAI21X1_512
timestamp 1515882711
transform 1 0 7880 0 -1 2210
box 0 0 64 200
use FILL  FILL_BUFX4_314
timestamp 1515882711
transform 1 0 7944 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_314
timestamp 1515882711
transform 1 0 7960 0 -1 2210
box 0 0 64 200
use FILL  FILL_11_1
timestamp 1515882711
transform -1 0 8040 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_2
timestamp 1515882711
transform -1 0 8056 0 -1 2210
box 0 0 16 200
use FILL  FILL_BUFX4_68
timestamp 1515882711
transform -1 0 24 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_68
timestamp 1515882711
transform -1 0 88 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_261
timestamp 1515882711
transform -1 0 104 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_261
timestamp 1515882711
transform -1 0 296 0 1 1810
box 0 0 192 200
use FILL  FILL_BUFX4_215
timestamp 1515882711
transform -1 0 312 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_215
timestamp 1515882711
transform -1 0 376 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_226
timestamp 1515882711
transform 1 0 376 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_226
timestamp 1515882711
transform 1 0 392 0 1 1810
box 0 0 192 200
use FILL  FILL_AOI21X1_58
timestamp 1515882711
transform 1 0 584 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_58
timestamp 1515882711
transform 1 0 600 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_134
timestamp 1515882711
transform -1 0 712 0 1 1810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_259
timestamp 1515882711
transform 1 0 712 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_259
timestamp 1515882711
transform 1 0 728 0 1 1810
box 0 0 192 200
use FILL  FILL_BUFX4_183
timestamp 1515882711
transform -1 0 936 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_0
timestamp 1515882711
transform -1 0 952 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1515882711
transform -1 0 968 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_183
timestamp 1515882711
transform -1 0 1032 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_211
timestamp 1515882711
transform 1 0 1032 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_211
timestamp 1515882711
transform 1 0 1048 0 1 1810
box 0 0 192 200
use FILL  FILL_AOI21X1_44
timestamp 1515882711
transform 1 0 1240 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_44
timestamp 1515882711
transform 1 0 1256 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_120
timestamp 1515882711
transform -1 0 1368 0 1 1810
box 0 0 48 200
use FILL  FILL_BUFX4_157
timestamp 1515882711
transform 1 0 1368 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_157
timestamp 1515882711
transform 1 0 1384 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_277
timestamp 1515882711
transform -1 0 1464 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_277
timestamp 1515882711
transform -1 0 1528 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_408
timestamp 1515882711
transform -1 0 1592 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_35
timestamp 1515882711
transform -1 0 1608 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_35
timestamp 1515882711
transform -1 0 1672 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_114
timestamp 1515882711
transform -1 0 1720 0 1 1810
box 0 0 48 200
use FILL  FILL_AOI21X1_38
timestamp 1515882711
transform -1 0 1736 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_38
timestamp 1515882711
transform -1 0 1800 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_205
timestamp 1515882711
transform 1 0 1800 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_205
timestamp 1515882711
transform 1 0 1816 0 1 1810
box 0 0 192 200
use FILL  FILL_9_1_0
timestamp 1515882711
transform -1 0 2024 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1515882711
transform -1 0 2040 0 1 1810
box 0 0 16 200
use FILL  FILL_AOI21X1_55
timestamp 1515882711
transform -1 0 2056 0 1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_55
timestamp 1515882711
transform -1 0 2120 0 1 1810
box 0 0 64 200
use FILL  FILL_INVX8_1
timestamp 1515882711
transform 1 0 2120 0 1 1810
box 0 0 16 200
use INVX8  INVX8_1
timestamp 1515882711
transform 1 0 2136 0 1 1810
box 0 0 80 200
use FILL  FILL_BUFX4_168
timestamp 1515882711
transform -1 0 2232 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_168
timestamp 1515882711
transform -1 0 2296 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_190
timestamp 1515882711
transform 1 0 2296 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_190
timestamp 1515882711
transform 1 0 2312 0 1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_164
timestamp 1515882711
transform -1 0 2392 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_164
timestamp 1515882711
transform -1 0 2440 0 1 1810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_12
timestamp 1515882711
transform 1 0 2440 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1515882711
transform 1 0 2456 0 1 1810
box 0 0 192 200
use FILL  FILL_INVX1_66
timestamp 1515882711
transform 1 0 2648 0 1 1810
box 0 0 16 200
use INVX1  INVX1_66
timestamp 1515882711
transform 1 0 2664 0 1 1810
box 0 0 32 200
use FILL  FILL_INVX8_12
timestamp 1515882711
transform -1 0 2712 0 1 1810
box 0 0 16 200
use INVX8  INVX8_12
timestamp 1515882711
transform -1 0 2792 0 1 1810
box 0 0 80 200
use FILL  FILL_BUFX4_237
timestamp 1515882711
transform -1 0 2808 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_237
timestamp 1515882711
transform -1 0 2872 0 1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_191
timestamp 1515882711
transform 1 0 2872 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_191
timestamp 1515882711
transform 1 0 2888 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_199
timestamp 1515882711
transform -1 0 3000 0 1 1810
box 0 0 64 200
use FILL  FILL_9_2_0
timestamp 1515882711
transform -1 0 3016 0 1 1810
box 0 0 16 200
use FILL  FILL_9_2_1
timestamp 1515882711
transform -1 0 3032 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_359
timestamp 1515882711
transform -1 0 3096 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_46
timestamp 1515882711
transform 1 0 3096 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_46
timestamp 1515882711
transform 1 0 3112 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_202
timestamp 1515882711
transform 1 0 3176 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_147
timestamp 1515882711
transform -1 0 3288 0 1 1810
box 0 0 48 200
use FILL  FILL_NAND2X1_195
timestamp 1515882711
transform -1 0 3304 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_195
timestamp 1515882711
transform -1 0 3352 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_2
timestamp 1515882711
transform 1 0 3352 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_80
timestamp 1515882711
transform 1 0 3416 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_41
timestamp 1515882711
transform -1 0 3528 0 1 1810
box 0 0 48 200
use FILL  FILL_NAND2X1_322
timestamp 1515882711
transform -1 0 3544 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_322
timestamp 1515882711
transform -1 0 3592 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_78
timestamp 1515882711
transform -1 0 3656 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_233
timestamp 1515882711
transform 1 0 3656 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_233
timestamp 1515882711
transform 1 0 3672 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_161
timestamp 1515882711
transform 1 0 3736 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_161
timestamp 1515882711
transform 1 0 3752 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_43
timestamp 1515882711
transform 1 0 3816 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_43
timestamp 1515882711
transform 1 0 3832 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_411
timestamp 1515882711
transform 1 0 3896 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_210
timestamp 1515882711
transform 1 0 3960 0 1 1810
box 0 0 64 200
use FILL  FILL_9_3_0
timestamp 1515882711
transform -1 0 4040 0 1 1810
box 0 0 16 200
use FILL  FILL_9_3_1
timestamp 1515882711
transform -1 0 4056 0 1 1810
box 0 0 16 200
use NOR2X1  NOR2X1_67
timestamp 1515882711
transform -1 0 4104 0 1 1810
box 0 0 48 200
use FILL  FILL_NAND2X1_350
timestamp 1515882711
transform -1 0 4120 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_350
timestamp 1515882711
transform -1 0 4168 0 1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_211
timestamp 1515882711
transform 1 0 4168 0 1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_36
timestamp 1515882711
transform 1 0 4232 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_300
timestamp 1515882711
transform -1 0 4312 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_300
timestamp 1515882711
transform -1 0 4376 0 1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_49
timestamp 1515882711
transform -1 0 4392 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_49
timestamp 1515882711
transform -1 0 4440 0 1 1810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_86
timestamp 1515882711
transform 1 0 4440 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_86
timestamp 1515882711
transform 1 0 4456 0 1 1810
box 0 0 192 200
use FILL  FILL_NAND2X1_67
timestamp 1515882711
transform 1 0 4648 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_67
timestamp 1515882711
transform 1 0 4664 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_86
timestamp 1515882711
transform -1 0 4776 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_304
timestamp 1515882711
transform -1 0 4792 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_304
timestamp 1515882711
transform -1 0 4856 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_49
timestamp 1515882711
transform 1 0 4856 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_49
timestamp 1515882711
transform 1 0 4872 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_246
timestamp 1515882711
transform -1 0 4952 0 1 1810
box 0 0 16 200
use FILL  FILL_9_4_0
timestamp 1515882711
transform -1 0 4968 0 1 1810
box 0 0 16 200
use FILL  FILL_9_4_1
timestamp 1515882711
transform -1 0 4984 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_246
timestamp 1515882711
transform -1 0 5176 0 1 1810
box 0 0 192 200
use FILL  FILL_NAND2X1_279
timestamp 1515882711
transform 1 0 5176 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_279
timestamp 1515882711
transform 1 0 5192 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_246
timestamp 1515882711
transform -1 0 5304 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_48
timestamp 1515882711
transform 1 0 5304 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_48
timestamp 1515882711
transform 1 0 5320 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_223
timestamp 1515882711
transform 1 0 5384 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_223
timestamp 1515882711
transform 1 0 5400 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_281
timestamp 1515882711
transform 1 0 5464 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_281
timestamp 1515882711
transform 1 0 5480 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_145
timestamp 1515882711
transform 1 0 5544 0 1 1810
box 0 0 48 200
use NOR3X1  NOR3X1_12
timestamp 1515882711
transform 1 0 5592 0 1 1810
box 0 0 128 200
use FILL  FILL_DFFPOSX1_68
timestamp 1515882711
transform -1 0 5736 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_68
timestamp 1515882711
transform -1 0 5928 0 1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_423
timestamp 1515882711
transform -1 0 5992 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_457
timestamp 1515882711
transform 1 0 5992 0 1 1810
box 0 0 64 200
use FILL  FILL_9_5_0
timestamp 1515882711
transform -1 0 6072 0 1 1810
box 0 0 16 200
use FILL  FILL_9_5_1
timestamp 1515882711
transform -1 0 6088 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_406
timestamp 1515882711
transform -1 0 6136 0 1 1810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_317
timestamp 1515882711
transform -1 0 6152 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_317
timestamp 1515882711
transform -1 0 6344 0 1 1810
box 0 0 192 200
use FILL  FILL_DFFPOSX1_332
timestamp 1515882711
transform -1 0 6360 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_332
timestamp 1515882711
transform -1 0 6552 0 1 1810
box 0 0 192 200
use FILL  FILL_BUFX4_8
timestamp 1515882711
transform -1 0 6568 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_8
timestamp 1515882711
transform -1 0 6632 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_358
timestamp 1515882711
transform -1 0 6696 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_198
timestamp 1515882711
transform -1 0 6760 0 1 1810
box 0 0 64 200
use FILL  FILL_MUX2X1_37
timestamp 1515882711
transform 1 0 6760 0 1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_37
timestamp 1515882711
transform 1 0 6776 0 1 1810
box 0 0 96 200
use NAND2X1  NAND2X1_435
timestamp 1515882711
transform 1 0 6872 0 1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_438
timestamp 1515882711
transform 1 0 6920 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_490
timestamp 1515882711
transform -1 0 7032 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_312
timestamp 1515882711
transform -1 0 7048 0 1 1810
box 0 0 16 200
use FILL  FILL_9_6_0
timestamp 1515882711
transform -1 0 7064 0 1 1810
box 0 0 16 200
use FILL  FILL_9_6_1
timestamp 1515882711
transform -1 0 7080 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_312
timestamp 1515882711
transform -1 0 7272 0 1 1810
box 0 0 192 200
use FILL  FILL_BUFX4_194
timestamp 1515882711
transform 1 0 7272 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_194
timestamp 1515882711
transform 1 0 7288 0 1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_270
timestamp 1515882711
transform 1 0 7352 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_270
timestamp 1515882711
transform 1 0 7368 0 1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_289
timestamp 1515882711
transform 1 0 7432 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_289
timestamp 1515882711
transform 1 0 7448 0 1 1810
box 0 0 48 200
use FILL  FILL_BUFX4_271
timestamp 1515882711
transform 1 0 7496 0 1 1810
box 0 0 16 200
use BUFX4  BUFX4_271
timestamp 1515882711
transform 1 0 7512 0 1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_266
timestamp 1515882711
transform 1 0 7576 0 1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_266
timestamp 1515882711
transform 1 0 7592 0 1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_4
timestamp 1515882711
transform 1 0 7640 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_5
timestamp 1515882711
transform -1 0 7768 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_511
timestamp 1515882711
transform 1 0 7768 0 1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_291
timestamp 1515882711
transform -1 0 7848 0 1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_291
timestamp 1515882711
transform -1 0 8040 0 1 1810
box 0 0 192 200
use FILL  FILL_10_1
timestamp 1515882711
transform 1 0 8040 0 1 1810
box 0 0 16 200
use NOR2X1  NOR2X1_81
timestamp 1515882711
transform -1 0 56 0 -1 1810
box 0 0 48 200
use FILL  FILL_AOI21X1_5
timestamp 1515882711
transform -1 0 72 0 -1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_5
timestamp 1515882711
transform -1 0 136 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_31
timestamp 1515882711
transform -1 0 200 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_30
timestamp 1515882711
transform 1 0 200 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_32
timestamp 1515882711
transform -1 0 328 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_207
timestamp 1515882711
transform 1 0 328 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_209
timestamp 1515882711
transform -1 0 456 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_208
timestamp 1515882711
transform 1 0 456 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1515882711
transform -1 0 584 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_10
timestamp 1515882711
transform 1 0 584 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_79
timestamp 1515882711
transform 1 0 648 0 -1 1810
box 0 0 48 200
use FILL  FILL_AOI21X1_3
timestamp 1515882711
transform -1 0 712 0 -1 1810
box 0 0 16 200
use AOI21X1  AOI21X1_3
timestamp 1515882711
transform -1 0 776 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_171
timestamp 1515882711
transform 1 0 776 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_171
timestamp 1515882711
transform 1 0 792 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_186
timestamp 1515882711
transform 1 0 856 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_0_0
timestamp 1515882711
transform 1 0 920 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1515882711
transform 1 0 936 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_187
timestamp 1515882711
transform 1 0 952 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_185
timestamp 1515882711
transform 1 0 1016 0 -1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_144
timestamp 1515882711
transform 1 0 1080 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_144
timestamp 1515882711
transform 1 0 1096 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_205
timestamp 1515882711
transform -1 0 1208 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_409
timestamp 1515882711
transform -1 0 1272 0 -1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_40
timestamp 1515882711
transform -1 0 1400 0 -1 1810
box 0 0 128 200
use NAND3X1  NAND3X1_28
timestamp 1515882711
transform 1 0 1400 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_316
timestamp 1515882711
transform -1 0 1528 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_27
timestamp 1515882711
transform 1 0 1528 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_315
timestamp 1515882711
transform -1 0 1656 0 -1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_18
timestamp 1515882711
transform 1 0 1656 0 -1 1810
box 0 0 128 200
use NAND3X1  NAND3X1_5
timestamp 1515882711
transform -1 0 1848 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_6
timestamp 1515882711
transform -1 0 1912 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_183
timestamp 1515882711
transform -1 0 1976 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_1_0
timestamp 1515882711
transform 1 0 1976 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1515882711
transform 1 0 1992 0 -1 1810
box 0 0 16 200
use NOR2X1  NOR2X1_131
timestamp 1515882711
transform 1 0 2008 0 -1 1810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_222
timestamp 1515882711
transform -1 0 2072 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_222
timestamp 1515882711
transform -1 0 2264 0 -1 1810
box 0 0 192 200
use NAND3X1  NAND3X1_182
timestamp 1515882711
transform 1 0 2264 0 -1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_158
timestamp 1515882711
transform -1 0 2344 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_158
timestamp 1515882711
transform -1 0 2392 0 -1 1810
box 0 0 48 200
use FILL  FILL_NAND2X1_162
timestamp 1515882711
transform -1 0 2408 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_162
timestamp 1515882711
transform -1 0 2456 0 -1 1810
box 0 0 48 200
use FILL  FILL_NAND2X1_147
timestamp 1515882711
transform 1 0 2456 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_147
timestamp 1515882711
transform 1 0 2472 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_162
timestamp 1515882711
transform -1 0 2584 0 -1 1810
box 0 0 64 200
use FILL  FILL_INVX2_28
timestamp 1515882711
transform -1 0 2600 0 -1 1810
box 0 0 16 200
use INVX2  INVX2_28
timestamp 1515882711
transform -1 0 2632 0 -1 1810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_178
timestamp 1515882711
transform -1 0 2648 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_178
timestamp 1515882711
transform -1 0 2840 0 -1 1810
box 0 0 192 200
use FILL  FILL_NAND2X1_376
timestamp 1515882711
transform 1 0 2840 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_376
timestamp 1515882711
transform 1 0 2856 0 -1 1810
box 0 0 48 200
use FILL  FILL_NAND2X1_206
timestamp 1515882711
transform 1 0 2904 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_206
timestamp 1515882711
transform 1 0 2920 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_2_0
timestamp 1515882711
transform -1 0 2984 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_2_1
timestamp 1515882711
transform -1 0 3000 0 -1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_443
timestamp 1515882711
transform -1 0 3064 0 -1 1810
box 0 0 64 200
use FILL  FILL_INVX1_89
timestamp 1515882711
transform -1 0 3080 0 -1 1810
box 0 0 16 200
use INVX1  INVX1_89
timestamp 1515882711
transform -1 0 3112 0 -1 1810
box 0 0 32 200
use FILL  FILL_DFFPOSX1_350
timestamp 1515882711
transform -1 0 3128 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_350
timestamp 1515882711
transform -1 0 3320 0 -1 1810
box 0 0 192 200
use FILL  FILL_BUFX4_61
timestamp 1515882711
transform 1 0 3320 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_61
timestamp 1515882711
transform 1 0 3336 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_13
timestamp 1515882711
transform -1 0 3464 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_81
timestamp 1515882711
transform -1 0 3528 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_18
timestamp 1515882711
transform 1 0 3528 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_18
timestamp 1515882711
transform 1 0 3544 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_174
timestamp 1515882711
transform 1 0 3608 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_174
timestamp 1515882711
transform 1 0 3624 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_251
timestamp 1515882711
transform 1 0 3688 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_251
timestamp 1515882711
transform 1 0 3704 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_252
timestamp 1515882711
transform -1 0 3784 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_252
timestamp 1515882711
transform -1 0 3848 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_253
timestamp 1515882711
transform 1 0 3848 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_253
timestamp 1515882711
transform 1 0 3864 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_67
timestamp 1515882711
transform -1 0 3992 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_3_0
timestamp 1515882711
transform 1 0 3992 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_3_1
timestamp 1515882711
transform 1 0 4008 0 -1 1810
box 0 0 16 200
use NAND3X1  NAND3X1_69
timestamp 1515882711
transform 1 0 4024 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_247
timestamp 1515882711
transform 1 0 4088 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_245
timestamp 1515882711
transform 1 0 4152 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_213
timestamp 1515882711
transform 1 0 4216 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_214
timestamp 1515882711
transform -1 0 4344 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_354
timestamp 1515882711
transform -1 0 4408 0 -1 1810
box 0 0 64 200
use FILL  FILL_INVX1_86
timestamp 1515882711
transform -1 0 4424 0 -1 1810
box 0 0 16 200
use INVX1  INVX1_86
timestamp 1515882711
transform -1 0 4456 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_69
timestamp 1515882711
transform -1 0 4520 0 -1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_69
timestamp 1515882711
transform -1 0 4536 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_69
timestamp 1515882711
transform -1 0 4728 0 -1 1810
box 0 0 192 200
use FILL  FILL_INVX1_85
timestamp 1515882711
transform 1 0 4728 0 -1 1810
box 0 0 16 200
use INVX1  INVX1_85
timestamp 1515882711
transform 1 0 4744 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_353
timestamp 1515882711
transform 1 0 4776 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_77
timestamp 1515882711
transform -1 0 4856 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_77
timestamp 1515882711
transform -1 0 4920 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_324
timestamp 1515882711
transform 1 0 4920 0 -1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_309
timestamp 1515882711
transform -1 0 5000 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_309
timestamp 1515882711
transform -1 0 5048 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_4_0
timestamp 1515882711
transform 1 0 5048 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_4_1
timestamp 1515882711
transform 1 0 5064 0 -1 1810
box 0 0 16 200
use FILL  FILL_NAND2X1_310
timestamp 1515882711
transform 1 0 5080 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_310
timestamp 1515882711
transform 1 0 5096 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_68
timestamp 1515882711
transform 1 0 5144 0 -1 1810
box 0 0 64 200
use FILL  FILL_NAND2X1_90
timestamp 1515882711
transform -1 0 5224 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_90
timestamp 1515882711
transform -1 0 5272 0 -1 1810
box 0 0 48 200
use FILL  FILL_DFFPOSX1_33
timestamp 1515882711
transform -1 0 5288 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_33
timestamp 1515882711
transform -1 0 5480 0 -1 1810
box 0 0 192 200
use NOR2X1  NOR2X1_40
timestamp 1515882711
transform 1 0 5480 0 -1 1810
box 0 0 48 200
use OAI22X1  OAI22X1_1
timestamp 1515882711
transform 1 0 5528 0 -1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_143
timestamp 1515882711
transform -1 0 5656 0 -1 1810
box 0 0 48 200
use FILL  FILL_MUX2X1_1
timestamp 1515882711
transform 1 0 5656 0 -1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_1
timestamp 1515882711
transform 1 0 5672 0 -1 1810
box 0 0 96 200
use NAND2X1  NAND2X1_402
timestamp 1515882711
transform 1 0 5768 0 -1 1810
box 0 0 48 200
use FILL  FILL_MUX2X1_42
timestamp 1515882711
transform -1 0 5832 0 -1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_42
timestamp 1515882711
transform -1 0 5928 0 -1 1810
box 0 0 96 200
use FILL  FILL_DFFPOSX1_315
timestamp 1515882711
transform -1 0 5944 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_315
timestamp 1515882711
transform -1 0 6136 0 -1 1810
box 0 0 192 200
use FILL  FILL_8_5_0
timestamp 1515882711
transform 1 0 6136 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_5_1
timestamp 1515882711
transform 1 0 6152 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_404
timestamp 1515882711
transform 1 0 6168 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_434
timestamp 1515882711
transform -1 0 6280 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_70
timestamp 1515882711
transform 1 0 6280 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_70
timestamp 1515882711
transform 1 0 6296 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_72
timestamp 1515882711
transform -1 0 6376 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_72
timestamp 1515882711
transform -1 0 6440 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_421
timestamp 1515882711
transform 1 0 6440 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_475
timestamp 1515882711
transform -1 0 6552 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_6
timestamp 1515882711
transform 1 0 6552 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_6
timestamp 1515882711
transform 1 0 6568 0 -1 1810
box 0 0 64 200
use FILL  FILL_BUFX4_208
timestamp 1515882711
transform -1 0 6648 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_208
timestamp 1515882711
transform -1 0 6712 0 -1 1810
box 0 0 64 200
use FILL  FILL_MUX2X1_27
timestamp 1515882711
transform -1 0 6728 0 -1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_27
timestamp 1515882711
transform -1 0 6824 0 -1 1810
box 0 0 96 200
use FILL  FILL_DFFPOSX1_308
timestamp 1515882711
transform -1 0 6840 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_308
timestamp 1515882711
transform -1 0 7032 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_487
timestamp 1515882711
transform -1 0 7096 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_6_0
timestamp 1515882711
transform 1 0 7096 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_6_1
timestamp 1515882711
transform 1 0 7112 0 -1 1810
box 0 0 16 200
use FILL  FILL_DFFPOSX1_296
timestamp 1515882711
transform 1 0 7128 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_296
timestamp 1515882711
transform 1 0 7144 0 -1 1810
box 0 0 192 200
use OAI21X1  OAI21X1_16
timestamp 1515882711
transform 1 0 7336 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_15
timestamp 1515882711
transform -1 0 7464 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_497
timestamp 1515882711
transform 1 0 7464 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_496
timestamp 1515882711
transform 1 0 7528 0 -1 1810
box 0 0 64 200
use FILL  FILL_DFFPOSX1_268
timestamp 1515882711
transform -1 0 7608 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_268
timestamp 1515882711
transform -1 0 7800 0 -1 1810
box 0 0 192 200
use FILL  FILL_DFFPOSX1_289
timestamp 1515882711
transform 1 0 7800 0 -1 1810
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_289
timestamp 1515882711
transform 1 0 7816 0 -1 1810
box 0 0 192 200
use FILL  FILL_9_1
timestamp 1515882711
transform -1 0 8024 0 -1 1810
box 0 0 16 200
use FILL  FILL_9_2
timestamp 1515882711
transform -1 0 8040 0 -1 1810
box 0 0 16 200
use FILL  FILL_9_3
timestamp 1515882711
transform -1 0 8056 0 -1 1810
box 0 0 16 200
use FILL  FILL_DFFPOSX1_256
timestamp 1515882711
transform 1 0 8 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_256
timestamp 1515882711
transform 1 0 24 0 1 1410
box 0 0 192 200
use FILL  FILL_BUFX4_139
timestamp 1515882711
transform 1 0 216 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_139
timestamp 1515882711
transform 1 0 232 0 1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_138
timestamp 1515882711
transform 1 0 296 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_138
timestamp 1515882711
transform 1 0 312 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_29
timestamp 1515882711
transform 1 0 376 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_206
timestamp 1515882711
transform 1 0 440 0 1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_60
timestamp 1515882711
transform -1 0 520 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_60
timestamp 1515882711
transform -1 0 584 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1515882711
transform 1 0 584 0 1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_58
timestamp 1515882711
transform -1 0 664 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_58
timestamp 1515882711
transform -1 0 728 0 1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_175
timestamp 1515882711
transform -1 0 744 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_175
timestamp 1515882711
transform -1 0 808 0 1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_167
timestamp 1515882711
transform -1 0 824 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_167
timestamp 1515882711
transform -1 0 1016 0 1 1410
box 0 0 192 200
use FILL  FILL_7_0_0
timestamp 1515882711
transform 1 0 1016 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1515882711
transform 1 0 1032 0 1 1410
box 0 0 16 200
use FILL  FILL_BUFX4_20
timestamp 1515882711
transform 1 0 1048 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_20
timestamp 1515882711
transform 1 0 1064 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_160
timestamp 1515882711
transform -1 0 1192 0 1 1410
box 0 0 64 200
use FILL  FILL_INVX2_12
timestamp 1515882711
transform -1 0 1208 0 1 1410
box 0 0 16 200
use INVX2  INVX2_12
timestamp 1515882711
transform -1 0 1240 0 1 1410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_176
timestamp 1515882711
transform -1 0 1256 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_176
timestamp 1515882711
transform -1 0 1448 0 1 1410
box 0 0 192 200
use FILL  FILL_INVX2_24
timestamp 1515882711
transform -1 0 1464 0 1 1410
box 0 0 16 200
use INVX2  INVX2_24
timestamp 1515882711
transform -1 0 1496 0 1 1410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_243
timestamp 1515882711
transform -1 0 1512 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_243
timestamp 1515882711
transform -1 0 1704 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_191
timestamp 1515882711
transform 1 0 1704 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_175
timestamp 1515882711
transform -1 0 1784 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_175
timestamp 1515882711
transform -1 0 1832 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_295
timestamp 1515882711
transform -1 0 1896 0 1 1410
box 0 0 64 200
use FILL  FILL_7_1_0
timestamp 1515882711
transform -1 0 1912 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1515882711
transform -1 0 1928 0 1 1410
box 0 0 16 200
use NOR3X1  NOR3X1_14
timestamp 1515882711
transform -1 0 2056 0 1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_296
timestamp 1515882711
transform -1 0 2120 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_400
timestamp 1515882711
transform -1 0 2184 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_399
timestamp 1515882711
transform 1 0 2184 0 1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_38
timestamp 1515882711
transform 1 0 2248 0 1 1410
box 0 0 128 200
use FILL  FILL_NAND2X1_313
timestamp 1515882711
transform -1 0 2392 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_313
timestamp 1515882711
transform -1 0 2440 0 1 1410
box 0 0 48 200
use FILL  FILL_INVX2_21
timestamp 1515882711
transform -1 0 2456 0 1 1410
box 0 0 16 200
use INVX2  INVX2_21
timestamp 1515882711
transform -1 0 2488 0 1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_188
timestamp 1515882711
transform 1 0 2488 0 1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_241
timestamp 1515882711
transform -1 0 2568 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_241
timestamp 1515882711
transform -1 0 2760 0 1 1410
box 0 0 192 200
use FILL  FILL_BUFX4_228
timestamp 1515882711
transform 1 0 2760 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_228
timestamp 1515882711
transform 1 0 2776 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_378
timestamp 1515882711
transform 1 0 2840 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_378
timestamp 1515882711
transform 1 0 2856 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_447
timestamp 1515882711
transform -1 0 2968 0 1 1410
box 0 0 64 200
use FILL  FILL_INVX1_11
timestamp 1515882711
transform -1 0 2984 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_0
timestamp 1515882711
transform -1 0 3000 0 1 1410
box 0 0 16 200
use FILL  FILL_7_2_1
timestamp 1515882711
transform -1 0 3016 0 1 1410
box 0 0 16 200
use INVX1  INVX1_11
timestamp 1515882711
transform -1 0 3048 0 1 1410
box 0 0 32 200
use FILL  FILL_DFFPOSX1_352
timestamp 1515882711
transform -1 0 3064 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_352
timestamp 1515882711
transform -1 0 3256 0 1 1410
box 0 0 192 200
use FILL  FILL_BUFX4_289
timestamp 1515882711
transform -1 0 3272 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_289
timestamp 1515882711
transform -1 0 3336 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_36
timestamp 1515882711
transform 1 0 3336 0 1 1410
box 0 0 48 200
use FILL  FILL_INVX1_88
timestamp 1515882711
transform -1 0 3400 0 1 1410
box 0 0 16 200
use INVX1  INVX1_88
timestamp 1515882711
transform -1 0 3432 0 1 1410
box 0 0 32 200
use FILL  FILL_NAND2X1_321
timestamp 1515882711
transform 1 0 3432 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_321
timestamp 1515882711
transform 1 0 3448 0 1 1410
box 0 0 48 200
use FILL  FILL_BUFX4_181
timestamp 1515882711
transform 1 0 3496 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_181
timestamp 1515882711
transform 1 0 3512 0 1 1410
box 0 0 64 200
use FILL  FILL_INVX8_10
timestamp 1515882711
transform -1 0 3592 0 1 1410
box 0 0 16 200
use INVX8  INVX8_10
timestamp 1515882711
transform -1 0 3672 0 1 1410
box 0 0 80 200
use FILL  FILL_BUFX4_41
timestamp 1515882711
transform -1 0 3688 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_41
timestamp 1515882711
transform -1 0 3752 0 1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_42
timestamp 1515882711
transform 1 0 3752 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_42
timestamp 1515882711
transform 1 0 3768 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_425
timestamp 1515882711
transform 1 0 3832 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_244
timestamp 1515882711
transform 1 0 3896 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_311
timestamp 1515882711
transform 1 0 3960 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_311
timestamp 1515882711
transform 1 0 3976 0 1 1410
box 0 0 48 200
use FILL  FILL_7_3_0
timestamp 1515882711
transform -1 0 4040 0 1 1410
box 0 0 16 200
use FILL  FILL_7_3_1
timestamp 1515882711
transform -1 0 4056 0 1 1410
box 0 0 16 200
use NOR2X1  NOR2X1_74
timestamp 1515882711
transform -1 0 4104 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_356
timestamp 1515882711
transform -1 0 4120 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_356
timestamp 1515882711
transform -1 0 4168 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_317
timestamp 1515882711
transform -1 0 4184 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_317
timestamp 1515882711
transform -1 0 4232 0 1 1410
box 0 0 48 200
use FILL  FILL_INVX1_91
timestamp 1515882711
transform 1 0 4232 0 1 1410
box 0 0 16 200
use INVX1  INVX1_91
timestamp 1515882711
transform 1 0 4248 0 1 1410
box 0 0 32 200
use FILL  FILL_BUFX2_5
timestamp 1515882711
transform 1 0 4280 0 1 1410
box 0 0 16 200
use BUFX2  BUFX2_5
timestamp 1515882711
transform 1 0 4296 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_318
timestamp 1515882711
transform 1 0 4344 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_318
timestamp 1515882711
transform 1 0 4360 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_319
timestamp 1515882711
transform 1 0 4408 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_319
timestamp 1515882711
transform 1 0 4424 0 1 1410
box 0 0 48 200
use FILL  FILL_BUFX4_198
timestamp 1515882711
transform 1 0 4472 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_198
timestamp 1515882711
transform 1 0 4488 0 1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_65
timestamp 1515882711
transform -1 0 4568 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_65
timestamp 1515882711
transform -1 0 4760 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_65
timestamp 1515882711
transform 1 0 4760 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_45
timestamp 1515882711
transform -1 0 4840 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_45
timestamp 1515882711
transform -1 0 4888 0 1 1410
box 0 0 48 200
use FILL  FILL_INVX1_70
timestamp 1515882711
transform 1 0 4888 0 1 1410
box 0 0 16 200
use INVX1  INVX1_70
timestamp 1515882711
transform 1 0 4904 0 1 1410
box 0 0 32 200
use FILL  FILL_NAND2X1_287
timestamp 1515882711
transform 1 0 4936 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_287
timestamp 1515882711
transform 1 0 4952 0 1 1410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_30
timestamp 1515882711
transform -1 0 5016 0 1 1410
box 0 0 16 200
use FILL  FILL_7_4_0
timestamp 1515882711
transform -1 0 5032 0 1 1410
box 0 0 16 200
use FILL  FILL_7_4_1
timestamp 1515882711
transform -1 0 5048 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_30
timestamp 1515882711
transform -1 0 5240 0 1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_35
timestamp 1515882711
transform 1 0 5240 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_57
timestamp 1515882711
transform 1 0 5304 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_57
timestamp 1515882711
transform 1 0 5320 0 1 1410
box 0 0 48 200
use FILL  FILL_BUFX4_266
timestamp 1515882711
transform -1 0 5384 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_266
timestamp 1515882711
transform -1 0 5448 0 1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_81
timestamp 1515882711
transform 1 0 5448 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_81
timestamp 1515882711
transform 1 0 5464 0 1 1410
box 0 0 192 200
use FILL  FILL_NAND2X1_62
timestamp 1515882711
transform 1 0 5656 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_62
timestamp 1515882711
transform 1 0 5672 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_81
timestamp 1515882711
transform -1 0 5784 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_33
timestamp 1515882711
transform 1 0 5784 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_33
timestamp 1515882711
transform 1 0 5800 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_53
timestamp 1515882711
transform -1 0 5912 0 1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_104
timestamp 1515882711
transform -1 0 5928 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_104
timestamp 1515882711
transform -1 0 6120 0 1 1410
box 0 0 192 200
use FILL  FILL_7_5_0
timestamp 1515882711
transform 1 0 6120 0 1 1410
box 0 0 16 200
use FILL  FILL_7_5_1
timestamp 1515882711
transform 1 0 6136 0 1 1410
box 0 0 16 200
use FILL  FILL_NAND2X1_86
timestamp 1515882711
transform 1 0 6152 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_86
timestamp 1515882711
transform 1 0 6168 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_104
timestamp 1515882711
transform -1 0 6280 0 1 1410
box 0 0 64 200
use OAI22X1  OAI22X1_8
timestamp 1515882711
transform 1 0 6280 0 1 1410
box 0 0 80 200
use NOR2X1  NOR2X1_73
timestamp 1515882711
transform -1 0 6408 0 1 1410
box 0 0 48 200
use FILL  FILL_MUX2X1_41
timestamp 1515882711
transform -1 0 6424 0 1 1410
box 0 0 16 200
use MUX2X1  MUX2X1_41
timestamp 1515882711
transform -1 0 6520 0 1 1410
box 0 0 96 200
use FILL  FILL_NAND2X1_105
timestamp 1515882711
transform -1 0 6536 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_105
timestamp 1515882711
transform -1 0 6584 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_402
timestamp 1515882711
transform 1 0 6584 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_344
timestamp 1515882711
transform -1 0 6664 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_344
timestamp 1515882711
transform -1 0 6712 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_267
timestamp 1515882711
transform 1 0 6712 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_267
timestamp 1515882711
transform 1 0 6728 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_351
timestamp 1515882711
transform -1 0 6792 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_351
timestamp 1515882711
transform -1 0 6840 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_291
timestamp 1515882711
transform 1 0 6840 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_291
timestamp 1515882711
transform 1 0 6856 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_424
timestamp 1515882711
transform 1 0 6904 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_306
timestamp 1515882711
transform -1 0 6984 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_306
timestamp 1515882711
transform -1 0 7032 0 1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_355
timestamp 1515882711
transform -1 0 7048 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_355
timestamp 1515882711
transform -1 0 7096 0 1 1410
box 0 0 48 200
use FILL  FILL_7_6_0
timestamp 1515882711
transform 1 0 7096 0 1 1410
box 0 0 16 200
use FILL  FILL_7_6_1
timestamp 1515882711
transform 1 0 7112 0 1 1410
box 0 0 16 200
use FILL  FILL_NAND2X1_119
timestamp 1515882711
transform 1 0 7128 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_119
timestamp 1515882711
transform 1 0 7144 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_134
timestamp 1515882711
transform -1 0 7256 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_327
timestamp 1515882711
transform -1 0 7320 0 1 1410
box 0 0 64 200
use FILL  FILL_INVX1_71
timestamp 1515882711
transform -1 0 7336 0 1 1410
box 0 0 16 200
use INVX1  INVX1_71
timestamp 1515882711
transform -1 0 7368 0 1 1410
box 0 0 32 200
use FILL  FILL_NAND2X1_305
timestamp 1515882711
transform 1 0 7368 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_305
timestamp 1515882711
transform 1 0 7384 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_348
timestamp 1515882711
transform -1 0 7496 0 1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_284
timestamp 1515882711
transform 1 0 7496 0 1 1410
box 0 0 16 200
use BUFX4  BUFX4_284
timestamp 1515882711
transform 1 0 7512 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_297
timestamp 1515882711
transform -1 0 7640 0 1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_196
timestamp 1515882711
transform -1 0 7656 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_196
timestamp 1515882711
transform -1 0 7704 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_152
timestamp 1515882711
transform 1 0 7704 0 1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_152
timestamp 1515882711
transform -1 0 7784 0 1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_152
timestamp 1515882711
transform -1 0 7976 0 1 1410
box 0 0 192 200
use FILL  FILL_NAND2X1_251
timestamp 1515882711
transform -1 0 7992 0 1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_251
timestamp 1515882711
transform -1 0 8040 0 1 1410
box 0 0 48 200
use FILL  FILL_8_1
timestamp 1515882711
transform 1 0 8040 0 1 1410
box 0 0 16 200
use NOR2X1  NOR2X1_76
timestamp 1515882711
transform -1 0 56 0 -1 1410
box 0 0 48 200
use FILL  FILL_AOI21X1_64
timestamp 1515882711
transform -1 0 72 0 -1 1410
box 0 0 16 200
use AOI21X1  AOI21X1_64
timestamp 1515882711
transform -1 0 136 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_63
timestamp 1515882711
transform -1 0 200 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_64
timestamp 1515882711
transform -1 0 264 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_65
timestamp 1515882711
transform -1 0 328 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_62
timestamp 1515882711
transform 1 0 328 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_242
timestamp 1515882711
transform 1 0 392 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_240
timestamp 1515882711
transform 1 0 456 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_241
timestamp 1515882711
transform 1 0 520 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_307
timestamp 1515882711
transform 1 0 584 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_306
timestamp 1515882711
transform 1 0 648 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_163
timestamp 1515882711
transform 1 0 712 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_162
timestamp 1515882711
transform -1 0 840 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_305
timestamp 1515882711
transform -1 0 904 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_94
timestamp 1515882711
transform 1 0 904 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_0_0
timestamp 1515882711
transform -1 0 968 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1515882711
transform -1 0 984 0 -1 1410
box 0 0 16 200
use FILL  FILL_AOI21X1_18
timestamp 1515882711
transform -1 0 1000 0 -1 1410
box 0 0 16 200
use AOI21X1  AOI21X1_18
timestamp 1515882711
transform -1 0 1064 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_355
timestamp 1515882711
transform -1 0 1128 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_195
timestamp 1515882711
transform -1 0 1192 0 -1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_27
timestamp 1515882711
transform -1 0 1320 0 -1 1410
box 0 0 128 200
use NAND3X1  NAND3X1_72
timestamp 1515882711
transform 1 0 1320 0 -1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1515882711
transform -1 0 1512 0 -1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_196
timestamp 1515882711
transform 1 0 1512 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_223
timestamp 1515882711
transform 1 0 1576 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_160
timestamp 1515882711
transform -1 0 1704 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_303
timestamp 1515882711
transform 1 0 1704 0 -1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_131
timestamp 1515882711
transform 1 0 1768 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_131
timestamp 1515882711
transform 1 0 1784 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_304
timestamp 1515882711
transform -1 0 1912 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_161
timestamp 1515882711
transform 1 0 1912 0 -1 1410
box 0 0 64 200
use FILL  FILL_6_1_0
timestamp 1515882711
transform -1 0 1992 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1515882711
transform -1 0 2008 0 -1 1410
box 0 0 16 200
use FILL  FILL_BUFX4_177
timestamp 1515882711
transform -1 0 2024 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_177
timestamp 1515882711
transform -1 0 2088 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_177
timestamp 1515882711
transform 1 0 2088 0 -1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_94
timestamp 1515882711
transform 1 0 2152 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_94
timestamp 1515882711
transform 1 0 2168 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_129
timestamp 1515882711
transform -1 0 2280 0 -1 1410
box 0 0 48 200
use FILL  FILL_AOI21X1_53
timestamp 1515882711
transform -1 0 2296 0 -1 1410
box 0 0 16 200
use AOI21X1  AOI21X1_53
timestamp 1515882711
transform -1 0 2360 0 -1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_220
timestamp 1515882711
transform -1 0 2376 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_220
timestamp 1515882711
transform -1 0 2568 0 -1 1410
box 0 0 192 200
use FILL  FILL_NAND2X1_173
timestamp 1515882711
transform -1 0 2584 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_173
timestamp 1515882711
transform -1 0 2632 0 -1 1410
box 0 0 48 200
use FILL  FILL_BUFX4_143
timestamp 1515882711
transform -1 0 2648 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_143
timestamp 1515882711
transform -1 0 2712 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1515882711
transform 1 0 2712 0 -1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_25
timestamp 1515882711
transform -1 0 2792 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_25
timestamp 1515882711
transform -1 0 2856 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_28
timestamp 1515882711
transform 1 0 2856 0 -1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_6
timestamp 1515882711
transform -1 0 2936 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_6
timestamp 1515882711
transform -1 0 2984 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_2_0
timestamp 1515882711
transform 1 0 2984 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_2_1
timestamp 1515882711
transform 1 0 3000 0 -1 1410
box 0 0 16 200
use FILL  FILL_DFFPOSX1_276
timestamp 1515882711
transform 1 0 3016 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_276
timestamp 1515882711
transform 1 0 3032 0 -1 1410
box 0 0 192 200
use FILL  FILL_BUFX4_285
timestamp 1515882711
transform -1 0 3240 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_285
timestamp 1515882711
transform -1 0 3304 0 -1 1410
box 0 0 64 200
use FILL  FILL_INVX1_90
timestamp 1515882711
transform 1 0 3304 0 -1 1410
box 0 0 16 200
use INVX1  INVX1_90
timestamp 1515882711
transform 1 0 3320 0 -1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_37
timestamp 1515882711
transform -1 0 3400 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_34
timestamp 1515882711
transform 1 0 3400 0 -1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_314
timestamp 1515882711
transform 1 0 3448 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_314
timestamp 1515882711
transform 1 0 3464 0 -1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_254
timestamp 1515882711
transform -1 0 3528 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_254
timestamp 1515882711
transform -1 0 3576 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_166
timestamp 1515882711
transform -1 0 3640 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_281
timestamp 1515882711
transform -1 0 3704 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_309
timestamp 1515882711
transform -1 0 3768 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_192
timestamp 1515882711
transform -1 0 3832 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_63
timestamp 1515882711
transform -1 0 3880 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_70
timestamp 1515882711
transform -1 0 3944 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_32
timestamp 1515882711
transform 1 0 3944 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_3_0
timestamp 1515882711
transform 1 0 3992 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_3_1
timestamp 1515882711
transform 1 0 4008 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_352
timestamp 1515882711
transform 1 0 4024 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_248
timestamp 1515882711
transform -1 0 4152 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_66
timestamp 1515882711
transform 1 0 4152 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_39
timestamp 1515882711
transform 1 0 4216 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_113
timestamp 1515882711
transform -1 0 4328 0 -1 1410
box 0 0 64 200
use BUFX2  BUFX2_45
timestamp 1515882711
transform -1 0 4376 0 -1 1410
box 0 0 48 200
use FILL  FILL_NAND2X1_345
timestamp 1515882711
transform -1 0 4392 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_345
timestamp 1515882711
transform -1 0 4440 0 -1 1410
box 0 0 48 200
use NAND3X1  NAND3X1_12
timestamp 1515882711
transform 1 0 4440 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_189
timestamp 1515882711
transform 1 0 4504 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_91
timestamp 1515882711
transform -1 0 4632 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_351
timestamp 1515882711
transform -1 0 4696 0 -1 1410
box 0 0 64 200
use FILL  FILL_INVX1_84
timestamp 1515882711
transform -1 0 4712 0 -1 1410
box 0 0 16 200
use INVX1  INVX1_84
timestamp 1515882711
transform -1 0 4744 0 -1 1410
box 0 0 32 200
use FILL  FILL_NAND2X1_30
timestamp 1515882711
transform 1 0 4744 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_30
timestamp 1515882711
transform 1 0 4760 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_51
timestamp 1515882711
transform -1 0 4872 0 -1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_51
timestamp 1515882711
transform -1 0 4888 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_51
timestamp 1515882711
transform -1 0 5080 0 -1 1410
box 0 0 192 200
use FILL  FILL_6_4_0
timestamp 1515882711
transform -1 0 5096 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_4_1
timestamp 1515882711
transform -1 0 5112 0 -1 1410
box 0 0 16 200
use FILL  FILL_BUFX4_24
timestamp 1515882711
transform -1 0 5128 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_24
timestamp 1515882711
transform -1 0 5192 0 -1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_18
timestamp 1515882711
transform 1 0 5192 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_18
timestamp 1515882711
transform 1 0 5208 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_112
timestamp 1515882711
transform 1 0 5400 0 -1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_334
timestamp 1515882711
transform -1 0 5480 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_334
timestamp 1515882711
transform -1 0 5528 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_303
timestamp 1515882711
transform -1 0 5592 0 -1 1410
box 0 0 64 200
use FILL  FILL_INVX1_58
timestamp 1515882711
transform -1 0 5608 0 -1 1410
box 0 0 16 200
use INVX1  INVX1_58
timestamp 1515882711
transform -1 0 5640 0 -1 1410
box 0 0 32 200
use FILL  FILL_NAND2X1_202
timestamp 1515882711
transform -1 0 5656 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_202
timestamp 1515882711
transform -1 0 5704 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_214
timestamp 1515882711
transform -1 0 5768 0 -1 1410
box 0 0 64 200
use FILL  FILL_INVX1_9
timestamp 1515882711
transform -1 0 5784 0 -1 1410
box 0 0 16 200
use INVX1  INVX1_9
timestamp 1515882711
transform -1 0 5816 0 -1 1410
box 0 0 32 200
use FILL  FILL_BUFX4_26
timestamp 1515882711
transform -1 0 5832 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_26
timestamp 1515882711
transform -1 0 5896 0 -1 1410
box 0 0 64 200
use FILL  FILL_BUFX4_162
timestamp 1515882711
transform 1 0 5896 0 -1 1410
box 0 0 16 200
use BUFX4  BUFX4_162
timestamp 1515882711
transform 1 0 5912 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_62
timestamp 1515882711
transform -1 0 6024 0 -1 1410
box 0 0 48 200
use FILL  FILL_DFFPOSX1_53
timestamp 1515882711
transform -1 0 6040 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_5_0
timestamp 1515882711
transform -1 0 6056 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_5_1
timestamp 1515882711
transform -1 0 6072 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_53
timestamp 1515882711
transform -1 0 6264 0 -1 1410
box 0 0 192 200
use NOR2X1  NOR2X1_31
timestamp 1515882711
transform 1 0 6264 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_30
timestamp 1515882711
transform -1 0 6360 0 -1 1410
box 0 0 48 200
use NOR3X1  NOR3X1_26
timestamp 1515882711
transform 1 0 6360 0 -1 1410
box 0 0 128 200
use OAI21X1  OAI21X1_122
timestamp 1515882711
transform 1 0 6488 0 -1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_122
timestamp 1515882711
transform 1 0 6552 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_122
timestamp 1515882711
transform 1 0 6568 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_298
timestamp 1515882711
transform -1 0 6824 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_415
timestamp 1515882711
transform -1 0 6888 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_328
timestamp 1515882711
transform -1 0 6952 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_349
timestamp 1515882711
transform 1 0 6952 0 -1 1410
box 0 0 64 200
use FILL  FILL_DFFPOSX1_134
timestamp 1515882711
transform -1 0 7032 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_6_0
timestamp 1515882711
transform -1 0 7048 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_6_1
timestamp 1515882711
transform -1 0 7064 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_134
timestamp 1515882711
transform -1 0 7256 0 -1 1410
box 0 0 192 200
use FILL  FILL_MUX2X1_43
timestamp 1515882711
transform 1 0 7256 0 -1 1410
box 0 0 16 200
use MUX2X1  MUX2X1_43
timestamp 1515882711
transform 1 0 7272 0 -1 1410
box 0 0 96 200
use FILL  FILL_DFFPOSX1_155
timestamp 1515882711
transform -1 0 7384 0 -1 1410
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_155
timestamp 1515882711
transform -1 0 7576 0 -1 1410
box 0 0 192 200
use OAI21X1  OAI21X1_155
timestamp 1515882711
transform 1 0 7576 0 -1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_141
timestamp 1515882711
transform 1 0 7640 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_141
timestamp 1515882711
transform 1 0 7656 0 -1 1410
box 0 0 48 200
use FILL  FILL_INVX1_54
timestamp 1515882711
transform -1 0 7720 0 -1 1410
box 0 0 16 200
use INVX1  INVX1_54
timestamp 1515882711
transform -1 0 7752 0 -1 1410
box 0 0 32 200
use FILL  FILL_NAND2X1_138
timestamp 1515882711
transform -1 0 7768 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_138
timestamp 1515882711
transform -1 0 7816 0 -1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_158
timestamp 1515882711
transform 1 0 7816 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_485
timestamp 1515882711
transform 1 0 7880 0 -1 1410
box 0 0 64 200
use FILL  FILL_NAND2X1_143
timestamp 1515882711
transform -1 0 7960 0 -1 1410
box 0 0 16 200
use NAND2X1  NAND2X1_143
timestamp 1515882711
transform -1 0 8008 0 -1 1410
box 0 0 48 200
use FILL  FILL_7_1
timestamp 1515882711
transform -1 0 8024 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_2
timestamp 1515882711
transform -1 0 8040 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_3
timestamp 1515882711
transform -1 0 8056 0 -1 1410
box 0 0 16 200
use NAND3X1  NAND3X1_278
timestamp 1515882711
transform -1 0 72 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_267
timestamp 1515882711
transform -1 0 136 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_289
timestamp 1515882711
transform -1 0 200 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_74
timestamp 1515882711
transform 1 0 200 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_75
timestamp 1515882711
transform 1 0 264 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_76
timestamp 1515882711
transform -1 0 392 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_243
timestamp 1515882711
transform -1 0 456 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_164
timestamp 1515882711
transform -1 0 520 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_165
timestamp 1515882711
transform -1 0 584 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_308
timestamp 1515882711
transform -1 0 648 0 1 1010
box 0 0 64 200
use FILL  FILL_AOI21X1_27
timestamp 1515882711
transform 1 0 648 0 1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_27
timestamp 1515882711
transform 1 0 664 0 1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_167
timestamp 1515882711
transform -1 0 744 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_167
timestamp 1515882711
transform -1 0 808 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_103
timestamp 1515882711
transform 1 0 808 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_71
timestamp 1515882711
transform -1 0 920 0 1 1010
box 0 0 64 200
use FILL  FILL_5_0_0
timestamp 1515882711
transform 1 0 920 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1515882711
transform 1 0 936 0 1 1010
box 0 0 16 200
use NAND3X1  NAND3X1_112
timestamp 1515882711
transform 1 0 952 0 1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_130
timestamp 1515882711
transform -1 0 1032 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_130
timestamp 1515882711
transform -1 0 1096 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_36
timestamp 1515882711
transform -1 0 1224 0 1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_391
timestamp 1515882711
transform 1 0 1224 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_356
timestamp 1515882711
transform 1 0 1288 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_9
timestamp 1515882711
transform -1 0 1480 0 1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_275
timestamp 1515882711
transform 1 0 1480 0 1 1010
box 0 0 64 200
use FILL  FILL_AOI21X1_36
timestamp 1515882711
transform 1 0 1544 0 1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_36
timestamp 1515882711
transform 1 0 1560 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_112
timestamp 1515882711
transform -1 0 1672 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_276
timestamp 1515882711
transform 1 0 1672 0 1 1010
box 0 0 64 200
use FILL  FILL_INVX2_19
timestamp 1515882711
transform -1 0 1752 0 1 1010
box 0 0 16 200
use INVX2  INVX2_19
timestamp 1515882711
transform -1 0 1784 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_392
timestamp 1515882711
transform 1 0 1784 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_186
timestamp 1515882711
transform 1 0 1848 0 1 1010
box 0 0 64 200
use FILL  FILL_INVX2_10
timestamp 1515882711
transform -1 0 1928 0 1 1010
box 0 0 16 200
use INVX2  INVX2_10
timestamp 1515882711
transform -1 0 1960 0 1 1010
box 0 0 32 200
use FILL  FILL_5_1_0
timestamp 1515882711
transform -1 0 1976 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1515882711
transform -1 0 1992 0 1 1010
box 0 0 16 200
use FILL  FILL_DFFPOSX1_230
timestamp 1515882711
transform -1 0 2008 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_230
timestamp 1515882711
transform -1 0 2200 0 1 1010
box 0 0 192 200
use FILL  FILL_INVX2_2
timestamp 1515882711
transform 1 0 2200 0 1 1010
box 0 0 16 200
use INVX2  INVX2_2
timestamp 1515882711
transform 1 0 2216 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_169
timestamp 1515882711
transform 1 0 2248 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_171
timestamp 1515882711
transform -1 0 2328 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_171
timestamp 1515882711
transform -1 0 2376 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_153
timestamp 1515882711
transform -1 0 2392 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_153
timestamp 1515882711
transform -1 0 2440 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_155
timestamp 1515882711
transform -1 0 2456 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_155
timestamp 1515882711
transform -1 0 2504 0 1 1010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_274
timestamp 1515882711
transform 1 0 2504 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_274
timestamp 1515882711
transform 1 0 2520 0 1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_4
timestamp 1515882711
transform 1 0 2712 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_4
timestamp 1515882711
transform 1 0 2728 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_280
timestamp 1515882711
transform 1 0 2776 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_299
timestamp 1515882711
transform -1 0 2904 0 1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_340
timestamp 1515882711
transform 1 0 2904 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_0
timestamp 1515882711
transform 1 0 2920 0 1 1010
box 0 0 16 200
use FILL  FILL_5_2_1
timestamp 1515882711
transform 1 0 2936 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_340
timestamp 1515882711
transform 1 0 2952 0 1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_247
timestamp 1515882711
transform 1 0 3144 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_247
timestamp 1515882711
transform 1 0 3160 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_271
timestamp 1515882711
transform -1 0 3272 0 1 1010
box 0 0 64 200
use FILL  FILL_INVX1_40
timestamp 1515882711
transform -1 0 3288 0 1 1010
box 0 0 16 200
use INVX1  INVX1_40
timestamp 1515882711
transform -1 0 3320 0 1 1010
box 0 0 32 200
use FILL  FILL_NAND2X1_366
timestamp 1515882711
transform 1 0 3320 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_366
timestamp 1515882711
transform 1 0 3336 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_433
timestamp 1515882711
transform -1 0 3448 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_21
timestamp 1515882711
transform 1 0 3448 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_21
timestamp 1515882711
transform 1 0 3464 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_42
timestamp 1515882711
transform -1 0 3576 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_394
timestamp 1515882711
transform 1 0 3576 0 1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_102
timestamp 1515882711
transform -1 0 3656 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_102
timestamp 1515882711
transform -1 0 3720 0 1 1010
box 0 0 64 200
use FILL  FILL_INVX1_46
timestamp 1515882711
transform -1 0 3736 0 1 1010
box 0 0 16 200
use INVX1  INVX1_46
timestamp 1515882711
transform -1 0 3768 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_282
timestamp 1515882711
transform -1 0 3832 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_403
timestamp 1515882711
transform 1 0 3832 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_9
timestamp 1515882711
transform -1 0 3944 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_188
timestamp 1515882711
transform -1 0 4008 0 1 1010
box 0 0 64 200
use FILL  FILL_5_3_0
timestamp 1515882711
transform 1 0 4008 0 1 1010
box 0 0 16 200
use FILL  FILL_5_3_1
timestamp 1515882711
transform 1 0 4024 0 1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_302
timestamp 1515882711
transform 1 0 4040 0 1 1010
box 0 0 64 200
use FILL  FILL_BUFX2_8
timestamp 1515882711
transform 1 0 4104 0 1 1010
box 0 0 16 200
use BUFX2  BUFX2_8
timestamp 1515882711
transform 1 0 4120 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_11
timestamp 1515882711
transform 1 0 4168 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_15
timestamp 1515882711
transform -1 0 4296 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_16
timestamp 1515882711
transform -1 0 4344 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_203
timestamp 1515882711
transform -1 0 4360 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_203
timestamp 1515882711
transform -1 0 4408 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_101
timestamp 1515882711
transform 1 0 4408 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_273
timestamp 1515882711
transform 1 0 4472 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_273
timestamp 1515882711
transform 1 0 4488 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_14
timestamp 1515882711
transform 1 0 4536 0 1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_191
timestamp 1515882711
transform 1 0 4600 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_325
timestamp 1515882711
transform -1 0 4680 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_325
timestamp 1515882711
transform -1 0 4728 0 1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_89
timestamp 1515882711
transform 1 0 4728 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_308
timestamp 1515882711
transform -1 0 4808 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_308
timestamp 1515882711
transform -1 0 4856 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_375
timestamp 1515882711
transform 1 0 4856 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_375
timestamp 1515882711
transform 1 0 4872 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_442
timestamp 1515882711
transform -1 0 4984 0 1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_100
timestamp 1515882711
transform -1 0 5000 0 1 1010
box 0 0 16 200
use FILL  FILL_5_4_0
timestamp 1515882711
transform -1 0 5016 0 1 1010
box 0 0 16 200
use FILL  FILL_5_4_1
timestamp 1515882711
transform -1 0 5032 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_100
timestamp 1515882711
transform -1 0 5096 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_124
timestamp 1515882711
transform 1 0 5096 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_124
timestamp 1515882711
transform 1 0 5112 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_90
timestamp 1515882711
transform -1 0 5224 0 1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_90
timestamp 1515882711
transform -1 0 5240 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_90
timestamp 1515882711
transform -1 0 5432 0 1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_201
timestamp 1515882711
transform 1 0 5432 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_201
timestamp 1515882711
transform 1 0 5448 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_168
timestamp 1515882711
transform -1 0 5560 0 1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_168
timestamp 1515882711
transform -1 0 5576 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_168
timestamp 1515882711
transform -1 0 5768 0 1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_60
timestamp 1515882711
transform 1 0 5768 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_60
timestamp 1515882711
transform 1 0 5784 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_78
timestamp 1515882711
transform -1 0 5896 0 1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_164
timestamp 1515882711
transform 1 0 5896 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_164
timestamp 1515882711
transform 1 0 5912 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_14
timestamp 1515882711
transform 1 0 5976 0 1 1010
box 0 0 48 200
use FILL  FILL_5_5_0
timestamp 1515882711
transform 1 0 6024 0 1 1010
box 0 0 16 200
use FILL  FILL_5_5_1
timestamp 1515882711
transform 1 0 6040 0 1 1010
box 0 0 16 200
use NOR3X1  NOR3X1_15
timestamp 1515882711
transform 1 0 6056 0 1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_15
timestamp 1515882711
transform 1 0 6184 0 1 1010
box 0 0 48 200
use NOR3X1  NOR3X1_21
timestamp 1515882711
transform 1 0 6232 0 1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_25
timestamp 1515882711
transform -1 0 6408 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_8
timestamp 1515882711
transform -1 0 6456 0 1 1010
box 0 0 48 200
use FILL  FILL_BUFX4_111
timestamp 1515882711
transform 1 0 6456 0 1 1010
box 0 0 16 200
use BUFX4  BUFX4_111
timestamp 1515882711
transform 1 0 6472 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_88
timestamp 1515882711
transform 1 0 6536 0 1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_71
timestamp 1515882711
transform -1 0 6616 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_71
timestamp 1515882711
transform -1 0 6664 0 1 1010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_88
timestamp 1515882711
transform 1 0 6664 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_88
timestamp 1515882711
transform 1 0 6680 0 1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_340
timestamp 1515882711
transform -1 0 6888 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_340
timestamp 1515882711
transform -1 0 6936 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_252
timestamp 1515882711
transform -1 0 6952 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_252
timestamp 1515882711
transform -1 0 7000 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_197
timestamp 1515882711
transform -1 0 7016 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_197
timestamp 1515882711
transform -1 0 7064 0 1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_324
timestamp 1515882711
transform -1 0 7080 0 1 1010
box 0 0 16 200
use FILL  FILL_5_6_0
timestamp 1515882711
transform -1 0 7096 0 1 1010
box 0 0 16 200
use FILL  FILL_5_6_1
timestamp 1515882711
transform -1 0 7112 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_324
timestamp 1515882711
transform -1 0 7160 0 1 1010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_140
timestamp 1515882711
transform -1 0 7176 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_140
timestamp 1515882711
transform -1 0 7368 0 1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_125
timestamp 1515882711
transform 1 0 7368 0 1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_125
timestamp 1515882711
transform 1 0 7384 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_140
timestamp 1515882711
transform -1 0 7496 0 1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_314
timestamp 1515882711
transform -1 0 7512 0 1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_314
timestamp 1515882711
transform -1 0 7704 0 1 1010
box 0 0 192 200
use NAND2X1  NAND2X1_440
timestamp 1515882711
transform 1 0 7704 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_493
timestamp 1515882711
transform -1 0 7816 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_155
timestamp 1515882711
transform 1 0 7816 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_207
timestamp 1515882711
transform -1 0 7928 0 1 1010
box 0 0 64 200
use FILL  FILL_INVX1_43
timestamp 1515882711
transform 1 0 7928 0 1 1010
box 0 0 16 200
use INVX1  INVX1_43
timestamp 1515882711
transform 1 0 7944 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_277
timestamp 1515882711
transform 1 0 7976 0 1 1010
box 0 0 64 200
use FILL  FILL_6_1
timestamp 1515882711
transform 1 0 8040 0 1 1010
box 0 0 16 200
use FILL  FILL_DFFPOSX1_248
timestamp 1515882711
transform -1 0 24 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_248
timestamp 1515882711
transform -1 0 216 0 -1 1010
box 0 0 192 200
use NAND3X1  NAND3X1_256
timestamp 1515882711
transform 1 0 216 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_2
timestamp 1515882711
transform 1 0 280 0 -1 1010
box 0 0 48 200
use FILL  FILL_AOI21X1_1
timestamp 1515882711
transform -1 0 344 0 -1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_1
timestamp 1515882711
transform -1 0 408 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_73
timestamp 1515882711
transform 1 0 408 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_214
timestamp 1515882711
transform -1 0 488 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_214
timestamp 1515882711
transform -1 0 552 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_150
timestamp 1515882711
transform -1 0 568 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_150
timestamp 1515882711
transform -1 0 632 0 -1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_194
timestamp 1515882711
transform 1 0 632 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_194
timestamp 1515882711
transform 1 0 648 0 -1 1010
box 0 0 192 200
use FILL  FILL_BUFX4_95
timestamp 1515882711
transform -1 0 856 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_95
timestamp 1515882711
transform -1 0 920 0 -1 1010
box 0 0 64 200
use FILL  FILL_4_0_0
timestamp 1515882711
transform -1 0 936 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1515882711
transform -1 0 952 0 -1 1010
box 0 0 16 200
use NAND3X1  NAND3X1_238
timestamp 1515882711
transform -1 0 1016 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_60
timestamp 1515882711
transform 1 0 1016 0 -1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_43
timestamp 1515882711
transform -1 0 1208 0 -1 1010
box 0 0 128 200
use OAI21X1  OAI21X1_421
timestamp 1515882711
transform -1 0 1272 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_422
timestamp 1515882711
transform -1 0 1336 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_345
timestamp 1515882711
transform -1 0 1400 0 -1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_25
timestamp 1515882711
transform 1 0 1400 0 -1 1010
box 0 0 128 200
use FILL  FILL_DFFPOSX1_203
timestamp 1515882711
transform 1 0 1528 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_203
timestamp 1515882711
transform 1 0 1544 0 -1 1010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_239
timestamp 1515882711
transform -1 0 1752 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_239
timestamp 1515882711
transform -1 0 1944 0 -1 1010
box 0 0 192 200
use FILL  FILL_BUFX4_140
timestamp 1515882711
transform -1 0 1960 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_0
timestamp 1515882711
transform -1 0 1976 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1515882711
transform -1 0 1992 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_140
timestamp 1515882711
transform -1 0 2056 0 -1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_185
timestamp 1515882711
transform 1 0 2056 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_185
timestamp 1515882711
transform 1 0 2072 0 -1 1010
box 0 0 192 200
use FILL  FILL_BUFX4_316
timestamp 1515882711
transform -1 0 2280 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_316
timestamp 1515882711
transform -1 0 2344 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_33
timestamp 1515882711
transform -1 0 2392 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_38
timestamp 1515882711
transform 1 0 2392 0 -1 1010
box 0 0 48 200
use FILL  FILL_INVX1_87
timestamp 1515882711
transform 1 0 2440 0 -1 1010
box 0 0 16 200
use INVX1  INVX1_87
timestamp 1515882711
transform 1 0 2456 0 -1 1010
box 0 0 32 200
use FILL  FILL_AND2X2_8
timestamp 1515882711
transform 1 0 2488 0 -1 1010
box 0 0 16 200
use AND2X2  AND2X2_8
timestamp 1515882711
transform 1 0 2504 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_105
timestamp 1515882711
transform -1 0 2584 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_105
timestamp 1515882711
transform -1 0 2648 0 -1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_316
timestamp 1515882711
transform 1 0 2648 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_316
timestamp 1515882711
transform 1 0 2664 0 -1 1010
box 0 0 48 200
use FILL  FILL_BUFX4_3
timestamp 1515882711
transform -1 0 2728 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_3
timestamp 1515882711
transform -1 0 2792 0 -1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_269
timestamp 1515882711
transform -1 0 2808 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_269
timestamp 1515882711
transform -1 0 2856 0 -1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_253
timestamp 1515882711
transform 1 0 2856 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_253
timestamp 1515882711
transform 1 0 2872 0 -1 1010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_341
timestamp 1515882711
transform 1 0 2920 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_0
timestamp 1515882711
transform 1 0 2936 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_2_1
timestamp 1515882711
transform 1 0 2952 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_341
timestamp 1515882711
transform 1 0 2968 0 -1 1010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_42
timestamp 1515882711
transform 1 0 3160 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_42
timestamp 1515882711
transform 1 0 3176 0 -1 1010
box 0 0 192 200
use FILL  FILL_NAND2X1_367
timestamp 1515882711
transform 1 0 3368 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_367
timestamp 1515882711
transform 1 0 3384 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_435
timestamp 1515882711
transform -1 0 3496 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_221
timestamp 1515882711
transform -1 0 3560 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_170
timestamp 1515882711
transform -1 0 3624 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_59
timestamp 1515882711
transform -1 0 3672 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_44
timestamp 1515882711
transform 1 0 3672 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_88
timestamp 1515882711
transform 1 0 3736 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_90
timestamp 1515882711
transform 1 0 3800 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_313
timestamp 1515882711
transform -1 0 3928 0 -1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_258
timestamp 1515882711
transform -1 0 3944 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_258
timestamp 1515882711
transform -1 0 3992 0 -1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_341
timestamp 1515882711
transform -1 0 4008 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_0
timestamp 1515882711
transform -1 0 4024 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_3_1
timestamp 1515882711
transform -1 0 4040 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_341
timestamp 1515882711
transform -1 0 4088 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_167
timestamp 1515882711
transform 1 0 4088 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_310
timestamp 1515882711
transform 1 0 4152 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_150
timestamp 1515882711
transform -1 0 4264 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_45
timestamp 1515882711
transform 1 0 4264 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_222
timestamp 1515882711
transform 1 0 4328 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_43
timestamp 1515882711
transform -1 0 4440 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_92
timestamp 1515882711
transform -1 0 4504 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_163
timestamp 1515882711
transform 1 0 4504 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_163
timestamp 1515882711
transform 1 0 4520 0 -1 1010
box 0 0 64 200
use FILL  FILL_DFFPOSX1_349
timestamp 1515882711
transform -1 0 4600 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_349
timestamp 1515882711
transform -1 0 4792 0 -1 1010
box 0 0 192 200
use FILL  FILL_BUFX4_290
timestamp 1515882711
transform -1 0 4808 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_290
timestamp 1515882711
transform -1 0 4872 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_268
timestamp 1515882711
transform 1 0 4872 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_268
timestamp 1515882711
transform 1 0 4888 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_213
timestamp 1515882711
transform -1 0 5016 0 -1 1010
box 0 0 64 200
use FILL  FILL_INVX1_8
timestamp 1515882711
transform -1 0 5032 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_4_0
timestamp 1515882711
transform -1 0 5048 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_4_1
timestamp 1515882711
transform -1 0 5064 0 -1 1010
box 0 0 16 200
use INVX1  INVX1_8
timestamp 1515882711
transform -1 0 5096 0 -1 1010
box 0 0 32 200
use FILL  FILL_NAND2X1_200
timestamp 1515882711
transform -1 0 5112 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_200
timestamp 1515882711
transform -1 0 5160 0 -1 1010
box 0 0 48 200
use FILL  FILL_BUFX4_288
timestamp 1515882711
transform 1 0 5160 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_288
timestamp 1515882711
transform 1 0 5176 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_283
timestamp 1515882711
transform -1 0 5304 0 -1 1010
box 0 0 64 200
use FILL  FILL_INVX1_47
timestamp 1515882711
transform -1 0 5320 0 -1 1010
box 0 0 16 200
use INVX1  INVX1_47
timestamp 1515882711
transform -1 0 5352 0 -1 1010
box 0 0 32 200
use FILL  FILL_NAND2X1_255
timestamp 1515882711
transform 1 0 5352 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_255
timestamp 1515882711
transform 1 0 5368 0 -1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_271
timestamp 1515882711
transform 1 0 5416 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_271
timestamp 1515882711
transform 1 0 5432 0 -1 1010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_78
timestamp 1515882711
transform -1 0 5496 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_78
timestamp 1515882711
transform -1 0 5688 0 -1 1010
box 0 0 192 200
use FILL  FILL_BUFX4_104
timestamp 1515882711
transform 1 0 5688 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_104
timestamp 1515882711
transform 1 0 5704 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_286
timestamp 1515882711
transform 1 0 5768 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_286
timestamp 1515882711
transform 1 0 5784 0 -1 1010
box 0 0 64 200
use FILL  FILL_BUFX4_85
timestamp 1515882711
transform 1 0 5848 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_85
timestamp 1515882711
transform 1 0 5864 0 -1 1010
box 0 0 64 200
use OAI22X1  OAI22X1_3
timestamp 1515882711
transform -1 0 6008 0 -1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_23
timestamp 1515882711
transform -1 0 6056 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_5_0
timestamp 1515882711
transform -1 0 6072 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_5_1
timestamp 1515882711
transform -1 0 6088 0 -1 1010
box 0 0 16 200
use OAI22X1  OAI22X1_6
timestamp 1515882711
transform -1 0 6168 0 -1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_69
timestamp 1515882711
transform -1 0 6216 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_42
timestamp 1515882711
transform 1 0 6216 0 -1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_9
timestamp 1515882711
transform -1 0 6344 0 -1 1010
box 0 0 80 200
use NOR3X1  NOR3X1_10
timestamp 1515882711
transform -1 0 6472 0 -1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_7
timestamp 1515882711
transform -1 0 6520 0 -1 1010
box 0 0 48 200
use OAI22X1  OAI22X1_16
timestamp 1515882711
transform -1 0 6600 0 -1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_58
timestamp 1515882711
transform -1 0 6648 0 -1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_149
timestamp 1515882711
transform -1 0 6696 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_393
timestamp 1515882711
transform 1 0 6696 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_278
timestamp 1515882711
transform 1 0 6760 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_362
timestamp 1515882711
transform 1 0 6824 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_208
timestamp 1515882711
transform 1 0 6888 0 -1 1010
box 0 0 64 200
use FILL  FILL_MUX2X1_45
timestamp 1515882711
transform -1 0 6968 0 -1 1010
box 0 0 16 200
use MUX2X1  MUX2X1_45
timestamp 1515882711
transform -1 0 7064 0 -1 1010
box 0 0 96 200
use FILL  FILL_4_6_0
timestamp 1515882711
transform 1 0 7064 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_6_1
timestamp 1515882711
transform 1 0 7080 0 -1 1010
box 0 0 16 200
use OAI21X1  OAI21X1_132
timestamp 1515882711
transform 1 0 7096 0 -1 1010
box 0 0 64 200
use FILL  FILL_NAND2X1_117
timestamp 1515882711
transform -1 0 7176 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_117
timestamp 1515882711
transform -1 0 7224 0 -1 1010
box 0 0 48 200
use FILL  FILL_NAND2X1_108
timestamp 1515882711
transform -1 0 7240 0 -1 1010
box 0 0 16 200
use NAND2X1  NAND2X1_108
timestamp 1515882711
transform -1 0 7288 0 -1 1010
box 0 0 48 200
use FILL  FILL_DFFPOSX1_125
timestamp 1515882711
transform -1 0 7304 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_125
timestamp 1515882711
transform -1 0 7496 0 -1 1010
box 0 0 192 200
use FILL  FILL_BUFX4_306
timestamp 1515882711
transform 1 0 7496 0 -1 1010
box 0 0 16 200
use BUFX4  BUFX4_306
timestamp 1515882711
transform 1 0 7512 0 -1 1010
box 0 0 64 200
use FILL  FILL_INVX1_82
timestamp 1515882711
transform -1 0 7592 0 -1 1010
box 0 0 16 200
use INVX1  INVX1_82
timestamp 1515882711
transform -1 0 7624 0 -1 1010
box 0 0 32 200
use FILL  FILL_DFFPOSX1_150
timestamp 1515882711
transform 1 0 7624 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_150
timestamp 1515882711
transform 1 0 7640 0 -1 1010
box 0 0 192 200
use FILL  FILL_DFFPOSX1_158
timestamp 1515882711
transform 1 0 7832 0 -1 1010
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_158
timestamp 1515882711
transform 1 0 7848 0 -1 1010
box 0 0 192 200
use FILL  FILL_5_1
timestamp 1515882711
transform -1 0 8056 0 -1 1010
box 0 0 16 200
use FILL  FILL_DFFPOSX1_159
timestamp 1515882711
transform 1 0 8 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_159
timestamp 1515882711
transform 1 0 24 0 1 610
box 0 0 192 200
use NOR2X1  NOR2X1_85
timestamp 1515882711
transform 1 0 216 0 1 610
box 0 0 48 200
use FILL  FILL_AOI21X1_9
timestamp 1515882711
transform -1 0 280 0 1 610
box 0 0 16 200
use AOI21X1  AOI21X1_9
timestamp 1515882711
transform -1 0 344 0 1 610
box 0 0 64 200
use FILL  FILL_AOI21X1_24
timestamp 1515882711
transform 1 0 344 0 1 610
box 0 0 16 200
use AOI21X1  AOI21X1_24
timestamp 1515882711
transform 1 0 360 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_99
timestamp 1515882711
transform -1 0 472 0 1 610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_173
timestamp 1515882711
transform -1 0 488 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_173
timestamp 1515882711
transform -1 0 680 0 1 610
box 0 0 192 200
use FILL  FILL_AOI21X1_43
timestamp 1515882711
transform 1 0 680 0 1 610
box 0 0 16 200
use AOI21X1  AOI21X1_43
timestamp 1515882711
transform 1 0 696 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_119
timestamp 1515882711
transform -1 0 808 0 1 610
box 0 0 48 200
use FILL  FILL_AOI21X1_41
timestamp 1515882711
transform 1 0 808 0 1 610
box 0 0 16 200
use AOI21X1  AOI21X1_41
timestamp 1515882711
transform 1 0 824 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_117
timestamp 1515882711
transform -1 0 936 0 1 610
box 0 0 48 200
use FILL  FILL_3_0_0
timestamp 1515882711
transform -1 0 952 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1515882711
transform -1 0 968 0 1 610
box 0 0 16 200
use NAND3X1  NAND3X1_38
timestamp 1515882711
transform -1 0 1032 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_215
timestamp 1515882711
transform -1 0 1096 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_325
timestamp 1515882711
transform -1 0 1160 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_413
timestamp 1515882711
transform -1 0 1224 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_239
timestamp 1515882711
transform -1 0 1288 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_61
timestamp 1515882711
transform 1 0 1288 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_347
timestamp 1515882711
transform -1 0 1416 0 1 610
box 0 0 64 200
use FILL  FILL_BUFX4_4
timestamp 1515882711
transform -1 0 1432 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_4
timestamp 1515882711
transform -1 0 1496 0 1 610
box 0 0 64 200
use FILL  FILL_BUFX4_292
timestamp 1515882711
transform -1 0 1512 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_292
timestamp 1515882711
transform -1 0 1576 0 1 610
box 0 0 64 200
use FILL  FILL_INVX2_7
timestamp 1515882711
transform -1 0 1592 0 1 610
box 0 0 16 200
use INVX2  INVX2_7
timestamp 1515882711
transform -1 0 1624 0 1 610
box 0 0 32 200
use FILL  FILL_DFFPOSX1_191
timestamp 1515882711
transform -1 0 1640 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_191
timestamp 1515882711
transform -1 0 1832 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_174
timestamp 1515882711
transform 1 0 1832 0 1 610
box 0 0 64 200
use FILL  FILL_INVX2_4
timestamp 1515882711
transform -1 0 1912 0 1 610
box 0 0 16 200
use INVX2  INVX2_4
timestamp 1515882711
transform -1 0 1944 0 1 610
box 0 0 32 200
use FILL  FILL_DFFPOSX1_187
timestamp 1515882711
transform -1 0 1960 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_0
timestamp 1515882711
transform -1 0 1976 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1515882711
transform -1 0 1992 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_187
timestamp 1515882711
transform -1 0 2184 0 1 610
box 0 0 192 200
use OAI21X1  OAI21X1_171
timestamp 1515882711
transform 1 0 2184 0 1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_10
timestamp 1515882711
transform 1 0 2248 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_10
timestamp 1515882711
transform 1 0 2264 0 1 610
box 0 0 192 200
use FILL  FILL_INVX1_55
timestamp 1515882711
transform 1 0 2456 0 1 610
box 0 0 16 200
use INVX1  INVX1_55
timestamp 1515882711
transform 1 0 2472 0 1 610
box 0 0 32 200
use FILL  FILL_INVX8_18
timestamp 1515882711
transform -1 0 2520 0 1 610
box 0 0 16 200
use INVX8  INVX8_18
timestamp 1515882711
transform -1 0 2600 0 1 610
box 0 0 80 200
use OAI21X1  OAI21X1_455
timestamp 1515882711
transform 1 0 2600 0 1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_266
timestamp 1515882711
transform 1 0 2664 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_266
timestamp 1515882711
transform 1 0 2680 0 1 610
box 0 0 192 200
use FILL  FILL_INVX1_44
timestamp 1515882711
transform 1 0 2872 0 1 610
box 0 0 16 200
use INVX1  INVX1_44
timestamp 1515882711
transform 1 0 2888 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_209
timestamp 1515882711
transform 1 0 2920 0 1 610
box 0 0 64 200
use FILL  FILL_3_2_0
timestamp 1515882711
transform 1 0 2984 0 1 610
box 0 0 16 200
use FILL  FILL_3_2_1
timestamp 1515882711
transform 1 0 3000 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_447
timestamp 1515882711
transform 1 0 3016 0 1 610
box 0 0 48 200
use FILL  FILL_NAND2X1_373
timestamp 1515882711
transform 1 0 3064 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_373
timestamp 1515882711
transform 1 0 3080 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_440
timestamp 1515882711
transform -1 0 3192 0 1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_347
timestamp 1515882711
transform 1 0 3192 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_347
timestamp 1515882711
transform 1 0 3208 0 1 610
box 0 0 192 200
use FILL  FILL_NAND2X1_293
timestamp 1515882711
transform -1 0 3416 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_293
timestamp 1515882711
transform -1 0 3464 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_330
timestamp 1515882711
transform -1 0 3528 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_416
timestamp 1515882711
transform -1 0 3592 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_331
timestamp 1515882711
transform 1 0 3592 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_70
timestamp 1515882711
transform -1 0 3704 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_363
timestamp 1515882711
transform 1 0 3704 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_211
timestamp 1515882711
transform 1 0 3768 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_26
timestamp 1515882711
transform -1 0 3880 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_312
timestamp 1515882711
transform -1 0 3944 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_169
timestamp 1515882711
transform -1 0 4008 0 1 610
box 0 0 64 200
use FILL  FILL_3_3_0
timestamp 1515882711
transform -1 0 4024 0 1 610
box 0 0 16 200
use FILL  FILL_3_3_1
timestamp 1515882711
transform -1 0 4040 0 1 610
box 0 0 16 200
use FILL  FILL_NAND2X1_296
timestamp 1515882711
transform -1 0 4056 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_296
timestamp 1515882711
transform -1 0 4104 0 1 610
box 0 0 48 200
use NAND3X1  NAND3X1_47
timestamp 1515882711
transform 1 0 4104 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_225
timestamp 1515882711
transform -1 0 4232 0 1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_352
timestamp 1515882711
transform -1 0 4248 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_352
timestamp 1515882711
transform -1 0 4296 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_210
timestamp 1515882711
transform -1 0 4360 0 1 610
box 0 0 64 200
use FILL  FILL_INVX1_7
timestamp 1515882711
transform -1 0 4376 0 1 610
box 0 0 16 200
use INVX1  INVX1_7
timestamp 1515882711
transform -1 0 4408 0 1 610
box 0 0 32 200
use FILL  FILL_NAND2X1_199
timestamp 1515882711
transform 1 0 4408 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_199
timestamp 1515882711
transform 1 0 4424 0 1 610
box 0 0 48 200
use FILL  FILL_BUFX2_12
timestamp 1515882711
transform 1 0 4472 0 1 610
box 0 0 16 200
use BUFX2  BUFX2_12
timestamp 1515882711
transform 1 0 4488 0 1 610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_334
timestamp 1515882711
transform -1 0 4552 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_334
timestamp 1515882711
transform -1 0 4744 0 1 610
box 0 0 192 200
use FILL  FILL_NAND2X1_360
timestamp 1515882711
transform 1 0 4744 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_360
timestamp 1515882711
transform 1 0 4760 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_284
timestamp 1515882711
transform -1 0 4872 0 1 610
box 0 0 64 200
use FILL  FILL_INVX1_48
timestamp 1515882711
transform -1 0 4888 0 1 610
box 0 0 16 200
use INVX1  INVX1_48
timestamp 1515882711
transform -1 0 4920 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_71
timestamp 1515882711
transform 1 0 4920 0 1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_52
timestamp 1515882711
transform -1 0 5000 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_52
timestamp 1515882711
transform -1 0 5048 0 1 610
box 0 0 48 200
use FILL  FILL_3_4_0
timestamp 1515882711
transform -1 0 5064 0 1 610
box 0 0 16 200
use FILL  FILL_3_4_1
timestamp 1515882711
transform -1 0 5080 0 1 610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_71
timestamp 1515882711
transform -1 0 5096 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_71
timestamp 1515882711
transform -1 0 5288 0 1 610
box 0 0 192 200
use FILL  FILL_NAND2X1_256
timestamp 1515882711
transform -1 0 5304 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_256
timestamp 1515882711
transform -1 0 5352 0 1 610
box 0 0 48 200
use FILL  FILL_BUFX4_293
timestamp 1515882711
transform -1 0 5368 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_293
timestamp 1515882711
transform -1 0 5432 0 1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_13
timestamp 1515882711
transform 1 0 5432 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_13
timestamp 1515882711
transform 1 0 5448 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_503
timestamp 1515882711
transform -1 0 5560 0 1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_26
timestamp 1515882711
transform -1 0 5576 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_26
timestamp 1515882711
transform -1 0 5768 0 1 610
box 0 0 192 200
use FILL  FILL_BUFX4_303
timestamp 1515882711
transform 1 0 5768 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_303
timestamp 1515882711
transform 1 0 5784 0 1 610
box 0 0 64 200
use FILL  FILL_MUX2X1_25
timestamp 1515882711
transform 1 0 5848 0 1 610
box 0 0 16 200
use MUX2X1  MUX2X1_25
timestamp 1515882711
transform 1 0 5864 0 1 610
box 0 0 96 200
use FILL  FILL_NAND2X1_103
timestamp 1515882711
transform -1 0 5976 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_103
timestamp 1515882711
transform -1 0 6024 0 1 610
box 0 0 48 200
use FILL  FILL_MUX2X1_35
timestamp 1515882711
transform 1 0 6024 0 1 610
box 0 0 16 200
use FILL  FILL_3_5_0
timestamp 1515882711
transform 1 0 6040 0 1 610
box 0 0 16 200
use FILL  FILL_3_5_1
timestamp 1515882711
transform 1 0 6056 0 1 610
box 0 0 16 200
use MUX2X1  MUX2X1_35
timestamp 1515882711
transform 1 0 6072 0 1 610
box 0 0 96 200
use FILL  FILL_NAND2X1_99
timestamp 1515882711
transform 1 0 6168 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_99
timestamp 1515882711
transform 1 0 6184 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_418
timestamp 1515882711
transform 1 0 6232 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_415
timestamp 1515882711
transform 1 0 6280 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_473
timestamp 1515882711
transform -1 0 6392 0 1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_329
timestamp 1515882711
transform -1 0 6408 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_329
timestamp 1515882711
transform -1 0 6600 0 1 610
box 0 0 192 200
use FILL  FILL_MUX2X1_36
timestamp 1515882711
transform 1 0 6600 0 1 610
box 0 0 16 200
use MUX2X1  MUX2X1_36
timestamp 1515882711
transform 1 0 6616 0 1 610
box 0 0 96 200
use FILL  FILL_MUX2X1_44
timestamp 1515882711
transform 1 0 6712 0 1 610
box 0 0 16 200
use MUX2X1  MUX2X1_44
timestamp 1515882711
transform 1 0 6728 0 1 610
box 0 0 96 200
use NOR2X1  NOR2X1_148
timestamp 1515882711
transform -1 0 6872 0 1 610
box 0 0 48 200
use NOR3X1  NOR3X1_34
timestamp 1515882711
transform 1 0 6872 0 1 610
box 0 0 128 200
use FILL  FILL_BUFX4_197
timestamp 1515882711
transform 1 0 7000 0 1 610
box 0 0 16 200
use BUFX4  BUFX4_197
timestamp 1515882711
transform 1 0 7016 0 1 610
box 0 0 64 200
use FILL  FILL_3_6_0
timestamp 1515882711
transform -1 0 7096 0 1 610
box 0 0 16 200
use FILL  FILL_3_6_1
timestamp 1515882711
transform -1 0 7112 0 1 610
box 0 0 16 200
use FILL  FILL_NAND2X1_323
timestamp 1515882711
transform -1 0 7128 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_323
timestamp 1515882711
transform -1 0 7176 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_268
timestamp 1515882711
transform -1 0 7240 0 1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_112
timestamp 1515882711
transform -1 0 7256 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_112
timestamp 1515882711
transform -1 0 7448 0 1 610
box 0 0 192 200
use FILL  FILL_DFFPOSX1_132
timestamp 1515882711
transform 1 0 7448 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_132
timestamp 1515882711
transform 1 0 7464 0 1 610
box 0 0 192 200
use FILL  FILL_MUX2X1_20
timestamp 1515882711
transform 1 0 7656 0 1 610
box 0 0 16 200
use MUX2X1  MUX2X1_20
timestamp 1515882711
transform 1 0 7672 0 1 610
box 0 0 96 200
use NAND2X1  NAND2X1_425
timestamp 1515882711
transform 1 0 7768 0 1 610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_306
timestamp 1515882711
transform 1 0 7816 0 1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_306
timestamp 1515882711
transform 1 0 7832 0 1 610
box 0 0 192 200
use FILL  FILL_4_1
timestamp 1515882711
transform 1 0 8024 0 1 610
box 0 0 16 200
use FILL  FILL_4_2
timestamp 1515882711
transform 1 0 8040 0 1 610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_160
timestamp 1515882711
transform 1 0 8 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_160
timestamp 1515882711
transform 1 0 24 0 -1 610
box 0 0 192 200
use NAND3X1  NAND3X1_46
timestamp 1515882711
transform 1 0 216 0 -1 610
box 0 0 64 200
use FILL  FILL_AOI21X1_10
timestamp 1515882711
transform 1 0 280 0 -1 610
box 0 0 16 200
use AOI21X1  AOI21X1_10
timestamp 1515882711
transform 1 0 296 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_86
timestamp 1515882711
transform 1 0 360 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_87
timestamp 1515882711
transform -1 0 472 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_84
timestamp 1515882711
transform 1 0 472 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_43
timestamp 1515882711
transform -1 0 600 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_40
timestamp 1515882711
transform 1 0 600 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_217
timestamp 1515882711
transform 1 0 664 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_210
timestamp 1515882711
transform 1 0 728 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_210
timestamp 1515882711
transform 1 0 744 0 -1 610
box 0 0 192 200
use FILL  FILL_2_0_0
timestamp 1515882711
transform 1 0 936 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1515882711
transform 1 0 952 0 -1 610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_208
timestamp 1515882711
transform 1 0 968 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_208
timestamp 1515882711
transform 1 0 984 0 -1 610
box 0 0 192 200
use NOR3X1  NOR3X1_41
timestamp 1515882711
transform -1 0 1304 0 -1 610
box 0 0 128 200
use OAI21X1  OAI21X1_414
timestamp 1515882711
transform -1 0 1368 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_326
timestamp 1515882711
transform -1 0 1432 0 -1 610
box 0 0 64 200
use NOR3X1  NOR3X1_20
timestamp 1515882711
transform 1 0 1432 0 -1 610
box 0 0 128 200
use NOR3X1  NOR3X1_28
timestamp 1515882711
transform -1 0 1688 0 -1 610
box 0 0 128 200
use OAI21X1  OAI21X1_360
timestamp 1515882711
transform -1 0 1752 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_83
timestamp 1515882711
transform 1 0 1752 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_361
timestamp 1515882711
transform -1 0 1880 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_206
timestamp 1515882711
transform -1 0 1944 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_159
timestamp 1515882711
transform -1 0 1960 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_0
timestamp 1515882711
transform -1 0 1976 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1515882711
transform -1 0 1992 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_159
timestamp 1515882711
transform -1 0 2040 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_205
timestamp 1515882711
transform -1 0 2104 0 -1 610
box 0 0 64 200
use NOR3X1  NOR3X1_23
timestamp 1515882711
transform 1 0 2104 0 -1 610
box 0 0 128 200
use FILL  FILL_BUFX4_319
timestamp 1515882711
transform -1 0 2248 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_319
timestamp 1515882711
transform -1 0 2312 0 -1 610
box 0 0 64 200
use FILL  FILL_BUFX4_302
timestamp 1515882711
transform -1 0 2328 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_302
timestamp 1515882711
transform -1 0 2392 0 -1 610
box 0 0 64 200
use BUFX2  BUFX2_51
timestamp 1515882711
transform -1 0 2440 0 -1 610
box 0 0 48 200
use FILL  FILL_BUFX2_11
timestamp 1515882711
transform -1 0 2456 0 -1 610
box 0 0 16 200
use BUFX2  BUFX2_11
timestamp 1515882711
transform -1 0 2504 0 -1 610
box 0 0 48 200
use FILL  FILL_NAND2X1_391
timestamp 1515882711
transform 1 0 2504 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_391
timestamp 1515882711
transform 1 0 2520 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_459
timestamp 1515882711
transform -1 0 2632 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_387
timestamp 1515882711
transform -1 0 2648 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_387
timestamp 1515882711
transform -1 0 2696 0 -1 610
box 0 0 48 200
use FILL  FILL_DFFPOSX1_14
timestamp 1515882711
transform 1 0 2696 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_14
timestamp 1515882711
transform 1 0 2712 0 -1 610
box 0 0 192 200
use FILL  FILL_INVX1_72
timestamp 1515882711
transform 1 0 2904 0 -1 610
box 0 0 16 200
use INVX1  INVX1_72
timestamp 1515882711
transform 1 0 2920 0 -1 610
box 0 0 32 200
use FILL  FILL_NAND2X1_198
timestamp 1515882711
transform -1 0 2968 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_0
timestamp 1515882711
transform -1 0 2984 0 -1 610
box 0 0 16 200
use FILL  FILL_2_2_1
timestamp 1515882711
transform -1 0 3000 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_198
timestamp 1515882711
transform -1 0 3048 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_18
timestamp 1515882711
transform -1 0 3112 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_385
timestamp 1515882711
transform 1 0 3112 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_385
timestamp 1515882711
transform 1 0 3128 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_453
timestamp 1515882711
transform 1 0 3176 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_8
timestamp 1515882711
transform 1 0 3240 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1515882711
transform 1 0 3256 0 -1 610
box 0 0 192 200
use FILL  FILL_NAND2X1_292
timestamp 1515882711
transform -1 0 3464 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_292
timestamp 1515882711
transform -1 0 3512 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_329
timestamp 1515882711
transform -1 0 3576 0 -1 610
box 0 0 64 200
use FILL  FILL_BUFX4_63
timestamp 1515882711
transform -1 0 3592 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_63
timestamp 1515882711
transform -1 0 3656 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_22
timestamp 1515882711
transform -1 0 3672 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_22
timestamp 1515882711
transform -1 0 3720 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_43
timestamp 1515882711
transform -1 0 3784 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_43
timestamp 1515882711
transform -1 0 3800 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_43
timestamp 1515882711
transform -1 0 3992 0 -1 610
box 0 0 192 200
use FILL  FILL_2_3_0
timestamp 1515882711
transform -1 0 4008 0 -1 610
box 0 0 16 200
use FILL  FILL_2_3_1
timestamp 1515882711
transform -1 0 4024 0 -1 610
box 0 0 16 200
use NAND3X1  NAND3X1_226
timestamp 1515882711
transform -1 0 4088 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_48
timestamp 1515882711
transform -1 0 4152 0 -1 610
box 0 0 64 200
use FILL  FILL_INVX1_73
timestamp 1515882711
transform -1 0 4168 0 -1 610
box 0 0 16 200
use INVX1  INVX1_73
timestamp 1515882711
transform -1 0 4200 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_124
timestamp 1515882711
transform -1 0 4264 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_28
timestamp 1515882711
transform 1 0 4264 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_28
timestamp 1515882711
transform 1 0 4280 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_49
timestamp 1515882711
transform -1 0 4392 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_49
timestamp 1515882711
transform -1 0 4408 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_49
timestamp 1515882711
transform -1 0 4600 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_300
timestamp 1515882711
transform 1 0 4600 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_270
timestamp 1515882711
transform -1 0 4680 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_270
timestamp 1515882711
transform -1 0 4728 0 -1 610
box 0 0 48 200
use FILL  FILL_INVX1_57
timestamp 1515882711
transform -1 0 4744 0 -1 610
box 0 0 16 200
use INVX1  INVX1_57
timestamp 1515882711
transform -1 0 4776 0 -1 610
box 0 0 32 200
use OAI21X1  OAI21X1_427
timestamp 1515882711
transform -1 0 4840 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_45
timestamp 1515882711
transform -1 0 4856 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_45
timestamp 1515882711
transform -1 0 5048 0 -1 610
box 0 0 192 200
use FILL  FILL_2_4_0
timestamp 1515882711
transform 1 0 5048 0 -1 610
box 0 0 16 200
use FILL  FILL_2_4_1
timestamp 1515882711
transform 1 0 5064 0 -1 610
box 0 0 16 200
use FILL  FILL_NAND2X1_25
timestamp 1515882711
transform 1 0 5080 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_25
timestamp 1515882711
transform 1 0 5096 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_45
timestamp 1515882711
transform -1 0 5208 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_15
timestamp 1515882711
transform 1 0 5208 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_15
timestamp 1515882711
transform 1 0 5224 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_36
timestamp 1515882711
transform -1 0 5336 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_304
timestamp 1515882711
transform 1 0 5336 0 -1 610
box 0 0 64 200
use FILL  FILL_BUFX4_64
timestamp 1515882711
transform -1 0 5416 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_64
timestamp 1515882711
transform -1 0 5480 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_272
timestamp 1515882711
transform -1 0 5496 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_272
timestamp 1515882711
transform -1 0 5544 0 -1 610
box 0 0 48 200
use FILL  FILL_BUFX4_106
timestamp 1515882711
transform -1 0 5560 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_106
timestamp 1515882711
transform -1 0 5624 0 -1 610
box 0 0 64 200
use FILL  FILL_NAND2X1_41
timestamp 1515882711
transform 1 0 5624 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_41
timestamp 1515882711
transform 1 0 5640 0 -1 610
box 0 0 48 200
use OAI21X1  OAI21X1_61
timestamp 1515882711
transform 1 0 5688 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_61
timestamp 1515882711
transform 1 0 5752 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_61
timestamp 1515882711
transform 1 0 5768 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_120
timestamp 1515882711
transform -1 0 6024 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_120
timestamp 1515882711
transform -1 0 6040 0 -1 610
box 0 0 16 200
use FILL  FILL_2_5_0
timestamp 1515882711
transform -1 0 6056 0 -1 610
box 0 0 16 200
use FILL  FILL_2_5_1
timestamp 1515882711
transform -1 0 6072 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_120
timestamp 1515882711
transform -1 0 6264 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_117
timestamp 1515882711
transform -1 0 6328 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_469
timestamp 1515882711
transform -1 0 6392 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_117
timestamp 1515882711
transform 1 0 6392 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_117
timestamp 1515882711
transform 1 0 6408 0 -1 610
box 0 0 192 200
use FILL  FILL_BUFX4_12
timestamp 1515882711
transform 1 0 6600 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_12
timestamp 1515882711
transform 1 0 6616 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_326
timestamp 1515882711
transform 1 0 6680 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_326
timestamp 1515882711
transform 1 0 6696 0 -1 610
box 0 0 192 200
use FILL  FILL_BUFX4_107
timestamp 1515882711
transform 1 0 6888 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_107
timestamp 1515882711
transform 1 0 6904 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_401
timestamp 1515882711
transform 1 0 6968 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_400
timestamp 1515882711
transform -1 0 7080 0 -1 610
box 0 0 48 200
use FILL  FILL_2_6_0
timestamp 1515882711
transform -1 0 7096 0 -1 610
box 0 0 16 200
use FILL  FILL_2_6_1
timestamp 1515882711
transform -1 0 7112 0 -1 610
box 0 0 16 200
use FILL  FILL_DFFPOSX1_46
timestamp 1515882711
transform -1 0 7128 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_46
timestamp 1515882711
transform -1 0 7320 0 -1 610
box 0 0 192 200
use OAI21X1  OAI21X1_115
timestamp 1515882711
transform 1 0 7320 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_115
timestamp 1515882711
transform 1 0 7384 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_115
timestamp 1515882711
transform 1 0 7400 0 -1 610
box 0 0 192 200
use FILL  FILL_BUFX4_65
timestamp 1515882711
transform -1 0 7608 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_65
timestamp 1515882711
transform -1 0 7672 0 -1 610
box 0 0 64 200
use FILL  FILL_BUFX4_66
timestamp 1515882711
transform 1 0 7672 0 -1 610
box 0 0 16 200
use BUFX4  BUFX4_66
timestamp 1515882711
transform 1 0 7688 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_477
timestamp 1515882711
transform 1 0 7752 0 -1 610
box 0 0 64 200
use FILL  FILL_DFFPOSX1_299
timestamp 1515882711
transform 1 0 7816 0 -1 610
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_299
timestamp 1515882711
transform 1 0 7832 0 -1 610
box 0 0 192 200
use FILL  FILL_3_1
timestamp 1515882711
transform -1 0 8040 0 -1 610
box 0 0 16 200
use FILL  FILL_3_2
timestamp 1515882711
transform -1 0 8056 0 -1 610
box 0 0 16 200
use NAND3X1  NAND3X1_68
timestamp 1515882711
transform -1 0 72 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_57
timestamp 1515882711
transform -1 0 136 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_79
timestamp 1515882711
transform -1 0 200 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_85
timestamp 1515882711
transform 1 0 200 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_86
timestamp 1515882711
transform 1 0 264 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_42
timestamp 1515882711
transform -1 0 392 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_219
timestamp 1515882711
transform 1 0 392 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_220
timestamp 1515882711
transform -1 0 520 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_41
timestamp 1515882711
transform -1 0 584 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_218
timestamp 1515882711
transform 1 0 584 0 1 210
box 0 0 64 200
use FILL  FILL_AOI21X1_28
timestamp 1515882711
transform 1 0 648 0 1 210
box 0 0 16 200
use AOI21X1  AOI21X1_28
timestamp 1515882711
transform 1 0 664 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_104
timestamp 1515882711
transform -1 0 776 0 1 210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_227
timestamp 1515882711
transform -1 0 792 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_227
timestamp 1515882711
transform -1 0 984 0 1 210
box 0 0 192 200
use FILL  FILL_1_0_0
timestamp 1515882711
transform -1 0 1000 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1515882711
transform -1 0 1016 0 1 210
box 0 0 16 200
use NAND3X1  NAND3X1_24
timestamp 1515882711
transform -1 0 1080 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_82
timestamp 1515882711
transform 1 0 1080 0 1 210
box 0 0 64 200
use FILL  FILL_AOI21X1_61
timestamp 1515882711
transform 1 0 1144 0 1 210
box 0 0 16 200
use AOI21X1  AOI21X1_61
timestamp 1515882711
transform 1 0 1160 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_137
timestamp 1515882711
transform -1 0 1272 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_216
timestamp 1515882711
transform -1 0 1336 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_39
timestamp 1515882711
transform 1 0 1336 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_35
timestamp 1515882711
transform -1 0 1464 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_121
timestamp 1515882711
transform 1 0 1464 0 1 210
box 0 0 48 200
use FILL  FILL_AOI21X1_46
timestamp 1515882711
transform -1 0 1528 0 1 210
box 0 0 16 200
use AOI21X1  AOI21X1_46
timestamp 1515882711
transform -1 0 1592 0 1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_231
timestamp 1515882711
transform -1 0 1608 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_231
timestamp 1515882711
transform -1 0 1800 0 1 210
box 0 0 192 200
use FILL  FILL_INVX2_11
timestamp 1515882711
transform 1 0 1800 0 1 210
box 0 0 16 200
use INVX2  INVX2_11
timestamp 1515882711
transform 1 0 1816 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_178
timestamp 1515882711
transform 1 0 1848 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_163
timestamp 1515882711
transform -1 0 1928 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_163
timestamp 1515882711
transform -1 0 1976 0 1 210
box 0 0 48 200
use FILL  FILL_1_1_0
timestamp 1515882711
transform 1 0 1976 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1515882711
transform 1 0 1992 0 1 210
box 0 0 16 200
use FILL  FILL_NAND2X1_145
timestamp 1515882711
transform 1 0 2008 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_145
timestamp 1515882711
transform 1 0 2024 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_161
timestamp 1515882711
transform -1 0 2136 0 1 210
box 0 0 64 200
use FILL  FILL_INVX2_23
timestamp 1515882711
transform -1 0 2152 0 1 210
box 0 0 16 200
use INVX2  INVX2_23
timestamp 1515882711
transform -1 0 2184 0 1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_177
timestamp 1515882711
transform -1 0 2200 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_177
timestamp 1515882711
transform -1 0 2392 0 1 210
box 0 0 192 200
use FILL  FILL_BUFX4_165
timestamp 1515882711
transform -1 0 2408 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_165
timestamp 1515882711
transform -1 0 2472 0 1 210
box 0 0 64 200
use FILL  FILL_INVX8_8
timestamp 1515882711
transform 1 0 2472 0 1 210
box 0 0 16 200
use INVX8  INVX8_8
timestamp 1515882711
transform 1 0 2488 0 1 210
box 0 0 80 200
use FILL  FILL_BUFX4_229
timestamp 1515882711
transform -1 0 2584 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_229
timestamp 1515882711
transform -1 0 2648 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_377
timestamp 1515882711
transform 1 0 2648 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_377
timestamp 1515882711
transform 1 0 2664 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_444
timestamp 1515882711
transform -1 0 2776 0 1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_351
timestamp 1515882711
transform 1 0 2776 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_351
timestamp 1515882711
transform 1 0 2792 0 1 210
box 0 0 192 200
use FILL  FILL_1_2_0
timestamp 1515882711
transform -1 0 3000 0 1 210
box 0 0 16 200
use FILL  FILL_1_2_1
timestamp 1515882711
transform -1 0 3016 0 1 210
box 0 0 16 200
use FILL  FILL_INVX1_6
timestamp 1515882711
transform -1 0 3032 0 1 210
box 0 0 16 200
use INVX1  INVX1_6
timestamp 1515882711
transform -1 0 3064 0 1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_280
timestamp 1515882711
transform -1 0 3080 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_280
timestamp 1515882711
transform -1 0 3272 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_31
timestamp 1515882711
transform -1 0 3336 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_9
timestamp 1515882711
transform -1 0 3352 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_9
timestamp 1515882711
transform -1 0 3400 0 1 210
box 0 0 48 200
use FILL  FILL_BUFX4_15
timestamp 1515882711
transform -1 0 3416 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_15
timestamp 1515882711
transform -1 0 3480 0 1 210
box 0 0 64 200
use FILL  FILL_INVX8_11
timestamp 1515882711
transform 1 0 3480 0 1 210
box 0 0 16 200
use INVX8  INVX8_11
timestamp 1515882711
transform 1 0 3496 0 1 210
box 0 0 80 200
use FILL  FILL_BUFX2_32
timestamp 1515882711
transform 1 0 3576 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_32
timestamp 1515882711
transform 1 0 3592 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_350
timestamp 1515882711
transform -1 0 3704 0 1 210
box 0 0 64 200
use FILL  FILL_BUFX2_26
timestamp 1515882711
transform 1 0 3704 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_26
timestamp 1515882711
transform 1 0 3720 0 1 210
box 0 0 48 200
use FILL  FILL_BUFX2_3
timestamp 1515882711
transform -1 0 3784 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_3
timestamp 1515882711
transform -1 0 3832 0 1 210
box 0 0 48 200
use FILL  FILL_NAND2X1_11
timestamp 1515882711
transform 1 0 3832 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_11
timestamp 1515882711
transform 1 0 3848 0 1 210
box 0 0 48 200
use FILL  FILL_BUFX2_18
timestamp 1515882711
transform 1 0 3896 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_18
timestamp 1515882711
transform 1 0 3912 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_33
timestamp 1515882711
transform -1 0 4024 0 1 210
box 0 0 64 200
use FILL  FILL_1_3_0
timestamp 1515882711
transform 1 0 4024 0 1 210
box 0 0 16 200
use FILL  FILL_1_3_1
timestamp 1515882711
transform 1 0 4040 0 1 210
box 0 0 16 200
use FILL  FILL_BUFX2_6
timestamp 1515882711
transform 1 0 4056 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_6
timestamp 1515882711
transform 1 0 4072 0 1 210
box 0 0 48 200
use FILL  FILL_BUFX2_24
timestamp 1515882711
transform 1 0 4120 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_24
timestamp 1515882711
transform 1 0 4136 0 1 210
box 0 0 48 200
use FILL  FILL_BUFX2_10
timestamp 1515882711
transform -1 0 4200 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_10
timestamp 1515882711
transform -1 0 4248 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_84
timestamp 1515882711
transform 1 0 4248 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_65
timestamp 1515882711
transform -1 0 4328 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_65
timestamp 1515882711
transform -1 0 4376 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_332
timestamp 1515882711
transform -1 0 4440 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_294
timestamp 1515882711
transform 1 0 4440 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_294
timestamp 1515882711
transform 1 0 4456 0 1 210
box 0 0 48 200
use FILL  FILL_NAND2X1_257
timestamp 1515882711
transform 1 0 4504 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_257
timestamp 1515882711
transform 1 0 4520 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_224
timestamp 1515882711
transform 1 0 4568 0 1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_344
timestamp 1515882711
transform -1 0 4648 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_344
timestamp 1515882711
transform -1 0 4840 0 1 210
box 0 0 192 200
use FILL  FILL_NAND2X1_370
timestamp 1515882711
transform 1 0 4840 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_370
timestamp 1515882711
transform 1 0 4856 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_437
timestamp 1515882711
transform -1 0 4968 0 1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_63
timestamp 1515882711
transform 1 0 4968 0 1 210
box 0 0 16 200
use FILL  FILL_1_4_0
timestamp 1515882711
transform 1 0 4984 0 1 210
box 0 0 16 200
use FILL  FILL_1_4_1
timestamp 1515882711
transform 1 0 5000 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_63
timestamp 1515882711
transform 1 0 5016 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_63
timestamp 1515882711
transform 1 0 5208 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_43
timestamp 1515882711
transform -1 0 5288 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_43
timestamp 1515882711
transform -1 0 5336 0 1 210
box 0 0 48 200
use FILL  FILL_INVX1_59
timestamp 1515882711
transform 1 0 5336 0 1 210
box 0 0 16 200
use INVX1  INVX1_59
timestamp 1515882711
transform 1 0 5352 0 1 210
box 0 0 32 200
use FILL  FILL_NAND2X1_224
timestamp 1515882711
transform -1 0 5400 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_224
timestamp 1515882711
transform -1 0 5448 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_190
timestamp 1515882711
transform -1 0 5512 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_333
timestamp 1515882711
transform -1 0 5576 0 1 210
box 0 0 64 200
use FILL  FILL_INVX1_75
timestamp 1515882711
transform -1 0 5592 0 1 210
box 0 0 16 200
use INVX1  INVX1_75
timestamp 1515882711
transform -1 0 5624 0 1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_190
timestamp 1515882711
transform -1 0 5640 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_190
timestamp 1515882711
transform -1 0 5832 0 1 210
box 0 0 192 200
use FILL  FILL_BUFX4_204
timestamp 1515882711
transform 1 0 5832 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_204
timestamp 1515882711
transform 1 0 5848 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_295
timestamp 1515882711
transform 1 0 5912 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_295
timestamp 1515882711
transform 1 0 5928 0 1 210
box 0 0 48 200
use FILL  FILL_BUFX4_28
timestamp 1515882711
transform 1 0 5976 0 1 210
box 0 0 16 200
use BUFX4  BUFX4_28
timestamp 1515882711
transform 1 0 5992 0 1 210
box 0 0 64 200
use FILL  FILL_1_5_0
timestamp 1515882711
transform 1 0 6056 0 1 210
box 0 0 16 200
use FILL  FILL_1_5_1
timestamp 1515882711
transform 1 0 6072 0 1 210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_13
timestamp 1515882711
transform 1 0 6088 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1515882711
transform 1 0 6104 0 1 210
box 0 0 192 200
use FILL  FILL_MUX2X1_26
timestamp 1515882711
transform -1 0 6312 0 1 210
box 0 0 16 200
use MUX2X1  MUX2X1_26
timestamp 1515882711
transform -1 0 6408 0 1 210
box 0 0 96 200
use FILL  FILL_DFFPOSX1_102
timestamp 1515882711
transform 1 0 6408 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_102
timestamp 1515882711
transform 1 0 6424 0 1 210
box 0 0 192 200
use OAI21X1  OAI21X1_102
timestamp 1515882711
transform 1 0 6616 0 1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_84
timestamp 1515882711
transform 1 0 6680 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_84
timestamp 1515882711
transform 1 0 6696 0 1 210
box 0 0 48 200
use FILL  FILL_MUX2X1_19
timestamp 1515882711
transform -1 0 6760 0 1 210
box 0 0 16 200
use MUX2X1  MUX2X1_19
timestamp 1515882711
transform -1 0 6856 0 1 210
box 0 0 96 200
use FILL  FILL_MUX2X1_18
timestamp 1515882711
transform 1 0 6856 0 1 210
box 0 0 16 200
use MUX2X1  MUX2X1_18
timestamp 1515882711
transform 1 0 6872 0 1 210
box 0 0 96 200
use FILL  FILL_NAND2X1_97
timestamp 1515882711
transform 1 0 6968 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_97
timestamp 1515882711
transform 1 0 6984 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_467
timestamp 1515882711
transform 1 0 7032 0 1 210
box 0 0 64 200
use FILL  FILL_1_6_0
timestamp 1515882711
transform -1 0 7112 0 1 210
box 0 0 16 200
use FILL  FILL_1_6_1
timestamp 1515882711
transform -1 0 7128 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_413
timestamp 1515882711
transform -1 0 7176 0 1 210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_324
timestamp 1515882711
transform -1 0 7192 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_324
timestamp 1515882711
transform -1 0 7384 0 1 210
box 0 0 192 200
use FILL  FILL_MUX2X1_34
timestamp 1515882711
transform -1 0 7400 0 1 210
box 0 0 16 200
use MUX2X1  MUX2X1_34
timestamp 1515882711
transform -1 0 7496 0 1 210
box 0 0 96 200
use FILL  FILL_NAND2X1_89
timestamp 1515882711
transform 1 0 7496 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_89
timestamp 1515882711
transform 1 0 7512 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_106
timestamp 1515882711
transform -1 0 7624 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_405
timestamp 1515882711
transform 1 0 7624 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_446
timestamp 1515882711
transform -1 0 7736 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_142
timestamp 1515882711
transform 1 0 7736 0 1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_142
timestamp 1515882711
transform 1 0 7800 0 1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_142
timestamp 1515882711
transform 1 0 7816 0 1 210
box 0 0 192 200
use FILL  FILL_2_1
timestamp 1515882711
transform 1 0 8008 0 1 210
box 0 0 16 200
use FILL  FILL_2_2
timestamp 1515882711
transform 1 0 8024 0 1 210
box 0 0 16 200
use FILL  FILL_2_3
timestamp 1515882711
transform 1 0 8040 0 1 210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_249
timestamp 1515882711
transform -1 0 24 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_249
timestamp 1515882711
transform -1 0 216 0 -1 210
box 0 0 192 200
use NOR2X1  NOR2X1_13
timestamp 1515882711
transform -1 0 264 0 -1 210
box 0 0 48 200
use FILL  FILL_AOI21X1_12
timestamp 1515882711
transform -1 0 280 0 -1 210
box 0 0 16 200
use AOI21X1  AOI21X1_12
timestamp 1515882711
transform -1 0 344 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_82
timestamp 1515882711
transform -1 0 392 0 -1 210
box 0 0 48 200
use FILL  FILL_AOI21X1_6
timestamp 1515882711
transform -1 0 408 0 -1 210
box 0 0 16 200
use AOI21X1  AOI21X1_6
timestamp 1515882711
transform -1 0 472 0 -1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_262
timestamp 1515882711
transform 1 0 472 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_262
timestamp 1515882711
transform 1 0 488 0 -1 210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_195
timestamp 1515882711
transform 1 0 680 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_195
timestamp 1515882711
transform 1 0 696 0 -1 210
box 0 0 192 200
use FILL  FILL_AOI21X1_59
timestamp 1515882711
transform 1 0 888 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_0
timestamp 1515882711
transform 1 0 904 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1515882711
transform 1 0 920 0 -1 210
box 0 0 16 200
use AOI21X1  AOI21X1_59
timestamp 1515882711
transform 1 0 936 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_135
timestamp 1515882711
transform 1 0 1000 0 -1 210
box 0 0 48 200
use FILL  FILL_BUFX4_16
timestamp 1515882711
transform -1 0 1064 0 -1 210
box 0 0 16 200
use BUFX4  BUFX4_16
timestamp 1515882711
transform -1 0 1128 0 -1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_229
timestamp 1515882711
transform 1 0 1128 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_229
timestamp 1515882711
transform 1 0 1144 0 -1 210
box 0 0 192 200
use FILL  FILL_INVX2_25
timestamp 1515882711
transform -1 0 1352 0 -1 210
box 0 0 16 200
use INVX2  INVX2_25
timestamp 1515882711
transform -1 0 1384 0 -1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_244
timestamp 1515882711
transform -1 0 1400 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_244
timestamp 1515882711
transform -1 0 1592 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_192
timestamp 1515882711
transform 1 0 1592 0 -1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_176
timestamp 1515882711
transform -1 0 1672 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_176
timestamp 1515882711
transform -1 0 1720 0 -1 210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_213
timestamp 1515882711
transform -1 0 1736 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_213
timestamp 1515882711
transform -1 0 1928 0 -1 210
box 0 0 192 200
use FILL  FILL_INVX2_27
timestamp 1515882711
transform -1 0 1944 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_0
timestamp 1515882711
transform -1 0 1960 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1515882711
transform -1 0 1976 0 -1 210
box 0 0 16 200
use INVX2  INVX2_27
timestamp 1515882711
transform -1 0 2008 0 -1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_247
timestamp 1515882711
transform -1 0 2024 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_247
timestamp 1515882711
transform -1 0 2216 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_194
timestamp 1515882711
transform 1 0 2216 0 -1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_178
timestamp 1515882711
transform -1 0 2296 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_178
timestamp 1515882711
transform -1 0 2344 0 -1 210
box 0 0 48 200
use FILL  FILL_INVX2_9
timestamp 1515882711
transform -1 0 2360 0 -1 210
box 0 0 16 200
use INVX2  INVX2_9
timestamp 1515882711
transform -1 0 2392 0 -1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_193
timestamp 1515882711
transform -1 0 2408 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_193
timestamp 1515882711
transform -1 0 2600 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_176
timestamp 1515882711
transform 1 0 2600 0 -1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_161
timestamp 1515882711
transform -1 0 2680 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_161
timestamp 1515882711
transform -1 0 2728 0 -1 210
box 0 0 48 200
use FILL  FILL_INVX8_6
timestamp 1515882711
transform 1 0 2728 0 -1 210
box 0 0 16 200
use INVX8  INVX8_6
timestamp 1515882711
transform 1 0 2744 0 -1 210
box 0 0 80 200
use FILL  FILL_INVX8_3
timestamp 1515882711
transform 1 0 2824 0 -1 210
box 0 0 16 200
use INVX8  INVX8_3
timestamp 1515882711
transform 1 0 2840 0 -1 210
box 0 0 80 200
use FILL  FILL_NAND2X1_393
timestamp 1515882711
transform 1 0 2920 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_393
timestamp 1515882711
transform 1 0 2936 0 -1 210
box 0 0 48 200
use FILL  FILL_0_2_0
timestamp 1515882711
transform -1 0 3000 0 -1 210
box 0 0 16 200
use FILL  FILL_0_2_1
timestamp 1515882711
transform -1 0 3016 0 -1 210
box 0 0 16 200
use OAI21X1  OAI21X1_461
timestamp 1515882711
transform -1 0 3080 0 -1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_16
timestamp 1515882711
transform 1 0 3080 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1515882711
transform 1 0 3096 0 -1 210
box 0 0 192 200
use FILL  FILL_INVX1_83
timestamp 1515882711
transform 1 0 3288 0 -1 210
box 0 0 16 200
use INVX1  INVX1_83
timestamp 1515882711
transform 1 0 3304 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_49
timestamp 1515882711
transform -1 0 3384 0 -1 210
box 0 0 48 200
use FILL  FILL_BUFX2_9
timestamp 1515882711
transform -1 0 3400 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_9
timestamp 1515882711
transform -1 0 3448 0 -1 210
box 0 0 48 200
use FILL  FILL_NAND2X1_307
timestamp 1515882711
transform -1 0 3464 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_307
timestamp 1515882711
transform -1 0 3512 0 -1 210
box 0 0 48 200
use FILL  FILL_BUFX2_1
timestamp 1515882711
transform 1 0 3512 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_1
timestamp 1515882711
transform 1 0 3528 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_33
timestamp 1515882711
transform -1 0 3624 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_41
timestamp 1515882711
transform 1 0 3624 0 -1 210
box 0 0 48 200
use FILL  FILL_BUFX4_202
timestamp 1515882711
transform 1 0 3672 0 -1 210
box 0 0 16 200
use BUFX4  BUFX4_202
timestamp 1515882711
transform 1 0 3688 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_64
timestamp 1515882711
transform 1 0 3752 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_43
timestamp 1515882711
transform 1 0 3800 0 -1 210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_282
timestamp 1515882711
transform -1 0 3864 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_282
timestamp 1515882711
transform -1 0 4056 0 -1 210
box 0 0 192 200
use FILL  FILL_0_3_0
timestamp 1515882711
transform -1 0 4072 0 -1 210
box 0 0 16 200
use FILL  FILL_0_3_1
timestamp 1515882711
transform -1 0 4088 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_48
timestamp 1515882711
transform -1 0 4136 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_57
timestamp 1515882711
transform -1 0 4184 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_46
timestamp 1515882711
transform -1 0 4232 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_62
timestamp 1515882711
transform -1 0 4280 0 -1 210
box 0 0 48 200
use FILL  FILL_BUFX2_20
timestamp 1515882711
transform 1 0 4280 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_20
timestamp 1515882711
transform 1 0 4296 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_59
timestamp 1515882711
transform 1 0 4344 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_50
timestamp 1515882711
transform 1 0 4392 0 -1 210
box 0 0 48 200
use FILL  FILL_INVX1_74
timestamp 1515882711
transform -1 0 4456 0 -1 210
box 0 0 16 200
use INVX1  INVX1_74
timestamp 1515882711
transform -1 0 4488 0 -1 210
box 0 0 32 200
use FILL  FILL_DFFPOSX1_84
timestamp 1515882711
transform 1 0 4488 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_84
timestamp 1515882711
transform 1 0 4504 0 -1 210
box 0 0 192 200
use BUFX2  BUFX2_34
timestamp 1515882711
transform -1 0 4744 0 -1 210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_224
timestamp 1515882711
transform -1 0 4760 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_224
timestamp 1515882711
transform -1 0 4952 0 -1 210
box 0 0 192 200
use FILL  FILL_BUFX4_27
timestamp 1515882711
transform 1 0 4952 0 -1 210
box 0 0 16 200
use BUFX4  BUFX4_27
timestamp 1515882711
transform 1 0 4968 0 -1 210
box 0 0 64 200
use FILL  FILL_0_4_0
timestamp 1515882711
transform -1 0 5048 0 -1 210
box 0 0 16 200
use FILL  FILL_0_4_1
timestamp 1515882711
transform -1 0 5064 0 -1 210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_36
timestamp 1515882711
transform -1 0 5080 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_36
timestamp 1515882711
transform -1 0 5272 0 -1 210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_28
timestamp 1515882711
transform 1 0 5272 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_28
timestamp 1515882711
transform 1 0 5288 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_13
timestamp 1515882711
transform 1 0 5480 0 -1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_35
timestamp 1515882711
transform 1 0 5544 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_35
timestamp 1515882711
transform 1 0 5560 0 -1 210
box 0 0 48 200
use FILL  FILL_NAND2X1_47
timestamp 1515882711
transform 1 0 5608 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_47
timestamp 1515882711
transform 1 0 5624 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_66
timestamp 1515882711
transform -1 0 5736 0 -1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_66
timestamp 1515882711
transform -1 0 5752 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_66
timestamp 1515882711
transform -1 0 5944 0 -1 210
box 0 0 192 200
use FILL  FILL_NAND2X1_68
timestamp 1515882711
transform -1 0 5960 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_68
timestamp 1515882711
transform -1 0 6008 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_46
timestamp 1515882711
transform -1 0 6072 0 -1 210
box 0 0 64 200
use FILL  FILL_0_5_0
timestamp 1515882711
transform -1 0 6088 0 -1 210
box 0 0 16 200
use FILL  FILL_0_5_1
timestamp 1515882711
transform -1 0 6104 0 -1 210
box 0 0 16 200
use FILL  FILL_DFFPOSX1_31
timestamp 1515882711
transform -1 0 6120 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_31
timestamp 1515882711
transform -1 0 6312 0 -1 210
box 0 0 192 200
use OAI21X1  OAI21X1_368
timestamp 1515882711
transform 1 0 6312 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_396
timestamp 1515882711
transform -1 0 6424 0 -1 210
box 0 0 48 200
use FILL  FILL_BUFX4_14
timestamp 1515882711
transform -1 0 6440 0 -1 210
box 0 0 16 200
use BUFX4  BUFX4_14
timestamp 1515882711
transform -1 0 6504 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_98
timestamp 1515882711
transform 1 0 6504 0 -1 210
box 0 0 64 200
use FILL  FILL_NAND2X1_81
timestamp 1515882711
transform -1 0 6584 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_81
timestamp 1515882711
transform -1 0 6632 0 -1 210
box 0 0 48 200
use FILL  FILL_DFFPOSX1_98
timestamp 1515882711
transform 1 0 6632 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_98
timestamp 1515882711
transform 1 0 6648 0 -1 210
box 0 0 192 200
use FILL  FILL_NAND2X1_78
timestamp 1515882711
transform -1 0 6856 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_78
timestamp 1515882711
transform -1 0 6904 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_96
timestamp 1515882711
transform -1 0 6968 0 -1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_96
timestamp 1515882711
transform -1 0 6984 0 -1 210
box 0 0 16 200
use FILL  FILL_0_6_0
timestamp 1515882711
transform -1 0 7000 0 -1 210
box 0 0 16 200
use FILL  FILL_0_6_1
timestamp 1515882711
transform -1 0 7016 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_96
timestamp 1515882711
transform -1 0 7208 0 -1 210
box 0 0 192 200
use FILL  FILL_NAND2X1_394
timestamp 1515882711
transform 1 0 7208 0 -1 210
box 0 0 16 200
use NAND2X1  NAND2X1_394
timestamp 1515882711
transform 1 0 7224 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_346
timestamp 1515882711
transform -1 0 7336 0 -1 210
box 0 0 64 200
use FILL  FILL_DFFPOSX1_342
timestamp 1515882711
transform 1 0 7336 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_342
timestamp 1515882711
transform 1 0 7352 0 -1 210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_106
timestamp 1515882711
transform -1 0 7560 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_106
timestamp 1515882711
transform -1 0 7752 0 -1 210
box 0 0 192 200
use FILL  FILL_DFFPOSX1_316
timestamp 1515882711
transform -1 0 7768 0 -1 210
box 0 0 16 200
use DFFPOSX1  DFFPOSX1_316
timestamp 1515882711
transform -1 0 7960 0 -1 210
box 0 0 192 200
use FILL  FILL_INVX1_5
timestamp 1515882711
transform -1 0 7976 0 -1 210
box 0 0 16 200
use INVX1  INVX1_5
timestamp 1515882711
transform -1 0 8008 0 -1 210
box 0 0 32 200
use FILL  FILL_1_1
timestamp 1515882711
transform -1 0 8024 0 -1 210
box 0 0 16 200
use FILL  FILL_1_2
timestamp 1515882711
transform -1 0 8040 0 -1 210
box 0 0 16 200
use FILL  FILL_1_3
timestamp 1515882711
transform -1 0 8056 0 -1 210
box 0 0 16 200
<< labels >>
flabel space 1156 42 1164 136 6 FreeSans 48 0 0 0 vdd
port 0 nsew
flabel space 2180 42 2188 136 6 FreeSans 48 0 0 0 gnd
port 1 nsew
flabel metal3 -48 1740 -48 1740 7 FreeSans 48 0 0 0 REG_D<0>
port 2 nsew
flabel metal2 2656 -40 2656 -40 7 FreeSans 48 270 0 0 REG_D<1>
port 3 nsew
flabel metal2 2880 -40 2880 -40 7 FreeSans 48 270 0 0 REG_D<2>
port 4 nsew
flabel metal2 2272 5660 2272 5660 3 FreeSans 48 90 0 0 REG_D<3>
port 5 nsew
flabel metal2 2208 5660 2208 5660 3 FreeSans 48 90 0 0 REG_D<4>
port 6 nsew
flabel metal3 -48 4320 -48 4320 7 FreeSans 48 0 0 0 REG_D<5>
port 7 nsew
flabel metal2 2320 5660 2320 5660 3 FreeSans 48 90 0 0 REG_D<6>
port 8 nsew
flabel metal2 1680 5660 1680 5660 3 FreeSans 48 90 0 0 REG_D<7>
port 9 nsew
flabel metal2 2992 -40 2992 -40 7 FreeSans 48 270 0 0 REG_D<8>
port 10 nsew
flabel metal2 1840 5660 1840 5660 3 FreeSans 48 90 0 0 REG_D<9>
port 11 nsew
flabel metal2 2848 -40 2848 -40 7 FreeSans 48 270 0 0 REG_D<10>
port 12 nsew
flabel metal2 2816 5660 2816 5660 3 FreeSans 48 90 0 0 REG_D<11>
port 13 nsew
flabel metal2 1824 -40 1824 -40 7 FreeSans 48 270 0 0 REG_D<12>
port 14 nsew
flabel metal2 2000 -40 2000 -40 7 FreeSans 48 270 0 0 REG_D<13>
port 15 nsew
flabel metal2 2688 5660 2688 5660 3 FreeSans 48 90 0 0 REG_D<14>
port 16 nsew
flabel metal2 2944 -40 2944 -40 7 FreeSans 48 270 0 0 REG_D<15>
port 17 nsew
flabel metal2 3536 -40 3536 -40 7 FreeSans 48 270 0 0 REG_RF1<0>
port 18 nsew
flabel metal2 3488 -40 3488 -40 7 FreeSans 48 270 0 0 REG_RF1<1>
port 19 nsew
flabel metal2 2704 -40 2704 -40 7 FreeSans 48 270 0 0 REG_RF1<2>
port 20 nsew
flabel metal2 2528 -40 2528 -40 7 FreeSans 48 270 0 0 REG_RF1<3>
port 21 nsew
flabel metal3 -48 3160 -48 3160 7 FreeSans 48 0 0 0 REG_RF2<0>
port 22 nsew
flabel metal3 -48 3120 -48 3120 7 FreeSans 48 0 0 0 REG_RF2<1>
port 23 nsew
flabel metal3 -48 2920 -48 2920 7 FreeSans 48 0 0 0 REG_RF2<2>
port 24 nsew
flabel metal3 -48 2960 -48 2960 7 FreeSans 48 0 0 0 REG_RF2<3>
port 25 nsew
flabel metal3 8112 3060 8112 3060 3 FreeSans 48 0 0 0 REG_RFD<0>
port 26 nsew
flabel metal3 8112 3100 8112 3100 3 FreeSans 48 0 0 0 REG_RFD<1>
port 27 nsew
flabel metal3 8112 3140 8112 3140 3 FreeSans 48 0 0 0 REG_RFD<2>
port 28 nsew
flabel metal3 8112 3220 8112 3220 3 FreeSans 48 0 0 0 REG_RFD<3>
port 29 nsew
flabel metal3 -48 1120 -48 1120 7 FreeSans 48 0 0 0 REG_R1<0>
port 30 nsew
flabel metal3 -48 320 -48 320 7 FreeSans 48 0 0 0 REG_R1<1>
port 31 nsew
flabel metal3 -48 2360 -48 2360 7 FreeSans 48 0 0 0 REG_R1<2>
port 32 nsew
flabel metal3 -48 4720 -48 4720 7 FreeSans 48 0 0 0 REG_R1<3>
port 33 nsew
flabel metal3 -48 4360 -48 4360 7 FreeSans 48 0 0 0 REG_R1<4>
port 34 nsew
flabel metal3 -48 4120 -48 4120 7 FreeSans 48 0 0 0 REG_R1<5>
port 35 nsew
flabel metal3 -48 3380 -48 3380 7 FreeSans 48 0 0 0 REG_R1<6>
port 36 nsew
flabel metal3 -48 4760 -48 4760 7 FreeSans 48 0 0 0 REG_R1<7>
port 37 nsew
flabel metal3 -48 1300 -48 1300 7 FreeSans 48 0 0 0 REG_R1<8>
port 38 nsew
flabel metal3 -48 3300 -48 3300 7 FreeSans 48 0 0 0 REG_R1<9>
port 39 nsew
flabel metal3 -48 1520 -48 1520 7 FreeSans 48 0 0 0 REG_R1<10>
port 40 nsew
flabel metal3 -48 3340 -48 3340 7 FreeSans 48 0 0 0 REG_R1<11>
port 41 nsew
flabel metal3 -48 1700 -48 1700 7 FreeSans 48 0 0 0 REG_R1<12>
port 42 nsew
flabel metal2 592 -40 592 -40 7 FreeSans 48 270 0 0 REG_R1<13>
port 43 nsew
flabel metal3 -48 4400 -48 4400 7 FreeSans 48 0 0 0 REG_R1<14>
port 44 nsew
flabel metal3 -48 1340 -48 1340 7 FreeSans 48 0 0 0 REG_R1<15>
port 45 nsew
flabel metal3 8112 3180 8112 3180 3 FreeSans 48 0 0 0 REG_Write
port 46 nsew
flabel metal2 3712 -40 3712 -40 7 FreeSans 48 270 0 0 REG_Interrupt_flag
port 47 nsew
flabel metal2 1808 5660 1808 5660 3 FreeSans 48 90 0 0 clk
port 48 nsew
flabel space 3904 5660 3904 5660 3 FreeSans 48 90 0 0 rst
port 49 nsew
flabel metal2 3584 -40 3584 -40 7 FreeSans 48 270 0 0 REG_A<0>
port 50 nsew
flabel metal2 4704 -40 4704 -40 7 FreeSans 48 270 0 0 REG_A<1>
port 51 nsew
flabel metal3 -48 2320 -48 2320 7 FreeSans 48 0 0 0 REG_A<2>
port 52 nsew
flabel metal2 4192 5660 4192 5660 3 FreeSans 48 90 0 0 REG_A<3>
port 53 nsew
flabel metal2 3328 5660 3328 5660 3 FreeSans 48 90 0 0 REG_A<4>
port 54 nsew
flabel metal3 -48 3520 -48 3520 7 FreeSans 48 0 0 0 REG_A<5>
port 55 nsew
flabel metal2 2928 5660 2928 5660 3 FreeSans 48 90 0 0 REG_A<6>
port 56 nsew
flabel metal2 2880 5660 2880 5660 3 FreeSans 48 90 0 0 REG_A<7>
port 57 nsew
flabel metal2 3664 -40 3664 -40 7 FreeSans 48 270 0 0 REG_A<8>
port 58 nsew
flabel metal2 3184 5660 3184 5660 3 FreeSans 48 90 0 0 REG_A<9>
port 59 nsew
flabel metal2 3840 -40 3840 -40 7 FreeSans 48 270 0 0 REG_A<10>
port 60 nsew
flabel metal3 -48 3720 -48 3720 7 FreeSans 48 0 0 0 REG_A<11>
port 61 nsew
flabel metal2 4336 -40 4336 -40 7 FreeSans 48 270 0 0 REG_A<12>
port 62 nsew
flabel metal2 4192 -40 4192 -40 7 FreeSans 48 270 0 0 REG_A<13>
port 63 nsew
flabel metal2 4144 5660 4144 5660 3 FreeSans 48 90 0 0 REG_A<14>
port 64 nsew
flabel metal2 4096 -40 4096 -40 7 FreeSans 48 270 0 0 REG_A<15>
port 65 nsew
flabel metal2 3344 -40 3344 -40 7 FreeSans 48 270 0 0 REG_B<0>
port 66 nsew
flabel metal2 4432 -40 4432 -40 7 FreeSans 48 270 0 0 REG_B<1>
port 67 nsew
flabel metal2 2416 -40 2416 -40 7 FreeSans 48 270 0 0 REG_B<2>
port 68 nsew
flabel metal2 3936 5660 3936 5660 3 FreeSans 48 90 0 0 REG_B<3>
port 69 nsew
flabel metal2 3792 5660 3792 5660 3 FreeSans 48 90 0 0 REG_B<4>
port 70 nsew
flabel metal3 -48 3560 -48 3560 7 FreeSans 48 0 0 0 REG_B<5>
port 71 nsew
flabel metal2 3104 5660 3104 5660 3 FreeSans 48 90 0 0 REG_B<6>
port 72 nsew
flabel metal2 2976 5660 2976 5660 3 FreeSans 48 90 0 0 REG_B<7>
port 73 nsew
flabel metal2 4144 -40 4144 -40 7 FreeSans 48 270 0 0 REG_B<8>
port 74 nsew
flabel metal2 3024 5660 3024 5660 3 FreeSans 48 90 0 0 REG_B<9>
port 75 nsew
flabel metal2 4384 -40 4384 -40 7 FreeSans 48 270 0 0 REG_B<10>
port 76 nsew
flabel metal2 3232 5660 3232 5660 3 FreeSans 48 90 0 0 REG_B<11>
port 77 nsew
flabel metal2 4240 5660 4240 5660 3 FreeSans 48 90 0 0 REG_B<12>
port 78 nsew
flabel metal2 4240 -40 4240 -40 7 FreeSans 48 270 0 0 REG_B<13>
port 79 nsew
flabel metal2 3856 5660 3856 5660 3 FreeSans 48 90 0 0 REG_B<14>
port 80 nsew
flabel metal2 3792 -40 3792 -40 7 FreeSans 48 270 0 0 REG_B<15>
port 81 nsew
<< end >>
