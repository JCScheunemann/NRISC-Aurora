module NRISC_ULA (ULA_A, ULA_B, ULA_ctrl, ULA_OUT, ULA_flags);

input [15:0] ULA_A;
input [15:0] ULA_B;
input [3:0] ULA_ctrl;
output [15:0] ULA_OUT;
output [2:0] ULA_flags;

wire vdd = 1'b1;
wire gnd = 1'b0;

AND2X2 AND2X2_1 ( .A(ULA_A[15]), .B(ULA_B[15]), .Y(_455_) );
AND2X2 AND2X2_2 ( .A(_167_), .B(_129_), .Y(_518__2_) );
AND2X2 AND2X2_3 ( .A(_499_), .B(_500_), .Y(_501_) );
AND2X2 AND2X2_4 ( .A(_101_), .B(_487__bF_buf2), .Y(_231_) );
AND2X2 AND2X2_5 ( .A(ULA_B_0_bF_buf0), .B(ULA_B_1_bF_buf4), .Y(_502_) );
AND2X2 AND2X2_6 ( .A(_30_), .B(_32_), .Y(_33_) );
AND2X2 AND2X2_7 ( .A(_63_), .B(_486_), .Y(_518__0_) );
AND2X2 AND2X2_8 ( .A(_212_), .B(_491_), .Y(_224_) );
AND2X2 AND2X2_9 ( .A(ULA_A[5]), .B(ULA_B[5]), .Y(_237_) );
AND2X2 AND2X2_10 ( .A(_283_), .B(_491_), .Y(_295_) );
AND2X2 AND2X2_11 ( .A(_237_), .B(_491_), .Y(_249_) );
AND2X2 AND2X2_12 ( .A(_484__bF_buf2), .B(_457_), .Y(_459_) );
AND2X2 AND2X2_13 ( .A(ULA_A[6]), .B(ULA_B[6]), .Y(_261_) );
AND2X2 AND2X2_14 ( .A(_261_), .B(_491_), .Y(_272_) );
AND2X2 AND2X2_15 ( .A(ULA_A[7]), .B(ULA_B[7]), .Y(_283_) );
AND2X2 AND2X2_16 ( .A(_484__bF_buf3), .B(_309_), .Y(_310_) );
AND2X2 AND2X2_17 ( .A(_484__bF_buf1), .B(_336_), .Y(_337_) );
AND2X2 AND2X2_18 ( .A(_478_), .B(_480__bF_buf2), .Y(_481_) );
AND2X2 AND2X2_19 ( .A(_484__bF_buf3), .B(_354_), .Y(_355_) );
AND2X2 AND2X2_20 ( .A(ULA_A[12]), .B(ULA_B[12]), .Y(_392_) );
AND2X2 AND2X2_21 ( .A(ULA_A[13]), .B(ULA_B[13]), .Y(_411_) );
AND2X2 AND2X2_22 ( .A(ULA_ctrl[2]), .B(ULA_ctrl[1]), .Y(_446_) );
AND2X2 AND2X2_23 ( .A(ULA_ctrl[1]), .B(ULA_ctrl[3]), .Y(_482_) );
AOI21X1 AOI21X1_1 ( .A(ULA_ctrl_0_bF_buf4), .B(_420_), .C(_484__bF_buf3), .Y(_421_) );
AOI21X1 AOI21X1_2 ( .A(_314_), .B(_315_), .C(_487__bF_buf1), .Y(_386_) );
AOI21X1 AOI21X1_3 ( .A(_387_), .B(_381_), .C(_311_), .Y(_388_) );
AOI21X1 AOI21X1_4 ( .A(_258_), .B(_260_), .C(_269_), .Y(_270_) );
AOI21X1 AOI21X1_5 ( .A(_65_), .B(_478_), .C(_1_), .Y(_390_) );
AOI21X1 AOI21X1_6 ( .A(ULA_ctrl_0_bF_buf0), .B(_426_), .C(_484__bF_buf0), .Y(_485_) );
AOI21X1 AOI21X1_7 ( .A(_208_), .B(_304_), .C(_395_), .Y(_396_) );
AOI21X1 AOI21X1_8 ( .A(_22_), .B(_48_), .C(_210_), .Y(_211_) );
AOI21X1 AOI21X1_9 ( .A(ULA_ctrl_0_bF_buf2), .B(_398_), .C(_484__bF_buf0), .Y(_399_) );
AOI21X1 AOI21X1_10 ( .A(_365_), .B(ULA_B_1_bF_buf0), .C(_27_), .Y(_407_) );
AOI21X1 AOI21X1_11 ( .A(_402_), .B(_408_), .C(_311_), .Y(_409_) );
AOI21X1 AOI21X1_12 ( .A(ULA_ctrl_0_bF_buf3), .B(_339_), .C(_484__bF_buf0), .Y(_340_) );
AOI21X1 AOI21X1_13 ( .A(ULA_ctrl_0_bF_buf0), .B(_416_), .C(_484__bF_buf2), .Y(_417_) );
AOI21X1 AOI21X1_14 ( .A(_498_), .B(ULA_A[14]), .C(ULA_B_1_bF_buf4), .Y(_424_) );
AOI21X1 AOI21X1_15 ( .A(_481_), .B(_432_), .C(_436_), .Y(_437_) );
AOI21X1 AOI21X1_16 ( .A(_37_), .B(_282_), .C(_292_), .Y(_293_) );
AOI21X1 AOI21X1_17 ( .A(_442_), .B(_303_), .C(_440_), .Y(_443_) );
AOI21X1 AOI21X1_18 ( .A(ULA_B_1_bF_buf3), .B(_405_), .C(_175_), .Y(_449_) );
AOI21X1 AOI21X1_19 ( .A(_450_), .B(_38__bF_buf3), .C(ULA_B_2_bF_buf4), .Y(_451_) );
AOI21X1 AOI21X1_20 ( .A(ULA_ctrl_0_bF_buf2), .B(_461_), .C(_484__bF_buf1), .Y(_462_) );
AOI21X1 AOI21X1_21 ( .A(_486_), .B(_63_), .C(_518__3_), .Y(_466_) );
AOI21X1 AOI21X1_22 ( .A(_488_), .B(_22_), .C(_491_), .Y(_23_) );
AOI21X1 AOI21X1_23 ( .A(ULA_ctrl_0_bF_buf1), .B(_357_), .C(_484__bF_buf2), .Y(_358_) );
AOI21X1 AOI21X1_24 ( .A(_22_), .B(_45_), .C(_49_), .Y(_50_) );
AOI21X1 AOI21X1_25 ( .A(_51_), .B(_37_), .C(_61_), .Y(_62_) );
AOI21X1 AOI21X1_26 ( .A(_46_), .B(_105_), .C(_109_), .Y(_110_) );
AOI21X1 AOI21X1_27 ( .A(_117_), .B(_120_), .C(_67_), .Y(_121_) );
AOI21X1 AOI21X1_28 ( .A(_110_), .B(_104_), .C(_122_), .Y(_123_) );
AOI21X1 AOI21X1_29 ( .A(_46_), .B(_152_), .C(_155_), .Y(_156_) );
AOI21X1 AOI21X1_30 ( .A(_156_), .B(_150_), .C(_165_), .Y(_166_) );
AOI21X1 AOI21X1_31 ( .A(_38__bF_buf1), .B(_70_), .C(_185_), .Y(_186_) );
AOI21X1 AOI21X1_32 ( .A(_184_), .B(_190_), .C(_199_), .Y(_200_) );
AOI21X1 AOI21X1_33 ( .A(_1_), .B(_204_), .C(_205_), .Y(_206_) );
AOI21X1 AOI21X1_34 ( .A(_40_), .B(_39_), .C(ULA_B_2_bF_buf4), .Y(_208_) );
AOI21X1 AOI21X1_35 ( .A(_211_), .B(_209_), .C(_221_), .Y(_222_) );
AOI21X1 AOI21X1_36 ( .A(_232_), .B(ULA_B[3]), .C(_235_), .Y(_236_) );
AOI21X1 AOI21X1_37 ( .A(_236_), .B(_37_), .C(_246_), .Y(_247_) );
AOI21X1 AOI21X1_38 ( .A(_3_), .B(_424_), .C(_425_), .Y(_427_) );
AOI21X1 AOI21X1_39 ( .A(_147_), .B(_46_), .C(_259_), .Y(_260_) );
AOI21X1 AOI21X1_40 ( .A(_297_), .B(_298_), .C(_299_), .Y(_300_) );
AOI21X1 AOI21X1_41 ( .A(_314_), .B(_315_), .C(_27_), .Y(_316_) );
AOI21X1 AOI21X1_42 ( .A(ULA_ctrl_0_bF_buf0), .B(_321_), .C(_484__bF_buf2), .Y(_322_) );
AOI21X1 AOI21X1_43 ( .A(_167_), .B(_129_), .C(_518__1_), .Y(_471_) );
AOI21X1 AOI21X1_44 ( .A(_327_), .B(_328_), .C(_27_), .Y(_329_) );
AOI21X1 AOI21X1_45 ( .A(_183_), .B(_304_), .C(_374_), .Y(_375_) );
AOI21X1 AOI21X1_46 ( .A(_429_), .B(_423_), .C(_311_), .Y(_430_) );
AOI21X1 AOI21X1_47 ( .A(ULA_ctrl_0_bF_buf4), .B(_377_), .C(_484__bF_buf1), .Y(_378_) );
AOI21X1 AOI21X1_48 ( .A(ULA_ctrl_0_bF_buf3), .B(_127_), .C(_484__bF_buf2), .Y(_128_) );
AOI21X1 AOI21X1_49 ( .A(_383_), .B(_384_), .C(ULA_B_2_bF_buf0), .Y(_385_) );
AOI22X1 AOI22X1_1 ( .A(_458_), .B(_479_), .C(_420_), .D(_434_), .Y(_435_) );
AOI22X1 AOI22X1_2 ( .A(_446_), .B(_479_), .C(_447_), .D(_482_), .Y(_483_) );
AOI22X1 AOI22X1_3 ( .A(_67_), .B(_124_), .C(_123_), .D(_97_), .Y(_518__1_) );
AOI22X1 AOI22X1_4 ( .A(ULA_B_2_bF_buf1), .B(_175_), .C(_497_), .D(_176_), .Y(_177_) );
AOI22X1 AOI22X1_5 ( .A(_67_), .B(_201_), .C(_200_), .D(_179_), .Y(_518__3_) );
AOI22X1 AOI22X1_6 ( .A(ULA_B[3]), .B(_257_), .C(_22_), .D(_152_), .Y(_258_) );
AOI22X1 AOI22X1_7 ( .A(_490_), .B(_494_), .C(_24_), .D(_29_), .Y(_389_) );
AOI22X1 AOI22X1_8 ( .A(_406_), .B(_407_), .C(_46_), .D(_403_), .Y(_408_) );
AOI22X1 AOI22X1_9 ( .A(_410_), .B(_412_), .C(_304_), .D(_231_), .Y(_413_) );
BUFX4 BUFX4_1 ( .A(_487_), .Y(_487__bF_buf1) );
BUFX4 BUFX4_2 ( .A(_518__2_), .Y(_518__2_) );
BUFX4 BUFX4_3 ( .A(_518__3_), .Y(_518__3_) );
BUFX4 BUFX4_4 ( .A(_518__4_), .Y(_518__4_) );
BUFX4 BUFX4_5 ( .A(_518__5_), .Y(_518__5_) );
BUFX4 BUFX4_6 ( .A(_518__6_), .Y(_518__6_) );
BUFX4 BUFX4_7 ( .A(_518__7_), .Y(_518__7_) );
BUFX4 BUFX4_8 ( .A(_518__8_), .Y(_518__8_) );
BUFX4 BUFX4_9 ( .A(_518__9_), .Y(_518__9_) );
BUFX4 BUFX4_10 ( .A(_518__10_), .Y(_518__10_) );
BUFX4 BUFX4_11 ( .A(_518__11_), .Y(_518__11_) );
BUFX4 BUFX4_12 ( .A(_484_), .Y(_484__bF_buf0) );
BUFX4 BUFX4_13 ( .A(_518__12_), .Y(_518__12_) );
BUFX4 BUFX4_14 ( .A(_518__13_), .Y(_518__13_) );
BUFX4 BUFX4_15 ( .A(_484_), .Y(_484__bF_buf1) );
BUFX4 BUFX4_16 ( .A(_518__14_), .Y(_518__14_) );
BUFX4 BUFX4_17 ( .A(_518__15_), .Y(_518__15_) );
BUFX4 BUFX4_18 ( .A(_519__0_), .Y(_519__0_) );
BUFX4 BUFX4_19 ( .A(_519__1_), .Y(_519__1_) );
BUFX4 BUFX4_20 ( .A(_519__2_), .Y(_519__2_) );
BUFX2 BUFX2_1 ( .A(_518__0_), .Y(_518__0_) );
BUFX2 BUFX2_2 ( .A(_518__1_), .Y(_518__1_) );
BUFX4 BUFX4_21 ( .A(_480_), .Y(_480__bF_buf3) );
BUFX2 BUFX2_3 ( .A(_518__2_), .Y(_518__2_) );
BUFX2 BUFX2_4 ( .A(_518__3_), .Y(_518__3_) );
BUFX2 BUFX2_5 ( .A(_518__4_), .Y(_518__4_) );
BUFX2 BUFX2_6 ( .A(_518__5_), .Y(_518__5_) );
BUFX2 BUFX2_7 ( .A(_518__6_), .Y(_518__6_) );
BUFX2 BUFX2_8 ( .A(_518__7_), .Y(_518__7_) );
BUFX2 BUFX2_9 ( .A(_518__8_), .Y(_518__8_) );
BUFX2 BUFX2_10 ( .A(_518__9_), .Y(_518__9_) );
BUFX2 BUFX2_11 ( .A(_518__10_), .Y(_518__10_) );
BUFX2 BUFX2_12 ( .A(_518__11_), .Y(_518__11_) );
BUFX4 BUFX4_22 ( .A(_480_), .Y(_480__bF_buf2) );
BUFX2 BUFX2_13 ( .A(_518__12_), .Y(_518__12_) );
BUFX2 BUFX2_14 ( .A(_518__13_), .Y(_518__13_) );
BUFX2 BUFX2_15 ( .A(_518__14_), .Y(_518__14_) );
BUFX2 BUFX2_16 ( .A(_518__15_), .Y(_518__15_) );
BUFX2 BUFX2_17 ( .A(_519__0_), .Y(_519__0_) );
BUFX2 BUFX2_18 ( .A(_519__1_), .Y(_519__1_) );
BUFX2 BUFX2_19 ( .A(_519__2_), .Y(_519__2_) );
BUFX4 BUFX4_23 ( .A(_480_), .Y(_480__bF_buf1) );
BUFX4 BUFX4_24 ( .A(_480_), .Y(_480__bF_buf0) );
BUFX4 BUFX4_25 ( .A(_487_), .Y(_487__bF_buf0) );
BUFX4 BUFX4_26 ( .A(_518__0_), .Y(_518__0_) );
BUFX4 BUFX4_27 ( .A(_518__1_), .Y(_518__1_) );
BUFX4 BUFX4_28 ( .A(_518__15_), .Y(_518__15_) );
BUFX4 BUFX4_29 ( .A(_518__8_), .Y(_518__8_) );
BUFX4 BUFX4_30 ( .A(_484_), .Y(_484__bF_buf2) );
BUFX4 BUFX4_31 ( .A(_38_), .Y(_38__bF_buf4) );
BUFX4 BUFX4_32 ( .A(_38_), .Y(_38__bF_buf3) );
BUFX4 BUFX4_33 ( .A(_518__1_), .Y(_518__1_) );
BUFX4 BUFX4_34 ( .A(_38_), .Y(_38__bF_buf2) );
BUFX4 BUFX4_35 ( .A(_519__0_), .Y(_519__0_) );
BUFX4 BUFX4_36 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf5) );
BUFX4 BUFX4_37 ( .A(_38_), .Y(_38__bF_buf1) );
BUFX4 BUFX4_38 ( .A(_38_), .Y(_38__bF_buf0) );
BUFX4 BUFX4_39 ( .A(ULA_B[2]), .Y(ULA_B_2_bF_buf4) );
BUFX4 BUFX4_40 ( .A(_518__8_), .Y(_518__8_) );
BUFX4 BUFX4_41 ( .A(_518__2_), .Y(_518__2_) );
BUFX4 BUFX4_42 ( .A(_518__3_), .Y(_518__3_) );
BUFX4 BUFX4_43 ( .A(_519__1_), .Y(_519__1_) );
BUFX4 BUFX4_44 ( .A(_518__9_), .Y(_518__9_) );
BUFX4 BUFX4_45 ( .A(_518__10_), .Y(_518__10_) );
BUFX4 BUFX4_46 ( .A(_518__11_), .Y(_518__11_) );
BUFX4 BUFX4_47 ( .A(_518__12_), .Y(_518__12_) );
BUFX4 BUFX4_48 ( .A(_518__13_), .Y(_518__13_) );
BUFX4 BUFX4_49 ( .A(_518__14_), .Y(_518__14_) );
BUFX4 BUFX4_50 ( .A(_518__15_), .Y(_518__15_) );
BUFX4 BUFX4_51 ( .A(_519__0_), .Y(_519__0_) );
BUFX4 BUFX4_52 ( .A(_518__0_), .Y(_518__0_) );
BUFX4 BUFX4_53 ( .A(_518__9_), .Y(_518__9_) );
BUFX4 BUFX4_54 ( .A(_519__1_), .Y(_519__1_) );
BUFX4 BUFX4_55 ( .A(_519__2_), .Y(_519__2_) );
BUFX4 BUFX4_56 ( .A(_518__10_), .Y(_518__10_) );
BUFX4 BUFX4_57 ( .A(_518__11_), .Y(_518__11_) );
BUFX4 BUFX4_58 ( .A(_518__12_), .Y(_518__12_) );
BUFX4 BUFX4_59 ( .A(_518__13_), .Y(_518__13_) );
BUFX4 BUFX4_60 ( .A(_518__14_), .Y(_518__14_) );
BUFX4 BUFX4_61 ( .A(_518__1_), .Y(_518__1_) );
BUFX4 BUFX4_62 ( .A(_519__2_), .Y(_519__2_) );
BUFX4 BUFX4_63 ( .A(_518__1_), .Y(_518__1_) );
BUFX4 BUFX4_64 ( .A(_518__0_), .Y(_518__0_) );
BUFX4 BUFX4_65 ( .A(gnd), .Y(_519__0_) );
BUFX4 BUFX4_66 ( .A(_518__4_), .Y(_518__4_) );
BUFX4 BUFX4_67 ( .A(_518__5_), .Y(_518__5_) );
BUFX4 BUFX4_68 ( .A(_518__6_), .Y(_518__6_) );
BUFX4 BUFX4_69 ( .A(_518__7_), .Y(_518__7_) );
BUFX4 BUFX4_70 ( .A(_518__8_), .Y(_518__8_) );
BUFX4 BUFX4_71 ( .A(_518__9_), .Y(_518__9_) );
BUFX4 BUFX4_72 ( .A(_518__10_), .Y(_518__10_) );
BUFX4 BUFX4_73 ( .A(_518__2_), .Y(_518__2_) );
BUFX4 BUFX4_74 ( .A(_518__2_), .Y(_518__2_) );
BUFX4 BUFX4_75 ( .A(_518__10_), .Y(_518__10_) );
BUFX4 BUFX4_76 ( .A(_518__11_), .Y(_518__11_) );
BUFX4 BUFX4_77 ( .A(_518__3_), .Y(_518__3_) );
BUFX4 BUFX4_78 ( .A(zero), .Y(_519__1_) );
BUFX4 BUFX4_79 ( .A(_518__12_), .Y(_518__12_) );
BUFX4 BUFX4_80 ( .A(_518__13_), .Y(_518__13_) );
BUFX4 BUFX4_81 ( .A(_518__14_), .Y(_518__14_) );
BUFX4 BUFX4_82 ( .A(_518__15_), .Y(_518__15_) );
BUFX4 BUFX4_83 ( .A(_519__0_), .Y(_519__0_) );
BUFX4 BUFX4_84 ( .A(_519__1_), .Y(_519__1_) );
BUFX4 BUFX4_85 ( .A(_518__3_), .Y(_518__3_) );
BUFX4 BUFX4_86 ( .A(_518__3_), .Y(_518__3_) );
BUFX4 BUFX4_87 ( .A(_519__2_), .Y(_519__2_) );
BUFX4 BUFX4_88 ( .A(_518__4_), .Y(_518__4_) );
BUFX4 BUFX4_89 ( .A(_518__5_), .Y(_518__5_) );
BUFX4 BUFX4_90 ( .A(_518__6_), .Y(_518__6_) );
BUFX4 BUFX4_91 ( .A(_518__1_), .Y(_518__1_) );
BUFX4 BUFX4_92 ( .A(_518__7_), .Y(_518__7_) );
BUFX4 BUFX4_93 ( .A(_518__8_), .Y(_518__8_) );
BUFX4 BUFX4_94 ( .A(_518__11_), .Y(_518__11_) );
BUFX4 BUFX4_95 ( .A(_518__12_), .Y(_518__12_) );
BUFX4 BUFX4_96 ( .A(_518__4_), .Y(_518__4_) );
BUFX4 BUFX4_97 ( .A(_518__13_), .Y(_518__13_) );
BUFX4 BUFX4_98 ( .A(_518__4_), .Y(_518__4_) );
BUFX4 BUFX4_99 ( .A(_518__14_), .Y(_518__14_) );
BUFX4 BUFX4_100 ( .A(_518__15_), .Y(_518__15_) );
BUFX4 BUFX4_101 ( .A(_518__0_), .Y(_518__0_) );
BUFX4 BUFX4_102 ( .A(ULA_B[2]), .Y(ULA_B_2_bF_buf3) );
BUFX4 BUFX4_103 ( .A(ULA_B[2]), .Y(ULA_B_2_bF_buf2) );
BUFX4 BUFX4_104 ( .A(_undef), .Y(_519__2_) );
BUFX4 BUFX4_105 ( .A(ULA_B[2]), .Y(ULA_B_2_bF_buf1) );
BUFX4 BUFX4_106 ( .A(ULA_B[2]), .Y(ULA_B_2_bF_buf0) );
BUFX4 BUFX4_107 ( .A(_518__5_), .Y(_518__5_) );
BUFX4 BUFX4_108 ( .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf2) );
BUFX4 BUFX4_109 ( .A(_504_), .Y(_504__bF_buf4) );
BUFX4 BUFX4_110 ( .A(_518__5_), .Y(_518__5_) );
BUFX4 BUFX4_111 ( .A(_504_), .Y(_504__bF_buf3) );
BUFX4 BUFX4_112 ( .A(_504_), .Y(_504__bF_buf2) );
BUFX4 BUFX4_113 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf4) );
BUFX4 BUFX4_114 ( .A(_504_), .Y(_504__bF_buf1) );
BUFX4 BUFX4_115 ( .A(_518__2_), .Y(_518__2_) );
BUFX4 BUFX4_116 ( .A(_504_), .Y(_504__bF_buf0) );
BUFX4 BUFX4_117 ( .A(_518__9_), .Y(_518__9_) );
BUFX4 BUFX4_118 ( .A(_518__6_), .Y(_518__6_) );
BUFX4 BUFX4_119 ( .A(ULA_B[1]), .Y(ULA_B_1_bF_buf4) );
BUFX4 BUFX4_120 ( .A(ULA_B[1]), .Y(ULA_B_1_bF_buf3) );
BUFX4 BUFX4_121 ( .A(ULA_B[1]), .Y(ULA_B_1_bF_buf2) );
BUFX4 BUFX4_122 ( .A(_518__6_), .Y(_518__6_) );
BUFX4 BUFX4_123 ( .A(ULA_B[1]), .Y(ULA_B_1_bF_buf1) );
BUFX4 BUFX4_124 ( .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf1) );
BUFX4 BUFX4_125 ( .A(ULA_B[1]), .Y(ULA_B_1_bF_buf0) );
BUFX4 BUFX4_126 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf3) );
BUFX4 BUFX4_127 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf2) );
BUFX4 BUFX4_128 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf1) );
BUFX4 BUFX4_129 ( .A(_518__7_), .Y(_518__7_) );
BUFX4 BUFX4_130 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf6) );
BUFX4 BUFX4_131 ( .A(_518__0_), .Y(_518__0_) );
BUFX4 BUFX4_132 ( .A(ULA_B[0]), .Y(ULA_B_0_bF_buf0) );
BUFX4 BUFX4_133 ( .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf4) );
BUFX4 BUFX4_134 ( .A(_518__7_), .Y(_518__7_) );
BUFX4 BUFX4_135 ( .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf3) );
BUFX4 BUFX4_136 ( .A(ULA_ctrl[0]), .Y(ULA_ctrl_0_bF_buf0) );
BUFX4 BUFX4_137 ( .A(_487_), .Y(_487__bF_buf3) );
BUFX4 BUFX4_138 ( .A(_487_), .Y(_487__bF_buf2) );
BUFX4 BUFX4_139 ( .A(_484_), .Y(_484__bF_buf3) );
INVX1 INVX1_1 ( .A(_66_), .Y(_432_) );
INVX1 INVX1_2 ( .A(_231_), .Y(_232_) );
INVX1 INVX1_3 ( .A(_37_), .Y(_259_) );
INVX2 INVX2_1 ( .A(_119_), .Y(_120_) );
INVX1 INVX1_4 ( .A(ULA_A[6]), .Y(_513_) );
INVX1 INVX1_5 ( .A(ULA_B[8]), .Y(_306_) );
INVX2 INVX2_2 ( .A(_311_), .Y(_312_) );
INVX2 INVX2_3 ( .A(ULA_A[9]), .Y(_86_) );
INVX1 INVX1_6 ( .A(_307_), .Y(_321_) );
INVX1 INVX1_7 ( .A(ULA_B[9]), .Y(_333_) );
INVX1 INVX1_8 ( .A(_478_), .Y(_441_) );
INVX1 INVX1_9 ( .A(ULA_A[0]), .Y(_157_) );
INVX1 INVX1_10 ( .A(_334_), .Y(_339_) );
INVX1 INVX1_11 ( .A(_52_), .Y(_434_) );
INVX1 INVX1_12 ( .A(ULA_B[10]), .Y(_351_) );
INVX1 INVX1_13 ( .A(ULA_A[2]), .Y(_125_) );
INVX1 INVX1_14 ( .A(_352_), .Y(_357_) );
INVX1 INVX1_15 ( .A(ULA_A[12]), .Y(_2_) );
INVX1 INVX1_16 ( .A(ULA_B[11]), .Y(_370_) );
INVX1 INVX1_17 ( .A(_371_), .Y(_377_) );
INVX2 INVX2_4 ( .A(ULA_A[4]), .Y(_509_) );
INVX1 INVX1_18 ( .A(_392_), .Y(_398_) );
INVX1 INVX1_19 ( .A(_79_), .Y(_170_) );
INVX1 INVX1_20 ( .A(_455_), .Y(_461_) );
INVX1 INVX1_21 ( .A(ULA_A[13]), .Y(_404_) );
INVX1 INVX1_22 ( .A(_411_), .Y(_416_) );
INVX1 INVX1_23 ( .A(_4_), .Y(_5_) );
INVX2 INVX2_5 ( .A(ULA_A[10]), .Y(_15_) );
INVX1 INVX1_24 ( .A(_35_), .Y(_36_) );
INVX1 INVX1_25 ( .A(_467_), .Y(_469_) );
INVX2 INVX2_6 ( .A(ULA_ctrl[1]), .Y(_477_) );
INVX1 INVX1_26 ( .A(ULA_A[14]), .Y(_6_) );
INVX2 INVX2_7 ( .A(ULA_A[8]), .Y(_11_) );
INVX1 INVX1_27 ( .A(ULA_A[7]), .Y(_77_) );
INVX1 INVX1_28 ( .A(_88_), .Y(_89_) );
INVX1 INVX1_29 ( .A(_13_), .Y(_14_) );
INVX1 INVX1_30 ( .A(_426_), .Y(_53_) );
INVX1 INVX1_31 ( .A(_57_), .Y(_58_) );
INVX1 INVX1_32 ( .A(ULA_A[5]), .Y(_73_) );
INVX1 INVX1_33 ( .A(_126_), .Y(_127_) );
INVX1 INVX1_34 ( .A(_75_), .Y(_76_) );
INVX1 INVX1_35 ( .A(ULA_A[11]), .Y(_90_) );
INVX1 INVX1_36 ( .A(_70_), .Y(_107_) );
INVX1 INVX1_37 ( .A(ULA_A[1]), .Y(_111_) );
INVX1 INVX1_38 ( .A(_274_), .Y(_440_) );
INVX1 INVX1_39 ( .A(_116_), .Y(_117_) );
INVX1 INVX1_40 ( .A(_495_), .Y(_130_) );
INVX1 INVX1_41 ( .A(_511_), .Y(_512_) );
INVX1 INVX1_42 ( .A(_515_), .Y(_133_) );
INVX1 INVX1_43 ( .A(_17_), .Y(_140_) );
INVX1 INVX1_44 ( .A(ULA_A[15]), .Y(_174_) );
INVX1 INVX1_45 ( .A(_175_), .Y(_180_) );
INVX1 INVX1_46 ( .A(ULA_B[4]), .Y(_25_) );
INVX1 INVX1_47 ( .A(_19_), .Y(_204_) );
INVX2 INVX2_8 ( .A(ULA_ctrl[3]), .Y(_479_) );
INVX2 INVX2_9 ( .A(ULA_B_0_bF_buf2), .Y(_498_) );
INVX2 INVX2_10 ( .A(ULA_A[3]), .Y(_505_) );
INVX4 INVX4_1 ( .A(_303_), .Y(_304_) );
INVX4 INVX4_2 ( .A(ULA_ctrl[2]), .Y(_447_) );
INVX4 INVX4_3 ( .A(ULA_ctrl_0_bF_buf2), .Y(_491_) );
INVX8 INVX8_1 ( .A(ULA_B[3]), .Y(_492_) );
INVX4 INVX4_4 ( .A(_46_), .Y(_47_) );
INVX8 INVX8_2 ( .A(_439_), .Y(_518__14_) );
INVX8 INVX8_3 ( .A(_464_), .Y(_518__15_) );
INVX8 INVX8_4 ( .A(ULA_B_2_bF_buf2), .Y(_487_) );
INVX8 INVX8_5 ( .A(ULA_B_1_bF_buf1), .Y(_38_) );
INVX8 INVX8_6 ( .A(_324_), .Y(_518__8_) );
INVX8 INVX8_7 ( .A(_342_), .Y(_518__9_) );
INVX8 INVX8_8 ( .A(_360_), .Y(_518__10_) );
INVX8 INVX8_9 ( .A(_380_), .Y(_518__11_) );
INVX8 INVX8_10 ( .A(_401_), .Y(_518__12_) );
INVX8 INVX8_11 ( .A(_419_), .Y(_518__13_) );
MUX2X1 MUX2X1_1 ( .A(_507_), .B(_501_), .S(_504__bF_buf4), .Y(_508_) );
MUX2X1 MUX2X1_2 ( .A(_217_), .B(_159_), .S(_38__bF_buf4), .Y(_218_) );
MUX2X1 MUX2X1_3 ( .A(_242_), .B(_192_), .S(_38__bF_buf2), .Y(_243_) );
MUX2X1 MUX2X1_4 ( .A(ULA_A[2]), .B(ULA_A[1]), .S(ULA_B_0_bF_buf4), .Y(_68_) );
MUX2X1 MUX2X1_5 ( .A(_265_), .B(_217_), .S(_38__bF_buf1), .Y(_266_) );
MUX2X1 MUX2X1_6 ( .A(_345_), .B(_313_), .S(_38__bF_buf0), .Y(_346_) );
MUX2X1 MUX2X1_7 ( .A(_94_), .B(_85_), .S(_497_), .Y(_95_) );
MUX2X1 MUX2X1_8 ( .A(ULA_A[10]), .B(ULA_A[11]), .S(ULA_B_0_bF_buf4), .Y(_365_) );
MUX2X1 MUX2X1_9 ( .A(_10_), .B(_19_), .S(_1_), .Y(_20_) );
MUX2X1 MUX2X1_10 ( .A(_0_), .B(_20_), .S(_495_), .Y(_21_) );
MUX2X1 MUX2X1_11 ( .A(_501_), .B(_507_), .S(_38__bF_buf1), .Y(_45_) );
MUX2X1 MUX2X1_12 ( .A(ULA_A[15]), .B(ULA_A[14]), .S(ULA_B_0_bF_buf4), .Y(_138_) );
MUX2X1 MUX2X1_13 ( .A(_515_), .B(_511_), .S(ULA_B_1_bF_buf2), .Y(_48_) );
MUX2X1 MUX2X1_14 ( .A(_81_), .B(_72_), .S(_1_), .Y(_82_) );
MUX2X1 MUX2X1_15 ( .A(_84_), .B(_98_), .S(_504__bF_buf4), .Y(_176_) );
MUX2X1 MUX2X1_16 ( .A(ULA_A[14]), .B(ULA_A[13]), .S(ULA_B_0_bF_buf4), .Y(_84_) );
MUX2X1 MUX2X1_17 ( .A(_82_), .B(_95_), .S(_495_), .Y(_96_) );
MUX2X1 MUX2X1_18 ( .A(ULA_A[12]), .B(ULA_A[11]), .S(ULA_B_0_bF_buf6), .Y(_98_) );
MUX2X1 MUX2X1_19 ( .A(_79_), .B(_75_), .S(ULA_B_1_bF_buf2), .Y(_105_) );
MUX2X1 MUX2X1_20 ( .A(_135_), .B(_132_), .S(_1_), .Y(_136_) );
MUX2X1 MUX2X1_21 ( .A(_17_), .B(_4_), .S(_38__bF_buf2), .Y(_147_) );
MUX2X1 MUX2X1_22 ( .A(ULA_A[4]), .B(ULA_A[5]), .S(ULA_B_0_bF_buf2), .Y(_287_) );
MUX2X1 MUX2X1_23 ( .A(_172_), .B(_169_), .S(_1_), .Y(_173_) );
MUX2X1 MUX2X1_24 ( .A(_173_), .B(_177_), .S(_495_), .Y(_178_) );
MUX2X1 MUX2X1_25 ( .A(_508_), .B(_517_), .S(_497_), .Y(_0_) );
MUX2X1 MUX2X1_26 ( .A(_98_), .B(_84_), .S(_38__bF_buf3), .Y(_181_) );
MUX2X1 MUX2X1_27 ( .A(_192_), .B(_115_), .S(_38__bF_buf0), .Y(_193_) );
NAND2X1 NAND2X1_1 ( .A(_390_), .B(_389_), .Y(_431_) );
NAND2X1 NAND2X1_2 ( .A(_487__bF_buf1), .B(_364_), .Y(_444_) );
NAND2X1 NAND2X1_3 ( .A(_38__bF_buf3), .B(_13_), .Y(_301_) );
NAND2X1 NAND2X1_4 ( .A(ULA_B_0_bF_buf2), .B(ULA_A[7]), .Y(_514_) );
NAND2X1 NAND2X1_5 ( .A(_57_), .B(_35_), .Y(_303_) );
NAND2X1 NAND2X1_6 ( .A(_478_), .B(_480__bF_buf0), .Y(_64_) );
NAND2X1 NAND2X1_7 ( .A(ULA_B_0_bF_buf3), .B(ULA_A[4]), .Y(_69_) );
NAND2X1 NAND2X1_8 ( .A(_391_), .B(_396_), .Y(_397_) );
NAND2X1 NAND2X1_9 ( .A(_70_), .B(_504__bF_buf2), .Y(_71_) );
NAND2X1 NAND2X1_10 ( .A(ULA_B_0_bF_buf1), .B(ULA_A[1]), .Y(_500_) );
NAND2X1 NAND2X1_11 ( .A(ULA_B_0_bF_buf1), .B(ULA_A[6]), .Y(_74_) );
NAND2X1 NAND2X1_12 ( .A(ULA_B_0_bF_buf6), .B(ULA_A[8]), .Y(_78_) );
NAND2X1 NAND2X1_13 ( .A(_369_), .B(_375_), .Y(_376_) );
NAND2X1 NAND2X1_14 ( .A(_79_), .B(_504__bF_buf0), .Y(_80_) );
NAND2X1 NAND2X1_15 ( .A(_515_), .B(_504__bF_buf3), .Y(_516_) );
NAND2X1 NAND2X1_16 ( .A(ULA_B_0_bF_buf3), .B(ULA_A[10]), .Y(_87_) );
NAND2X1 NAND2X1_17 ( .A(ULA_B_0_bF_buf1), .B(ULA_A[12]), .Y(_91_) );
NAND2X1 NAND2X1_18 ( .A(_304_), .B(_103_), .Y(_332_) );
NAND2X1 NAND2X1_19 ( .A(_92_), .B(_504__bF_buf2), .Y(_93_) );
NAND2X1 NAND2X1_20 ( .A(ULA_B_2_bF_buf3), .B(_367_), .Y(_453_) );
NAND2X1 NAND2X1_21 ( .A(_33_), .B(_96_), .Y(_97_) );
NAND2X1 NAND2X1_22 ( .A(ULA_B_1_bF_buf2), .B(_265_), .Y(_315_) );
NAND2X1 NAND2X1_23 ( .A(ULA_B_1_bF_buf0), .B(_98_), .Y(_99_) );
NAND2X1 NAND2X1_24 ( .A(_327_), .B(_328_), .Y(_403_) );
NAND2X1 NAND2X1_25 ( .A(ULA_B_2_bF_buf0), .B(_101_), .Y(_102_) );
NAND2X1 NAND2X1_26 ( .A(_25_), .B(_118_), .Y(_311_) );
NAND2X1 NAND2X1_27 ( .A(_57_), .B(_118_), .Y(_119_) );
NAND2X1 NAND2X1_28 ( .A(_38__bF_buf2), .B(_382_), .Y(_383_) );
NAND2X1 NAND2X1_29 ( .A(_114_), .B(_121_), .Y(_122_) );
NAND2X1 NAND2X1_30 ( .A(_511_), .B(_504__bF_buf0), .Y(_131_) );
NAND2X1 NAND2X1_31 ( .A(ULA_B_1_bF_buf4), .B(_287_), .Y(_363_) );
NAND2X1 NAND2X1_32 ( .A(_13_), .B(_504__bF_buf3), .Y(_134_) );
NAND2X1 NAND2X1_33 ( .A(_4_), .B(_504__bF_buf0), .Y(_141_) );
NAND2X1 NAND2X1_34 ( .A(_38__bF_buf1), .B(_326_), .Y(_327_) );
NAND2X1 NAND2X1_35 ( .A(_487__bF_buf3), .B(_147_), .Y(_148_) );
NAND2X1 NAND2X1_36 ( .A(ULA_B[3]), .B(_149_), .Y(_150_) );
NAND2X1 NAND2X1_37 ( .A(ULA_A[0]), .B(_498_), .Y(_499_) );
NAND2X1 NAND2X1_38 ( .A(_464_), .B(_360_), .Y(_473_) );
NAND2X1 NAND2X1_39 ( .A(_38__bF_buf1), .B(_133_), .Y(_151_) );
NAND2X1 NAND2X1_40 ( .A(ULA_A[14]), .B(ULA_B[14]), .Y(_420_) );
NAND2X1 NAND2X1_41 ( .A(_161_), .B(_120_), .Y(_162_) );
NAND2X1 NAND2X1_42 ( .A(ULA_B_1_bF_buf2), .B(_345_), .Y(_384_) );
NAND2X1 NAND2X1_43 ( .A(_166_), .B(_145_), .Y(_167_) );
NAND2X1 NAND2X1_44 ( .A(_38__bF_buf4), .B(_365_), .Y(_366_) );
NAND2X1 NAND2X1_45 ( .A(_75_), .B(_504__bF_buf3), .Y(_168_) );
NAND2X1 NAND2X1_46 ( .A(ULA_B_1_bF_buf1), .B(_288_), .Y(_328_) );
NAND2X1 NAND2X1_47 ( .A(_88_), .B(_504__bF_buf1), .Y(_171_) );
NAND2X1 NAND2X1_48 ( .A(_38__bF_buf2), .B(_313_), .Y(_314_) );
NAND2X1 NAND2X1_49 ( .A(_33_), .B(_178_), .Y(_179_) );
NAND2X1 NAND2X1_50 ( .A(_487__bF_buf1), .B(_181_), .Y(_182_) );
NAND2X1 NAND2X1_51 ( .A(ULA_B_1_bF_buf0), .B(_88_), .Y(_187_) );
NAND2X1 NAND2X1_52 ( .A(ULA_B_0_bF_buf1), .B(ULA_A[2]), .Y(_191_) );
NAND2X1 NAND2X1_53 ( .A(_120_), .B(_194_), .Y(_195_) );
NAND2X1 NAND2X1_54 ( .A(ULA_A[0]), .B(ULA_B_0_bF_buf6), .Y(_426_) );
NAND2X1 NAND2X1_55 ( .A(ULA_B_1_bF_buf3), .B(_491_), .Y(_503_) );
NAND2X1 NAND2X1_56 ( .A(ULA_B_0_bF_buf0), .B(ULA_A[13]), .Y(_3_) );
NAND2X1 NAND2X1_57 ( .A(ULA_B_0_bF_buf1), .B(ULA_A[11]), .Y(_16_) );
NAND2X1 NAND2X1_58 ( .A(_24_), .B(_29_), .Y(_30_) );
NAND2X1 NAND2X1_59 ( .A(ULA_B_1_bF_buf0), .B(_8_), .Y(_40_) );
NAND2X1 NAND2X1_60 ( .A(_497_), .B(_10_), .Y(_202_) );
NAND2X1 NAND2X1_61 ( .A(ULA_B_0_bF_buf6), .B(ULA_A[3]), .Y(_216_) );
NAND2X1 NAND2X1_62 ( .A(_487__bF_buf3), .B(_218_), .Y(_219_) );
NAND2X1 NAND2X1_63 ( .A(_215_), .B(_219_), .Y(_220_) );
NAND2X1 NAND2X1_64 ( .A(_497_), .B(_85_), .Y(_226_) );
NAND2X1 NAND2X1_65 ( .A(_33_), .B(_229_), .Y(_230_) );
NAND2X1 NAND2X1_66 ( .A(_22_), .B(_105_), .Y(_233_) );
NAND2X1 NAND2X1_67 ( .A(_46_), .B(_100_), .Y(_234_) );
NAND2X1 NAND2X1_68 ( .A(_233_), .B(_234_), .Y(_235_) );
NAND2X1 NAND2X1_69 ( .A(_38__bF_buf3), .B(_115_), .Y(_240_) );
NAND2X1 NAND2X1_70 ( .A(ULA_B_1_bF_buf4), .B(_17_), .Y(_42_) );
NAND2X1 NAND2X1_71 ( .A(ULA_ctrl[1]), .B(ULA_ctrl[3]), .Y(_31_) );
NAND2X1 NAND2X1_72 ( .A(_17_), .B(_504__bF_buf4), .Y(_18_) );
NAND2X1 NAND2X1_73 ( .A(ULA_B_0_bF_buf5), .B(ULA_A[15]), .Y(_7_) );
NAND2X1 NAND2X1_74 ( .A(ULA_B_0_bF_buf6), .B(_505_), .Y(_506_) );
NAND2X1 NAND2X1_75 ( .A(_487__bF_buf0), .B(_488_), .Y(_489_) );
NAND2X1 NAND2X1_76 ( .A(ULA_B_2_bF_buf2), .B(_240_), .Y(_241_) );
NAND2X1 NAND2X1_77 ( .A(_487__bF_buf1), .B(_243_), .Y(_244_) );
NAND2X1 NAND2X1_78 ( .A(_241_), .B(_244_), .Y(_245_) );
NAND2X1 NAND2X1_79 ( .A(_497_), .B(_130_), .Y(_252_) );
NAND2X1 NAND2X1_80 ( .A(_33_), .B(_255_), .Y(_256_) );
NAND2X1 NAND2X1_81 ( .A(_451_), .B(_449_), .Y(_452_) );
NAND2X1 NAND2X1_82 ( .A(_487__bF_buf0), .B(_146_), .Y(_257_) );
NAND2X1 NAND2X1_83 ( .A(_33_), .B(_21_), .Y(_34_) );
NAND2X1 NAND2X1_84 ( .A(ULA_B_2_bF_buf1), .B(_160_), .Y(_264_) );
NAND2X1 NAND2X1_85 ( .A(ULA_B[4]), .B(_23_), .Y(_24_) );
NAND2X1 NAND2X1_86 ( .A(_487__bF_buf3), .B(_266_), .Y(_267_) );
NAND2X1 NAND2X1_87 ( .A(_8_), .B(_504__bF_buf1), .Y(_9_) );
NAND2X1 NAND2X1_88 ( .A(_264_), .B(_267_), .Y(_268_) );
NAND2X1 NAND2X1_89 ( .A(ULA_B_0_bF_buf4), .B(ULA_A[5]), .Y(_510_) );
NAND2X1 NAND2X1_90 ( .A(ULA_B[3]), .B(_274_), .Y(_275_) );
NAND2X1 NAND2X1_91 ( .A(_494_), .B(_490_), .Y(_495_) );
NAND2X1 NAND2X1_92 ( .A(_62_), .B(_34_), .Y(_63_) );
NAND2X1 NAND2X1_93 ( .A(_33_), .B(_278_), .Y(_279_) );
NAND2X1 NAND2X1_94 ( .A(_22_), .B(_188_), .Y(_280_) );
NAND2X1 NAND2X1_95 ( .A(_38__bF_buf2), .B(_4_), .Y(_39_) );
NAND2X1 NAND2X1_96 ( .A(_46_), .B(_181_), .Y(_281_) );
NAND2X1 NAND2X1_97 ( .A(ULA_B_2_bF_buf0), .B(_193_), .Y(_286_) );
NAND2X1 NAND2X1_98 ( .A(_25_), .B(_28_), .Y(_29_) );
NAND2X1 NAND2X1_99 ( .A(_38__bF_buf0), .B(_288_), .Y(_289_) );
NAND2X1 NAND2X1_100 ( .A(_1_), .B(_10_), .Y(_297_) );
NAND2X1 NAND2X1_101 ( .A(ULA_B_0_bF_buf3), .B(ULA_A[9]), .Y(_12_) );
NAND2X1 NAND2X1_102 ( .A(_497_), .B(_19_), .Y(_298_) );
NAND3X1 NAND3X1_1 ( .A(ULA_B[3]), .B(_264_), .C(_267_), .Y(_423_) );
NAND3X1 NAND3X1_2 ( .A(_484__bF_buf3), .B(_413_), .C(_414_), .Y(_415_) );
NAND3X1 NAND3X1_3 ( .A(_459_), .B(_454_), .C(_448_), .Y(_460_) );
NAND3X1 NAND3X1_4 ( .A(_487__bF_buf2), .B(_301_), .C(_42_), .Y(_302_) );
NAND3X1 NAND3X1_5 ( .A(_342_), .B(_439_), .C(_380_), .Y(_467_) );
NAND3X1 NAND3X1_6 ( .A(_483_), .B(_468_), .C(_481_), .Y(_484_) );
NAND3X1 NAND3X1_7 ( .A(_465_), .B(_466_), .C(_469_), .Y(_470_) );
NAND3X1 NAND3X1_8 ( .A(_250_), .B(_230_), .C(_247_), .Y(_518__5_) );
NAND3X1 NAND3X1_9 ( .A(_324_), .B(_401_), .C(_419_), .Y(_474_) );
NAND3X1 NAND3X1_10 ( .A(_471_), .B(_472_), .C(_475_), .Y(_476_) );
NAND3X1 NAND3X1_11 ( .A(ULA_ctrl_0_bF_buf3), .B(ULA_B[3]), .C(_489_), .Y(_490_) );
NAND3X1 NAND3X1_12 ( .A(_350_), .B(_355_), .C(_348_), .Y(_356_) );
NAND3X1 NAND3X1_13 ( .A(ULA_B_2_bF_buf2), .B(_39_), .C(_40_), .Y(_41_) );
NAND3X1 NAND3X1_14 ( .A(_441_), .B(_495_), .C(_30_), .Y(_442_) );
NAND3X1 NAND3X1_15 ( .A(ULA_ctrl[2]), .B(ULA_ctrl[1]), .C(_479_), .Y(_52_) );
NAND3X1 NAND3X1_16 ( .A(_304_), .B(_41_), .C(_302_), .Y(_305_) );
NAND3X1 NAND3X1_17 ( .A(ULA_ctrl[2]), .B(ULA_ctrl[3]), .C(_477_), .Y(_56_) );
NAND3X1 NAND3X1_18 ( .A(ULA_A[0]), .B(_493_), .C(_59_), .Y(_60_) );
NAND3X1 NAND3X1_19 ( .A(_65_), .B(_56_), .C(_483_), .Y(_66_) );
NAND3X1 NAND3X1_20 ( .A(ULA_B_1_bF_buf1), .B(ULA_A[15]), .C(_498_), .Y(_83_) );
NAND3X1 NAND3X1_21 ( .A(ULA_ctrl[3]), .B(_447_), .C(_477_), .Y(_478_) );
NAND3X1 NAND3X1_22 ( .A(_38__bF_buf3), .B(_487__bF_buf1), .C(_115_), .Y(_116_) );
NAND3X1 NAND3X1_23 ( .A(ULA_B[3]), .B(_215_), .C(_219_), .Y(_381_) );
NAND3X1 NAND3X1_24 ( .A(_484__bF_buf1), .B(_164_), .C(_162_), .Y(_165_) );
NAND3X1 NAND3X1_25 ( .A(_484__bF_buf0), .B(_198_), .C(_195_), .Y(_199_) );
NAND3X1 NAND3X1_26 ( .A(_270_), .B(_273_), .C(_256_), .Y(_518__6_) );
NAND3X1 NAND3X1_27 ( .A(_275_), .B(_281_), .C(_280_), .Y(_282_) );
NAND3X1 NAND3X1_28 ( .A(_55_), .B(_60_), .C(_484__bF_buf3), .Y(_61_) );
NAND3X1 NAND3X1_29 ( .A(_296_), .B(_293_), .C(_279_), .Y(_518__7_) );
NAND3X1 NAND3X1_30 ( .A(_286_), .B(_444_), .C(_445_), .Y(_448_) );
NAND3X1 NAND3X1_31 ( .A(_495_), .B(_32_), .C(_30_), .Y(_299_) );
NAND3X1 NAND3X1_32 ( .A(ULA_A[0]), .B(ULA_B[3]), .C(_493_), .Y(_317_) );
NAND3X1 NAND3X1_33 ( .A(_305_), .B(_310_), .C(_319_), .Y(_320_) );
NAND3X1 NAND3X1_34 ( .A(_222_), .B(_225_), .C(_207_), .Y(_518__4_) );
NAND3X1 NAND3X1_35 ( .A(_337_), .B(_331_), .C(_332_), .Y(_338_) );
NAND3X1 NAND3X1_36 ( .A(ULA_ctrl[2]), .B(_477_), .C(_479_), .Y(_480_) );
NAND3X1 NAND3X1_37 ( .A(_349_), .B(_304_), .C(_148_), .Y(_350_) );
NAND3X1 NAND3X1_38 ( .A(_10_), .B(_390_), .C(_389_), .Y(_391_) );
NAND3X1 NAND3X1_39 ( .A(_120_), .B(_452_), .C(_453_), .Y(_454_) );
NAND3X1 NAND3X1_40 ( .A(ULA_B[3]), .B(_241_), .C(_244_), .Y(_402_) );
NAND3X1 NAND3X1_41 ( .A(ULA_ctrl[2]), .B(ULA_ctrl[1]), .C(ULA_ctrl[3]), .Y(_65_) );
NAND3X1 NAND3X1_42 ( .A(_85_), .B(_390_), .C(_389_), .Y(_414_) );
NOR2X1 NOR2X1_1 ( .A(_487__bF_buf2), .B(_346_), .Y(_428_) );
NOR2X1 NOR2X1_2 ( .A(_299_), .B(_95_), .Y(_325_) );
NOR2X1 NOR2X1_3 ( .A(_86_), .B(_333_), .Y(_334_) );
NOR2X1 NOR2X1_4 ( .A(_495_), .B(_202_), .Y(_203_) );
NOR2X1 NOR2X1_5 ( .A(_299_), .B(_143_), .Y(_343_) );
NOR2X1 NOR2X1_6 ( .A(ULA_ctrl[2]), .B(_31_), .Y(_35_) );
NOR2X1 NOR2X1_7 ( .A(_15_), .B(_351_), .Y(_352_) );
NOR2X1 NOR2X1_8 ( .A(ULA_B_2_bF_buf3), .B(_160_), .Y(_161_) );
NOR2X1 NOR2X1_9 ( .A(_299_), .B(_177_), .Y(_361_) );
NOR2X1 NOR2X1_10 ( .A(_90_), .B(_370_), .Y(_371_) );
NOR2X1 NOR2X1_11 ( .A(_518__7_), .B(_518__4_), .Y(_465_) );
NOR2X1 NOR2X1_12 ( .A(_491_), .B(_261_), .Y(_271_) );
NOR2X1 NOR2X1_13 ( .A(_518__6_), .B(_518__5_), .Y(_472_) );
NOR2X1 NOR2X1_14 ( .A(ULA_A[14]), .B(ULA_B[14]), .Y(_433_) );
NOR2X1 NOR2X1_15 ( .A(_473_), .B(_474_), .Y(_475_) );
NOR2X1 NOR2X1_16 ( .A(_509_), .B(_25_), .Y(_212_) );
NOR2X1 NOR2X1_17 ( .A(_470_), .B(_476_), .Y(zero) );
NOR2X1 NOR2X1_18 ( .A(ULA_ctrl[1]), .B(_447_), .Y(_458_) );
NOR2X1 NOR2X1_19 ( .A(ULA_B[4]), .B(_36_), .Y(_37_) );
NOR2X1 NOR2X1_20 ( .A(ULA_B[3]), .B(_487__bF_buf2), .Y(_46_) );
NOR2X1 NOR2X1_21 ( .A(ULA_B_0_bF_buf5), .B(ULA_B_1_bF_buf2), .Y(_488_) );
NOR2X1 NOR2X1_22 ( .A(_47_), .B(_48_), .Y(_49_) );
NOR2X1 NOR2X1_23 ( .A(_174_), .B(_489_), .Y(_274_) );
NOR2X1 NOR2X1_24 ( .A(ULA_B[3]), .B(ULA_B[4]), .Y(_57_) );
NOR2X1 NOR2X1_25 ( .A(_56_), .B(_58_), .Y(_59_) );
NOR2X1 NOR2X1_26 ( .A(_111_), .B(_38__bF_buf4), .Y(_112_) );
NOR2X1 NOR2X1_27 ( .A(_125_), .B(_487__bF_buf0), .Y(_126_) );
NOR2X1 NOR2X1_28 ( .A(_64_), .B(_66_), .Y(_67_) );
NOR2X1 NOR2X1_29 ( .A(_130_), .B(_136_), .Y(_137_) );
NOR2X1 NOR2X1_30 ( .A(_495_), .B(_143_), .Y(_144_) );
NOR2X1 NOR2X1_31 ( .A(ULA_B_1_bF_buf4), .B(_138_), .Y(_146_) );
NOR2X1 NOR2X1_32 ( .A(_174_), .B(_26_), .Y(_175_) );
NOR2X1 NOR2X1_33 ( .A(_186_), .B(_189_), .Y(_190_) );
NOR2X1 NOR2X1_34 ( .A(ULA_B_1_bF_buf3), .B(_507_), .Y(_153_) );
NOR2X1 NOR2X1_35 ( .A(ULA_B_2_bF_buf0), .B(_193_), .Y(_194_) );
NOR2X1 NOR2X1_36 ( .A(_492_), .B(_311_), .Y(_445_) );
NOR2X1 NOR2X1_37 ( .A(_505_), .B(_492_), .Y(_196_) );
NOR2X1 NOR2X1_38 ( .A(_491_), .B(_212_), .Y(_223_) );
NOR2X1 NOR2X1_39 ( .A(_497_), .B(_94_), .Y(_227_) );
NOR2X1 NOR2X1_40 ( .A(_491_), .B(_237_), .Y(_248_) );
NOR2X1 NOR2X1_41 ( .A(ULA_B_2_bF_buf4), .B(ULA_B[3]), .Y(_22_) );
NOR2X1 NOR2X1_42 ( .A(_497_), .B(_142_), .Y(_253_) );
NOR2X1 NOR2X1_43 ( .A(_497_), .B(_176_), .Y(_276_) );
NOR2X1 NOR2X1_44 ( .A(_498_), .B(_6_), .Y(_450_) );
NOR2X1 NOR2X1_45 ( .A(_491_), .B(_283_), .Y(_294_) );
NOR2X1 NOR2X1_46 ( .A(ULA_B_1_bF_buf1), .B(_68_), .Y(_106_) );
NOR2X1 NOR2X1_47 ( .A(_11_), .B(_306_), .Y(_307_) );
NOR3X1 NOR3X1_1 ( .A(ULA_B_0_bF_buf4), .B(ULA_B_1_bF_buf1), .C(ULA_B_2_bF_buf1), .Y(_493_) );
NOR3X1 NOR3X1_2 ( .A(ULA_B_2_bF_buf3), .B(_492_), .C(_160_), .Y(_344_) );
NOR3X1 NOR3X1_3 ( .A(ULA_B_2_bF_buf1), .B(_492_), .C(_193_), .Y(_362_) );
OAI21X1 OAI21X1_1 ( .A(ULA_ctrl_0_bF_buf3), .B(_420_), .C(_421_), .Y(_422_) );
OAI21X1 OAI21X1_2 ( .A(ULA_B_0_bF_buf5), .B(_509_), .C(_216_), .Y(_217_) );
OAI21X1 OAI21X1_3 ( .A(ULA_B_1_bF_buf0), .B(_138_), .C(ULA_B_2_bF_buf2), .Y(_349_) );
OAI21X1 OAI21X1_4 ( .A(ULA_B_0_bF_buf0), .B(_90_), .C(_91_), .Y(_92_) );
OAI21X1 OAI21X1_5 ( .A(_487__bF_buf0), .B(_180_), .C(_182_), .Y(_183_) );
OAI21X1 OAI21X1_6 ( .A(_251_), .B(_431_), .C(_437_), .Y(_438_) );
OAI21X1 OAI21X1_7 ( .A(_504__bF_buf1), .B(_89_), .C(_93_), .Y(_94_) );
OAI21X1 OAI21X1_8 ( .A(_52_), .B(_307_), .C(_480__bF_buf0), .Y(_308_) );
OAI21X1 OAI21X1_9 ( .A(ULA_B_1_bF_buf4), .B(_88_), .C(_99_), .Y(_100_) );
OAI21X1 OAI21X1_10 ( .A(ULA_B_1_bF_buf3), .B(_84_), .C(_83_), .Y(_101_) );
OAI21X1 OAI21X1_11 ( .A(_119_), .B(_291_), .C(_285_), .Y(_292_) );
OAI21X1 OAI21X1_12 ( .A(ULA_B_2_bF_buf4), .B(_100_), .C(_102_), .Y(_103_) );
OAI21X1 OAI21X1_13 ( .A(_455_), .B(_52_), .C(_480__bF_buf3), .Y(_456_) );
OAI21X1 OAI21X1_14 ( .A(_38__bF_buf0), .B(_107_), .C(_22_), .Y(_108_) );
OAI21X1 OAI21X1_15 ( .A(_52_), .B(_352_), .C(_480__bF_buf2), .Y(_353_) );
OAI21X1 OAI21X1_16 ( .A(_106_), .B(_108_), .C(_37_), .Y(_109_) );
OAI21X1 OAI21X1_17 ( .A(_52_), .B(_112_), .C(_480__bF_buf3), .Y(_113_) );
OAI21X1 OAI21X1_18 ( .A(ULA_A[1]), .B(ULA_B_1_bF_buf0), .C(_113_), .Y(_114_) );
OAI21X1 OAI21X1_19 ( .A(_47_), .B(_218_), .C(_317_), .Y(_318_) );
OAI21X1 OAI21X1_20 ( .A(ULA_B_0_bF_buf5), .B(_111_), .C(_426_), .Y(_115_) );
OAI21X1 OAI21X1_21 ( .A(_447_), .B(_31_), .C(_56_), .Y(_118_) );
OAI21X1 OAI21X1_22 ( .A(_430_), .B(_438_), .C(_422_), .Y(_439_) );
OAI21X1 OAI21X1_23 ( .A(ULA_A[8]), .B(ULA_B[8]), .C(_308_), .Y(_309_) );
OAI21X1 OAI21X1_24 ( .A(_119_), .B(_220_), .C(_214_), .Y(_221_) );
OAI21X1 OAI21X1_25 ( .A(ULA_B_0_bF_buf0), .B(_15_), .C(_16_), .Y(_17_) );
OAI21X1 OAI21X1_26 ( .A(ULA_ctrl_0_bF_buf2), .B(_127_), .C(_128_), .Y(_129_) );
OAI21X1 OAI21X1_27 ( .A(ULA_A[10]), .B(ULA_B[10]), .C(_353_), .Y(_354_) );
OAI21X1 OAI21X1_28 ( .A(_504__bF_buf4), .B(_507_), .C(_131_), .Y(_132_) );
OAI21X1 OAI21X1_29 ( .A(_504__bF_buf2), .B(_133_), .C(_134_), .Y(_135_) );
OAI21X1 OAI21X1_30 ( .A(_504__bF_buf1), .B(_138_), .C(_1_), .Y(_139_) );
OAI21X1 OAI21X1_31 ( .A(_504__bF_buf4), .B(_140_), .C(_141_), .Y(_142_) );
OAI21X1 OAI21X1_32 ( .A(_1_), .B(_142_), .C(_139_), .Y(_143_) );
OAI21X1 OAI21X1_33 ( .A(_38__bF_buf2), .B(_76_), .C(_22_), .Y(_185_) );
OAI21X1 OAI21X1_34 ( .A(_144_), .B(_137_), .C(_33_), .Y(_145_) );
OAI21X1 OAI21X1_35 ( .A(ULA_B_0_bF_buf1), .B(_77_), .C(_74_), .Y(_288_) );
OAI21X1 OAI21X1_36 ( .A(_487__bF_buf2), .B(_146_), .C(_148_), .Y(_149_) );
OAI21X1 OAI21X1_37 ( .A(_38__bF_buf0), .B(_13_), .C(_151_), .Y(_152_) );
OAI21X1 OAI21X1_38 ( .A(_504__bF_buf3), .B(_14_), .C(_18_), .Y(_19_) );
OAI21X1 OAI21X1_39 ( .A(ULA_ctrl_0_bF_buf0), .B(_357_), .C(_358_), .Y(_359_) );
OAI21X1 OAI21X1_40 ( .A(_38__bF_buf4), .B(_512_), .C(_22_), .Y(_154_) );
OAI21X1 OAI21X1_41 ( .A(ULA_A[15]), .B(ULA_B[15]), .C(_456_), .Y(_457_) );
OAI21X1 OAI21X1_42 ( .A(ULA_B_1_bF_buf4), .B(_170_), .C(_187_), .Y(_188_) );
OAI21X1 OAI21X1_43 ( .A(_47_), .B(_188_), .C(_37_), .Y(_189_) );
OAI21X1 OAI21X1_44 ( .A(ULA_B_0_bF_buf0), .B(_505_), .C(_191_), .Y(_192_) );
OAI21X1 OAI21X1_45 ( .A(_52_), .B(_196_), .C(_480__bF_buf1), .Y(_197_) );
OAI21X1 OAI21X1_46 ( .A(_223_), .B(_224_), .C(_67_), .Y(_225_) );
OAI21X1 OAI21X1_47 ( .A(ULA_B_0_bF_buf0), .B(_11_), .C(_514_), .Y(_313_) );
OAI21X1 OAI21X1_48 ( .A(ULA_A[3]), .B(ULA_B[3]), .C(_197_), .Y(_198_) );
OAI21X1 OAI21X1_49 ( .A(_1_), .B(_517_), .C(_495_), .Y(_205_) );
OAI21X1 OAI21X1_50 ( .A(_203_), .B(_206_), .C(_33_), .Y(_207_) );
OAI21X1 OAI21X1_51 ( .A(_447_), .B(_31_), .C(_478_), .Y(_32_) );
OAI21X1 OAI21X1_52 ( .A(_1_), .B(_81_), .C(_495_), .Y(_228_) );
OAI21X1 OAI21X1_53 ( .A(_237_), .B(_52_), .C(_480__bF_buf3), .Y(_238_) );
OAI21X1 OAI21X1_54 ( .A(ULA_A[5]), .B(ULA_B[5]), .C(_238_), .Y(_239_) );
OAI21X1 OAI21X1_55 ( .A(ULA_ctrl_0_bF_buf4), .B(_426_), .C(_485_), .Y(_486_) );
OAI21X1 OAI21X1_56 ( .A(_343_), .B(_356_), .C(_359_), .Y(_360_) );
OAI21X1 OAI21X1_57 ( .A(ULA_B_0_bF_buf4), .B(_73_), .C(_69_), .Y(_242_) );
OAI21X1 OAI21X1_58 ( .A(_119_), .B(_245_), .C(_239_), .Y(_246_) );
OAI21X1 OAI21X1_59 ( .A(_248_), .B(_249_), .C(_67_), .Y(_250_) );
OAI21X1 OAI21X1_60 ( .A(_460_), .B(_443_), .C(_463_), .Y(_464_) );
OAI21X1 OAI21X1_61 ( .A(ULA_B_1_bF_buf3), .B(_288_), .C(_363_), .Y(_364_) );
OAI21X1 OAI21X1_62 ( .A(_153_), .B(_154_), .C(_37_), .Y(_155_) );
OAI21X1 OAI21X1_63 ( .A(_1_), .B(_135_), .C(_495_), .Y(_254_) );
OAI21X1 OAI21X1_64 ( .A(ULA_B_1_bF_buf3), .B(_14_), .C(_42_), .Y(_43_) );
OAI21X1 OAI21X1_65 ( .A(_261_), .B(_52_), .C(_480__bF_buf2), .Y(_262_) );
OAI21X1 OAI21X1_66 ( .A(ULA_A[6]), .B(ULA_B[6]), .C(_262_), .Y(_263_) );
OAI21X1 OAI21X1_67 ( .A(_26_), .B(_27_), .C(ULA_ctrl_0_bF_buf0), .Y(_28_) );
OAI21X1 OAI21X1_68 ( .A(ULA_B_0_bF_buf3), .B(_513_), .C(_510_), .Y(_265_) );
OAI21X1 OAI21X1_69 ( .A(_119_), .B(_268_), .C(_263_), .Y(_269_) );
OAI21X1 OAI21X1_70 ( .A(_271_), .B(_272_), .C(_67_), .Y(_273_) );
OAI21X1 OAI21X1_71 ( .A(ULA_ctrl_0_bF_buf4), .B(_321_), .C(_322_), .Y(_323_) );
OAI21X1 OAI21X1_72 ( .A(_1_), .B(_172_), .C(_495_), .Y(_277_) );
OAI21X1 OAI21X1_73 ( .A(_427_), .B(_428_), .C(_492_), .Y(_429_) );
OAI21X1 OAI21X1_74 ( .A(_276_), .B(_277_), .C(_275_), .Y(_278_) );
OAI21X1 OAI21X1_75 ( .A(_283_), .B(_52_), .C(_480__bF_buf1), .Y(_284_) );
OAI21X1 OAI21X1_76 ( .A(ULA_B_0_bF_buf3), .B(_157_), .C(ULA_B_1_bF_buf2), .Y(_158_) );
OAI21X1 OAI21X1_77 ( .A(ULA_B_2_bF_buf1), .B(_43_), .C(_41_), .Y(_44_) );
OAI21X1 OAI21X1_78 ( .A(_47_), .B(_43_), .C(_37_), .Y(_210_) );
OAI21X1 OAI21X1_79 ( .A(ULA_A[7]), .B(ULA_B[7]), .C(_284_), .Y(_285_) );
OAI21X1 OAI21X1_80 ( .A(_300_), .B(_320_), .C(_323_), .Y(_324_) );
OAI21X1 OAI21X1_81 ( .A(ULA_B_0_bF_buf6), .B(_86_), .C(_78_), .Y(_326_) );
OAI21X1 OAI21X1_82 ( .A(_329_), .B(_330_), .C(_312_), .Y(_331_) );
OAI21X1 OAI21X1_83 ( .A(_52_), .B(_334_), .C(_480__bF_buf3), .Y(_335_) );
OAI21X1 OAI21X1_84 ( .A(ULA_A[9]), .B(ULA_B[9]), .C(_335_), .Y(_336_) );
OAI21X1 OAI21X1_85 ( .A(_38__bF_buf3), .B(_326_), .C(_366_), .Y(_367_) );
OAI21X1 OAI21X1_86 ( .A(_446_), .B(_458_), .C(ULA_ctrl[3]), .Y(_468_) );
OAI21X1 OAI21X1_87 ( .A(ULA_ctrl_0_bF_buf2), .B(_339_), .C(_340_), .Y(_341_) );
OAI21X1 OAI21X1_88 ( .A(_325_), .B(_338_), .C(_341_), .Y(_342_) );
OAI21X1 OAI21X1_89 ( .A(_316_), .B(_318_), .C(_312_), .Y(_319_) );
OAI21X1 OAI21X1_90 ( .A(ULA_B_0_bF_buf5), .B(_15_), .C(_12_), .Y(_345_) );
OAI21X1 OAI21X1_91 ( .A(ULA_B_1_bF_buf1), .B(_159_), .C(_158_), .Y(_160_) );
OAI21X1 OAI21X1_92 ( .A(_362_), .B(_368_), .C(_312_), .Y(_369_) );
OAI21X1 OAI21X1_93 ( .A(_52_), .B(_371_), .C(_480__bF_buf1), .Y(_372_) );
OAI21X1 OAI21X1_94 ( .A(ULA_A[11]), .B(ULA_B[11]), .C(_372_), .Y(_373_) );
OAI21X1 OAI21X1_95 ( .A(ULA_B_0_bF_buf3), .B(ULA_B_1_bF_buf0), .C(ULA_ctrl_0_bF_buf1), .Y(_496_) );
OAI21X1 OAI21X1_96 ( .A(_492_), .B(_44_), .C(_50_), .Y(_51_) );
OAI21X1 OAI21X1_97 ( .A(_64_), .B(_66_), .C(_373_), .Y(_374_) );
OAI21X1 OAI21X1_98 ( .A(ULA_ctrl_0_bF_buf3), .B(_377_), .C(_378_), .Y(_379_) );
OAI21X1 OAI21X1_99 ( .A(_361_), .B(_376_), .C(_379_), .Y(_380_) );
OAI21X1 OAI21X1_100 ( .A(_52_), .B(_212_), .C(_480__bF_buf0), .Y(_213_) );
OAI21X1 OAI21X1_101 ( .A(ULA_B_0_bF_buf3), .B(_2_), .C(_16_), .Y(_382_) );
OAI21X1 OAI21X1_102 ( .A(_53_), .B(_52_), .C(_480__bF_buf1), .Y(_54_) );
OAI21X1 OAI21X1_103 ( .A(_38__bF_buf4), .B(_287_), .C(_289_), .Y(_290_) );
OAI21X1 OAI21X1_104 ( .A(_385_), .B(_386_), .C(_492_), .Y(_387_) );
OAI21X1 OAI21X1_105 ( .A(_52_), .B(_126_), .C(_480__bF_buf2), .Y(_163_) );
OAI21X1 OAI21X1_106 ( .A(_392_), .B(_52_), .C(_480__bF_buf0), .Y(_393_) );
OAI21X1 OAI21X1_107 ( .A(ULA_A[12]), .B(ULA_B[12]), .C(_393_), .Y(_394_) );
OAI21X1 OAI21X1_108 ( .A(ULA_B_0_bF_buf2), .B(_125_), .C(_500_), .Y(_159_) );
OAI21X1 OAI21X1_109 ( .A(_64_), .B(_66_), .C(_394_), .Y(_395_) );
OAI21X1 OAI21X1_110 ( .A(ULA_ctrl_0_bF_buf1), .B(_398_), .C(_399_), .Y(_400_) );
OAI21X1 OAI21X1_111 ( .A(ULA_A[4]), .B(ULA_B[4]), .C(_213_), .Y(_214_) );
OAI21X1 OAI21X1_112 ( .A(_388_), .B(_397_), .C(_400_), .Y(_401_) );
OAI21X1 OAI21X1_113 ( .A(_502_), .B(_496_), .C(_503_), .Y(_504_) );
OAI21X1 OAI21X1_114 ( .A(ULA_B_0_bF_buf2), .B(_404_), .C(_91_), .Y(_405_) );
OAI21X1 OAI21X1_115 ( .A(_504__bF_buf0), .B(_170_), .C(_171_), .Y(_172_) );
OAI21X1 OAI21X1_116 ( .A(_411_), .B(_52_), .C(_480__bF_buf3), .Y(_412_) );
OAI21X1 OAI21X1_117 ( .A(ULA_ctrl_0_bF_buf4), .B(_416_), .C(_417_), .Y(_418_) );
OAI21X1 OAI21X1_118 ( .A(ULA_B_2_bF_buf4), .B(_290_), .C(_286_), .Y(_291_) );
OAI21X1 OAI21X1_119 ( .A(ULA_A[2]), .B(ULA_B_2_bF_buf2), .C(_163_), .Y(_164_) );
OAI21X1 OAI21X1_120 ( .A(_347_), .B(_344_), .C(_312_), .Y(_348_) );
OAI21X1 OAI21X1_121 ( .A(_409_), .B(_415_), .C(_418_), .Y(_419_) );
OAI21X1 OAI21X1_122 ( .A(ULA_ctrl_0_bF_buf1), .B(_461_), .C(_462_), .Y(_463_) );
OAI21X1 OAI21X1_123 ( .A(ULA_B_0_bF_buf5), .B(ULA_A[2]), .C(_506_), .Y(_507_) );
OAI21X1 OAI21X1_124 ( .A(ULA_B_0_bF_buf3), .B(_509_), .C(_510_), .Y(_511_) );
OAI21X1 OAI21X1_125 ( .A(ULA_B_0_bF_buf1), .B(_513_), .C(_514_), .Y(_515_) );
OAI21X1 OAI21X1_126 ( .A(_504__bF_buf2), .B(_512_), .C(_516_), .Y(_517_) );
OAI21X1 OAI21X1_127 ( .A(ULA_B_0_bF_buf6), .B(_2_), .C(_3_), .Y(_4_) );
OAI21X1 OAI21X1_128 ( .A(ULA_A[0]), .B(ULA_B_0_bF_buf5), .C(_54_), .Y(_55_) );
OAI21X1 OAI21X1_129 ( .A(_38__bF_buf4), .B(_382_), .C(_487__bF_buf3), .Y(_425_) );
OAI21X1 OAI21X1_130 ( .A(ULA_B_0_bF_buf4), .B(_6_), .C(_7_), .Y(_8_) );
OAI21X1 OAI21X1_131 ( .A(_504__bF_buf0), .B(_5_), .C(_9_), .Y(_10_) );
OAI21X1 OAI21X1_132 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
OAI21X1 OAI21X1_133 ( .A(ULA_B_1_bF_buf3), .B(_499_), .C(ULA_B_2_bF_buf3), .Y(_215_) );
OAI21X1 OAI21X1_134 ( .A(ULA_B_0_bF_buf2), .B(_11_), .C(_12_), .Y(_13_) );
OAI21X1 OAI21X1_135 ( .A(_294_), .B(_295_), .C(_67_), .Y(_296_) );
OAI21X1 OAI21X1_136 ( .A(ULA_B_0_bF_buf2), .B(_505_), .C(_69_), .Y(_70_) );
OAI21X1 OAI21X1_137 ( .A(_504__bF_buf1), .B(_68_), .C(_71_), .Y(_72_) );
OAI21X1 OAI21X1_138 ( .A(ULA_B_0_bF_buf0), .B(_73_), .C(_74_), .Y(_75_) );
OAI21X1 OAI21X1_139 ( .A(ULA_B_0_bF_buf5), .B(_77_), .C(_78_), .Y(_79_) );
OAI21X1 OAI21X1_140 ( .A(_504__bF_buf2), .B(_107_), .C(_168_), .Y(_169_) );
OAI21X1 OAI21X1_141 ( .A(_504__bF_buf4), .B(_76_), .C(_80_), .Y(_81_) );
OAI21X1 OAI21X1_142 ( .A(_84_), .B(_504__bF_buf3), .C(_83_), .Y(_85_) );
OAI21X1 OAI21X1_143 ( .A(ULA_B_0_bF_buf2), .B(_86_), .C(_87_), .Y(_88_) );
OAI22X1 OAI22X1_1 ( .A(_433_), .B(_435_), .C(_303_), .D(_257_), .Y(_436_) );
OAI22X1 OAI22X1_2 ( .A(_495_), .B(_226_), .C(_227_), .D(_228_), .Y(_229_) );
OAI22X1 OAI22X1_3 ( .A(_251_), .B(_252_), .C(_253_), .D(_254_), .Y(_255_) );
OAI22X1 OAI22X1_4 ( .A(_492_), .B(_116_), .C(_47_), .D(_243_), .Y(_330_) );
OAI22X1 OAI22X1_5 ( .A(_27_), .B(_346_), .C(_47_), .D(_266_), .Y(_347_) );
OAI22X1 OAI22X1_6 ( .A(_27_), .B(_367_), .C(_47_), .D(_364_), .Y(_368_) );
OR2X2 OR2X2_1 ( .A(ULA_B_0_bF_buf6), .B(ULA_B_1_bF_buf2), .Y(_26_) );
OR2X2 OR2X2_2 ( .A(ULA_B_2_bF_buf3), .B(ULA_B[3]), .Y(_27_) );
OR2X2 OR2X2_3 ( .A(_103_), .B(_492_), .Y(_104_) );
OR2X2 OR2X2_4 ( .A(_183_), .B(_492_), .Y(_184_) );
OR2X2 OR2X2_5 ( .A(_208_), .B(_492_), .Y(_209_) );
OR2X2 OR2X2_6 ( .A(_504__bF_buf3), .B(_138_), .Y(_251_) );
OR2X2 OR2X2_7 ( .A(_405_), .B(ULA_B_1_bF_buf1), .Y(_406_) );
OR2X2 OR2X2_8 ( .A(ULA_A[13]), .B(ULA_B[13]), .Y(_410_) );
XNOR2X1 XNOR2X1_1 ( .A(_496_), .B(_487__bF_buf3), .Y(_497_) );
XNOR2X1 XNOR2X1_2 ( .A(_496_), .B(ULA_B_2_bF_buf0), .Y(_1_) );
XNOR2X1 XNOR2X1_3 ( .A(_112_), .B(ULA_ctrl_0_bF_buf4), .Y(_124_) );
XNOR2X1 XNOR2X1_4 ( .A(_196_), .B(ULA_ctrl_0_bF_buf1), .Y(_201_) );
BUFX2 BUFX2_20 ( .A(_518__0_), .Y(ULA_OUT[0]) );
BUFX2 BUFX2_21 ( .A(_518__1_), .Y(ULA_OUT[1]) );
BUFX2 BUFX2_22 ( .A(_518__2_), .Y(ULA_OUT[2]) );
BUFX2 BUFX2_23 ( .A(_518__3_), .Y(ULA_OUT[3]) );
BUFX2 BUFX2_24 ( .A(_518__4_), .Y(ULA_OUT[4]) );
BUFX2 BUFX2_25 ( .A(_518__5_), .Y(ULA_OUT[5]) );
BUFX2 BUFX2_26 ( .A(_518__6_), .Y(ULA_OUT[6]) );
BUFX2 BUFX2_27 ( .A(_518__7_), .Y(ULA_OUT[7]) );
BUFX2 BUFX2_28 ( .A(_518__8_), .Y(ULA_OUT[8]) );
BUFX2 BUFX2_29 ( .A(_518__9_), .Y(ULA_OUT[9]) );
BUFX2 BUFX2_30 ( .A(_518__10_), .Y(ULA_OUT[10]) );
BUFX2 BUFX2_31 ( .A(_518__11_), .Y(ULA_OUT[11]) );
BUFX2 BUFX2_32 ( .A(_518__12_), .Y(ULA_OUT[12]) );
BUFX2 BUFX2_33 ( .A(_518__13_), .Y(ULA_OUT[13]) );
BUFX2 BUFX2_34 ( .A(_518__14_), .Y(ULA_OUT[14]) );
BUFX2 BUFX2_35 ( .A(_518__15_), .Y(ULA_OUT[15]) );
BUFX2 BUFX2_36 ( .A(_519__0_), .Y(ULA_flags[0]) );
BUFX2 BUFX2_37 ( .A(_519__1_), .Y(ULA_flags[1]) );
BUFX2 BUFX2_38 ( .A(_519__2_), .Y(ULA_flags[2]) );
endmodule
