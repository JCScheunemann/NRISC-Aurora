module NRISC_REGs ( gnd, vdd, REG_D, REG_RF1, REG_RF2, REG_RFD, REG_R1, REG_Write, REG_Interrupt_flag, clk, rst, REG_A, REG_B);

input gnd, vdd;
input REG_Write;
input REG_Interrupt_flag;
input clk;
input rst;
input [15:0] REG_D;
input [3:0] REG_RF1;
input [3:0] REG_RF2;
input [3:0] REG_RFD;
input [15:0] REG_R1;
output [15:0] REG_A;
output [15:0] REG_B;

AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_1626_), .B(_500_), .Y(_501_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_500_), .Y(_518_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_1680_), .B(_500_), .Y(_536_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_500_), .Y(_568_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_1717_), .Y(_585_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_500_), .Y(_603_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(REG_RF2[3]), .Y(_673_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(REG_RF1[3]), .Y(_1294_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_1623_), .Y(_1604_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf0), .B(_501__bF_buf0), .C(_502_), .Y(_224_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf0), .B(_501__bF_buf2), .C(_511_), .Y(_233_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf3), .B(_501__bF_buf1), .C(_512_), .Y(_234_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf0), .B(_501__bF_buf4), .C(_513_), .Y(_235_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf3), .B(_501__bF_buf1), .C(_514_), .Y(_236_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf0), .B(_501__bF_buf0), .C(_515_), .Y(_237_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf3), .B(_501__bF_buf3), .C(_516_), .Y(_238_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf0), .B(_501__bF_buf4), .C(_517_), .Y(_239_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf0), .B(_518__bF_buf1), .C(_519_), .Y(_240_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf3), .B(_518__bF_buf1), .C(_520_), .Y(_241_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_518__bF_buf4), .C(_521_), .Y(_242_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf3), .B(_501__bF_buf0), .C(_503_), .Y(_225_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf3), .B(_518__bF_buf2), .C(_522_), .Y(_243_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf0), .B(_518__bF_buf3), .C(_523_), .Y(_244_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf3), .B(_518__bF_buf3), .C(_524_), .Y(_245_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf3), .B(_518__bF_buf4), .C(_525_), .Y(_246_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf3), .B(_518__bF_buf2), .C(_526_), .Y(_247_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf2), .B(_518__bF_buf0), .C(_527_), .Y(_248_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf0), .B(_518__bF_buf0), .C(_528_), .Y(_249_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf3), .B(_518__bF_buf4), .C(_529_), .Y(_250_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf0), .B(_518__bF_buf0), .C(_530_), .Y(_251_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf3), .B(_518__bF_buf0), .C(_531_), .Y(_252_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_501__bF_buf2), .C(_504_), .Y(_226_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf0), .B(_518__bF_buf1), .C(_532_), .Y(_253_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf3), .B(_518__bF_buf2), .C(_533_), .Y(_254_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf0), .B(_518__bF_buf3), .C(_534_), .Y(_255_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf0), .B(_568__bF_buf3), .C(_569_), .Y(_272_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf3), .B(_568__bF_buf3), .C(_570_), .Y(_273_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_568__bF_buf2), .C(_571_), .Y(_274_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf3), .B(_568__bF_buf4), .C(_572_), .Y(_275_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf0), .B(_568__bF_buf1), .C(_573_), .Y(_276_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf3), .B(_568__bF_buf1), .C(_574_), .Y(_277_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf3), .B(_568__bF_buf1), .C(_575_), .Y(_278_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf3), .B(_501__bF_buf3), .C(_505_), .Y(_227_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf3), .B(_568__bF_buf4), .C(_576_), .Y(_279_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf2), .B(_568__bF_buf0), .C(_577_), .Y(_280_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf0), .B(_568__bF_buf1), .C(_578_), .Y(_281_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf3), .B(_568__bF_buf0), .C(_579_), .Y(_282_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf0), .B(_568__bF_buf2), .C(_580_), .Y(_283_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf3), .B(_568__bF_buf0), .C(_581_), .Y(_284_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf0), .B(_568__bF_buf3), .C(_582_), .Y(_285_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf3), .B(_568__bF_buf4), .C(_583_), .Y(_286_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf0), .B(_568__bF_buf3), .C(_584_), .Y(_287_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf0), .B(_585__bF_buf2), .C(_586_), .Y(_288_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf0), .B(_501__bF_buf4), .C(_506_), .Y(_228_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf3), .B(_585__bF_buf0), .C(_587_), .Y(_289_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_585__bF_buf1), .C(_588_), .Y(_290_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf3), .B(_585__bF_buf3), .C(_589_), .Y(_291_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf0), .B(_585__bF_buf4), .C(_590_), .Y(_292_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf3), .B(_585__bF_buf4), .C(_591_), .Y(_293_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf3), .B(_585__bF_buf4), .C(_592_), .Y(_294_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf3), .B(_585__bF_buf3), .C(_593_), .Y(_295_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf2), .B(_585__bF_buf1), .C(_594_), .Y(_296_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf0), .B(_585__bF_buf4), .C(_595_), .Y(_297_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf3), .B(_585__bF_buf1), .C(_596_), .Y(_298_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf3), .B(_501__bF_buf4), .C(_507_), .Y(_229_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf0), .B(_585__bF_buf2), .C(_597_), .Y(_299_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf3), .B(_585__bF_buf2), .C(_598_), .Y(_300_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf0), .B(_585__bF_buf0), .C(_599_), .Y(_301_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf3), .B(_585__bF_buf3), .C(_600_), .Y(_302_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf0), .B(_585__bF_buf0), .C(_601_), .Y(_303_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf3), .B(_501__bF_buf2), .C(_508_), .Y(_230_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf3), .B(_501__bF_buf3), .C(_509_), .Y(_231_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf2), .B(_501__bF_buf1), .C(_510_), .Y(_232_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_1748__0_), .Y(_1748__0_) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_1748__9_), .Y(_1748__9_) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_1748__10_), .Y(_1748__10_) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_1748__11_), .Y(_1748__11_) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_1748__12_), .Y(_1748__12_) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_1748__13_), .Y(_1748__13_) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_1748__14_), .Y(_1748__14_) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_1748__15_), .Y(_1748__15_) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_1749__0_), .Y(_1749__0_) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_1749__1_), .Y(_1749__1_) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_1749__2_), .Y(_1749__2_) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_1748__1_), .Y(_1748__1_) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_1749__3_), .Y(_1749__3_) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_1749__4_), .Y(_1749__4_) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_1749__5_), .Y(_1749__5_) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_1749__6_), .Y(_1749__6_) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_1749__7_), .Y(_1749__7_) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_1749__8_), .Y(_1749__8_) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_1749__9_), .Y(_1749__9_) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_1749__10_), .Y(_1749__10_) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_1749__11_), .Y(_1749__11_) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_1749__12_), .Y(_1749__12_) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_1748__2_), .Y(_1748__2_) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_1749__13_), .Y(_1749__13_) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1749__14_), .Y(_1749__14_) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_1749__15_), .Y(_1749__15_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_1748__3_), .Y(_1748__3_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_1748__4_), .Y(_1748__4_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1748__5_), .Y(_1748__5_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_1748__6_), .Y(_1748__6_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_1748__7_), .Y(_1748__7_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_1748__8_), .Y(_1748__8_) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_397_), .Y(_397__bF_buf2) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf8) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf7) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf6) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf5) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf4) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf3) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf2) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf1) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf0) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .Y(_1653__bF_buf3) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_397_), .Y(_397__bF_buf1) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .Y(_1653__bF_buf2) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .Y(_1653__bF_buf1) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .Y(_1653__bF_buf0) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf6) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf5) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf4) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf3) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf2) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf1) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .Y(_1268__bF_buf0) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(_397_), .Y(_397__bF_buf0) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .Y(_1647__bF_buf3) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .Y(_1647__bF_buf2) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .Y(_1647__bF_buf1) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .Y(_1647__bF_buf0) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .Y(_1641__bF_buf3) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .Y(_1641__bF_buf2) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .Y(_1641__bF_buf1) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .Y(_1641__bF_buf0) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf3) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf2) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf6) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf1) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .Y(_1735__bF_buf0) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf6) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf5) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf4) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf3) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf2) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf1) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1294__bF_buf0) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf4) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf5) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf3) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf2) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf1) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_414_), .Y(_414__bF_buf0) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .Y(_1635__bF_buf3) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .Y(_1635__bF_buf2) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .Y(_1635__bF_buf1) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .Y(_1635__bF_buf0) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf6) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf5) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf4) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf4) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf3) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf2) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf1) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_640__bF_buf0) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .Y(_1629__bF_buf3) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .Y(_1629__bF_buf2) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .Y(_1629__bF_buf1) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .Y(_1629__bF_buf0) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf4) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf3) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf3) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf2) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf1) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1699__bF_buf0) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .Y(_1661__bF_buf4) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .Y(_1661__bF_buf3) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .Y(_1661__bF_buf2) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .Y(_1661__bF_buf1) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .Y(_1661__bF_buf0) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .Y(_1655__bF_buf3) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf2) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .Y(_1655__bF_buf2) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .Y(_1655__bF_buf1) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .Y(_1655__bF_buf0) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(_431_), .Y(_431__bF_buf4) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(_431_), .Y(_431__bF_buf3) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(_431_), .Y(_431__bF_buf2) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(_431_), .Y(_431__bF_buf1) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(_431_), .Y(_431__bF_buf0) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .Y(_1649__bF_buf3) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .Y(_1649__bF_buf2) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf1) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .Y(_1649__bF_buf1) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .Y(_1649__bF_buf0) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .Y(_1264__bF_buf4) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .Y(_1264__bF_buf3) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .Y(_1264__bF_buf2) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .Y(_1264__bF_buf1) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .Y(_1264__bF_buf0) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(_1587__bF_buf4) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(_1587__bF_buf3) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(_1587__bF_buf2) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(_644_), .Y(_644__bF_buf0) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(_1587__bF_buf1) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(_1587__bF_buf0) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .Y(_1643__bF_buf3) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .Y(_1643__bF_buf2) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .Y(_1643__bF_buf1) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .Y(_1643__bF_buf0) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1681__bF_buf4) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1681__bF_buf3) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1681__bF_buf2) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1681__bF_buf1) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_585__bF_buf4) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1681__bF_buf0) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .Y(_1637__bF_buf3) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .Y(_1637__bF_buf2) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .Y(_1637__bF_buf1) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .Y(_1637__bF_buf0) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(_448_), .Y(_448__bF_buf4) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(_448_), .Y(_448__bF_buf3) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(_448_), .Y(_448__bF_buf2) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(_448_), .Y(_448__bF_buf1) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(_448_), .Y(_448__bF_buf0) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_585__bF_buf3) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf3) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf2) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf1) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1631__bF_buf0) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_636__bF_buf4) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_636__bF_buf3) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_636__bF_buf2) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_636__bF_buf1) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(_636_), .Y(_636__bF_buf0) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(_501_), .Y(_501__bF_buf4) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_585__bF_buf2) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_501_), .Y(_501__bF_buf3) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_501_), .Y(_501__bF_buf2) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_501_), .Y(_501__bF_buf1) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_501_), .Y(_501__bF_buf0) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_536_), .Y(_536__bF_buf4) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_536_), .Y(_536__bF_buf3) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_536_), .Y(_536__bF_buf2) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(_536_), .Y(_536__bF_buf1) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(_536_), .Y(_536__bF_buf0) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .Y(_1278__bF_buf5) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_585__bF_buf1) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .Y(_1278__bF_buf4) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .Y(_1278__bF_buf3) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .Y(_1278__bF_buf2) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .Y(_1278__bF_buf1) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .Y(_1278__bF_buf0) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .Y(_1622__bF_buf3) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .Y(_1622__bF_buf2) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .Y(_1622__bF_buf1) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .Y(_1622__bF_buf0) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(_380_), .Y(_380__bF_buf4) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_585__bF_buf0) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(_380_), .Y(_380__bF_buf3) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(_380_), .Y(_380__bF_buf2) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(_380_), .Y(_380__bF_buf1) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_380_), .Y(_380__bF_buf0) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .Y(_1657__bF_buf3) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .Y(_1657__bF_buf2) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .Y(_1657__bF_buf1) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .Y(_1657__bF_buf0) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_568_), .Y(_568__bF_buf4) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_568_), .Y(_568__bF_buf3) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_603_), .Y(_603__bF_buf4) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_568_), .Y(_568__bF_buf2) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_568_), .Y(_568__bF_buf1) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_568_), .Y(_568__bF_buf0) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .Y(_1275__bF_buf4) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .Y(_1275__bF_buf3) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .Y(_1275__bF_buf2) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .Y(_1275__bF_buf1) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .Y(_1275__bF_buf0) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf6) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf5) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_603_), .Y(_603__bF_buf3) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf4) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf3) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf2) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf1) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .Y(_1272__bF_buf0) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .Y(_1651__bF_buf3) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .Y(_1651__bF_buf2) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .Y(_1651__bF_buf1) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .Y(_1651__bF_buf0) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(_465_), .Y(_465__bF_buf4) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(_603_), .Y(_603__bF_buf2) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(_465_), .Y(_465__bF_buf3) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_465_), .Y(_465__bF_buf2) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_465_), .Y(_465__bF_buf1) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_465_), .Y(_465__bF_buf0) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf13) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf12) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf11) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf10) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf9) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf8) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(_603_), .Y(_603__bF_buf1) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf7) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf6) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf5) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf4) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf3) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf2) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf1) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag), .Y(REG_Interrupt_flag_bF_buf0) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf4) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf3) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_603_), .Y(_603__bF_buf0) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf2) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf1) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_518_), .Y(_518__bF_buf0) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .Y(_1645__bF_buf3) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .Y(_1645__bF_buf2) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .Y(_1645__bF_buf1) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .Y(_1645__bF_buf0) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_650__bF_buf5) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_650__bF_buf4) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_650__bF_buf3) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .Y(_1633__bF_buf3) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_650__bF_buf2) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_650__bF_buf1) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_650__bF_buf0) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .Y(_1604__bF_buf4) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .Y(_1604__bF_buf3) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .Y(_1604__bF_buf2) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .Y(_1604__bF_buf1) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .Y(_1604__bF_buf0) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(_362_), .Y(_362__bF_buf4) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(_362_), .Y(_362__bF_buf3) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .Y(_1633__bF_buf2) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(_362_), .Y(_362__bF_buf2) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(_362_), .Y(_362__bF_buf1) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(_362_), .Y(_362__bF_buf0) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_647__bF_buf4) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_647__bF_buf3) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_647__bF_buf2) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_647__bF_buf1) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(_647_), .Y(_647__bF_buf0) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .Y(_1639__bF_buf3) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .Y(_1639__bF_buf2) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .Y(_1633__bF_buf1) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .Y(_1639__bF_buf1) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .Y(_1639__bF_buf0) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .Y(_1633__bF_buf0) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf6) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf5) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf4) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf3) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf2) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf1) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(_673_), .Y(_673__bF_buf0) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(_482_), .Y(_482__bF_buf4) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(_482_), .Y(_482__bF_buf3) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_482_), .Y(_482__bF_buf2) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_482_), .Y(_482__bF_buf1) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_482_), .Y(_482__bF_buf0) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .Y(_1627__bF_buf4) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .Y(_1627__bF_buf3) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .Y(_1627__bF_buf2) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .Y(_1627__bF_buf1) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .Y(_1627__bF_buf0) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .Y(_1718__bF_buf4) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .Y(_1718__bF_buf3) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .Y(_1718__bF_buf2) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .Y(_1718__bF_buf1) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(_1718_), .Y(_1718__bF_buf0) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_1621__bF_buf3) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_1621__bF_buf2) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_1621__bF_buf1) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_1621__bF_buf0) );
BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf48) );
BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf47) );
BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf46) );
BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf45) );
BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf44) );
BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf43) );
BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf42) );
BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf41) );
BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf40) );
BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf39) );
BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf38) );
BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf37) );
BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf36) );
BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf35) );
BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf34) );
BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf33) );
BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf32) );
BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf31) );
BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf30) );
BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf29) );
BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(_397_), .Y(_397__bF_buf4) );
BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28) );
BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf27) );
BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf26) );
BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf25) );
BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf24) );
BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf23) );
BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf22) );
BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf21) );
BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf20) );
BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf19) );
BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(_397_), .Y(_397__bF_buf3) );
BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf18) );
BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf17) );
BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf16) );
BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf15) );
BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf14) );
BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf13) );
BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf12) );
BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf11) );
BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf10) );
BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf9) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_32_), .Q(FIRQ_REGS_4__0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_41_), .Q(FIRQ_REGS_4__9_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_339_), .Q(FIRQ_REGS_0__3_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_340_), .Q(FIRQ_REGS_0__4_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_341_), .Q(FIRQ_REGS_0__5_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_342_), .Q(FIRQ_REGS_0__6_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_343_), .Q(FIRQ_REGS_0__7_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_344_), .Q(FIRQ_REGS_0__8_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_345_), .Q(FIRQ_REGS_0__9_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_346_), .Q(FIRQ_REGS_0__10_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_347_), .Q(FIRQ_REGS_0__11_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_348_), .Q(FIRQ_REGS_0__12_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_42_), .Q(FIRQ_REGS_4__10_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_349_), .Q(FIRQ_REGS_0__13_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_350_), .Q(FIRQ_REGS_0__14_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_351_), .Q(FIRQ_REGS_0__15_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0_), .Q(FIRQ_REGS_2__0_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_1_), .Q(FIRQ_REGS_2__1_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_2_), .Q(FIRQ_REGS_2__2_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3_), .Q(FIRQ_REGS_2__3_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_4_), .Q(FIRQ_REGS_2__4_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_5_), .Q(FIRQ_REGS_2__5_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_6_), .Q(FIRQ_REGS_2__6_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_43_), .Q(FIRQ_REGS_4__11_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_7_), .Q(FIRQ_REGS_2__7_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_8_), .Q(FIRQ_REGS_2__8_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_9_), .Q(FIRQ_REGS_2__9_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10_), .Q(FIRQ_REGS_2__10_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_11_), .Q(FIRQ_REGS_2__11_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_12_), .Q(FIRQ_REGS_2__12_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_13_), .Q(FIRQ_REGS_2__13_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_14_), .Q(FIRQ_REGS_2__14_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_15_), .Q(FIRQ_REGS_2__15_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_112_), .Q(USR_REGS_1__0_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_44_), .Q(FIRQ_REGS_4__12_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_113_), .Q(USR_REGS_1__1_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_114_), .Q(USR_REGS_1__2_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_115_), .Q(USR_REGS_1__3_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_116_), .Q(USR_REGS_1__4_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_117_), .Q(USR_REGS_1__5_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_118_), .Q(USR_REGS_1__6_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_119_), .Q(USR_REGS_1__7_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_120_), .Q(USR_REGS_1__8_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_121_), .Q(USR_REGS_1__9_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_122_), .Q(USR_REGS_1__10_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_45_), .Q(FIRQ_REGS_4__13_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_123_), .Q(USR_REGS_1__11_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_124_), .Q(USR_REGS_1__12_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_125_), .Q(USR_REGS_1__13_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_126_), .Q(USR_REGS_1__14_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_127_), .Q(USR_REGS_1__15_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_128_), .Q(USR_REGS_2__0_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_129_), .Q(USR_REGS_2__1_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_130_), .Q(USR_REGS_2__2_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_131_), .Q(USR_REGS_2__3_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_132_), .Q(USR_REGS_2__4_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_46_), .Q(FIRQ_REGS_4__14_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_133_), .Q(USR_REGS_2__5_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_134_), .Q(USR_REGS_2__6_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_135_), .Q(USR_REGS_2__7_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_136_), .Q(USR_REGS_2__8_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_137_), .Q(USR_REGS_2__9_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_138_), .Q(USR_REGS_2__10_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_139_), .Q(USR_REGS_2__11_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_140_), .Q(USR_REGS_2__12_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_141_), .Q(USR_REGS_2__13_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_142_), .Q(USR_REGS_2__14_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_47_), .Q(FIRQ_REGS_4__15_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_143_), .Q(USR_REGS_2__15_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_144_), .Q(USR_REGS_3__0_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_145_), .Q(USR_REGS_3__1_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_146_), .Q(USR_REGS_3__2_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_147_), .Q(USR_REGS_3__3_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_148_), .Q(USR_REGS_3__4_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_149_), .Q(USR_REGS_3__5_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_150_), .Q(USR_REGS_3__6_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_151_), .Q(USR_REGS_3__7_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_152_), .Q(USR_REGS_3__8_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_16_), .Q(FIRQ_REGS_3__0_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_153_), .Q(USR_REGS_3__9_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_154_), .Q(USR_REGS_3__10_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_155_), .Q(USR_REGS_3__11_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_156_), .Q(USR_REGS_3__12_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_157_), .Q(USR_REGS_3__13_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_158_), .Q(USR_REGS_3__14_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_159_), .Q(USR_REGS_3__15_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_160_), .Q(USR_REGS_4__0_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_161_), .Q(USR_REGS_4__1_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_162_), .Q(USR_REGS_4__2_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_17_), .Q(FIRQ_REGS_3__1_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_163_), .Q(USR_REGS_4__3_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_164_), .Q(USR_REGS_4__4_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_165_), .Q(USR_REGS_4__5_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_166_), .Q(USR_REGS_4__6_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_167_), .Q(USR_REGS_4__7_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_168_), .Q(USR_REGS_4__8_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_169_), .Q(USR_REGS_4__9_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_170_), .Q(USR_REGS_4__10_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_171_), .Q(USR_REGS_4__11_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_172_), .Q(USR_REGS_4__12_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_18_), .Q(FIRQ_REGS_3__2_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_173_), .Q(USR_REGS_4__13_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_174_), .Q(USR_REGS_4__14_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_175_), .Q(USR_REGS_4__15_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_176_), .Q(USR_REGS_5__0_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_177_), .Q(USR_REGS_5__1_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_178_), .Q(USR_REGS_5__2_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_179_), .Q(USR_REGS_5__3_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_180_), .Q(USR_REGS_5__4_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_181_), .Q(USR_REGS_5__5_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_182_), .Q(USR_REGS_5__6_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_33_), .Q(FIRQ_REGS_4__1_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_19_), .Q(FIRQ_REGS_3__3_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_183_), .Q(USR_REGS_5__7_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_184_), .Q(USR_REGS_5__8_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_185_), .Q(USR_REGS_5__9_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_186_), .Q(USR_REGS_5__10_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_187_), .Q(USR_REGS_5__11_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_188_), .Q(USR_REGS_5__12_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_189_), .Q(USR_REGS_5__13_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_190_), .Q(USR_REGS_5__14_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_191_), .Q(USR_REGS_5__15_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_192_), .Q(USR_REGS_6__0_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_20_), .Q(FIRQ_REGS_3__4_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_193_), .Q(USR_REGS_6__1_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_194_), .Q(USR_REGS_6__2_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_195_), .Q(USR_REGS_6__3_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_196_), .Q(USR_REGS_6__4_) );
DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_197_), .Q(USR_REGS_6__5_) );
DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_198_), .Q(USR_REGS_6__6_) );
DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_199_), .Q(USR_REGS_6__7_) );
DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_200_), .Q(USR_REGS_6__8_) );
DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_201_), .Q(USR_REGS_6__9_) );
DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_202_), .Q(USR_REGS_6__10_) );
DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_21_), .Q(FIRQ_REGS_3__5_) );
DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_203_), .Q(USR_REGS_6__11_) );
DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_204_), .Q(USR_REGS_6__12_) );
DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_205_), .Q(USR_REGS_6__13_) );
DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_206_), .Q(USR_REGS_6__14_) );
DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_207_), .Q(USR_REGS_6__15_) );
DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_208_), .Q(USR_REGS_7__0_) );
DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_209_), .Q(USR_REGS_7__1_) );
DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_210_), .Q(USR_REGS_7__2_) );
DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_211_), .Q(USR_REGS_7__3_) );
DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_212_), .Q(USR_REGS_7__4_) );
DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_22_), .Q(FIRQ_REGS_3__6_) );
DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_213_), .Q(USR_REGS_7__5_) );
DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_214_), .Q(USR_REGS_7__6_) );
DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_215_), .Q(USR_REGS_7__7_) );
DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_216_), .Q(USR_REGS_7__8_) );
DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_217_), .Q(USR_REGS_7__9_) );
DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_218_), .Q(USR_REGS_7__10_) );
DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_219_), .Q(USR_REGS_7__11_) );
DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_220_), .Q(USR_REGS_7__12_) );
DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_221_), .Q(USR_REGS_7__13_) );
DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_222_), .Q(USR_REGS_7__14_) );
DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_23_), .Q(FIRQ_REGS_3__7_) );
DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_223_), .Q(USR_REGS_7__15_) );
DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_240_), .Q(REGS_3__0_) );
DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_241_), .Q(REGS_3__1_) );
DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_242_), .Q(REGS_3__2_) );
DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_243_), .Q(REGS_3__3_) );
DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_244_), .Q(REGS_3__4_) );
DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_245_), .Q(REGS_3__5_) );
DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_246_), .Q(REGS_3__6_) );
DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_247_), .Q(REGS_3__7_) );
DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_248_), .Q(REGS_3__8_) );
DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_24_), .Q(FIRQ_REGS_3__8_) );
DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_249_), .Q(REGS_3__9_) );
DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_250_), .Q(REGS_3__10_) );
DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_251_), .Q(REGS_3__11_) );
DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_252_), .Q(REGS_3__12_) );
DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_253_), .Q(REGS_3__13_) );
DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_254_), .Q(REGS_3__14_) );
DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_255_), .Q(REGS_3__15_) );
DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_256_), .Q(REGS_4__0_) );
DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_257_), .Q(REGS_4__1_) );
DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_258_), .Q(REGS_4__2_) );
DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_25_), .Q(FIRQ_REGS_3__9_) );
DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_259_), .Q(REGS_4__3_) );
DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_260_), .Q(REGS_4__4_) );
DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_261_), .Q(REGS_4__5_) );
DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_262_), .Q(REGS_4__6_) );
DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_263_), .Q(REGS_4__7_) );
DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_264_), .Q(REGS_4__8_) );
DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_265_), .Q(REGS_4__9_) );
DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_266_), .Q(REGS_4__10_) );
DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_267_), .Q(REGS_4__11_) );
DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_268_), .Q(REGS_4__12_) );
DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_26_), .Q(FIRQ_REGS_3__10_) );
DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_269_), .Q(REGS_4__13_) );
DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_270_), .Q(REGS_4__14_) );
DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_271_), .Q(REGS_4__15_) );
DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_272_), .Q(REGS_5__0_) );
DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_273_), .Q(REGS_5__1_) );
DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_274_), .Q(REGS_5__2_) );
DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_275_), .Q(REGS_5__3_) );
DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_276_), .Q(REGS_5__4_) );
DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_277_), .Q(REGS_5__5_) );
DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_278_), .Q(REGS_5__6_) );
DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_27_), .Q(FIRQ_REGS_3__11_) );
DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_279_), .Q(REGS_5__7_) );
DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_280_), .Q(REGS_5__8_) );
DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_281_), .Q(REGS_5__9_) );
DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_282_), .Q(REGS_5__10_) );
DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_283_), .Q(REGS_5__11_) );
DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_284_), .Q(REGS_5__12_) );
DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_285_), .Q(REGS_5__13_) );
DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_286_), .Q(REGS_5__14_) );
DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_287_), .Q(REGS_5__15_) );
DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_288_), .Q(REGS_6__0_) );
DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_28_), .Q(FIRQ_REGS_3__12_) );
DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_289_), .Q(REGS_6__1_) );
DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_290_), .Q(REGS_6__2_) );
DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_291_), .Q(REGS_6__3_) );
DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_292_), .Q(REGS_6__4_) );
DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_293_), .Q(REGS_6__5_) );
DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_294_), .Q(REGS_6__6_) );
DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_295_), .Q(REGS_6__7_) );
DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_296_), .Q(REGS_6__8_) );
DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_297_), .Q(REGS_6__9_) );
DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_298_), .Q(REGS_6__10_) );
DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_34_), .Q(FIRQ_REGS_4__2_) );
DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_29_), .Q(FIRQ_REGS_3__13_) );
DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_299_), .Q(REGS_6__11_) );
DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_300_), .Q(REGS_6__12_) );
DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_301_), .Q(REGS_6__13_) );
DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_302_), .Q(REGS_6__14_) );
DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_303_), .Q(REGS_6__15_) );
DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_304_), .Q(REGS_7__0_) );
DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_305_), .Q(REGS_7__1_) );
DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_306_), .Q(REGS_7__2_) );
DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_307_), .Q(REGS_7__3_) );
DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_308_), .Q(REGS_7__4_) );
DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_30_), .Q(FIRQ_REGS_3__14_) );
DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_309_), .Q(REGS_7__5_) );
DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_310_), .Q(REGS_7__6_) );
DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_311_), .Q(REGS_7__7_) );
DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_312_), .Q(REGS_7__8_) );
DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_313_), .Q(REGS_7__9_) );
DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_314_), .Q(REGS_7__10_) );
DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_315_), .Q(REGS_7__11_) );
DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_316_), .Q(REGS_7__12_) );
DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_317_), .Q(REGS_7__13_) );
DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_318_), .Q(REGS_7__14_) );
DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_31_), .Q(FIRQ_REGS_3__15_) );
DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_319_), .Q(REGS_7__15_) );
DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_224_), .Q(REGS_2__0_) );
DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_225_), .Q(REGS_2__1_) );
DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_226_), .Q(REGS_2__2_) );
DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_227_), .Q(REGS_2__3_) );
DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_228_), .Q(REGS_2__4_) );
DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_229_), .Q(REGS_2__5_) );
DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_230_), .Q(REGS_2__6_) );
DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_231_), .Q(REGS_2__7_) );
DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_232_), .Q(REGS_2__8_) );
DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_80_), .Q(FIRQ_REGS_7__0_) );
DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_233_), .Q(REGS_2__9_) );
DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_234_), .Q(REGS_2__10_) );
DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_235_), .Q(REGS_2__11_) );
DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_236_), .Q(REGS_2__12_) );
DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_237_), .Q(REGS_2__13_) );
DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_238_), .Q(REGS_2__14_) );
DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_239_), .Q(REGS_2__15_) );
DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_96_), .Q(USR_REGS_0__0_) );
DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_97_), .Q(USR_REGS_0__1_) );
DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_98_), .Q(USR_REGS_0__2_) );
DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_81_), .Q(FIRQ_REGS_7__1_) );
DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_99_), .Q(USR_REGS_0__3_) );
DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_100_), .Q(USR_REGS_0__4_) );
DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_101_), .Q(USR_REGS_0__5_) );
DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_102_), .Q(USR_REGS_0__6_) );
DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_103_), .Q(USR_REGS_0__7_) );
DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_104_), .Q(USR_REGS_0__8_) );
DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_105_), .Q(USR_REGS_0__9_) );
DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_106_), .Q(USR_REGS_0__10_) );
DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_107_), .Q(USR_REGS_0__11_) );
DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_108_), .Q(USR_REGS_0__12_) );
DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_82_), .Q(FIRQ_REGS_7__2_) );
DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_109_), .Q(USR_REGS_0__13_) );
DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_110_), .Q(USR_REGS_0__14_) );
DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_111_), .Q(USR_REGS_0__15_) );
DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_83_), .Q(FIRQ_REGS_7__3_) );
DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_84_), .Q(FIRQ_REGS_7__4_) );
DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_85_), .Q(FIRQ_REGS_7__5_) );
DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_86_), .Q(FIRQ_REGS_7__6_) );
DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_35_), .Q(FIRQ_REGS_4__3_) );
DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_87_), .Q(FIRQ_REGS_7__7_) );
DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_88_), .Q(FIRQ_REGS_7__8_) );
DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_89_), .Q(FIRQ_REGS_7__9_) );
DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_90_), .Q(FIRQ_REGS_7__10_) );
DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_91_), .Q(FIRQ_REGS_7__11_) );
DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_92_), .Q(FIRQ_REGS_7__12_) );
DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_93_), .Q(FIRQ_REGS_7__13_) );
DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_94_), .Q(FIRQ_REGS_7__14_) );
DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_95_), .Q(FIRQ_REGS_7__15_) );
DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_64_), .Q(FIRQ_REGS_6__0_) );
DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_36_), .Q(FIRQ_REGS_4__4_) );
DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_65_), .Q(FIRQ_REGS_6__1_) );
DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_66_), .Q(FIRQ_REGS_6__2_) );
DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_67_), .Q(FIRQ_REGS_6__3_) );
DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_68_), .Q(FIRQ_REGS_6__4_) );
DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_69_), .Q(FIRQ_REGS_6__5_) );
DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_70_), .Q(FIRQ_REGS_6__6_) );
DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_71_), .Q(FIRQ_REGS_6__7_) );
DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_72_), .Q(FIRQ_REGS_6__8_) );
DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_73_), .Q(FIRQ_REGS_6__9_) );
DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_74_), .Q(FIRQ_REGS_6__10_) );
DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_37_), .Q(FIRQ_REGS_4__5_) );
DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_75_), .Q(FIRQ_REGS_6__11_) );
DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_76_), .Q(FIRQ_REGS_6__12_) );
DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_77_), .Q(FIRQ_REGS_6__13_) );
DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_78_), .Q(FIRQ_REGS_6__14_) );
DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_79_), .Q(FIRQ_REGS_6__15_) );
DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_48_), .Q(FIRQ_REGS_5__0_) );
DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_49_), .Q(FIRQ_REGS_5__1_) );
DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_50_), .Q(FIRQ_REGS_5__2_) );
DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_51_), .Q(FIRQ_REGS_5__3_) );
DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_52_), .Q(FIRQ_REGS_5__4_) );
DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_38_), .Q(FIRQ_REGS_4__6_) );
DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_53_), .Q(FIRQ_REGS_5__5_) );
DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_54_), .Q(FIRQ_REGS_5__6_) );
DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_55_), .Q(FIRQ_REGS_5__7_) );
DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_56_), .Q(FIRQ_REGS_5__8_) );
DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_57_), .Q(FIRQ_REGS_5__9_) );
DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_58_), .Q(FIRQ_REGS_5__10_) );
DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_59_), .Q(FIRQ_REGS_5__11_) );
DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_60_), .Q(FIRQ_REGS_5__12_) );
DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_61_), .Q(FIRQ_REGS_5__13_) );
DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_62_), .Q(FIRQ_REGS_5__14_) );
DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_39_), .Q(FIRQ_REGS_4__7_) );
DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_63_), .Q(FIRQ_REGS_5__15_) );
DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_320_), .Q(FIRQ_REGS_1__0_) );
DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_321_), .Q(FIRQ_REGS_1__1_) );
DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_322_), .Q(FIRQ_REGS_1__2_) );
DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_323_), .Q(FIRQ_REGS_1__3_) );
DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_324_), .Q(FIRQ_REGS_1__4_) );
DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_325_), .Q(FIRQ_REGS_1__5_) );
DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_326_), .Q(FIRQ_REGS_1__6_) );
DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_327_), .Q(FIRQ_REGS_1__7_) );
DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_328_), .Q(FIRQ_REGS_1__8_) );
DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_40_), .Q(FIRQ_REGS_4__8_) );
DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_329_), .Q(FIRQ_REGS_1__9_) );
DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_330_), .Q(FIRQ_REGS_1__10_) );
DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_331_), .Q(FIRQ_REGS_1__11_) );
DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_332_), .Q(FIRQ_REGS_1__12_) );
DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_333_), .Q(FIRQ_REGS_1__13_) );
DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_334_), .Q(FIRQ_REGS_1__14_) );
DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_335_), .Q(FIRQ_REGS_1__15_) );
DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_336_), .Q(FIRQ_REGS_0__0_) );
DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_337_), .Q(FIRQ_REGS_0__1_) );
DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_338_), .Q(FIRQ_REGS_0__2_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[2]), .Y(_1624_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__0_), .Y(_678_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__0_), .Y(_683_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__0_), .Y(_687_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__1_), .Y(_707_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__1_), .Y(_713_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__1_), .Y(_716_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__1_), .Y(_721_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__1_), .Y(_725_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__2_), .Y(_745_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__2_), .Y(_751_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[1]), .Y(_1678_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__2_), .Y(_754_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__2_), .Y(_759_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__2_), .Y(_763_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__3_), .Y(_783_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__3_), .Y(_789_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__3_), .Y(_792_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__3_), .Y(_797_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__3_), .Y(_801_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__4_), .Y(_821_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__4_), .Y(_827_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .Y(_1736_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__4_), .Y(_830_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__4_), .Y(_835_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__4_), .Y(_839_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__5_), .Y(_859_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__5_), .Y(_865_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__5_), .Y(_868_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__5_), .Y(_873_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__5_), .Y(_877_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__6_), .Y(_897_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__6_), .Y(_903_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[2]), .Y(_635_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__6_), .Y(_906_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__6_), .Y(_911_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__6_), .Y(_915_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__7_), .Y(_935_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__7_), .Y(_941_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__7_), .Y(_944_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__7_), .Y(_949_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__7_), .Y(_953_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__8_), .Y(_973_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__8_), .Y(_979_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[0]), .Y(_639_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__8_), .Y(_982_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__8_), .Y(_987_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__8_), .Y(_991_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__9_), .Y(_1011_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__9_), .Y(_1017_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__9_), .Y(_1020_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__9_), .Y(_1025_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__9_), .Y(_1029_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__10_), .Y(_1049_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__10_), .Y(_1055_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[1]), .Y(_643_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__10_), .Y(_1058_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__10_), .Y(_1063_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__10_), .Y(_1067_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__11_), .Y(_1087_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__11_), .Y(_1093_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__11_), .Y(_1096_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__11_), .Y(_1101_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__11_), .Y(_1105_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__12_), .Y(_1125_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__12_), .Y(_1131_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_656_), .Y(_657_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__12_), .Y(_1134_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__12_), .Y(_1139_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__12_), .Y(_1143_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__13_), .Y(_1163_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__13_), .Y(_1169_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__13_), .Y(_1172_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__13_), .Y(_1177_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__13_), .Y(_1181_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__14_), .Y(_1201_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__14_), .Y(_1207_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__0_), .Y(_667_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__14_), .Y(_1210_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__14_), .Y(_1215_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__14_), .Y(_1219_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__15_), .Y(_1239_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__15_), .Y(_1245_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__15_), .Y(_1248_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__15_), .Y(_1253_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__15_), .Y(_1257_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[2]), .Y(_1263_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[0]), .Y(_1267_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_0__0_), .Y(_675_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[1]), .Y(_1271_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .Y(_1285_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[0]), .Y(_1659_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__8_), .Y(_552_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__9_), .Y(_554_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__10_), .Y(_556_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__11_), .Y(_558_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__12_), .Y(_560_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__13_), .Y(_562_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__14_), .Y(_564_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__15_), .Y(_566_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__0_), .Y(_602_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__1_), .Y(_605_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__0_), .Y(_535_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__2_), .Y(_607_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__3_), .Y(_609_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__4_), .Y(_611_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__5_), .Y(_613_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__6_), .Y(_615_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__7_), .Y(_617_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__8_), .Y(_619_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__9_), .Y(_621_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__10_), .Y(_623_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__11_), .Y(_625_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__1_), .Y(_538_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__12_), .Y(_627_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__13_), .Y(_629_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__14_), .Y(_631_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(REGS_7__15_), .Y(_633_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__2_), .Y(_540_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__3_), .Y(_542_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__4_), .Y(_544_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__5_), .Y(_546_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__6_), .Y(_548_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(REGS_4__7_), .Y(_550_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_1622__bF_buf0), .Y(_1623_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(REG_D[0]), .Y(_1621_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(REG_D[9]), .Y(_1645_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(REG_D[10]), .Y(_1647_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(REG_D[11]), .Y(_1649_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(REG_D[12]), .Y(_1651_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(REG_D[13]), .Y(_1653_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(REG_D[14]), .Y(_1655_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(REG_D[15]), .Y(_1657_) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(_646_), .Y(_647_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .Y(_1275_) );
INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(REG_D[1]), .Y(_1629_) );
INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(REG_D[2]), .Y(_1631_) );
INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(REG_D[3]), .Y(_1633_) );
INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(REG_D[4]), .Y(_1635_) );
INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(REG_D[5]), .Y(_1637_) );
INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(REG_D[6]), .Y(_1639_) );
INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(REG_D[7]), .Y(_1641_) );
INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(REG_D[8]), .Y(_1643_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__0_), .B(USR_REGS_5__0_), .S(REG_Interrupt_flag_bF_buf1), .Y(_659_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__3_), .B(USR_REGS_5__3_), .S(REG_Interrupt_flag_bF_buf8), .Y(_778_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__3_), .B(USR_REGS_4__3_), .S(REG_Interrupt_flag_bF_buf8), .Y(_780_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__3_), .B(USR_REGS_6__3_), .S(REG_Interrupt_flag_bF_buf8), .Y(_782_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__4_), .B(USR_REGS_5__4_), .S(REG_Interrupt_flag_bF_buf13), .Y(_816_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__4_), .B(USR_REGS_4__4_), .S(REG_Interrupt_flag_bF_buf13), .Y(_818_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__4_), .B(USR_REGS_6__4_), .S(REG_Interrupt_flag_bF_buf13), .Y(_820_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__5_), .B(USR_REGS_5__5_), .S(REG_Interrupt_flag_bF_buf8), .Y(_854_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__5_), .B(USR_REGS_4__5_), .S(REG_Interrupt_flag_bF_buf6), .Y(_856_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__5_), .B(USR_REGS_6__5_), .S(REG_Interrupt_flag_bF_buf9), .Y(_858_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__6_), .B(USR_REGS_5__6_), .S(REG_Interrupt_flag_bF_buf8), .Y(_892_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__0_), .B(USR_REGS_4__0_), .S(REG_Interrupt_flag_bF_buf1), .Y(_662_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__6_), .B(USR_REGS_4__6_), .S(REG_Interrupt_flag_bF_buf8), .Y(_894_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__6_), .B(USR_REGS_6__6_), .S(REG_Interrupt_flag_bF_buf8), .Y(_896_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__7_), .B(USR_REGS_5__7_), .S(REG_Interrupt_flag_bF_buf13), .Y(_930_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__7_), .B(USR_REGS_4__7_), .S(REG_Interrupt_flag_bF_buf13), .Y(_932_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__7_), .B(USR_REGS_6__7_), .S(REG_Interrupt_flag_bF_buf8), .Y(_934_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__8_), .B(USR_REGS_5__8_), .S(REG_Interrupt_flag_bF_buf5), .Y(_968_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__8_), .B(USR_REGS_4__8_), .S(REG_Interrupt_flag_bF_buf5), .Y(_970_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__8_), .B(USR_REGS_6__8_), .S(REG_Interrupt_flag_bF_buf11), .Y(_972_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__9_), .B(USR_REGS_5__9_), .S(REG_Interrupt_flag_bF_buf8), .Y(_1006_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__9_), .B(USR_REGS_4__9_), .S(REG_Interrupt_flag_bF_buf13), .Y(_1008_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__0_), .B(USR_REGS_6__0_), .S(REG_Interrupt_flag_bF_buf0), .Y(_665_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__9_), .B(USR_REGS_6__9_), .S(REG_Interrupt_flag_bF_buf9), .Y(_1010_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__10_), .B(USR_REGS_5__10_), .S(REG_Interrupt_flag_bF_buf5), .Y(_1044_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__10_), .B(USR_REGS_4__10_), .S(REG_Interrupt_flag_bF_buf5), .Y(_1046_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__10_), .B(USR_REGS_6__10_), .S(REG_Interrupt_flag_bF_buf11), .Y(_1048_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__11_), .B(USR_REGS_5__11_), .S(REG_Interrupt_flag_bF_buf9), .Y(_1082_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__11_), .B(USR_REGS_4__11_), .S(REG_Interrupt_flag_bF_buf9), .Y(_1084_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__11_), .B(USR_REGS_6__11_), .S(REG_Interrupt_flag_bF_buf9), .Y(_1086_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__12_), .B(USR_REGS_5__12_), .S(REG_Interrupt_flag_bF_buf1), .Y(_1120_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__12_), .B(USR_REGS_4__12_), .S(REG_Interrupt_flag_bF_buf1), .Y(_1122_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__12_), .B(USR_REGS_6__12_), .S(REG_Interrupt_flag_bF_buf1), .Y(_1124_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__1_), .B(USR_REGS_5__1_), .S(REG_Interrupt_flag_bF_buf11), .Y(_702_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__13_), .B(USR_REGS_5__13_), .S(REG_Interrupt_flag_bF_buf5), .Y(_1158_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__13_), .B(USR_REGS_4__13_), .S(REG_Interrupt_flag_bF_buf5), .Y(_1160_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__13_), .B(USR_REGS_6__13_), .S(REG_Interrupt_flag_bF_buf1), .Y(_1162_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__14_), .B(USR_REGS_5__14_), .S(REG_Interrupt_flag_bF_buf8), .Y(_1196_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__14_), .B(USR_REGS_4__14_), .S(REG_Interrupt_flag_bF_buf8), .Y(_1198_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__14_), .B(USR_REGS_6__14_), .S(REG_Interrupt_flag_bF_buf8), .Y(_1200_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__15_), .B(USR_REGS_5__15_), .S(REG_Interrupt_flag_bF_buf1), .Y(_1234_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__15_), .B(USR_REGS_4__15_), .S(REG_Interrupt_flag_bF_buf1), .Y(_1236_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__15_), .B(USR_REGS_6__15_), .S(REG_Interrupt_flag_bF_buf11), .Y(_1238_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__1_), .B(USR_REGS_4__1_), .S(REG_Interrupt_flag_bF_buf5), .Y(_704_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__1_), .B(USR_REGS_6__1_), .S(REG_Interrupt_flag_bF_buf11), .Y(_706_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__2_), .B(USR_REGS_5__2_), .S(REG_Interrupt_flag_bF_buf1), .Y(_740_) );
MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__2_), .B(USR_REGS_4__2_), .S(REG_Interrupt_flag_bF_buf0), .Y(_742_) );
MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__2_), .B(USR_REGS_6__2_), .S(REG_Interrupt_flag_bF_buf0), .Y(_744_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[1]), .B(_1624_), .Y(_1625_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__7_), .B(_1627__bF_buf2), .Y(_1642_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__7_), .B(_362__bF_buf0), .Y(_370_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__8_), .B(_362__bF_buf1), .Y(_371_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__9_), .B(_362__bF_buf0), .Y(_372_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__10_), .B(_362__bF_buf1), .Y(_373_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__11_), .B(_362__bF_buf3), .Y(_374_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__12_), .B(_362__bF_buf2), .Y(_375_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__13_), .B(_362__bF_buf4), .Y(_376_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__14_), .B(_362__bF_buf0), .Y(_377_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__15_), .B(_362__bF_buf4), .Y(_378_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_379_), .Y(_380_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__8_), .B(_1627__bF_buf0), .Y(_1644_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__0_), .B(_380__bF_buf2), .Y(_381_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__1_), .B(_380__bF_buf3), .Y(_382_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__2_), .B(_380__bF_buf2), .Y(_383_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__3_), .B(_380__bF_buf4), .Y(_384_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__4_), .B(_380__bF_buf4), .Y(_385_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__5_), .B(_380__bF_buf2), .Y(_386_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__6_), .B(_380__bF_buf4), .Y(_387_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__7_), .B(_380__bF_buf0), .Y(_388_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__8_), .B(_380__bF_buf0), .Y(_389_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__9_), .B(_380__bF_buf4), .Y(_390_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__9_), .B(_1627__bF_buf4), .Y(_1646_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__10_), .B(_380__bF_buf3), .Y(_391_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__11_), .B(_380__bF_buf1), .Y(_392_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__12_), .B(_380__bF_buf2), .Y(_393_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__13_), .B(_380__bF_buf0), .Y(_394_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__14_), .B(_380__bF_buf1), .Y(_395_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_1__15_), .B(_380__bF_buf3), .Y(_396_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_1626_), .Y(_397_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__0_), .B(_397__bF_buf4), .Y(_398_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__1_), .B(_397__bF_buf3), .Y(_399_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__2_), .B(_397__bF_buf4), .Y(_400_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__10_), .B(_1627__bF_buf0), .Y(_1648_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__3_), .B(_397__bF_buf1), .Y(_401_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__4_), .B(_397__bF_buf2), .Y(_402_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__5_), .B(_397__bF_buf2), .Y(_403_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__6_), .B(_397__bF_buf1), .Y(_404_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__7_), .B(_397__bF_buf4), .Y(_405_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__8_), .B(_397__bF_buf0), .Y(_406_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__9_), .B(_397__bF_buf3), .Y(_407_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__10_), .B(_397__bF_buf0), .Y(_408_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__11_), .B(_397__bF_buf1), .Y(_409_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__12_), .B(_397__bF_buf3), .Y(_410_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__11_), .B(_1627__bF_buf4), .Y(_1650_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__13_), .B(_397__bF_buf0), .Y(_411_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__14_), .B(_397__bF_buf2), .Y(_412_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_2__15_), .B(_397__bF_buf4), .Y(_413_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_1660_), .Y(_414_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__0_), .B(_414__bF_buf3), .Y(_415_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__1_), .B(_414__bF_buf1), .Y(_416_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__2_), .B(_414__bF_buf3), .Y(_417_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__3_), .B(_414__bF_buf0), .Y(_418_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__4_), .B(_414__bF_buf4), .Y(_419_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__5_), .B(_414__bF_buf3), .Y(_420_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__12_), .B(_1627__bF_buf1), .Y(_1652_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__6_), .B(_414__bF_buf0), .Y(_421_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__7_), .B(_414__bF_buf4), .Y(_422_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__8_), .B(_414__bF_buf2), .Y(_423_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__9_), .B(_414__bF_buf0), .Y(_424_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__10_), .B(_414__bF_buf2), .Y(_425_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__11_), .B(_414__bF_buf3), .Y(_426_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__12_), .B(_414__bF_buf2), .Y(_427_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__13_), .B(_414__bF_buf1), .Y(_428_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__14_), .B(_414__bF_buf4), .Y(_429_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_3__15_), .B(_414__bF_buf1), .Y(_430_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__13_), .B(_1627__bF_buf0), .Y(_1654_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_1680_), .Y(_431_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__0_), .B(_431__bF_buf4), .Y(_432_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__1_), .B(_431__bF_buf1), .Y(_433_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__2_), .B(_431__bF_buf1), .Y(_434_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__3_), .B(_431__bF_buf3), .Y(_435_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__4_), .B(_431__bF_buf0), .Y(_436_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__5_), .B(_431__bF_buf3), .Y(_437_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__6_), .B(_431__bF_buf3), .Y(_438_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__7_), .B(_431__bF_buf0), .Y(_439_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__8_), .B(_431__bF_buf2), .Y(_440_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__14_), .B(_1627__bF_buf4), .Y(_1656_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__9_), .B(_431__bF_buf0), .Y(_441_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__10_), .B(_431__bF_buf2), .Y(_442_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__11_), .B(_431__bF_buf4), .Y(_443_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__12_), .B(_431__bF_buf4), .Y(_444_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__13_), .B(_431__bF_buf2), .Y(_445_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__14_), .B(_431__bF_buf3), .Y(_446_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_4__15_), .B(_431__bF_buf1), .Y(_447_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_1698_), .Y(_448_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__0_), .B(_448__bF_buf0), .Y(_449_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__1_), .B(_448__bF_buf3), .Y(_450_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__15_), .B(_1627__bF_buf1), .Y(_1658_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__2_), .B(_448__bF_buf4), .Y(_451_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__3_), .B(_448__bF_buf2), .Y(_452_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__4_), .B(_448__bF_buf2), .Y(_453_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__5_), .B(_448__bF_buf0), .Y(_454_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__6_), .B(_448__bF_buf1), .Y(_455_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__7_), .B(_448__bF_buf2), .Y(_456_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__8_), .B(_448__bF_buf3), .Y(_457_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__9_), .B(_448__bF_buf1), .Y(_458_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__10_), .B(_448__bF_buf4), .Y(_459_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__11_), .B(_448__bF_buf0), .Y(_460_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1660_), .Y(_1661_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__12_), .B(_448__bF_buf0), .Y(_461_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__13_), .B(_448__bF_buf4), .Y(_462_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__14_), .B(_448__bF_buf1), .Y(_463_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_5__15_), .B(_448__bF_buf3), .Y(_464_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(_359_), .Y(_465_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__0_), .B(_465__bF_buf1), .Y(_466_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__1_), .B(_465__bF_buf0), .Y(_467_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__2_), .B(_465__bF_buf2), .Y(_468_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__3_), .B(_465__bF_buf4), .Y(_469_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__4_), .B(_465__bF_buf3), .Y(_470_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1626_), .Y(_1627_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__0_), .B(_1661__bF_buf1), .Y(_1662_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__5_), .B(_465__bF_buf3), .Y(_471_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__6_), .B(_465__bF_buf4), .Y(_472_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__7_), .B(_465__bF_buf3), .Y(_473_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__8_), .B(_465__bF_buf0), .Y(_474_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__9_), .B(_465__bF_buf2), .Y(_475_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__10_), .B(_465__bF_buf1), .Y(_476_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__11_), .B(_465__bF_buf4), .Y(_477_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__12_), .B(_465__bF_buf2), .Y(_478_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__13_), .B(_465__bF_buf1), .Y(_479_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__14_), .B(_465__bF_buf3), .Y(_480_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__1_), .B(_1661__bF_buf0), .Y(_1663_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_6__15_), .B(_465__bF_buf0), .Y(_481_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_1736_), .Y(_482_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__0_), .B(_482__bF_buf3), .Y(_483_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__1_), .B(_482__bF_buf4), .Y(_484_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__2_), .B(_482__bF_buf3), .Y(_485_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__3_), .B(_482__bF_buf0), .Y(_486_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__4_), .B(_482__bF_buf0), .Y(_487_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__5_), .B(_482__bF_buf1), .Y(_488_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__6_), .B(_482__bF_buf1), .Y(_489_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__7_), .B(_482__bF_buf1), .Y(_490_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__2_), .B(_1661__bF_buf3), .Y(_1664_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__8_), .B(_482__bF_buf4), .Y(_491_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__9_), .B(_482__bF_buf3), .Y(_492_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__10_), .B(_482__bF_buf2), .Y(_493_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__11_), .B(_482__bF_buf0), .Y(_494_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__12_), .B(_482__bF_buf2), .Y(_495_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__13_), .B(_482__bF_buf2), .Y(_496_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__14_), .B(_482__bF_buf3), .Y(_497_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_7__15_), .B(_482__bF_buf4), .Y(_498_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(REG_D[0]), .B(_536__bF_buf2), .Y(_537_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(REG_D[1]), .B(_536__bF_buf4), .Y(_539_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__3_), .B(_1661__bF_buf4), .Y(_1665_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(REG_D[2]), .B(_536__bF_buf1), .Y(_541_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(REG_D[3]), .B(_536__bF_buf0), .Y(_543_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(REG_D[4]), .B(_536__bF_buf0), .Y(_545_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(REG_D[5]), .B(_536__bF_buf0), .Y(_547_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(REG_D[6]), .B(_536__bF_buf3), .Y(_549_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(REG_D[7]), .B(_536__bF_buf3), .Y(_551_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(REG_D[8]), .B(_536__bF_buf1), .Y(_553_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(REG_D[9]), .B(_536__bF_buf3), .Y(_555_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(REG_D[10]), .B(_536__bF_buf1), .Y(_557_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(REG_D[11]), .B(_536__bF_buf2), .Y(_559_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__4_), .B(_1661__bF_buf2), .Y(_1666_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(REG_D[12]), .B(_536__bF_buf1), .Y(_561_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(REG_D[13]), .B(_536__bF_buf4), .Y(_563_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(REG_D[14]), .B(_536__bF_buf3), .Y(_565_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(REG_D[15]), .B(_536__bF_buf4), .Y(_567_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(REG_D[0]), .B(_603__bF_buf2), .Y(_604_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(REG_D[1]), .B(_603__bF_buf4), .Y(_606_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(REG_D[2]), .B(_603__bF_buf2), .Y(_608_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(REG_D[3]), .B(_603__bF_buf0), .Y(_610_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(REG_D[4]), .B(_603__bF_buf0), .Y(_612_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(REG_D[5]), .B(_603__bF_buf1), .Y(_614_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__5_), .B(_1661__bF_buf2), .Y(_1667_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(REG_D[6]), .B(_603__bF_buf3), .Y(_616_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(REG_D[7]), .B(_603__bF_buf3), .Y(_618_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(REG_D[8]), .B(_603__bF_buf2), .Y(_620_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(REG_D[9]), .B(_603__bF_buf3), .Y(_622_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(REG_D[10]), .B(_603__bF_buf2), .Y(_624_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(REG_D[11]), .B(_603__bF_buf0), .Y(_626_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(REG_D[12]), .B(_603__bF_buf1), .Y(_628_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(REG_D[13]), .B(_603__bF_buf4), .Y(_630_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(REG_D[14]), .B(_603__bF_buf3), .Y(_632_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(REG_D[15]), .B(_603__bF_buf4), .Y(_634_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__6_), .B(_1661__bF_buf2), .Y(_1668_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_637_), .B(_636__bF_buf4), .Y(_638_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[1]), .B(REG_RF2[0]), .Y(_646_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf4), .B(_636__bF_buf1), .Y(_648_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[3]), .B(REG_RF2[2]), .Y(_656_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_640__bF_buf3), .Y(_658_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_637_), .B(_657_), .Y(_661_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_644__bF_buf0), .Y(_664_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(FIRQ_REGS_7__0_), .Y(_668_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_666_), .Y(_670_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_637_), .B(_673__bF_buf1), .Y(_674_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__7_), .B(_1661__bF_buf3), .Y(_1669_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(_675_), .Y(_676_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_1__0_), .Y(_679_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(FIRQ_REGS_3__0_), .Y(_684_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_2__0_), .Y(_688_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_690_), .Y(_691_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf11), .B(FIRQ_REGS_7__1_), .Y(_708_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_666_), .Y(_710_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(_713_), .Y(_714_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_1__1_), .Y(_717_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf5), .B(FIRQ_REGS_3__1_), .Y(_722_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__8_), .B(_1661__bF_buf1), .Y(_1670_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf1), .B(FIRQ_REGS_2__1_), .Y(_726_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_728_), .Y(_729_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(FIRQ_REGS_7__2_), .Y(_746_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_666_), .Y(_748_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(_751_), .Y(_752_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_1__2_), .Y(_755_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_3__2_), .Y(_760_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(FIRQ_REGS_2__2_), .Y(_764_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_766_), .Y(_767_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf8), .B(FIRQ_REGS_7__3_), .Y(_784_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__9_), .B(_1661__bF_buf4), .Y(_1671_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_666_), .Y(_786_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf13), .B(_789_), .Y(_790_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf13), .B(FIRQ_REGS_1__3_), .Y(_793_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf13), .B(FIRQ_REGS_3__3_), .Y(_798_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_2__3_), .Y(_802_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_804_), .Y(_805_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf9), .B(FIRQ_REGS_7__4_), .Y(_822_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_823_), .B(_666_), .Y(_824_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(_827_), .Y(_828_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf13), .B(FIRQ_REGS_1__4_), .Y(_831_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__0_), .B(_1627__bF_buf2), .Y(_1628_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__10_), .B(_1661__bF_buf0), .Y(_1672_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_3__4_), .Y(_836_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_2__4_), .Y(_840_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(_842_), .Y(_843_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf9), .B(FIRQ_REGS_7__5_), .Y(_860_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_861_), .B(_666_), .Y(_862_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(_865_), .Y(_866_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_1__5_), .Y(_869_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_3__5_), .Y(_874_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_2__5_), .Y(_878_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_880_), .Y(_881_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__11_), .B(_1661__bF_buf3), .Y(_1673_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf9), .B(FIRQ_REGS_7__6_), .Y(_898_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_666_), .Y(_900_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(_903_), .Y(_904_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_1__6_), .Y(_907_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_3__6_), .Y(_912_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_2__6_), .Y(_916_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_918_), .Y(_919_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf9), .B(FIRQ_REGS_7__7_), .Y(_936_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_666_), .Y(_938_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf13), .B(_941_), .Y(_942_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__12_), .B(_1661__bF_buf3), .Y(_1674_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(FIRQ_REGS_1__7_), .Y(_945_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_3__7_), .Y(_950_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_2__7_), .Y(_954_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_956_), .Y(_957_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf11), .B(FIRQ_REGS_7__8_), .Y(_974_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_666_), .Y(_976_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(_979_), .Y(_980_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(FIRQ_REGS_1__8_), .Y(_983_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf5), .B(FIRQ_REGS_3__8_), .Y(_988_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf5), .B(FIRQ_REGS_2__8_), .Y(_992_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__13_), .B(_1661__bF_buf0), .Y(_1675_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_994_), .Y(_995_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(FIRQ_REGS_7__9_), .Y(_1012_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_666_), .Y(_1014_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(_1017_), .Y(_1018_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(FIRQ_REGS_1__9_), .Y(_1021_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_3__9_), .Y(_1026_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(FIRQ_REGS_2__9_), .Y(_1030_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1032_), .Y(_1033_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf11), .B(FIRQ_REGS_7__10_), .Y(_1050_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_666_), .Y(_1052_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__14_), .B(_1661__bF_buf4), .Y(_1676_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(_1055_), .Y(_1056_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_1__10_), .Y(_1059_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf5), .B(FIRQ_REGS_3__10_), .Y(_1064_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf5), .B(FIRQ_REGS_2__10_), .Y(_1068_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1066_), .B(_1070_), .Y(_1071_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf9), .B(FIRQ_REGS_7__11_), .Y(_1088_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_666_), .Y(_1090_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(_1093_), .Y(_1094_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_1__11_), .Y(_1097_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf4), .B(FIRQ_REGS_3__11_), .Y(_1102_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_3__15_), .B(_1661__bF_buf1), .Y(_1677_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_2__11_), .Y(_1106_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_1108_), .Y(_1109_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(FIRQ_REGS_7__12_), .Y(_1126_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_666_), .Y(_1128_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(_1131_), .Y(_1132_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(FIRQ_REGS_1__12_), .Y(_1135_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf1), .B(FIRQ_REGS_3__12_), .Y(_1140_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_2__12_), .Y(_1144_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_1146_), .Y(_1147_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf11), .B(FIRQ_REGS_7__13_), .Y(_1164_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[2]), .B(_1678_), .Y(_1679_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_666_), .Y(_1166_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(_1169_), .Y(_1170_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(FIRQ_REGS_1__13_), .Y(_1173_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_3__13_), .Y(_1178_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf5), .B(FIRQ_REGS_2__13_), .Y(_1182_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(_1184_), .Y(_1185_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(FIRQ_REGS_7__14_), .Y(_1202_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_666_), .Y(_1204_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(_1207_), .Y(_1208_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_1__14_), .Y(_1211_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1680_), .Y(_1681_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf2), .B(FIRQ_REGS_3__14_), .Y(_1216_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf6), .B(FIRQ_REGS_2__14_), .Y(_1220_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1218_), .B(_1222_), .Y(_1223_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf11), .B(FIRQ_REGS_7__15_), .Y(_1240_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_666_), .Y(_1242_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(_1245_), .Y(_1246_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_1__15_), .Y(_1249_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_3__15_), .Y(_1254_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf10), .B(FIRQ_REGS_2__15_), .Y(_1258_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1260_), .Y(_1261_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__0_), .B(_1681__bF_buf4), .Y(_1682_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1264__bF_buf3), .Y(_1266_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[1]), .B(REG_RF1[0]), .Y(_1274_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf3), .B(_1264__bF_buf0), .Y(_1276_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[3]), .B(REG_RF1[2]), .Y(_1284_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1268__bF_buf5), .Y(_1286_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1285_), .Y(_1287_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1272__bF_buf3), .Y(_1289_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_1290_), .Y(_1291_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1294__bF_buf3), .Y(_1295_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1299_), .Y(_1300_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__1_), .B(_1681__bF_buf1), .Y(_1683_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_1290_), .Y(_1312_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_1318_), .Y(_1319_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_1290_), .Y(_1331_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1337_), .Y(_1338_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_1290_), .Y(_1350_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1355_), .B(_1356_), .Y(_1357_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_823_), .B(_1290_), .Y(_1369_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .B(_1375_), .Y(_1376_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_861_), .B(_1290_), .Y(_1388_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1393_), .B(_1394_), .Y(_1395_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__1_), .B(_1627__bF_buf1), .Y(_1630_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__2_), .B(_1681__bF_buf4), .Y(_1684_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_1290_), .Y(_1407_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1413_), .Y(_1414_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_1290_), .Y(_1426_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1431_), .B(_1432_), .Y(_1433_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_1290_), .Y(_1445_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1451_), .Y(_1452_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_1290_), .Y(_1464_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1470_), .Y(_1471_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1290_), .Y(_1483_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1489_), .Y(_1490_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__3_), .B(_1681__bF_buf0), .Y(_1685_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1290_), .Y(_1502_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .B(_1508_), .Y(_1509_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1290_), .Y(_1521_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_1527_), .Y(_1528_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1290_), .Y(_1540_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1546_), .Y(_1547_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_1290_), .Y(_1559_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1565_), .Y(_1566_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1290_), .Y(_1578_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1583_), .B(_1584_), .Y(_1585_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__4_), .B(_1681__bF_buf3), .Y(_1686_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_379_), .Y(_1587_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__0_), .B(_1587__bF_buf0), .Y(_1588_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__1_), .B(_1587__bF_buf2), .Y(_1589_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__2_), .B(_1587__bF_buf4), .Y(_1590_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__3_), .B(_1587__bF_buf3), .Y(_1591_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__4_), .B(_1587__bF_buf3), .Y(_1592_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__5_), .B(_1587__bF_buf3), .Y(_1593_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__6_), .B(_1587__bF_buf4), .Y(_1594_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__7_), .B(_1587__bF_buf1), .Y(_1595_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__8_), .B(_1587__bF_buf1), .Y(_1596_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__5_), .B(_1681__bF_buf4), .Y(_1687_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__9_), .B(_1587__bF_buf3), .Y(_1597_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__10_), .B(_1587__bF_buf2), .Y(_1598_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__11_), .B(_1587__bF_buf4), .Y(_1599_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__12_), .B(_1587__bF_buf0), .Y(_1600_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__13_), .B(_1587__bF_buf1), .Y(_1601_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__14_), .B(_1587__bF_buf0), .Y(_1602_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_1__15_), .B(_1587__bF_buf2), .Y(_1603_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(REG_D[0]), .B(_1604__bF_buf4), .Y(_1605_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(REG_D[1]), .B(_1604__bF_buf3), .Y(_1606_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(REG_D[2]), .B(_1604__bF_buf4), .Y(_1607_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__6_), .B(_1681__bF_buf0), .Y(_1688_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(REG_D[3]), .B(_1604__bF_buf1), .Y(_1608_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(REG_D[4]), .B(_1604__bF_buf1), .Y(_1609_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(REG_D[5]), .B(_1604__bF_buf0), .Y(_1610_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(REG_D[6]), .B(_1604__bF_buf0), .Y(_1611_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(REG_D[7]), .B(_1604__bF_buf1), .Y(_1612_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(REG_D[8]), .B(_1604__bF_buf3), .Y(_1613_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(REG_D[9]), .B(_1604__bF_buf2), .Y(_1614_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(REG_D[10]), .B(_1604__bF_buf4), .Y(_1615_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(REG_D[11]), .B(_1604__bF_buf2), .Y(_1616_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(REG_D[12]), .B(_1604__bF_buf0), .Y(_1617_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__7_), .B(_1681__bF_buf3), .Y(_1689_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(REG_D[13]), .B(_1604__bF_buf3), .Y(_1618_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(REG_D[14]), .B(_1604__bF_buf2), .Y(_1619_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(REG_D[15]), .B(_1604__bF_buf3), .Y(_1620_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__8_), .B(_1681__bF_buf1), .Y(_1690_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__9_), .B(_1681__bF_buf3), .Y(_1691_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__10_), .B(_1681__bF_buf2), .Y(_1692_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__11_), .B(_1681__bF_buf4), .Y(_1693_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__2_), .B(_1627__bF_buf2), .Y(_1632_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__12_), .B(_1681__bF_buf2), .Y(_1694_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__13_), .B(_1681__bF_buf1), .Y(_1695_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__14_), .B(_1681__bF_buf0), .Y(_1696_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_4__15_), .B(_1681__bF_buf2), .Y(_1697_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1698_), .Y(_1699_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__0_), .B(_1699__bF_buf0), .Y(_1700_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__1_), .B(_1699__bF_buf0), .Y(_1701_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__2_), .B(_1699__bF_buf2), .Y(_1702_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__3_), .B(_1699__bF_buf3), .Y(_1703_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__4_), .B(_1699__bF_buf3), .Y(_1704_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__3_), .B(_1627__bF_buf3), .Y(_1634_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__5_), .B(_1699__bF_buf4), .Y(_1705_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__6_), .B(_1699__bF_buf4), .Y(_1706_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__7_), .B(_1699__bF_buf3), .Y(_1707_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__8_), .B(_1699__bF_buf0), .Y(_1708_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__9_), .B(_1699__bF_buf4), .Y(_1709_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__10_), .B(_1699__bF_buf2), .Y(_1710_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__11_), .B(_1699__bF_buf1), .Y(_1711_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__12_), .B(_1699__bF_buf1), .Y(_1712_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__13_), .B(_1699__bF_buf2), .Y(_1713_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__14_), .B(_1699__bF_buf4), .Y(_1714_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__4_), .B(_1627__bF_buf3), .Y(_1636_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_5__15_), .B(_1699__bF_buf1), .Y(_1715_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[1]), .B(REG_RFD[2]), .Y(_1716_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1717_), .Y(_1718_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__0_), .B(_1718__bF_buf3), .Y(_1719_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__1_), .B(_1718__bF_buf2), .Y(_1720_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__2_), .B(_1718__bF_buf1), .Y(_1721_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__3_), .B(_1718__bF_buf0), .Y(_1722_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__4_), .B(_1718__bF_buf4), .Y(_1723_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__5_), .B(_1718__bF_buf4), .Y(_1724_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__6_), .B(_1718__bF_buf0), .Y(_1725_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__5_), .B(_1627__bF_buf3), .Y(_1638_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__7_), .B(_1718__bF_buf0), .Y(_1726_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__8_), .B(_1718__bF_buf2), .Y(_1727_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__9_), .B(_1718__bF_buf1), .Y(_1728_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__10_), .B(_1718__bF_buf3), .Y(_1729_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__11_), .B(_1718__bF_buf1), .Y(_1730_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__12_), .B(_1718__bF_buf1), .Y(_1731_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__13_), .B(_1718__bF_buf3), .Y(_1732_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__14_), .B(_1718__bF_buf4), .Y(_1733_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_6__15_), .B(_1718__bF_buf2), .Y(_1734_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1736_), .Y(_1737_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(FIRQ_REGS_2__6_), .B(_1627__bF_buf3), .Y(_1640_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[3]), .B(REG_Write), .Y(_358_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1678_), .B(_1624_), .Y(_360_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_361_), .Y(_362_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__0_), .B(_362__bF_buf4), .Y(_363_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__1_), .B(_362__bF_buf4), .Y(_364_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__2_), .B(_362__bF_buf1), .Y(_365_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__3_), .B(_362__bF_buf3), .Y(_366_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__4_), .B(_362__bF_buf3), .Y(_367_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__5_), .B(_362__bF_buf2), .Y(_368_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(USR_REGS_0__6_), .B(_362__bF_buf2), .Y(_369_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[3]), .B(REG_Write), .C(REG_Interrupt_flag_bF_buf0), .Y(_1622_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_689_), .C(_673__bF_buf4), .Y(_690_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf0), .B(_1031_), .C(_673__bF_buf1), .Y(_1032_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_1034_), .C(_1005_), .Y(_1749__9_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__10_), .B(_636__bF_buf2), .C(_640__bF_buf4), .Y(_1035_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__10_), .B(_636__bF_buf2), .C(_644__bF_buf6), .Y(_1037_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__10_), .B(_650__bF_buf3), .C(_647__bF_buf3), .Y(_1039_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[10]), .B(_650__bF_buf3), .C(_640__bF_buf4), .Y(_1040_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__10_), .B(_650__bF_buf3), .C(_644__bF_buf3), .Y(_1041_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1040_), .C(_1041_), .Y(_1042_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_1060_), .C(_673__bF_buf5), .Y(_1061_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf0), .B(_1065_), .C(_673__bF_buf3), .Y(_1066_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_692_), .C(_655_), .Y(_1749__0_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_1069_), .C(_673__bF_buf3), .Y(_1070_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1054_), .B(_1072_), .C(_1043_), .Y(_1749__10_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__11_), .B(_636__bF_buf1), .C(_640__bF_buf5), .Y(_1073_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__11_), .B(_636__bF_buf1), .C(_644__bF_buf4), .Y(_1075_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__11_), .B(_650__bF_buf4), .C(_647__bF_buf4), .Y(_1077_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[11]), .B(_650__bF_buf0), .C(_640__bF_buf6), .Y(_1078_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__11_), .B(_650__bF_buf0), .C(_644__bF_buf4), .Y(_1079_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1078_), .C(_1079_), .Y(_1080_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf0), .B(_1098_), .C(_673__bF_buf1), .Y(_1099_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_1103_), .C(_673__bF_buf1), .Y(_1104_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__1_), .B(_636__bF_buf3), .C(_640__bF_buf2), .Y(_693_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf0), .B(_1107_), .C(_673__bF_buf1), .Y(_1108_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .B(_1110_), .C(_1081_), .Y(_1749__11_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__12_), .B(_636__bF_buf2), .C(_640__bF_buf4), .Y(_1111_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__12_), .B(_636__bF_buf2), .C(_644__bF_buf6), .Y(_1113_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__12_), .B(_650__bF_buf3), .C(_647__bF_buf3), .Y(_1115_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[12]), .B(_650__bF_buf0), .C(_640__bF_buf4), .Y(_1116_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__12_), .B(_650__bF_buf0), .C(_644__bF_buf3), .Y(_1117_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1116_), .C(_1117_), .Y(_1118_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_1136_), .C(_673__bF_buf4), .Y(_1137_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf0), .B(_1141_), .C(_673__bF_buf4), .Y(_1142_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__1_), .B(_636__bF_buf3), .C(_644__bF_buf6), .Y(_695_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_1145_), .C(_673__bF_buf4), .Y(_1146_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1148_), .C(_1119_), .Y(_1749__12_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__13_), .B(_636__bF_buf3), .C(_640__bF_buf2), .Y(_1149_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__13_), .B(_636__bF_buf3), .C(_644__bF_buf6), .Y(_1151_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__13_), .B(_650__bF_buf2), .C(_647__bF_buf3), .Y(_1153_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[13]), .B(_650__bF_buf2), .C(_640__bF_buf2), .Y(_1154_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__13_), .B(_650__bF_buf2), .C(_644__bF_buf3), .Y(_1155_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1154_), .C(_1155_), .Y(_1156_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_1174_), .C(_673__bF_buf5), .Y(_1175_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf0), .B(_1179_), .C(_673__bF_buf3), .Y(_1180_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__1_), .B(_650__bF_buf0), .C(_647__bF_buf3), .Y(_697_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_1183_), .C(_673__bF_buf3), .Y(_1184_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1186_), .C(_1157_), .Y(_1749__13_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__14_), .B(_636__bF_buf0), .C(_640__bF_buf5), .Y(_1187_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__14_), .B(_636__bF_buf0), .C(_644__bF_buf1), .Y(_1189_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__14_), .B(_650__bF_buf5), .C(_647__bF_buf4), .Y(_1191_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[14]), .B(_650__bF_buf4), .C(_640__bF_buf6), .Y(_1192_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__14_), .B(_650__bF_buf4), .C(_644__bF_buf4), .Y(_1193_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(_1192_), .C(_1193_), .Y(_1194_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf3), .B(_1212_), .C(_673__bF_buf0), .Y(_1213_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_1217_), .C(_673__bF_buf2), .Y(_1218_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[1]), .B(_650__bF_buf2), .C(_640__bF_buf2), .Y(_698_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf0), .B(_1221_), .C(_673__bF_buf0), .Y(_1222_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1206_), .B(_1224_), .C(_1195_), .Y(_1749__14_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__15_), .B(_636__bF_buf3), .C(_640__bF_buf2), .Y(_1225_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__15_), .B(_636__bF_buf3), .C(_644__bF_buf6), .Y(_1227_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__15_), .B(_650__bF_buf2), .C(_647__bF_buf3), .Y(_1229_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[15]), .B(_650__bF_buf2), .C(_640__bF_buf2), .Y(_1230_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__15_), .B(_650__bF_buf2), .C(_644__bF_buf3), .Y(_1231_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .B(_1230_), .C(_1231_), .Y(_1232_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_1250_), .C(_673__bF_buf5), .Y(_1251_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf0), .B(_1255_), .C(_673__bF_buf5), .Y(_1256_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__1_), .B(_650__bF_buf2), .C(_644__bF_buf3), .Y(_699_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_1259_), .C(_673__bF_buf4), .Y(_1260_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1262_), .C(_1233_), .Y(_1749__15_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__0_), .B(_1264__bF_buf2), .C(_1268__bF_buf3), .Y(_1269_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__0_), .B(_1264__bF_buf3), .C(_1272__bF_buf6), .Y(_1273_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__0_), .B(_1278__bF_buf1), .C(_1275__bF_buf1), .Y(_1279_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[0]), .B(_1278__bF_buf5), .C(_1268__bF_buf0), .Y(_1280_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__0_), .B(_1278__bF_buf1), .C(_1272__bF_buf1), .Y(_1281_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1280_), .C(_1281_), .Y(_1282_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf4), .B(_680_), .C(_1294__bF_buf0), .Y(_1296_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_685_), .C(_1294__bF_buf3), .Y(_1298_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_698_), .C(_699_), .Y(_700_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf5), .B(_689_), .C(_1294__bF_buf3), .Y(_1299_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1301_), .C(_1283_), .Y(_1748__0_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__1_), .B(_1264__bF_buf2), .C(_1268__bF_buf3), .Y(_1302_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__1_), .B(_1264__bF_buf2), .C(_1272__bF_buf6), .Y(_1304_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__1_), .B(_1278__bF_buf5), .C(_1275__bF_buf1), .Y(_1306_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[1]), .B(_1278__bF_buf5), .C(_1268__bF_buf0), .Y(_1307_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__1_), .B(_1278__bF_buf5), .C(_1272__bF_buf1), .Y(_1308_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1307_), .C(_1308_), .Y(_1309_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf5), .B(_718_), .C(_1294__bF_buf3), .Y(_1315_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_723_), .C(_1294__bF_buf2), .Y(_1317_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_718_), .C(_673__bF_buf5), .Y(_719_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf3), .B(_727_), .C(_1294__bF_buf1), .Y(_1318_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1320_), .C(_1310_), .Y(_1748__1_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__2_), .B(_1264__bF_buf1), .C(_1268__bF_buf4), .Y(_1321_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__2_), .B(_1264__bF_buf1), .C(_1272__bF_buf5), .Y(_1323_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__2_), .B(_1278__bF_buf2), .C(_1275__bF_buf4), .Y(_1325_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[2]), .B(_1278__bF_buf2), .C(_1268__bF_buf0), .Y(_1326_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__2_), .B(_1278__bF_buf4), .C(_1272__bF_buf5), .Y(_1327_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1326_), .C(_1327_), .Y(_1328_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf4), .B(_756_), .C(_1294__bF_buf0), .Y(_1334_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf4), .B(_761_), .C(_1294__bF_buf0), .Y(_1336_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf0), .B(_723_), .C(_673__bF_buf3), .Y(_724_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf5), .B(_765_), .C(_1294__bF_buf0), .Y(_1337_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1333_), .B(_1339_), .C(_1329_), .Y(_1748__2_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__3_), .B(_1264__bF_buf4), .C(_1268__bF_buf6), .Y(_1340_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__3_), .B(_1264__bF_buf4), .C(_1272__bF_buf2), .Y(_1342_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__3_), .B(_1278__bF_buf0), .C(_1275__bF_buf3), .Y(_1344_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[3]), .B(_1278__bF_buf0), .C(_1268__bF_buf1), .Y(_1345_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__3_), .B(_1278__bF_buf0), .C(_1272__bF_buf4), .Y(_1346_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_1345_), .C(_1346_), .Y(_1347_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_794_), .C(_1294__bF_buf6), .Y(_1353_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf0), .B(_799_), .C(_1294__bF_buf4), .Y(_1355_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__0_), .B(_636__bF_buf3), .C(_640__bF_buf4), .Y(_641_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_727_), .C(_673__bF_buf5), .Y(_728_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_803_), .C(_1294__bF_buf4), .Y(_1356_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1358_), .C(_1348_), .Y(_1748__3_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__4_), .B(_1264__bF_buf0), .C(_1268__bF_buf6), .Y(_1359_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__4_), .B(_1264__bF_buf0), .C(_1272__bF_buf4), .Y(_1361_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__4_), .B(_1278__bF_buf0), .C(_1275__bF_buf3), .Y(_1363_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[4]), .B(_1278__bF_buf3), .C(_1268__bF_buf1), .Y(_1364_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__4_), .B(_1278__bF_buf3), .C(_1272__bF_buf4), .Y(_1365_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1364_), .C(_1365_), .Y(_1366_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_832_), .C(_1294__bF_buf6), .Y(_1372_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf0), .B(_837_), .C(_1294__bF_buf4), .Y(_1374_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_730_), .C(_701_), .Y(_1749__1_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_841_), .C(_1294__bF_buf4), .Y(_1375_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1371_), .B(_1377_), .C(_1367_), .Y(_1748__4_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__5_), .B(_1264__bF_buf0), .C(_1268__bF_buf1), .Y(_1378_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__5_), .B(_1264__bF_buf4), .C(_1272__bF_buf2), .Y(_1380_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__5_), .B(_1278__bF_buf3), .C(_1275__bF_buf3), .Y(_1382_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[5]), .B(_1278__bF_buf3), .C(_1268__bF_buf1), .Y(_1383_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__5_), .B(_1278__bF_buf3), .C(_1272__bF_buf4), .Y(_1384_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1383_), .C(_1384_), .Y(_1385_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf4), .B(_870_), .C(_1294__bF_buf0), .Y(_1391_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf4), .B(_875_), .C(_1294__bF_buf0), .Y(_1393_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__2_), .B(_636__bF_buf4), .C(_640__bF_buf0), .Y(_731_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf5), .B(_879_), .C(_1294__bF_buf0), .Y(_1394_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1396_), .C(_1386_), .Y(_1748__5_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__6_), .B(_1264__bF_buf4), .C(_1268__bF_buf6), .Y(_1397_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__6_), .B(_1264__bF_buf4), .C(_1272__bF_buf2), .Y(_1399_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__6_), .B(_1278__bF_buf4), .C(_1275__bF_buf4), .Y(_1401_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[6]), .B(_1278__bF_buf4), .C(_1268__bF_buf6), .Y(_1402_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__6_), .B(_1278__bF_buf4), .C(_1272__bF_buf2), .Y(_1403_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1401_), .B(_1402_), .C(_1403_), .Y(_1404_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_908_), .C(_1294__bF_buf6), .Y(_1410_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf0), .B(_913_), .C(_1294__bF_buf4), .Y(_1412_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__2_), .B(_636__bF_buf4), .C(_644__bF_buf2), .Y(_733_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_917_), .C(_1294__bF_buf4), .Y(_1413_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(_1415_), .C(_1405_), .Y(_1748__6_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__7_), .B(_1264__bF_buf0), .C(_1268__bF_buf1), .Y(_1416_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__7_), .B(_1264__bF_buf0), .C(_1272__bF_buf4), .Y(_1418_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__7_), .B(_1278__bF_buf0), .C(_1275__bF_buf3), .Y(_1420_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[7]), .B(_1278__bF_buf0), .C(_1268__bF_buf1), .Y(_1421_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__7_), .B(_1278__bF_buf0), .C(_1272__bF_buf4), .Y(_1422_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1421_), .C(_1422_), .Y(_1423_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_946_), .C(_1294__bF_buf5), .Y(_1429_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf4), .B(_951_), .C(_1294__bF_buf5), .Y(_1431_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__2_), .B(_650__bF_buf1), .C(_647__bF_buf1), .Y(_735_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_955_), .C(_1294__bF_buf5), .Y(_1432_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1428_), .B(_1434_), .C(_1424_), .Y(_1748__7_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__8_), .B(_1264__bF_buf3), .C(_1268__bF_buf3), .Y(_1435_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__8_), .B(_1264__bF_buf3), .C(_1272__bF_buf6), .Y(_1437_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__8_), .B(_1278__bF_buf1), .C(_1275__bF_buf1), .Y(_1439_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[8]), .B(_1278__bF_buf1), .C(_1268__bF_buf3), .Y(_1440_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__8_), .B(_1278__bF_buf1), .C(_1272__bF_buf6), .Y(_1441_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1440_), .C(_1441_), .Y(_1442_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf5), .B(_984_), .C(_1294__bF_buf3), .Y(_1448_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_989_), .C(_1294__bF_buf2), .Y(_1450_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[2]), .B(_650__bF_buf3), .C(_640__bF_buf0), .Y(_736_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf3), .B(_993_), .C(_1294__bF_buf2), .Y(_1451_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1453_), .C(_1443_), .Y(_1748__8_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__9_), .B(_1264__bF_buf1), .C(_1268__bF_buf6), .Y(_1454_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__9_), .B(_1264__bF_buf1), .C(_1272__bF_buf2), .Y(_1456_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__9_), .B(_1278__bF_buf4), .C(_1275__bF_buf4), .Y(_1458_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[9]), .B(_1278__bF_buf4), .C(_1268__bF_buf6), .Y(_1459_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__9_), .B(_1278__bF_buf4), .C(_1272__bF_buf5), .Y(_1460_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_1459_), .C(_1460_), .Y(_1461_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_1022_), .C(_1294__bF_buf6), .Y(_1467_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf0), .B(_1027_), .C(_1294__bF_buf6), .Y(_1469_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__2_), .B(_650__bF_buf1), .C(_644__bF_buf2), .Y(_737_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_1031_), .C(_1294__bF_buf5), .Y(_1470_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1472_), .C(_1462_), .Y(_1748__9_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__10_), .B(_1264__bF_buf3), .C(_1268__bF_buf4), .Y(_1473_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__10_), .B(_1264__bF_buf3), .C(_1272__bF_buf6), .Y(_1475_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__10_), .B(_1278__bF_buf2), .C(_1275__bF_buf4), .Y(_1477_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[10]), .B(_1278__bF_buf2), .C(_1268__bF_buf4), .Y(_1478_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__10_), .B(_1278__bF_buf2), .C(_1272__bF_buf5), .Y(_1479_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1477_), .B(_1478_), .C(_1479_), .Y(_1480_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf5), .B(_1060_), .C(_1294__bF_buf3), .Y(_1486_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_1065_), .C(_1294__bF_buf2), .Y(_1488_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_736_), .C(_737_), .Y(_738_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf3), .B(_1069_), .C(_1294__bF_buf2), .Y(_1489_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1485_), .B(_1491_), .C(_1481_), .Y(_1748__10_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__11_), .B(_1264__bF_buf1), .C(_1268__bF_buf0), .Y(_1492_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__11_), .B(_1264__bF_buf1), .C(_1272__bF_buf2), .Y(_1494_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__11_), .B(_1278__bF_buf4), .C(_1275__bF_buf3), .Y(_1496_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[11]), .B(_1278__bF_buf3), .C(_1268__bF_buf0), .Y(_1497_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__11_), .B(_1278__bF_buf5), .C(_1272__bF_buf1), .Y(_1498_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_1497_), .C(_1498_), .Y(_1499_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_1098_), .C(_1294__bF_buf5), .Y(_1505_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf0), .B(_1103_), .C(_1294__bF_buf5), .Y(_1507_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf0), .B(_756_), .C(_673__bF_buf6), .Y(_757_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_1107_), .C(_1294__bF_buf5), .Y(_1508_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1504_), .B(_1510_), .C(_1500_), .Y(_1748__11_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__12_), .B(_1264__bF_buf1), .C(_1268__bF_buf4), .Y(_1511_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__12_), .B(_1264__bF_buf3), .C(_1272__bF_buf6), .Y(_1513_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__12_), .B(_1278__bF_buf2), .C(_1275__bF_buf1), .Y(_1515_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[12]), .B(_1278__bF_buf2), .C(_1268__bF_buf0), .Y(_1516_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__12_), .B(_1278__bF_buf2), .C(_1272__bF_buf6), .Y(_1517_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .B(_1516_), .C(_1517_), .Y(_1518_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf5), .B(_1136_), .C(_1294__bF_buf1), .Y(_1524_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_1141_), .C(_1294__bF_buf1), .Y(_1526_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf1), .B(_761_), .C(_673__bF_buf6), .Y(_762_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf3), .B(_1145_), .C(_1294__bF_buf1), .Y(_1527_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1529_), .C(_1519_), .Y(_1748__12_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__13_), .B(_1264__bF_buf2), .C(_1268__bF_buf3), .Y(_1530_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__13_), .B(_1264__bF_buf2), .C(_1272__bF_buf1), .Y(_1532_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__13_), .B(_1278__bF_buf1), .C(_1275__bF_buf1), .Y(_1534_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[13]), .B(_1278__bF_buf1), .C(_1268__bF_buf3), .Y(_1535_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__13_), .B(_1278__bF_buf1), .C(_1272__bF_buf1), .Y(_1536_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1534_), .B(_1535_), .C(_1536_), .Y(_1537_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf5), .B(_1174_), .C(_1294__bF_buf3), .Y(_1543_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_1179_), .C(_1294__bF_buf2), .Y(_1545_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__0_), .B(_636__bF_buf2), .C(_644__bF_buf6), .Y(_645_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf2), .B(_765_), .C(_673__bF_buf6), .Y(_766_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf3), .B(_1183_), .C(_1294__bF_buf2), .Y(_1546_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1548_), .C(_1538_), .Y(_1748__13_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__14_), .B(_1264__bF_buf4), .C(_1268__bF_buf6), .Y(_1549_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__14_), .B(_1264__bF_buf4), .C(_1272__bF_buf2), .Y(_1551_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__14_), .B(_1278__bF_buf3), .C(_1275__bF_buf3), .Y(_1553_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[14]), .B(_1278__bF_buf0), .C(_1268__bF_buf1), .Y(_1554_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__14_), .B(_1278__bF_buf3), .C(_1272__bF_buf4), .Y(_1555_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1554_), .C(_1555_), .Y(_1556_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf2), .B(_1212_), .C(_1294__bF_buf6), .Y(_1562_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf0), .B(_1217_), .C(_1294__bF_buf6), .Y(_1564_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_768_), .C(_739_), .Y(_1749__2_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf0), .B(_1221_), .C(_1294__bF_buf4), .Y(_1565_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_1567_), .C(_1557_), .Y(_1748__14_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__15_), .B(_1264__bF_buf2), .C(_1268__bF_buf3), .Y(_1568_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__15_), .B(_1264__bF_buf2), .C(_1272__bF_buf1), .Y(_1570_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__15_), .B(_1278__bF_buf5), .C(_1275__bF_buf1), .Y(_1572_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[15]), .B(_1278__bF_buf5), .C(_1268__bF_buf0), .Y(_1573_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__15_), .B(_1278__bF_buf5), .C(_1272__bF_buf1), .Y(_1574_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_1573_), .C(_1574_), .Y(_1575_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1268__bF_buf5), .B(_1250_), .C(_1294__bF_buf1), .Y(_1581_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1275__bF_buf2), .B(_1255_), .C(_1294__bF_buf1), .Y(_1583_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__3_), .B(_636__bF_buf0), .C(_640__bF_buf5), .Y(_769_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1272__bF_buf3), .B(_1259_), .C(_1294__bF_buf1), .Y(_1584_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_1586_), .C(_1576_), .Y(_1748__15_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__3_), .B(_636__bF_buf0), .C(_644__bF_buf1), .Y(_771_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__3_), .B(_650__bF_buf5), .C(_647__bF_buf4), .Y(_773_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[3]), .B(_650__bF_buf5), .C(_640__bF_buf6), .Y(_774_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__3_), .B(_650__bF_buf5), .C(_644__bF_buf4), .Y(_775_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_774_), .C(_775_), .Y(_776_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf3), .B(_794_), .C(_673__bF_buf2), .Y(_795_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_799_), .C(_673__bF_buf2), .Y(_800_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__0_), .B(_650__bF_buf0), .C(_647__bF_buf3), .Y(_651_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf0), .B(_803_), .C(_673__bF_buf0), .Y(_804_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_806_), .C(_777_), .Y(_1749__3_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__4_), .B(_636__bF_buf1), .C(_640__bF_buf5), .Y(_807_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__4_), .B(_636__bF_buf1), .C(_644__bF_buf1), .Y(_809_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__4_), .B(_650__bF_buf5), .C(_647__bF_buf4), .Y(_811_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[4]), .B(_650__bF_buf4), .C(_640__bF_buf6), .Y(_812_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__4_), .B(_650__bF_buf4), .C(_644__bF_buf4), .Y(_813_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_812_), .C(_813_), .Y(_814_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf3), .B(_832_), .C(_673__bF_buf2), .Y(_833_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_837_), .C(_673__bF_buf0), .Y(_838_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[0]), .B(_650__bF_buf0), .C(_640__bF_buf2), .Y(_652_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf0), .B(_841_), .C(_673__bF_buf0), .Y(_842_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_826_), .B(_844_), .C(_815_), .Y(_1749__4_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__5_), .B(_636__bF_buf1), .C(_640__bF_buf5), .Y(_845_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__5_), .B(_636__bF_buf0), .C(_644__bF_buf1), .Y(_847_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__5_), .B(_650__bF_buf4), .C(_647__bF_buf4), .Y(_849_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[5]), .B(_650__bF_buf4), .C(_640__bF_buf6), .Y(_850_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__5_), .B(_650__bF_buf4), .C(_644__bF_buf4), .Y(_851_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_849_), .B(_850_), .C(_851_), .Y(_852_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf0), .B(_870_), .C(_673__bF_buf1), .Y(_871_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf1), .B(_875_), .C(_673__bF_buf6), .Y(_876_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__0_), .B(_650__bF_buf0), .C(_644__bF_buf3), .Y(_653_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf2), .B(_879_), .C(_673__bF_buf6), .Y(_880_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_882_), .C(_853_), .Y(_1749__5_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__6_), .B(_636__bF_buf4), .C(_640__bF_buf5), .Y(_883_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__6_), .B(_636__bF_buf4), .C(_644__bF_buf1), .Y(_885_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__6_), .B(_650__bF_buf1), .C(_647__bF_buf1), .Y(_887_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[6]), .B(_650__bF_buf1), .C(_640__bF_buf0), .Y(_888_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__6_), .B(_650__bF_buf1), .C(_644__bF_buf2), .Y(_889_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_887_), .B(_888_), .C(_889_), .Y(_890_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf3), .B(_908_), .C(_673__bF_buf2), .Y(_909_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_913_), .C(_673__bF_buf0), .Y(_914_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_652_), .C(_653_), .Y(_654_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf0), .B(_917_), .C(_673__bF_buf0), .Y(_918_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_920_), .C(_891_), .Y(_1749__6_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__7_), .B(_636__bF_buf1), .C(_640__bF_buf6), .Y(_921_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__7_), .B(_636__bF_buf0), .C(_644__bF_buf1), .Y(_923_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__7_), .B(_650__bF_buf5), .C(_647__bF_buf4), .Y(_925_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[7]), .B(_650__bF_buf5), .C(_640__bF_buf6), .Y(_926_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__7_), .B(_650__bF_buf5), .C(_644__bF_buf4), .Y(_927_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_926_), .C(_927_), .Y(_928_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf3), .B(_946_), .C(_673__bF_buf1), .Y(_947_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_951_), .C(_673__bF_buf6), .Y(_952_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_680_), .C(_673__bF_buf4), .Y(_681_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf2), .B(_955_), .C(_673__bF_buf6), .Y(_956_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_958_), .C(_929_), .Y(_1749__7_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__8_), .B(_636__bF_buf2), .C(_640__bF_buf4), .Y(_959_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__8_), .B(_636__bF_buf2), .C(_644__bF_buf6), .Y(_961_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__8_), .B(_650__bF_buf3), .C(_647__bF_buf3), .Y(_963_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[8]), .B(_650__bF_buf3), .C(_640__bF_buf4), .Y(_964_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__8_), .B(_650__bF_buf3), .C(_644__bF_buf3), .Y(_965_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_964_), .C(_965_), .Y(_966_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf1), .B(_984_), .C(_673__bF_buf5), .Y(_985_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf0), .B(_989_), .C(_673__bF_buf3), .Y(_990_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf1), .B(_685_), .C(_673__bF_buf4), .Y(_686_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_644__bF_buf5), .B(_993_), .C(_673__bF_buf3), .Y(_994_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_996_), .C(_967_), .Y(_1749__8_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__9_), .B(_636__bF_buf4), .C(_640__bF_buf5), .Y(_997_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__9_), .B(_636__bF_buf4), .C(_644__bF_buf1), .Y(_999_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__9_), .B(_650__bF_buf1), .C(_647__bF_buf1), .Y(_1001_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(REG_R1[9]), .B(_650__bF_buf1), .C(_640__bF_buf0), .Y(_1002_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__9_), .B(_650__bF_buf1), .C(_644__bF_buf2), .Y(_1003_) );
NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1002_), .C(_1003_), .Y(_1004_) );
NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_640__bF_buf3), .B(_1022_), .C(_673__bF_buf2), .Y(_1023_) );
NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_647__bF_buf2), .B(_1027_), .C(_673__bF_buf2), .Y(_1028_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[0]), .B(_1625_), .Y(_1626_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__0_), .B(_501__bF_buf0), .Y(_502_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_910_), .Y(_920_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_658_), .Y(_931_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_661_), .Y(_933_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_948_), .Y(_958_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_658_), .Y(_969_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_661_), .Y(_971_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_995_), .B(_986_), .Y(_996_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_658_), .Y(_1007_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_661_), .Y(_1009_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .B(_1024_), .Y(_1034_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__1_), .B(_501__bF_buf0), .Y(_503_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_658_), .Y(_1045_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_661_), .Y(_1047_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1062_), .Y(_1072_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1082_), .B(_658_), .Y(_1083_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_661_), .Y(_1085_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1109_), .B(_1100_), .Y(_1110_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1120_), .B(_658_), .Y(_1121_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_661_), .Y(_1123_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1138_), .Y(_1148_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .B(_658_), .Y(_1159_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__2_), .B(_501__bF_buf2), .Y(_504_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_661_), .Y(_1161_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1176_), .Y(_1186_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_658_), .Y(_1197_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_661_), .Y(_1199_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1214_), .Y(_1224_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_658_), .Y(_1235_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_661_), .Y(_1237_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1252_), .Y(_1262_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[3]), .B(_1263_), .Y(_1264_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[1]), .B(REG_RF1[0]), .Y(_1265_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__3_), .B(_501__bF_buf3), .Y(_505_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[1]), .B(_1267_), .Y(_1268_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[0]), .B(_1271_), .Y(_1272_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(REG_RF1[3]), .B(REG_RF1[2]), .Y(_1278_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1284_), .Y(_1290_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1288_), .Y(_1293_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1297_), .Y(_1301_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .B(_1311_), .Y(_1314_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1319_), .B(_1316_), .Y(_1320_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_1330_), .Y(_1333_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1335_), .Y(_1339_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__4_), .B(_501__bF_buf3), .Y(_506_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1351_), .B(_1349_), .Y(_1352_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1354_), .Y(_1358_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1368_), .Y(_1371_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .B(_1373_), .Y(_1377_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_1387_), .Y(_1390_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_1392_), .Y(_1396_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1406_), .Y(_1409_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1411_), .Y(_1415_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1427_), .B(_1425_), .Y(_1428_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1430_), .Y(_1434_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__5_), .B(_501__bF_buf4), .Y(_507_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1444_), .Y(_1447_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_1449_), .Y(_1453_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_1463_), .Y(_1466_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1468_), .Y(_1472_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_1482_), .Y(_1485_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1487_), .Y(_1491_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .B(_1501_), .Y(_1504_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .B(_1506_), .Y(_1510_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1520_), .Y(_1523_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1525_), .Y(_1529_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__6_), .B(_501__bF_buf2), .Y(_508_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1539_), .Y(_1542_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1544_), .Y(_1548_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .B(_1558_), .Y(_1561_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(_1563_), .Y(_1567_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1577_), .Y(_1580_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1582_), .Y(_1586_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__7_), .B(_501__bF_buf3), .Y(_509_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__8_), .B(_501__bF_buf1), .Y(_510_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__9_), .B(_501__bF_buf2), .Y(_511_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1625_), .Y(_1660_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__10_), .B(_501__bF_buf1), .Y(_512_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__11_), .B(_501__bF_buf4), .Y(_513_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__12_), .B(_501__bF_buf1), .Y(_514_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__13_), .B(_501__bF_buf0), .Y(_515_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__14_), .B(_501__bF_buf3), .Y(_516_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(REGS_2__15_), .B(_501__bF_buf4), .Y(_517_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__0_), .B(_518__bF_buf1), .Y(_519_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__1_), .B(_518__bF_buf1), .Y(_520_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__2_), .B(_518__bF_buf4), .Y(_521_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__3_), .B(_518__bF_buf2), .Y(_522_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[0]), .B(_1679_), .Y(_1680_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__4_), .B(_518__bF_buf3), .Y(_523_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__5_), .B(_518__bF_buf3), .Y(_524_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__6_), .B(_518__bF_buf4), .Y(_525_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__7_), .B(_518__bF_buf2), .Y(_526_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__8_), .B(_518__bF_buf0), .Y(_527_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__9_), .B(_518__bF_buf4), .Y(_528_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__10_), .B(_518__bF_buf4), .Y(_529_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__11_), .B(_518__bF_buf3), .Y(_530_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__12_), .B(_518__bF_buf0), .Y(_531_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__13_), .B(_518__bF_buf1), .Y(_532_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1679_), .Y(_1698_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__14_), .B(_518__bF_buf2), .Y(_533_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(REGS_3__15_), .B(_518__bF_buf3), .Y(_534_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__0_), .B(_568__bF_buf0), .Y(_569_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__1_), .B(_568__bF_buf3), .Y(_570_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__2_), .B(_568__bF_buf2), .Y(_571_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__3_), .B(_568__bF_buf4), .Y(_572_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__4_), .B(_568__bF_buf1), .Y(_573_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__5_), .B(_568__bF_buf4), .Y(_574_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__6_), .B(_568__bF_buf1), .Y(_575_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__7_), .B(_568__bF_buf4), .Y(_576_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[0]), .B(_1716_), .Y(_1717_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__8_), .B(_568__bF_buf0), .Y(_577_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__9_), .B(_568__bF_buf2), .Y(_578_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__10_), .B(_568__bF_buf0), .Y(_579_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__11_), .B(_568__bF_buf2), .Y(_580_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__12_), .B(_568__bF_buf2), .Y(_581_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__13_), .B(_568__bF_buf3), .Y(_582_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__14_), .B(_568__bF_buf4), .Y(_583_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(REGS_5__15_), .B(_568__bF_buf3), .Y(_584_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__0_), .B(_585__bF_buf2), .Y(_586_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__1_), .B(_585__bF_buf0), .Y(_587_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf0), .B(_358_), .Y(_359_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__2_), .B(_585__bF_buf1), .Y(_588_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__3_), .B(_585__bF_buf3), .Y(_589_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__4_), .B(_585__bF_buf3), .Y(_590_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__5_), .B(_585__bF_buf4), .Y(_591_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__6_), .B(_585__bF_buf4), .Y(_592_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__7_), .B(_585__bF_buf3), .Y(_593_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__8_), .B(_585__bF_buf1), .Y(_594_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__9_), .B(_585__bF_buf4), .Y(_595_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__10_), .B(_585__bF_buf1), .Y(_596_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__11_), .B(_585__bF_buf2), .Y(_597_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[0]), .B(_360_), .Y(_361_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__12_), .B(_585__bF_buf2), .Y(_598_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__13_), .B(_585__bF_buf0), .Y(_599_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__14_), .B(_585__bF_buf3), .Y(_600_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(REGS_6__15_), .B(_585__bF_buf0), .Y(_601_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[3]), .B(_635_), .Y(_636_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[1]), .B(REG_RF2[0]), .Y(_637_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[1]), .B(_639_), .Y(_640_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[0]), .B(_643_), .Y(_644_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(REG_RF2[3]), .B(REG_RF2[2]), .Y(_650_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_658_), .Y(_660_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_360_), .Y(_379_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_661_), .Y(_663_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_656_), .Y(_666_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_682_), .Y(_692_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_658_), .Y(_703_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_661_), .Y(_705_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_720_), .Y(_730_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_658_), .Y(_741_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_661_), .Y(_743_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_758_), .Y(_768_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_658_), .Y(_779_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[3]), .B(_499_), .Y(_500_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_661_), .Y(_781_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_796_), .Y(_806_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_658_), .Y(_817_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_661_), .Y(_819_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_834_), .Y(_844_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_658_), .Y(_855_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_661_), .Y(_857_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_872_), .Y(_882_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(_658_), .Y(_893_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_661_), .Y(_895_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_649_), .C(_654_), .Y(_655_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_819_), .C(_825_), .Y(_826_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_848_), .C(_852_), .Y(_853_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_857_), .C(_863_), .Y(_864_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_886_), .C(_890_), .Y(_891_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_895_), .C(_901_), .Y(_902_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_924_), .C(_928_), .Y(_929_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_933_), .C(_939_), .Y(_940_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(_962_), .C(_966_), .Y(_967_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_971_), .C(_977_), .Y(_978_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_1000_), .C(_1004_), .Y(_1005_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_663_), .C(_671_), .Y(_672_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .B(_1009_), .C(_1015_), .Y(_1016_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1036_), .B(_1038_), .C(_1042_), .Y(_1043_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1047_), .C(_1053_), .Y(_1054_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1076_), .C(_1080_), .Y(_1081_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1085_), .C(_1091_), .Y(_1092_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1114_), .C(_1118_), .Y(_1119_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1123_), .C(_1129_), .Y(_1130_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1152_), .C(_1156_), .Y(_1157_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1161_), .C(_1167_), .Y(_1168_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1190_), .C(_1194_), .Y(_1195_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_696_), .C(_700_), .Y(_701_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_1199_), .C(_1205_), .Y(_1206_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1228_), .C(_1232_), .Y(_1233_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1235_), .B(_1237_), .C(_1243_), .Y(_1244_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_1277_), .C(_1282_), .Y(_1283_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1305_), .C(_1309_), .Y(_1310_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(_1324_), .C(_1328_), .Y(_1329_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1343_), .C(_1347_), .Y(_1348_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1362_), .C(_1366_), .Y(_1367_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .B(_1381_), .C(_1385_), .Y(_1386_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1398_), .B(_1400_), .C(_1404_), .Y(_1405_) );
NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_705_), .C(_711_), .Y(_712_) );
NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1419_), .C(_1423_), .Y(_1424_) );
NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1438_), .C(_1442_), .Y(_1443_) );
NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1455_), .B(_1457_), .C(_1461_), .Y(_1462_) );
NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_1476_), .C(_1480_), .Y(_1481_) );
NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1495_), .C(_1499_), .Y(_1500_) );
NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1514_), .C(_1518_), .Y(_1519_) );
NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1533_), .C(_1537_), .Y(_1538_) );
NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_1552_), .C(_1556_), .Y(_1557_) );
NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1571_), .C(_1575_), .Y(_1576_) );
NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_734_), .C(_738_), .Y(_739_) );
NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_743_), .C(_749_), .Y(_750_) );
NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_772_), .C(_776_), .Y(_777_) );
NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_781_), .C(_787_), .Y(_788_) );
NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_810_), .C(_814_), .Y(_815_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf1), .B(_1627__bF_buf2), .C(_1628_), .Y(_0_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf1), .B(_1627__bF_buf4), .C(_1646_), .Y(_9_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1645__bF_buf1), .C(_1747_), .Y(_89_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_1622__bF_buf3), .C(FIRQ_REGS_7__10_), .Y(_352_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1647__bF_buf2), .C(_352_), .Y(_90_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_1622__bF_buf1), .C(FIRQ_REGS_7__11_), .Y(_353_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1649__bF_buf3), .C(_353_), .Y(_91_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_1622__bF_buf2), .C(FIRQ_REGS_7__12_), .Y(_354_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1651__bF_buf1), .C(_354_), .Y(_92_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_1622__bF_buf3), .C(FIRQ_REGS_7__13_), .Y(_355_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1653__bF_buf3), .C(_355_), .Y(_93_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_1622__bF_buf0), .C(FIRQ_REGS_7__14_), .Y(_356_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf1), .B(_1627__bF_buf0), .C(_1648_), .Y(_10_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1655__bF_buf2), .C(_356_), .Y(_94_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_1622__bF_buf3), .C(FIRQ_REGS_7__15_), .Y(_357_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1657__bF_buf1), .C(_357_), .Y(_95_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf1), .B(_362__bF_buf2), .C(_363_), .Y(_96_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf3), .B(_362__bF_buf4), .C(_364_), .Y(_97_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf2), .B(_362__bF_buf1), .C(_365_), .Y(_98_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf1), .B(_362__bF_buf3), .C(_366_), .Y(_99_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf1), .B(_362__bF_buf3), .C(_367_), .Y(_100_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf3), .B(_362__bF_buf2), .C(_368_), .Y(_101_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf3), .B(_362__bF_buf0), .C(_369_), .Y(_102_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf1), .B(_1627__bF_buf4), .C(_1650_), .Y(_11_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf3), .B(_362__bF_buf0), .C(_370_), .Y(_103_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf2), .B(_362__bF_buf1), .C(_371_), .Y(_104_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf2), .B(_362__bF_buf3), .C(_372_), .Y(_105_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf3), .B(_362__bF_buf1), .C(_373_), .Y(_106_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf2), .B(_362__bF_buf3), .C(_374_), .Y(_107_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf3), .B(_362__bF_buf2), .C(_375_), .Y(_108_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf1), .B(_362__bF_buf4), .C(_376_), .Y(_109_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf3), .B(_362__bF_buf0), .C(_377_), .Y(_110_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf2), .B(_362__bF_buf4), .C(_378_), .Y(_111_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf1), .B(_380__bF_buf2), .C(_381_), .Y(_112_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf2), .B(_1627__bF_buf1), .C(_1652_), .Y(_12_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf2), .B(_380__bF_buf3), .C(_382_), .Y(_113_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf1), .B(_380__bF_buf2), .C(_383_), .Y(_114_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf1), .B(_380__bF_buf4), .C(_384_), .Y(_115_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf1), .B(_380__bF_buf4), .C(_385_), .Y(_116_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf2), .B(_380__bF_buf1), .C(_386_), .Y(_117_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf2), .B(_380__bF_buf1), .C(_387_), .Y(_118_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf0), .B(_380__bF_buf0), .C(_388_), .Y(_119_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf1), .B(_380__bF_buf0), .C(_389_), .Y(_120_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf2), .B(_380__bF_buf4), .C(_390_), .Y(_121_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf1), .B(_380__bF_buf3), .C(_391_), .Y(_122_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf2), .B(_1627__bF_buf0), .C(_1654_), .Y(_13_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf2), .B(_380__bF_buf1), .C(_392_), .Y(_123_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf2), .B(_380__bF_buf3), .C(_393_), .Y(_124_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf1), .B(_380__bF_buf0), .C(_394_), .Y(_125_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf0), .B(_380__bF_buf1), .C(_395_), .Y(_126_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf2), .B(_380__bF_buf3), .C(_396_), .Y(_127_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf2), .B(_397__bF_buf4), .C(_398_), .Y(_128_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf1), .B(_397__bF_buf3), .C(_399_), .Y(_129_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf1), .B(_397__bF_buf3), .C(_400_), .Y(_130_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf1), .B(_397__bF_buf1), .C(_401_), .Y(_131_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf3), .B(_397__bF_buf2), .C(_402_), .Y(_132_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf2), .B(_1627__bF_buf4), .C(_1656_), .Y(_14_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf2), .B(_397__bF_buf2), .C(_403_), .Y(_133_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf0), .B(_397__bF_buf1), .C(_404_), .Y(_134_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf0), .B(_397__bF_buf4), .C(_405_), .Y(_135_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf1), .B(_397__bF_buf0), .C(_406_), .Y(_136_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf1), .B(_397__bF_buf3), .C(_407_), .Y(_137_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf1), .B(_397__bF_buf0), .C(_408_), .Y(_138_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf1), .B(_397__bF_buf1), .C(_409_), .Y(_139_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf2), .B(_397__bF_buf3), .C(_410_), .Y(_140_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf2), .B(_397__bF_buf0), .C(_411_), .Y(_141_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf0), .B(_397__bF_buf2), .C(_412_), .Y(_142_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf2), .B(_1627__bF_buf1), .C(_1658_), .Y(_15_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf2), .B(_397__bF_buf4), .C(_413_), .Y(_143_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf1), .B(_414__bF_buf3), .C(_415_), .Y(_144_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf2), .B(_414__bF_buf1), .C(_416_), .Y(_145_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf1), .B(_414__bF_buf3), .C(_417_), .Y(_146_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf1), .B(_414__bF_buf0), .C(_418_), .Y(_147_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf1), .B(_414__bF_buf4), .C(_419_), .Y(_148_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf2), .B(_414__bF_buf3), .C(_420_), .Y(_149_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf2), .B(_414__bF_buf0), .C(_421_), .Y(_150_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf2), .B(_414__bF_buf4), .C(_422_), .Y(_151_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf3), .B(_414__bF_buf2), .C(_423_), .Y(_152_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf1), .B(_1661__bF_buf1), .C(_1662_), .Y(_16_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf2), .B(_414__bF_buf0), .C(_424_), .Y(_153_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf2), .B(_414__bF_buf2), .C(_425_), .Y(_154_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf2), .B(_414__bF_buf4), .C(_426_), .Y(_155_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf1), .B(_414__bF_buf2), .C(_427_), .Y(_156_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf1), .B(_414__bF_buf1), .C(_428_), .Y(_157_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf0), .B(_414__bF_buf4), .C(_429_), .Y(_158_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf3), .B(_414__bF_buf1), .C(_430_), .Y(_159_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf2), .B(_431__bF_buf4), .C(_432_), .Y(_160_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf1), .B(_431__bF_buf1), .C(_433_), .Y(_161_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf3), .B(_431__bF_buf1), .C(_434_), .Y(_162_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf2), .B(_1661__bF_buf0), .C(_1663_), .Y(_17_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf2), .B(_431__bF_buf3), .C(_435_), .Y(_163_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf2), .B(_431__bF_buf0), .C(_436_), .Y(_164_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf1), .B(_431__bF_buf4), .C(_437_), .Y(_165_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf0), .B(_431__bF_buf3), .C(_438_), .Y(_166_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf1), .B(_431__bF_buf0), .C(_439_), .Y(_167_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf0), .B(_431__bF_buf2), .C(_440_), .Y(_168_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf3), .B(_431__bF_buf0), .C(_441_), .Y(_169_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf0), .B(_431__bF_buf2), .C(_442_), .Y(_170_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf1), .B(_431__bF_buf4), .C(_443_), .Y(_171_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf0), .B(_431__bF_buf4), .C(_444_), .Y(_172_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_1661__bF_buf3), .C(_1664_), .Y(_18_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf2), .B(_431__bF_buf2), .C(_445_), .Y(_173_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf1), .B(_431__bF_buf3), .C(_446_), .Y(_174_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf3), .B(_431__bF_buf1), .C(_447_), .Y(_175_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf2), .B(_448__bF_buf4), .C(_449_), .Y(_176_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf0), .B(_448__bF_buf3), .C(_450_), .Y(_177_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_448__bF_buf4), .C(_451_), .Y(_178_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf2), .B(_448__bF_buf2), .C(_452_), .Y(_179_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf1), .B(_448__bF_buf2), .C(_453_), .Y(_180_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf0), .B(_448__bF_buf0), .C(_454_), .Y(_181_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf1), .B(_448__bF_buf1), .C(_455_), .Y(_182_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf2), .B(_1627__bF_buf1), .C(_1630_), .Y(_1_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf2), .B(_1661__bF_buf4), .C(_1665_), .Y(_19_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf1), .B(_448__bF_buf2), .C(_456_), .Y(_183_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf0), .B(_448__bF_buf3), .C(_457_), .Y(_184_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf3), .B(_448__bF_buf1), .C(_458_), .Y(_185_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf0), .B(_448__bF_buf4), .C(_459_), .Y(_186_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf1), .B(_448__bF_buf0), .C(_460_), .Y(_187_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf0), .B(_448__bF_buf3), .C(_461_), .Y(_188_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf2), .B(_448__bF_buf4), .C(_462_), .Y(_189_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf1), .B(_448__bF_buf1), .C(_463_), .Y(_190_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf3), .B(_448__bF_buf3), .C(_464_), .Y(_191_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf3), .B(_465__bF_buf1), .C(_466_), .Y(_192_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf3), .B(_1661__bF_buf2), .C(_1666_), .Y(_20_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf1), .B(_465__bF_buf0), .C(_467_), .Y(_193_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf3), .B(_465__bF_buf2), .C(_468_), .Y(_194_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf0), .B(_465__bF_buf4), .C(_469_), .Y(_195_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf2), .B(_465__bF_buf3), .C(_470_), .Y(_196_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf1), .B(_465__bF_buf3), .C(_471_), .Y(_197_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf1), .B(_465__bF_buf4), .C(_472_), .Y(_198_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf1), .B(_465__bF_buf3), .C(_473_), .Y(_199_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf3), .B(_465__bF_buf0), .C(_474_), .Y(_200_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf1), .B(_465__bF_buf2), .C(_475_), .Y(_201_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf2), .B(_465__bF_buf1), .C(_476_), .Y(_202_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf2), .B(_1661__bF_buf2), .C(_1667_), .Y(_21_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf3), .B(_465__bF_buf4), .C(_477_), .Y(_203_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf0), .B(_465__bF_buf2), .C(_478_), .Y(_204_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf3), .B(_465__bF_buf1), .C(_479_), .Y(_205_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf1), .B(_465__bF_buf4), .C(_480_), .Y(_206_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf1), .B(_465__bF_buf0), .C(_481_), .Y(_207_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf3), .B(_482__bF_buf2), .C(_483_), .Y(_208_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf0), .B(_482__bF_buf4), .C(_484_), .Y(_209_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf3), .B(_482__bF_buf3), .C(_485_), .Y(_210_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf0), .B(_482__bF_buf0), .C(_486_), .Y(_211_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf3), .B(_482__bF_buf0), .C(_487_), .Y(_212_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf2), .B(_1661__bF_buf4), .C(_1668_), .Y(_22_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf1), .B(_482__bF_buf1), .C(_488_), .Y(_213_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf1), .B(_482__bF_buf1), .C(_489_), .Y(_214_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf2), .B(_482__bF_buf1), .C(_490_), .Y(_215_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf3), .B(_482__bF_buf4), .C(_491_), .Y(_216_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf1), .B(_482__bF_buf3), .C(_492_), .Y(_217_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf2), .B(_482__bF_buf2), .C(_493_), .Y(_218_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf3), .B(_482__bF_buf0), .C(_494_), .Y(_219_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf1), .B(_482__bF_buf4), .C(_495_), .Y(_220_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf3), .B(_482__bF_buf2), .C(_496_), .Y(_221_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf2), .B(_482__bF_buf3), .C(_497_), .Y(_222_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf2), .B(_1661__bF_buf2), .C(_1669_), .Y(_23_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf1), .B(_482__bF_buf4), .C(_498_), .Y(_223_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(REG_RFD[1]), .B(REG_RFD[2]), .C(REG_Write), .Y(_499_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536__bF_buf2), .C(_537_), .Y(_256_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_536__bF_buf4), .C(_539_), .Y(_257_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_536__bF_buf1), .C(_541_), .Y(_258_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_536__bF_buf0), .C(_543_), .Y(_259_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_536__bF_buf0), .C(_545_), .Y(_260_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_536__bF_buf2), .C(_547_), .Y(_261_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_536__bF_buf3), .C(_549_), .Y(_262_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_536__bF_buf0), .C(_551_), .Y(_263_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf1), .B(_1661__bF_buf1), .C(_1670_), .Y(_24_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_536__bF_buf1), .C(_553_), .Y(_264_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_536__bF_buf3), .C(_555_), .Y(_265_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_536__bF_buf4), .C(_557_), .Y(_266_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_536__bF_buf2), .C(_559_), .Y(_267_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_536__bF_buf2), .C(_561_), .Y(_268_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_536__bF_buf4), .C(_563_), .Y(_269_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_536__bF_buf3), .C(_565_), .Y(_270_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_536__bF_buf4), .C(_567_), .Y(_271_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_603__bF_buf4), .C(_604_), .Y(_304_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_603__bF_buf4), .C(_606_), .Y(_305_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf3), .B(_1661__bF_buf4), .C(_1671_), .Y(_25_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_603__bF_buf2), .C(_608_), .Y(_306_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_603__bF_buf0), .C(_610_), .Y(_307_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_603__bF_buf0), .C(_612_), .Y(_308_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_603__bF_buf1), .C(_614_), .Y(_309_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_603__bF_buf3), .C(_616_), .Y(_310_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_603__bF_buf3), .C(_618_), .Y(_311_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_603__bF_buf1), .C(_620_), .Y(_312_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_603__bF_buf1), .C(_622_), .Y(_313_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_603__bF_buf2), .C(_624_), .Y(_314_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_603__bF_buf0), .C(_626_), .Y(_315_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf1), .B(_1661__bF_buf0), .C(_1672_), .Y(_26_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_603__bF_buf1), .C(_628_), .Y(_316_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_603__bF_buf4), .C(_630_), .Y(_317_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_603__bF_buf3), .C(_632_), .Y(_318_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_603__bF_buf4), .C(_634_), .Y(_319_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_535_), .C(_641_), .Y(_642_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_602_), .C(_645_), .Y(_649_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(REG_Interrupt_flag_bF_buf0), .C(_668_), .Y(_669_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_665_), .C(_670_), .Y(_671_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(USR_REGS_0__0_), .C(_676_), .Y(_677_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(REG_Interrupt_flag_bF_buf3), .C(_679_), .Y(_680_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf2), .B(_1661__bF_buf3), .C(_1673_), .Y(_27_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_677_), .C(_681_), .Y(_682_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(REG_Interrupt_flag_bF_buf3), .C(_684_), .Y(_685_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(REG_Interrupt_flag_bF_buf3), .C(_688_), .Y(_689_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_538_), .C(_693_), .Y(_694_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_605_), .C(_695_), .Y(_696_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(REG_Interrupt_flag_bF_buf11), .C(_708_), .Y(_709_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_706_), .C(_710_), .Y(_711_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(USR_REGS_0__1_), .C(_714_), .Y(_715_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(REG_Interrupt_flag_bF_buf10), .C(_717_), .Y(_718_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_715_), .C(_719_), .Y(_720_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf2), .B(_1661__bF_buf3), .C(_1674_), .Y(_28_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(REG_Interrupt_flag_bF_buf10), .C(_722_), .Y(_723_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(REG_Interrupt_flag_bF_buf1), .C(_726_), .Y(_727_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_540_), .C(_731_), .Y(_732_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_607_), .C(_733_), .Y(_734_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(REG_Interrupt_flag_bF_buf0), .C(_746_), .Y(_747_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_744_), .C(_748_), .Y(_749_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(USR_REGS_0__2_), .C(_752_), .Y(_753_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(REG_Interrupt_flag_bF_buf4), .C(_755_), .Y(_756_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_753_), .C(_757_), .Y(_758_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(REG_Interrupt_flag_bF_buf4), .C(_760_), .Y(_761_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf1), .B(_1627__bF_buf2), .C(_1632_), .Y(_2_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf1), .B(_1661__bF_buf0), .C(_1675_), .Y(_29_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(REG_Interrupt_flag_bF_buf4), .C(_764_), .Y(_765_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_542_), .C(_769_), .Y(_770_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_609_), .C(_771_), .Y(_772_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(REG_Interrupt_flag_bF_buf8), .C(_784_), .Y(_785_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_782_), .C(_786_), .Y(_787_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__3_), .C(_790_), .Y(_791_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(REG_Interrupt_flag_bF_buf13), .C(_793_), .Y(_794_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_791_), .C(_795_), .Y(_796_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(REG_Interrupt_flag_bF_buf13), .C(_798_), .Y(_799_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(REG_Interrupt_flag_bF_buf6), .C(_802_), .Y(_803_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf0), .B(_1661__bF_buf4), .C(_1676_), .Y(_30_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_544_), .C(_807_), .Y(_808_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_611_), .C(_809_), .Y(_810_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(REG_Interrupt_flag_bF_buf9), .C(_822_), .Y(_823_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_820_), .C(_824_), .Y(_825_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__4_), .C(_828_), .Y(_829_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(REG_Interrupt_flag_bF_buf13), .C(_831_), .Y(_832_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_829_), .C(_833_), .Y(_834_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(REG_Interrupt_flag_bF_buf2), .C(_836_), .Y(_837_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(REG_Interrupt_flag_bF_buf2), .C(_840_), .Y(_841_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_546_), .C(_845_), .Y(_846_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf3), .B(_1661__bF_buf1), .C(_1677_), .Y(_31_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_613_), .C(_847_), .Y(_848_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(REG_Interrupt_flag_bF_buf9), .C(_860_), .Y(_861_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_858_), .C(_862_), .Y(_863_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__5_), .C(_866_), .Y(_867_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(REG_Interrupt_flag_bF_buf4), .C(_869_), .Y(_870_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_867_), .C(_871_), .Y(_872_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(REG_Interrupt_flag_bF_buf4), .C(_874_), .Y(_875_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(REG_Interrupt_flag_bF_buf4), .C(_878_), .Y(_879_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_548_), .C(_883_), .Y(_884_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_615_), .C(_885_), .Y(_886_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf2), .B(_1681__bF_buf4), .C(_1682_), .Y(_32_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_897_), .B(REG_Interrupt_flag_bF_buf8), .C(_898_), .Y(_899_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_896_), .C(_900_), .Y(_901_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__6_), .C(_904_), .Y(_905_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_906_), .B(REG_Interrupt_flag_bF_buf2), .C(_907_), .Y(_908_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_905_), .C(_909_), .Y(_910_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(REG_Interrupt_flag_bF_buf2), .C(_912_), .Y(_913_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_915_), .B(REG_Interrupt_flag_bF_buf6), .C(_916_), .Y(_917_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_550_), .C(_921_), .Y(_922_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_617_), .C(_923_), .Y(_924_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(REG_Interrupt_flag_bF_buf9), .C(_936_), .Y(_937_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf1), .B(_1681__bF_buf1), .C(_1683_), .Y(_33_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_934_), .C(_938_), .Y(_939_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf13), .B(USR_REGS_0__7_), .C(_942_), .Y(_943_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(REG_Interrupt_flag_bF_buf7), .C(_945_), .Y(_946_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_943_), .C(_947_), .Y(_948_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(REG_Interrupt_flag_bF_buf2), .C(_950_), .Y(_951_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_953_), .B(REG_Interrupt_flag_bF_buf4), .C(_954_), .Y(_955_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_552_), .C(_959_), .Y(_960_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_619_), .C(_961_), .Y(_962_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(REG_Interrupt_flag_bF_buf11), .C(_974_), .Y(_975_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_972_), .C(_976_), .Y(_977_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_1681__bF_buf4), .C(_1684_), .Y(_34_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(USR_REGS_0__8_), .C(_980_), .Y(_981_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(REG_Interrupt_flag_bF_buf3), .C(_983_), .Y(_984_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_981_), .C(_985_), .Y(_986_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(REG_Interrupt_flag_bF_buf5), .C(_988_), .Y(_989_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(REG_Interrupt_flag_bF_buf10), .C(_992_), .Y(_993_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_554_), .C(_997_), .Y(_998_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_621_), .C(_999_), .Y(_1000_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(REG_Interrupt_flag_bF_buf0), .C(_1012_), .Y(_1013_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1010_), .C(_1014_), .Y(_1015_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__9_), .C(_1018_), .Y(_1019_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf2), .B(_1681__bF_buf0), .C(_1685_), .Y(_35_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1020_), .B(REG_Interrupt_flag_bF_buf12), .C(_1021_), .Y(_1022_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1019_), .C(_1023_), .Y(_1024_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(REG_Interrupt_flag_bF_buf6), .C(_1026_), .Y(_1027_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(REG_Interrupt_flag_bF_buf6), .C(_1030_), .Y(_1031_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_556_), .C(_1035_), .Y(_1036_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_623_), .C(_1037_), .Y(_1038_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(REG_Interrupt_flag_bF_buf11), .C(_1050_), .Y(_1051_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1048_), .C(_1052_), .Y(_1053_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(USR_REGS_0__10_), .C(_1056_), .Y(_1057_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(REG_Interrupt_flag_bF_buf7), .C(_1059_), .Y(_1060_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf2), .B(_1681__bF_buf3), .C(_1686_), .Y(_36_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1057_), .C(_1061_), .Y(_1062_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(REG_Interrupt_flag_bF_buf1), .C(_1064_), .Y(_1065_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .B(REG_Interrupt_flag_bF_buf10), .C(_1068_), .Y(_1069_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_558_), .C(_1073_), .Y(_1074_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_625_), .C(_1075_), .Y(_1076_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1087_), .B(REG_Interrupt_flag_bF_buf9), .C(_1088_), .Y(_1089_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1086_), .C(_1090_), .Y(_1091_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__11_), .C(_1094_), .Y(_1095_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(REG_Interrupt_flag_bF_buf2), .C(_1097_), .Y(_1098_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1095_), .C(_1099_), .Y(_1100_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf0), .B(_1681__bF_buf3), .C(_1687_), .Y(_37_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .B(REG_Interrupt_flag_bF_buf4), .C(_1102_), .Y(_1103_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(REG_Interrupt_flag_bF_buf6), .C(_1106_), .Y(_1107_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_560_), .C(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_627_), .C(_1113_), .Y(_1114_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .B(REG_Interrupt_flag_bF_buf0), .C(_1126_), .Y(_1127_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1124_), .C(_1128_), .Y(_1129_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf3), .B(USR_REGS_0__12_), .C(_1132_), .Y(_1133_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1134_), .B(REG_Interrupt_flag_bF_buf3), .C(_1135_), .Y(_1136_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1133_), .C(_1137_), .Y(_1138_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(REG_Interrupt_flag_bF_buf1), .C(_1140_), .Y(_1141_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf0), .B(_1681__bF_buf0), .C(_1688_), .Y(_38_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(REG_Interrupt_flag_bF_buf1), .C(_1144_), .Y(_1145_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_562_), .C(_1149_), .Y(_1150_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_629_), .C(_1151_), .Y(_1152_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(REG_Interrupt_flag_bF_buf11), .C(_1164_), .Y(_1165_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1162_), .C(_1166_), .Y(_1167_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(USR_REGS_0__13_), .C(_1170_), .Y(_1171_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1172_), .B(REG_Interrupt_flag_bF_buf7), .C(_1173_), .Y(_1174_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1171_), .C(_1175_), .Y(_1176_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(REG_Interrupt_flag_bF_buf10), .C(_1178_), .Y(_1179_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(REG_Interrupt_flag_bF_buf5), .C(_1182_), .Y(_1183_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf1), .B(_1627__bF_buf3), .C(_1634_), .Y(_3_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf1), .B(_1681__bF_buf3), .C(_1689_), .Y(_39_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_564_), .C(_1187_), .Y(_1188_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_631_), .C(_1189_), .Y(_1190_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(REG_Interrupt_flag_bF_buf9), .C(_1202_), .Y(_1203_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1200_), .C(_1204_), .Y(_1205_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf12), .B(USR_REGS_0__14_), .C(_1208_), .Y(_1209_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1210_), .B(REG_Interrupt_flag_bF_buf6), .C(_1211_), .Y(_1212_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1209_), .C(_1213_), .Y(_1214_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(REG_Interrupt_flag_bF_buf2), .C(_1216_), .Y(_1217_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1219_), .B(REG_Interrupt_flag_bF_buf2), .C(_1220_), .Y(_1221_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_566_), .C(_1225_), .Y(_1226_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf0), .B(_1681__bF_buf1), .C(_1690_), .Y(_40_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_633_), .C(_1227_), .Y(_1228_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(REG_Interrupt_flag_bF_buf11), .C(_1240_), .Y(_1241_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_1238_), .C(_1242_), .Y(_1243_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(REG_Interrupt_flag_bF_buf7), .B(USR_REGS_0__15_), .C(_1246_), .Y(_1247_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(REG_Interrupt_flag_bF_buf10), .C(_1249_), .Y(_1250_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_1247_), .C(_1251_), .Y(_1252_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1253_), .B(REG_Interrupt_flag_bF_buf10), .C(_1254_), .Y(_1255_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1257_), .B(REG_Interrupt_flag_bF_buf10), .C(_1258_), .Y(_1259_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_535_), .C(_1269_), .Y(_1270_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_602_), .C(_1273_), .Y(_1277_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf2), .B(_1681__bF_buf3), .C(_1691_), .Y(_41_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_665_), .C(_1291_), .Y(_1292_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_677_), .C(_1296_), .Y(_1297_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_538_), .C(_1302_), .Y(_1303_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_605_), .C(_1304_), .Y(_1305_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_706_), .C(_1312_), .Y(_1313_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_715_), .C(_1315_), .Y(_1316_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_540_), .C(_1321_), .Y(_1322_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_607_), .C(_1323_), .Y(_1324_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_744_), .C(_1331_), .Y(_1332_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_753_), .C(_1334_), .Y(_1335_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf0), .B(_1681__bF_buf2), .C(_1692_), .Y(_42_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_542_), .C(_1340_), .Y(_1341_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_609_), .C(_1342_), .Y(_1343_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_782_), .C(_1350_), .Y(_1351_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_791_), .C(_1353_), .Y(_1354_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_544_), .C(_1359_), .Y(_1360_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_611_), .C(_1361_), .Y(_1362_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_820_), .C(_1369_), .Y(_1370_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_829_), .C(_1372_), .Y(_1373_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_546_), .C(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_613_), .C(_1380_), .Y(_1381_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf1), .B(_1681__bF_buf4), .C(_1693_), .Y(_43_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_858_), .C(_1388_), .Y(_1389_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_867_), .C(_1391_), .Y(_1392_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_548_), .C(_1397_), .Y(_1398_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_615_), .C(_1399_), .Y(_1400_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_896_), .C(_1407_), .Y(_1408_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_905_), .C(_1410_), .Y(_1411_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_550_), .C(_1416_), .Y(_1417_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_617_), .C(_1418_), .Y(_1419_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_934_), .C(_1426_), .Y(_1427_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_943_), .C(_1429_), .Y(_1430_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf0), .B(_1681__bF_buf2), .C(_1694_), .Y(_44_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_552_), .C(_1435_), .Y(_1436_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_619_), .C(_1437_), .Y(_1438_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_972_), .C(_1445_), .Y(_1446_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_981_), .C(_1448_), .Y(_1449_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_554_), .C(_1454_), .Y(_1455_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_621_), .C(_1456_), .Y(_1457_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1010_), .C(_1464_), .Y(_1465_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1019_), .C(_1467_), .Y(_1468_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_556_), .C(_1473_), .Y(_1474_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_623_), .C(_1475_), .Y(_1476_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf2), .B(_1681__bF_buf1), .C(_1695_), .Y(_45_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1048_), .C(_1483_), .Y(_1484_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1057_), .C(_1486_), .Y(_1487_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_558_), .C(_1492_), .Y(_1493_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_625_), .C(_1494_), .Y(_1495_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1086_), .C(_1502_), .Y(_1503_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1095_), .C(_1505_), .Y(_1506_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_560_), .C(_1511_), .Y(_1512_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_627_), .C(_1513_), .Y(_1514_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1124_), .C(_1521_), .Y(_1522_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1133_), .C(_1524_), .Y(_1525_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf1), .B(_1681__bF_buf0), .C(_1696_), .Y(_46_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_562_), .C(_1530_), .Y(_1531_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_629_), .C(_1532_), .Y(_1533_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1162_), .C(_1540_), .Y(_1541_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1171_), .C(_1543_), .Y(_1544_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_564_), .C(_1549_), .Y(_1550_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_631_), .C(_1551_), .Y(_1552_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1200_), .C(_1559_), .Y(_1560_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1209_), .C(_1562_), .Y(_1563_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_566_), .C(_1568_), .Y(_1569_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_633_), .C(_1570_), .Y(_1571_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf3), .B(_1681__bF_buf2), .C(_1697_), .Y(_47_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1238_), .C(_1578_), .Y(_1579_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1295_), .B(_1247_), .C(_1581_), .Y(_1582_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf2), .B(_1587__bF_buf0), .C(_1588_), .Y(_320_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf2), .B(_1587__bF_buf2), .C(_1589_), .Y(_321_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf1), .B(_1587__bF_buf4), .C(_1590_), .Y(_322_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf3), .B(_1587__bF_buf3), .C(_1591_), .Y(_323_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf1), .B(_1587__bF_buf3), .C(_1592_), .Y(_324_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf2), .B(_1587__bF_buf4), .C(_1593_), .Y(_325_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf2), .B(_1587__bF_buf4), .C(_1594_), .Y(_326_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf0), .B(_1587__bF_buf1), .C(_1595_), .Y(_327_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf3), .B(_1699__bF_buf0), .C(_1700_), .Y(_48_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf1), .B(_1587__bF_buf1), .C(_1596_), .Y(_328_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf2), .B(_1587__bF_buf3), .C(_1597_), .Y(_329_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf1), .B(_1587__bF_buf2), .C(_1598_), .Y(_330_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf2), .B(_1587__bF_buf4), .C(_1599_), .Y(_331_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf2), .B(_1587__bF_buf0), .C(_1600_), .Y(_332_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf1), .B(_1587__bF_buf1), .C(_1601_), .Y(_333_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf2), .B(_1587__bF_buf0), .C(_1602_), .Y(_334_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf2), .B(_1587__bF_buf2), .C(_1603_), .Y(_335_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_1604__bF_buf4), .C(_1605_), .Y(_336_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_1604__bF_buf3), .C(_1606_), .Y(_337_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf3), .B(_1627__bF_buf4), .C(_1636_), .Y(_4_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf0), .B(_1699__bF_buf0), .C(_1701_), .Y(_49_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_1604__bF_buf4), .C(_1607_), .Y(_338_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_1604__bF_buf1), .C(_1608_), .Y(_339_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_827_), .B(_1604__bF_buf1), .C(_1609_), .Y(_340_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_1604__bF_buf0), .C(_1610_), .Y(_341_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_1604__bF_buf0), .C(_1611_), .Y(_342_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1604__bF_buf1), .C(_1612_), .Y(_343_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_979_), .B(_1604__bF_buf4), .C(_1613_), .Y(_344_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .B(_1604__bF_buf2), .C(_1614_), .Y(_345_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1604__bF_buf4), .C(_1615_), .Y(_346_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1604__bF_buf2), .C(_1616_), .Y(_347_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf0), .B(_1699__bF_buf2), .C(_1702_), .Y(_50_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_1604__bF_buf0), .C(_1617_), .Y(_348_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1604__bF_buf3), .C(_1618_), .Y(_349_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1604__bF_buf2), .C(_1619_), .Y(_350_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .B(_1604__bF_buf3), .C(_1620_), .Y(_351_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf2), .B(_1699__bF_buf3), .C(_1703_), .Y(_51_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf2), .B(_1699__bF_buf3), .C(_1704_), .Y(_52_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf0), .B(_1699__bF_buf3), .C(_1705_), .Y(_53_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf1), .B(_1699__bF_buf4), .C(_1706_), .Y(_54_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf1), .B(_1699__bF_buf3), .C(_1707_), .Y(_55_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf0), .B(_1699__bF_buf0), .C(_1708_), .Y(_56_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf3), .B(_1699__bF_buf4), .C(_1709_), .Y(_57_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf0), .B(_1699__bF_buf2), .C(_1710_), .Y(_58_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf0), .B(_1627__bF_buf3), .C(_1638_), .Y(_5_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf3), .B(_1699__bF_buf1), .C(_1711_), .Y(_59_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf1), .B(_1699__bF_buf1), .C(_1712_), .Y(_60_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf3), .B(_1699__bF_buf2), .C(_1713_), .Y(_61_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf1), .B(_1699__bF_buf4), .C(_1714_), .Y(_62_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf1), .B(_1699__bF_buf1), .C(_1715_), .Y(_63_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_1621__bF_buf3), .B(_1718__bF_buf3), .C(_1719_), .Y(_64_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1629__bF_buf0), .B(_1718__bF_buf2), .C(_1720_), .Y(_65_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1631__bF_buf3), .B(_1718__bF_buf1), .C(_1721_), .Y(_66_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1633__bF_buf0), .B(_1718__bF_buf0), .C(_1722_), .Y(_67_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1635__bF_buf2), .B(_1718__bF_buf4), .C(_1723_), .Y(_68_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf2), .B(_1627__bF_buf3), .C(_1640_), .Y(_6_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_1637__bF_buf1), .B(_1718__bF_buf4), .C(_1724_), .Y(_69_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1639__bF_buf1), .B(_1718__bF_buf0), .C(_1725_), .Y(_70_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf2), .B(_1718__bF_buf0), .C(_1726_), .Y(_71_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf3), .B(_1718__bF_buf2), .C(_1727_), .Y(_72_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_1645__bF_buf3), .B(_1718__bF_buf1), .C(_1728_), .Y(_73_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1647__bF_buf2), .B(_1718__bF_buf3), .C(_1729_), .Y(_74_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1649__bF_buf3), .B(_1718__bF_buf4), .C(_1730_), .Y(_75_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1651__bF_buf1), .B(_1718__bF_buf3), .C(_1731_), .Y(_76_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_1653__bF_buf3), .B(_1718__bF_buf3), .C(_1732_), .Y(_77_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1655__bF_buf2), .B(_1718__bF_buf4), .C(_1733_), .Y(_78_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_1641__bF_buf0), .B(_1627__bF_buf2), .C(_1642_), .Y(_7_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1657__bF_buf1), .B(_1718__bF_buf2), .C(_1734_), .Y(_79_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_1622__bF_buf2), .C(FIRQ_REGS_7__0_), .Y(_1738_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1621__bF_buf3), .C(_1738_), .Y(_80_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_1622__bF_buf3), .C(FIRQ_REGS_7__1_), .Y(_1739_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1629__bF_buf1), .C(_1739_), .Y(_81_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_1622__bF_buf2), .C(FIRQ_REGS_7__2_), .Y(_1740_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1631__bF_buf3), .C(_1740_), .Y(_82_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_1622__bF_buf1), .C(FIRQ_REGS_7__3_), .Y(_1741_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1633__bF_buf0), .C(_1741_), .Y(_83_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_1622__bF_buf0), .C(FIRQ_REGS_7__4_), .Y(_1742_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_1643__bF_buf1), .B(_1627__bF_buf0), .C(_1644_), .Y(_8_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1635__bF_buf3), .C(_1742_), .Y(_84_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_1622__bF_buf1), .C(FIRQ_REGS_7__5_), .Y(_1743_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1637__bF_buf1), .C(_1743_), .Y(_85_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf2), .B(_1622__bF_buf0), .C(FIRQ_REGS_7__6_), .Y(_1744_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1639__bF_buf0), .C(_1744_), .Y(_86_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf1), .B(_1622__bF_buf1), .C(FIRQ_REGS_7__7_), .Y(_1745_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1641__bF_buf2), .C(_1745_), .Y(_87_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf3), .B(_1622__bF_buf3), .C(FIRQ_REGS_7__8_), .Y(_1746_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1643__bF_buf3), .C(_1746_), .Y(_88_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1735__bF_buf0), .B(_1622__bF_buf2), .C(FIRQ_REGS_7__9_), .Y(_1747_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_1287_), .C(_1286_), .D(_659_), .Y(_1288_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_1287_), .C(_1286_), .D(_1006_), .Y(_1463_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1287_), .C(_1286_), .D(_1044_), .Y(_1482_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1287_), .C(_1286_), .D(_1082_), .Y(_1501_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1287_), .C(_1286_), .D(_1120_), .Y(_1520_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1287_), .C(_1286_), .D(_1158_), .Y(_1539_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1287_), .C(_1286_), .D(_1196_), .Y(_1558_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1287_), .C(_1286_), .D(_1234_), .Y(_1577_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_1287_), .C(_1286_), .D(_702_), .Y(_1311_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_742_), .B(_1287_), .C(_1286_), .D(_740_), .Y(_1330_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_1287_), .C(_1286_), .D(_778_), .Y(_1349_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_1287_), .C(_1286_), .D(_816_), .Y(_1368_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_1287_), .C(_1286_), .D(_854_), .Y(_1387_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_1287_), .C(_1286_), .D(_892_), .Y(_1406_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_1287_), .C(_1286_), .D(_930_), .Y(_1425_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_1287_), .C(_1286_), .D(_968_), .Y(_1444_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_1716_), .B(_1659_), .Y(_1735_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_1748__0_), .Y(REG_A[0]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_1748__1_), .Y(REG_A[1]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_1748__2_), .Y(REG_A[2]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_1748__3_), .Y(REG_A[3]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_1748__4_), .Y(REG_A[4]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_1748__5_), .Y(REG_A[5]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_1748__6_), .Y(REG_A[6]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_1748__7_), .Y(REG_A[7]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_1748__8_), .Y(REG_A[8]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_1748__9_), .Y(REG_A[9]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_1748__10_), .Y(REG_A[10]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_1748__11_), .Y(REG_A[11]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_1748__12_), .Y(REG_A[12]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_1748__13_), .Y(REG_A[13]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_1748__14_), .Y(REG_A[14]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_1748__15_), .Y(REG_A[15]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_1749__0_), .Y(REG_B[0]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_1749__1_), .Y(REG_B[1]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_1749__2_), .Y(REG_B[2]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_1749__3_), .Y(REG_B[3]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_1749__4_), .Y(REG_B[4]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_1749__5_), .Y(REG_B[5]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_1749__6_), .Y(REG_B[6]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_1749__7_), .Y(REG_B[7]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_1749__8_), .Y(REG_B[8]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_1749__9_), .Y(REG_B[9]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_1749__10_), .Y(REG_B[10]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_1749__11_), .Y(REG_B[11]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_1749__12_), .Y(REG_B[12]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_1749__13_), .Y(REG_B[13]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_1749__14_), .Y(REG_B[14]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_1749__15_), .Y(REG_B[15]) );
endmodule
