magic
tech scmos
magscale 1 4
timestamp 1515334672
<< metal1 >>
rect 1976 2157 2003 2163
rect 2013 2157 2024 2163
rect 2120 2157 2163 2163
rect 2568 2156 2572 2164
rect 141 2137 152 2143
rect 237 2137 248 2143
rect 333 2137 344 2143
rect 637 2137 675 2143
rect 72 2117 83 2123
rect 552 2117 563 2123
rect 637 2123 643 2137
rect 808 2137 819 2143
rect 909 2137 947 2143
rect 1016 2137 1027 2143
rect 1112 2137 1139 2143
rect 1213 2137 1251 2143
rect 1400 2137 1411 2143
rect 1565 2137 1592 2143
rect 621 2117 643 2123
rect 952 2117 963 2123
rect 1277 2117 1331 2123
rect 1500 2117 1528 2123
rect 1500 2116 1508 2117
rect 1816 2117 1827 2123
rect 2029 2117 2040 2123
rect 2493 2117 2531 2123
rect 1181 2097 1192 2103
rect 2093 2097 2104 2103
rect 2317 2097 2328 2103
rect 2445 2097 2456 2103
rect 2797 2097 2808 2103
rect 2776 2077 2835 2083
rect 2877 2077 2904 2083
rect 1005 1937 1048 1943
rect 509 1917 547 1923
rect 61 1897 72 1903
rect 61 1883 67 1897
rect 141 1897 152 1903
rect 584 1897 595 1903
rect 717 1903 723 1923
rect 717 1897 755 1903
rect 45 1877 67 1883
rect 141 1877 152 1883
rect 301 1877 328 1883
rect 445 1877 467 1883
rect 989 1883 995 1923
rect 1032 1917 1048 1923
rect 1581 1897 1592 1903
rect 1757 1903 1763 1923
rect 1789 1917 1811 1923
rect 1757 1897 1795 1903
rect 2013 1903 2019 1923
rect 2840 1916 2844 1924
rect 2904 1916 2908 1924
rect 2968 1916 2972 1924
rect 1981 1897 2019 1903
rect 2333 1897 2344 1903
rect 2792 1897 2835 1903
rect 2888 1897 2899 1903
rect 2936 1897 2963 1903
rect 3101 1897 3139 1903
rect 968 1877 995 1883
rect 1064 1877 1075 1883
rect 1149 1877 1176 1883
rect 1192 1877 1203 1883
rect 1272 1877 1288 1883
rect 1528 1877 1555 1883
rect 1608 1877 1619 1883
rect 2536 1877 2579 1883
rect 2808 1877 2819 1883
rect 829 1857 851 1863
rect 948 1856 952 1864
rect 2413 1837 2424 1843
rect 3117 1757 3139 1763
rect 45 1737 56 1743
rect 733 1737 744 1743
rect 1048 1737 1080 1743
rect 1197 1737 1208 1743
rect 253 1717 264 1723
rect 376 1717 387 1723
rect 749 1717 787 1723
rect 749 1697 755 1717
rect 872 1717 883 1723
rect 920 1717 947 1723
rect 1197 1717 1203 1737
rect 2248 1737 2259 1743
rect 2461 1737 2472 1743
rect 2552 1737 2563 1743
rect 2941 1737 2952 1743
rect 1277 1717 1304 1723
rect 1421 1717 1432 1723
rect 1517 1717 1540 1723
rect 1532 1712 1540 1717
rect 1896 1717 1907 1723
rect 2077 1717 2120 1723
rect 2168 1717 2196 1723
rect 2188 1716 2196 1717
rect 2264 1717 2275 1723
rect 3021 1717 3059 1723
rect 1533 1697 1544 1703
rect 1656 1697 1667 1703
rect 1976 1696 1980 1704
rect 2696 1697 2707 1703
rect 3021 1697 3027 1717
rect 3144 1717 3155 1723
rect 3165 1717 3176 1723
rect 1613 1677 1688 1683
rect 2712 1677 2739 1683
rect 2104 1637 2131 1643
rect 3165 1557 3192 1563
rect 232 1497 243 1503
rect 312 1497 323 1503
rect 493 1497 504 1503
rect 493 1483 499 1497
rect 856 1497 883 1503
rect 1128 1497 1139 1503
rect 1213 1503 1219 1523
rect 1192 1497 1219 1503
rect 1309 1497 1320 1503
rect 1660 1503 1668 1508
rect 1629 1497 1668 1503
rect 1816 1497 1827 1503
rect 477 1477 499 1483
rect 616 1477 627 1483
rect 797 1477 851 1483
rect 845 1457 851 1477
rect 1208 1477 1235 1483
rect 1245 1477 1256 1483
rect 1821 1477 1827 1497
rect 2077 1497 2147 1503
rect 2248 1497 2275 1503
rect 2589 1497 2600 1503
rect 2701 1497 2739 1503
rect 2749 1497 2760 1503
rect 2941 1497 2952 1503
rect 2040 1477 2051 1483
rect 2621 1477 2648 1483
rect 2765 1477 2776 1483
rect 1405 1457 1427 1463
rect 2077 1457 2088 1463
rect 605 1337 616 1343
rect 24 1317 35 1323
rect 184 1317 211 1323
rect 344 1317 355 1323
rect 376 1317 387 1323
rect 589 1317 627 1323
rect 760 1317 771 1323
rect 925 1317 952 1323
rect 1325 1323 1331 1343
rect 2104 1337 2147 1343
rect 2381 1337 2392 1343
rect 2445 1337 2456 1343
rect 2664 1337 2675 1343
rect 2941 1337 2952 1343
rect 3080 1337 3091 1343
rect 1277 1317 1315 1323
rect 1325 1317 1352 1323
rect 1896 1317 1907 1323
rect 2093 1317 2104 1323
rect 2573 1317 2611 1323
rect 317 1297 339 1303
rect 1709 1297 1720 1303
rect 1912 1296 1916 1304
rect 2605 1297 2611 1317
rect 2808 1317 2819 1323
rect 2093 1237 2120 1243
rect 244 1116 248 1124
rect 152 1097 163 1103
rect 621 1097 659 1103
rect 1357 1097 1368 1103
rect 2013 1103 2019 1123
rect 2664 1116 2668 1124
rect 3101 1117 3112 1123
rect 1773 1097 1811 1103
rect 1965 1097 2003 1103
rect 2013 1097 2051 1103
rect 2189 1097 2232 1103
rect 2312 1097 2339 1103
rect 2621 1097 2632 1103
rect 125 1077 136 1083
rect 189 1077 200 1083
rect 573 1077 584 1083
rect 637 1077 648 1083
rect 637 1057 643 1077
rect 861 1077 872 1083
rect 989 1077 1032 1083
rect 1117 1077 1128 1083
rect 1245 1077 1256 1083
rect 1165 1057 1176 1063
rect 1245 1057 1251 1077
rect 1373 1077 1411 1083
rect 1533 1077 1544 1083
rect 1741 1077 1752 1083
rect 2536 1077 2547 1083
rect 2861 1077 2872 1083
rect 2957 1077 3011 1083
rect 3112 1077 3139 1083
rect 2269 1057 2307 1063
rect 2344 1057 2355 1063
rect 3181 1057 3192 1063
rect 504 957 515 963
rect 1341 957 1368 963
rect 1432 957 1443 963
rect 301 937 312 943
rect 573 937 584 943
rect 1165 937 1176 943
rect 1533 943 1539 963
rect 1592 957 1603 963
rect 1464 937 1507 943
rect 1533 937 1571 943
rect 2301 937 2339 943
rect 2360 937 2387 943
rect 2632 937 2643 943
rect 3016 937 3027 943
rect 3080 937 3091 943
rect 3181 937 3192 943
rect 104 917 115 923
rect 248 917 275 923
rect 333 917 387 923
rect 813 917 824 923
rect 1277 917 1304 923
rect 685 897 696 903
rect 1277 897 1283 917
rect 1645 917 1683 923
rect 1949 917 1987 923
rect 1864 896 1868 904
rect 1949 897 1955 917
rect 2264 917 2275 923
rect 3084 923 3092 928
rect 3069 917 3092 923
rect 2141 897 2152 903
rect 3181 757 3192 763
rect 125 717 163 723
rect 173 717 195 723
rect 328 697 371 703
rect 520 697 547 703
rect 1165 697 1203 703
rect 232 677 243 683
rect 872 677 883 683
rect 1197 677 1203 697
rect 1368 697 1379 703
rect 1389 697 1416 703
rect 1453 703 1459 723
rect 1837 717 1859 723
rect 1453 697 1491 703
rect 1773 697 1811 703
rect 2104 697 2131 703
rect 1512 677 1523 683
rect 2157 677 2168 683
rect 269 657 291 663
rect 989 657 1011 663
rect 1965 657 1992 663
rect 2157 657 2163 677
rect 2701 677 2712 683
rect 2792 677 2803 683
rect 3032 657 3043 663
rect 1597 637 1608 643
rect 1752 577 1774 583
rect 1976 577 2014 583
rect 1416 556 1420 564
rect 2916 556 2920 564
rect 77 537 99 543
rect 77 523 83 537
rect 461 537 472 543
rect 45 517 83 523
rect 157 517 184 523
rect 445 517 456 523
rect 973 523 979 543
rect 1549 537 1576 543
rect 1709 537 1768 543
rect 1805 537 1848 543
rect 2045 537 2147 543
rect 2552 537 2563 543
rect 936 517 979 523
rect 989 517 1016 523
rect 1048 517 1059 523
rect 1117 517 1155 523
rect 2461 517 2472 523
rect 2845 523 2851 543
rect 2888 537 2899 543
rect 2936 537 2963 543
rect 3181 537 3192 543
rect 2792 517 2851 523
rect 2861 517 2888 523
rect 285 497 296 503
rect 408 497 419 503
rect 1453 497 1464 503
rect 205 477 232 483
rect 1356 483 1364 488
rect 1320 477 1364 483
rect 141 303 147 323
rect 1933 317 1944 323
rect 2248 316 2252 324
rect 2360 316 2364 324
rect 2445 317 2456 323
rect 141 297 179 303
rect 317 297 339 303
rect 333 277 339 297
rect 845 297 883 303
rect 1645 297 1672 303
rect 1709 297 1763 303
rect 1848 297 1859 303
rect 2024 297 2035 303
rect 2541 297 2579 303
rect 397 277 435 283
rect 584 277 595 283
rect 2504 277 2515 283
rect 2600 277 2611 283
rect 2701 277 2712 283
rect 2968 277 2995 283
rect 840 256 844 264
rect 2088 257 2124 263
rect 2484 256 2488 264
rect 2786 236 2792 244
rect 1629 157 1640 163
rect 1816 157 1827 163
rect 2397 157 2408 163
rect 557 137 579 143
rect 1021 137 1064 143
rect 1245 137 1256 143
rect 1597 137 1608 143
rect 2285 137 2296 143
rect 2957 137 2984 143
rect 3181 137 3192 143
rect 1165 117 1203 123
rect 813 97 835 103
rect 904 97 915 103
rect 1197 97 1203 117
rect 1437 117 1448 123
rect 2040 117 2051 123
rect 2317 117 2339 123
rect 1220 96 1224 104
rect 1476 96 1480 104
rect 2580 96 2584 104
rect 2077 37 2104 43
<< m2contact >>
rect 2077 2202 2113 2218
rect 3080 2172 3096 2188
rect 40 2152 56 2168
rect 696 2152 712 2168
rect 776 2152 792 2168
rect 920 2152 936 2168
rect 1048 2152 1064 2168
rect 1176 2152 1192 2168
rect 1640 2152 1656 2168
rect 1912 2152 1928 2168
rect 2024 2152 2040 2168
rect 2104 2152 2120 2168
rect 2552 2152 2568 2168
rect 3032 2152 3048 2168
rect 3064 2154 3080 2170
rect 1352 2148 1368 2150
rect 152 2132 168 2148
rect 248 2132 264 2148
rect 344 2132 360 2148
rect 8 2112 24 2128
rect 56 2112 72 2128
rect 88 2112 104 2128
rect 136 2112 152 2128
rect 168 2112 200 2128
rect 232 2112 296 2128
rect 328 2112 344 2128
rect 360 2112 392 2128
rect 424 2112 440 2128
rect 472 2112 488 2128
rect 520 2112 552 2128
rect 568 2112 584 2128
rect 792 2132 808 2148
rect 1000 2132 1016 2148
rect 1096 2132 1112 2148
rect 1192 2132 1208 2148
rect 1304 2132 1320 2148
rect 1352 2134 1400 2148
rect 1368 2132 1400 2134
rect 1512 2132 1528 2148
rect 1592 2132 1608 2148
rect 2040 2132 2056 2148
rect 2168 2132 2184 2148
rect 2264 2132 2280 2148
rect 2296 2132 2312 2148
rect 2328 2132 2344 2148
rect 2392 2132 2408 2148
rect 2504 2132 2552 2148
rect 2584 2132 2600 2148
rect 2856 2132 2872 2148
rect 3096 2132 3112 2148
rect 664 2112 680 2128
rect 712 2112 760 2128
rect 808 2112 824 2128
rect 856 2112 904 2128
rect 936 2112 952 2128
rect 1016 2112 1032 2128
rect 1064 2112 1096 2128
rect 1144 2112 1160 2128
rect 1256 2112 1272 2128
rect 1352 2112 1368 2128
rect 1432 2112 1448 2128
rect 1528 2112 1544 2128
rect 1608 2112 1624 2128
rect 1656 2112 1688 2128
rect 1704 2112 1720 2128
rect 1800 2112 1816 2128
rect 1880 2112 1896 2128
rect 1944 2112 1960 2128
rect 2040 2112 2072 2128
rect 2184 2112 2200 2128
rect 2280 2112 2296 2128
rect 2344 2112 2360 2128
rect 2408 2112 2424 2128
rect 2616 2112 2632 2128
rect 2680 2112 2696 2128
rect 2760 2112 2776 2128
rect 2824 2112 2840 2128
rect 2904 2112 2920 2128
rect 2968 2112 2984 2128
rect 3048 2112 3064 2128
rect 3112 2112 3128 2128
rect 760 2092 776 2108
rect 984 2092 1000 2108
rect 1192 2092 1208 2108
rect 1224 2092 1240 2108
rect 1288 2092 1304 2108
rect 1688 2092 1704 2108
rect 1896 2092 1912 2108
rect 1928 2092 1944 2108
rect 2104 2092 2120 2108
rect 2328 2092 2344 2108
rect 2456 2092 2472 2108
rect 2552 2092 2568 2108
rect 2600 2092 2616 2108
rect 2664 2092 2680 2108
rect 2776 2092 2792 2108
rect 2808 2092 2824 2108
rect 2888 2092 2904 2108
rect 2952 2092 2968 2108
rect 600 2072 616 2088
rect 1720 2072 1736 2088
rect 1848 2072 1864 2088
rect 1960 2072 1976 2088
rect 2632 2072 2648 2088
rect 2696 2072 2712 2088
rect 2744 2072 2776 2088
rect 2904 2072 2936 2088
rect 2984 2072 3000 2088
rect 3016 2072 3032 2088
rect 408 2032 424 2048
rect 504 2032 520 2048
rect 952 2032 968 2048
rect 1560 2032 1576 2048
rect 1704 2032 1720 2048
rect 1768 2032 1784 2048
rect 2056 2032 2072 2048
rect 2232 2032 2248 2048
rect 2376 2032 2392 2048
rect 2408 2032 2424 2048
rect 2488 2032 2504 2048
rect 2616 2032 2632 2048
rect 2680 2032 2696 2048
rect 2728 2032 2744 2048
rect 2808 2032 2824 2048
rect 2904 2032 2920 2048
rect 2968 2032 2984 2048
rect 3144 2032 3160 2048
rect 1037 2002 1073 2018
rect 1224 1972 1240 1988
rect 1976 1972 1992 1988
rect 2328 1972 2344 1988
rect 2776 1972 2792 1988
rect 1048 1932 1064 1948
rect 1272 1932 1288 1948
rect 552 1912 568 1928
rect 692 1912 708 1928
rect 8 1892 24 1908
rect 72 1892 104 1908
rect 152 1892 200 1908
rect 232 1892 248 1908
rect 264 1892 280 1908
rect 344 1892 360 1908
rect 392 1892 424 1908
rect 472 1892 488 1908
rect 568 1892 584 1908
rect 632 1892 664 1908
rect 680 1892 696 1908
rect 728 1912 744 1928
rect 776 1892 792 1908
rect 840 1892 856 1908
rect 904 1892 920 1908
rect 968 1892 984 1908
rect 152 1872 168 1888
rect 328 1872 344 1888
rect 504 1872 536 1888
rect 664 1872 680 1888
rect 760 1872 776 1888
rect 792 1872 808 1888
rect 872 1872 888 1888
rect 920 1872 936 1888
rect 952 1872 968 1888
rect 1016 1912 1032 1928
rect 1048 1912 1064 1928
rect 1112 1912 1128 1928
rect 1304 1912 1320 1928
rect 1368 1912 1384 1928
rect 1080 1892 1096 1908
rect 1160 1892 1192 1908
rect 1240 1892 1256 1908
rect 1288 1892 1304 1908
rect 1320 1892 1336 1908
rect 1384 1892 1400 1908
rect 1416 1892 1432 1908
rect 1448 1892 1480 1908
rect 1592 1892 1608 1908
rect 1624 1892 1656 1908
rect 1720 1892 1736 1908
rect 1832 1892 1848 1908
rect 1864 1892 1880 1908
rect 1960 1892 1976 1908
rect 2136 1912 2152 1928
rect 2296 1912 2312 1928
rect 2744 1912 2760 1928
rect 2824 1912 2840 1928
rect 2856 1912 2872 1928
rect 2888 1912 2904 1928
rect 2920 1912 2936 1928
rect 2952 1912 2968 1928
rect 2984 1912 3016 1928
rect 3064 1912 3080 1928
rect 2040 1892 2056 1908
rect 2216 1892 2232 1908
rect 2344 1892 2360 1908
rect 2376 1892 2392 1908
rect 2488 1892 2504 1908
rect 2600 1892 2616 1908
rect 2632 1892 2648 1908
rect 2696 1892 2712 1908
rect 2776 1892 2792 1908
rect 2856 1892 2888 1908
rect 2920 1892 2936 1908
rect 3032 1892 3048 1908
rect 3080 1892 3096 1908
rect 3160 1892 3176 1908
rect 2248 1888 2264 1892
rect 1016 1872 1032 1888
rect 1048 1872 1064 1888
rect 1176 1872 1192 1888
rect 1224 1872 1240 1888
rect 1288 1872 1304 1888
rect 1336 1872 1352 1888
rect 1400 1872 1416 1888
rect 1432 1872 1448 1888
rect 1480 1872 1496 1888
rect 1512 1872 1528 1888
rect 1592 1872 1608 1888
rect 1656 1872 1672 1888
rect 1704 1872 1720 1888
rect 1768 1872 1784 1888
rect 1816 1872 1832 1888
rect 1848 1872 1864 1888
rect 1992 1872 2024 1888
rect 2056 1872 2072 1888
rect 2200 1872 2216 1888
rect 2232 1876 2264 1888
rect 2232 1872 2248 1876
rect 2344 1872 2376 1888
rect 2504 1872 2536 1888
rect 2616 1872 2632 1888
rect 2680 1872 2696 1888
rect 2792 1872 2808 1888
rect 2872 1872 2888 1888
rect 2936 1872 2952 1888
rect 3000 1872 3016 1888
rect 3048 1872 3064 1888
rect 3112 1872 3128 1888
rect 3176 1872 3192 1888
rect 424 1852 440 1868
rect 888 1852 904 1868
rect 952 1852 968 1868
rect 1128 1852 1144 1868
rect 1368 1852 1384 1868
rect 1512 1852 1528 1868
rect 1592 1852 1608 1868
rect 1688 1852 1704 1868
rect 1928 1852 1960 1868
rect 2104 1852 2136 1868
rect 2152 1852 2184 1868
rect 2504 1852 2520 1868
rect 216 1832 232 1848
rect 376 1832 392 1848
rect 616 1832 632 1848
rect 808 1832 824 1848
rect 1112 1832 1128 1848
rect 1496 1832 1512 1848
rect 1672 1832 1688 1848
rect 1752 1832 1768 1848
rect 1784 1832 1800 1848
rect 1896 1832 1912 1848
rect 1976 1832 1992 1848
rect 2184 1832 2200 1848
rect 2280 1832 2296 1848
rect 2424 1832 2440 1848
rect 2504 1832 2520 1848
rect 2664 1832 2680 1848
rect 2728 1832 2744 1848
rect 3128 1832 3144 1848
rect 2077 1802 2113 1818
rect 216 1772 232 1788
rect 568 1772 584 1788
rect 664 1772 680 1788
rect 1096 1772 1112 1788
rect 1224 1772 1240 1788
rect 1736 1772 1752 1788
rect 1848 1772 1864 1788
rect 2312 1772 2328 1788
rect 2792 1772 2808 1788
rect 2872 1772 2888 1788
rect 312 1752 328 1768
rect 1240 1752 1256 1768
rect 1720 1752 1736 1768
rect 1832 1752 1848 1768
rect 2040 1752 2056 1768
rect 2152 1752 2168 1768
rect 2328 1752 2344 1768
rect 2408 1752 2424 1768
rect 2680 1752 2696 1768
rect 2824 1752 2840 1768
rect 3096 1752 3112 1768
rect 56 1732 104 1748
rect 472 1732 488 1748
rect 712 1732 728 1748
rect 744 1732 776 1748
rect 792 1732 808 1748
rect 856 1732 872 1748
rect 904 1732 936 1748
rect 984 1732 1000 1748
rect 1032 1732 1048 1748
rect 1080 1732 1096 1748
rect 1112 1732 1128 1748
rect 1144 1732 1160 1748
rect 1176 1732 1192 1748
rect 8 1712 24 1728
rect 88 1712 104 1728
rect 136 1712 168 1728
rect 184 1712 200 1728
rect 232 1712 248 1728
rect 264 1712 296 1728
rect 328 1712 376 1728
rect 424 1712 456 1728
rect 504 1712 520 1728
rect 536 1712 552 1728
rect 584 1712 616 1728
rect 632 1712 648 1728
rect 680 1712 712 1728
rect 808 1712 824 1728
rect 856 1712 872 1728
rect 904 1712 920 1728
rect 1016 1712 1032 1728
rect 1128 1712 1144 1728
rect 1208 1732 1224 1748
rect 1256 1732 1272 1748
rect 1352 1732 1384 1748
rect 1880 1732 1896 1748
rect 1944 1732 1960 1748
rect 2024 1732 2040 1748
rect 2168 1732 2184 1748
rect 2232 1732 2248 1748
rect 2344 1732 2360 1748
rect 2472 1732 2488 1748
rect 2536 1732 2552 1748
rect 2600 1732 2616 1748
rect 2760 1732 2776 1748
rect 2952 1732 2984 1748
rect 3080 1732 3096 1748
rect 1208 1712 1224 1728
rect 1304 1712 1320 1728
rect 1336 1712 1352 1728
rect 1384 1712 1400 1728
rect 1432 1712 1464 1728
rect 1496 1712 1512 1728
rect 1544 1712 1560 1728
rect 1624 1712 1640 1728
rect 1672 1712 1688 1728
rect 1752 1712 1768 1728
rect 1800 1712 1816 1728
rect 1864 1712 1896 1728
rect 1960 1712 1976 1728
rect 2120 1712 2136 1728
rect 2152 1712 2168 1728
rect 2248 1712 2264 1728
rect 2360 1712 2376 1728
rect 2440 1712 2456 1728
rect 2488 1712 2504 1728
rect 2584 1712 2600 1728
rect 2616 1712 2632 1728
rect 2728 1712 2744 1728
rect 2840 1712 2856 1728
rect 2904 1712 2920 1728
rect 2984 1712 3000 1728
rect 840 1692 856 1708
rect 904 1692 920 1708
rect 968 1692 1000 1708
rect 1080 1692 1096 1708
rect 1144 1692 1160 1708
rect 1288 1692 1320 1708
rect 1544 1692 1560 1708
rect 1640 1692 1656 1708
rect 1816 1692 1832 1708
rect 1928 1692 1944 1708
rect 1960 1692 1976 1708
rect 1992 1692 2008 1708
rect 2296 1692 2312 1708
rect 2392 1692 2424 1708
rect 2520 1692 2536 1708
rect 2680 1692 2696 1708
rect 2792 1692 2808 1708
rect 3064 1712 3080 1728
rect 3128 1712 3144 1728
rect 3176 1712 3192 1728
rect 3032 1692 3048 1708
rect 408 1672 424 1688
rect 1560 1672 1576 1688
rect 1688 1672 1704 1688
rect 1784 1672 1800 1688
rect 2488 1672 2504 1688
rect 2648 1672 2664 1688
rect 2696 1672 2712 1688
rect 808 1652 824 1668
rect 776 1632 792 1648
rect 936 1632 952 1648
rect 1336 1632 1352 1648
rect 1480 1632 1496 1648
rect 1576 1632 1592 1648
rect 1624 1632 1640 1648
rect 1704 1632 1720 1648
rect 1768 1632 1784 1648
rect 1896 1632 1912 1648
rect 2008 1632 2024 1648
rect 2056 1632 2072 1648
rect 2088 1632 2104 1648
rect 2264 1632 2280 1648
rect 2360 1632 2376 1648
rect 2664 1632 2680 1648
rect 2744 1632 2760 1648
rect 2808 1632 2824 1648
rect 2984 1632 3000 1648
rect 1037 1602 1073 1618
rect 360 1572 376 1588
rect 552 1572 568 1588
rect 696 1572 712 1588
rect 3192 1552 3208 1568
rect 168 1532 184 1548
rect 1496 1532 1512 1548
rect 1688 1532 1704 1548
rect 2792 1532 2808 1548
rect 2984 1532 3000 1548
rect 1112 1512 1128 1528
rect 8 1492 24 1508
rect 72 1492 104 1508
rect 136 1492 152 1508
rect 216 1492 232 1508
rect 280 1492 312 1508
rect 328 1492 344 1508
rect 376 1492 392 1508
rect 440 1492 456 1508
rect 200 1472 216 1488
rect 232 1472 248 1488
rect 504 1492 536 1508
rect 568 1492 584 1508
rect 600 1492 616 1508
rect 664 1492 696 1508
rect 728 1492 744 1508
rect 760 1492 776 1508
rect 840 1492 856 1508
rect 952 1492 968 1508
rect 984 1492 1000 1508
rect 1016 1492 1032 1508
rect 1080 1492 1096 1508
rect 1112 1492 1128 1508
rect 1160 1492 1192 1508
rect 1464 1512 1480 1528
rect 1640 1512 1656 1528
rect 1720 1512 1736 1528
rect 1768 1512 1784 1528
rect 2168 1512 2200 1528
rect 2204 1512 2220 1528
rect 2248 1512 2264 1528
rect 2632 1512 2648 1528
rect 2712 1512 2728 1528
rect 2872 1512 2888 1528
rect 2952 1512 2968 1528
rect 1256 1492 1272 1508
rect 1320 1492 1336 1508
rect 1368 1492 1384 1508
rect 1448 1492 1464 1508
rect 1496 1492 1512 1508
rect 1528 1492 1544 1508
rect 1608 1492 1624 1508
rect 1672 1492 1688 1508
rect 1800 1492 1816 1508
rect 600 1472 616 1488
rect 424 1452 440 1468
rect 648 1452 664 1468
rect 856 1472 872 1488
rect 968 1472 984 1488
rect 1000 1472 1016 1488
rect 1064 1472 1080 1488
rect 1096 1472 1112 1488
rect 1192 1472 1208 1488
rect 1256 1472 1288 1488
rect 1512 1472 1528 1488
rect 1592 1472 1608 1488
rect 1752 1472 1768 1488
rect 1800 1472 1816 1488
rect 1944 1492 1992 1508
rect 2024 1492 2040 1508
rect 2216 1492 2248 1508
rect 2280 1492 2296 1508
rect 2376 1492 2392 1508
rect 2600 1492 2616 1508
rect 2760 1492 2776 1508
rect 2808 1492 2824 1508
rect 2840 1492 2856 1508
rect 2904 1492 2920 1508
rect 2952 1492 2968 1508
rect 2984 1492 3000 1508
rect 3128 1492 3144 1508
rect 2328 1488 2344 1492
rect 1912 1472 1928 1488
rect 2024 1472 2040 1488
rect 2120 1472 2136 1488
rect 2232 1472 2248 1488
rect 2296 1476 2344 1488
rect 2296 1472 2328 1476
rect 2424 1472 2440 1488
rect 2520 1472 2536 1488
rect 2600 1472 2616 1488
rect 2648 1472 2664 1488
rect 2680 1472 2696 1488
rect 2776 1472 2792 1488
rect 2824 1472 2840 1488
rect 2856 1472 2872 1488
rect 2888 1472 2904 1488
rect 3000 1472 3032 1488
rect 3112 1472 3128 1488
rect 856 1452 872 1468
rect 1144 1452 1160 1468
rect 1192 1452 1208 1468
rect 1304 1452 1320 1468
rect 1384 1452 1400 1468
rect 1432 1452 1448 1468
rect 1928 1452 1944 1468
rect 2008 1452 2024 1468
rect 2088 1452 2104 1468
rect 2408 1452 2424 1468
rect 2648 1452 2664 1468
rect 2776 1452 2792 1468
rect 40 1432 56 1448
rect 120 1432 136 1448
rect 168 1432 184 1448
rect 408 1432 424 1448
rect 632 1432 648 1448
rect 888 1432 904 1448
rect 1336 1432 1352 1448
rect 1560 1432 1576 1448
rect 1688 1432 1704 1448
rect 1736 1432 1752 1448
rect 1784 1432 1800 1448
rect 1864 1432 1880 1448
rect 1992 1432 2008 1448
rect 2168 1432 2184 1448
rect 2360 1432 2376 1448
rect 2392 1432 2408 1448
rect 2456 1432 2472 1448
rect 2552 1432 2568 1448
rect 2664 1432 2680 1448
rect 3080 1432 3096 1448
rect 2077 1402 2113 1418
rect 1192 1372 1208 1388
rect 1304 1372 1320 1388
rect 1736 1372 1752 1388
rect 2024 1372 2040 1388
rect 2776 1372 2792 1388
rect 120 1352 136 1368
rect 296 1352 312 1368
rect 728 1352 744 1368
rect 1176 1352 1192 1368
rect 1240 1352 1256 1368
rect 1720 1352 1736 1368
rect 1816 1352 1832 1368
rect 2040 1352 2072 1368
rect 2728 1352 2744 1368
rect 2760 1352 2776 1368
rect 184 1332 200 1348
rect 360 1332 376 1348
rect 616 1332 648 1348
rect 664 1332 680 1348
rect 1208 1332 1224 1348
rect 8 1312 24 1328
rect 72 1312 104 1328
rect 168 1312 184 1328
rect 216 1312 232 1328
rect 264 1312 280 1328
rect 328 1312 344 1328
rect 360 1312 376 1328
rect 392 1312 408 1328
rect 440 1312 456 1328
rect 488 1312 504 1328
rect 536 1312 568 1328
rect 680 1312 712 1328
rect 744 1312 760 1328
rect 776 1312 792 1328
rect 824 1312 840 1328
rect 856 1312 888 1328
rect 952 1312 984 1328
rect 1016 1312 1048 1328
rect 1096 1312 1112 1328
rect 1144 1312 1176 1328
rect 1224 1312 1240 1328
rect 1656 1332 1672 1348
rect 1704 1332 1720 1348
rect 1832 1332 1848 1348
rect 1880 1332 1896 1348
rect 1944 1332 1960 1348
rect 2088 1332 2104 1348
rect 2184 1332 2216 1348
rect 2248 1332 2264 1348
rect 2392 1332 2424 1348
rect 2456 1332 2472 1348
rect 2488 1332 2504 1348
rect 2536 1332 2552 1348
rect 2600 1332 2616 1348
rect 2648 1332 2664 1348
rect 2824 1332 2840 1348
rect 2872 1332 2888 1348
rect 2952 1332 2984 1348
rect 3064 1332 3080 1348
rect 1352 1312 1368 1328
rect 1400 1312 1432 1328
rect 1464 1312 1480 1328
rect 1512 1312 1528 1328
rect 1560 1312 1592 1328
rect 1608 1312 1624 1328
rect 1672 1312 1688 1328
rect 1784 1312 1800 1328
rect 1880 1312 1896 1328
rect 1960 1312 1976 1328
rect 1992 1312 2024 1328
rect 2104 1312 2120 1328
rect 2168 1312 2184 1328
rect 2232 1312 2248 1328
rect 2280 1312 2296 1328
rect 2344 1312 2376 1328
rect 2392 1312 2408 1328
rect 2456 1312 2472 1328
rect 2520 1312 2536 1328
rect 2552 1312 2568 1328
rect 136 1292 152 1308
rect 568 1292 584 1308
rect 1288 1292 1304 1308
rect 1480 1292 1496 1308
rect 1592 1292 1608 1308
rect 1720 1292 1736 1308
rect 1800 1292 1816 1308
rect 1896 1292 1912 1308
rect 1928 1292 1944 1308
rect 2136 1292 2152 1308
rect 2200 1292 2216 1308
rect 2264 1292 2280 1308
rect 2328 1292 2344 1308
rect 2584 1292 2600 1308
rect 2632 1312 2648 1328
rect 2680 1312 2696 1328
rect 2792 1312 2808 1328
rect 2840 1312 2856 1328
rect 2904 1312 2920 1328
rect 56 1272 72 1288
rect 1448 1272 1464 1288
rect 1624 1272 1640 1288
rect 1768 1272 1784 1288
rect 2296 1272 2312 1288
rect 1528 1252 1544 1268
rect 2408 1252 2424 1268
rect 104 1232 120 1248
rect 168 1232 184 1248
rect 248 1232 264 1248
rect 408 1232 424 1248
rect 504 1232 520 1248
rect 664 1232 680 1248
rect 792 1232 808 1248
rect 888 1232 904 1248
rect 984 1232 1000 1248
rect 1112 1232 1128 1248
rect 1272 1232 1288 1248
rect 1384 1232 1400 1248
rect 1464 1232 1480 1248
rect 1608 1232 1624 1248
rect 1784 1232 1800 1248
rect 1864 1232 1880 1248
rect 2120 1232 2136 1248
rect 2312 1232 2328 1248
rect 2712 1232 2728 1248
rect 2744 1232 2760 1248
rect 2936 1232 2952 1248
rect 3032 1232 3048 1248
rect 3144 1232 3160 1248
rect 1037 1202 1073 1218
rect 24 1172 40 1188
rect 2136 1172 2152 1188
rect 2424 1172 2440 1188
rect 3160 1172 3176 1188
rect 56 1132 72 1148
rect 440 1132 456 1148
rect 2120 1132 2136 1148
rect 216 1112 232 1128
rect 248 1112 264 1128
rect 328 1112 344 1128
rect 1320 1112 1336 1128
rect 1528 1112 1544 1128
rect 1704 1112 1720 1128
rect 1784 1112 1800 1128
rect 1864 1112 1880 1128
rect 88 1092 104 1108
rect 136 1092 152 1108
rect 248 1092 264 1108
rect 296 1092 328 1108
rect 344 1092 360 1108
rect 408 1092 424 1108
rect 536 1092 552 1108
rect 600 1092 616 1108
rect 696 1092 728 1108
rect 760 1092 776 1108
rect 808 1092 824 1108
rect 840 1092 856 1108
rect 904 1092 952 1108
rect 984 1092 1000 1108
rect 1048 1092 1080 1108
rect 1112 1092 1128 1108
rect 1176 1092 1208 1108
rect 1256 1092 1272 1108
rect 1304 1092 1320 1108
rect 1368 1092 1384 1108
rect 1400 1092 1416 1108
rect 1448 1092 1480 1108
rect 1496 1092 1512 1108
rect 1560 1092 1576 1108
rect 1608 1092 1656 1108
rect 2024 1112 2040 1128
rect 2152 1112 2168 1128
rect 2264 1112 2280 1128
rect 2504 1112 2520 1128
rect 2648 1112 2664 1128
rect 2680 1112 2696 1128
rect 2856 1112 2872 1128
rect 3112 1112 3128 1128
rect 2136 1092 2152 1108
rect 2232 1092 2248 1108
rect 2296 1092 2312 1108
rect 2408 1092 2424 1108
rect 2472 1092 2488 1108
rect 2568 1092 2584 1108
rect 2632 1092 2664 1108
rect 2712 1092 2728 1108
rect 2760 1092 2776 1108
rect 2824 1092 2840 1108
rect 2920 1092 2952 1108
rect 2984 1092 3000 1108
rect 3048 1092 3064 1108
rect 72 1072 88 1088
rect 136 1072 152 1088
rect 200 1072 216 1088
rect 264 1072 296 1088
rect 488 1072 504 1088
rect 520 1072 536 1088
rect 584 1072 600 1088
rect 472 1052 488 1068
rect 648 1072 664 1088
rect 760 1072 776 1088
rect 792 1072 808 1088
rect 872 1072 888 1088
rect 1032 1072 1048 1088
rect 1128 1072 1144 1088
rect 1208 1072 1224 1088
rect 664 1052 696 1068
rect 872 1052 888 1068
rect 1144 1052 1160 1068
rect 1176 1052 1192 1068
rect 1256 1072 1272 1088
rect 1288 1072 1304 1088
rect 1336 1072 1352 1088
rect 1480 1072 1496 1088
rect 1544 1072 1560 1088
rect 1656 1072 1672 1088
rect 1752 1072 1768 1088
rect 1816 1072 1832 1088
rect 1896 1072 1912 1088
rect 1944 1072 1960 1088
rect 1976 1072 1992 1088
rect 2056 1072 2072 1088
rect 2168 1072 2184 1088
rect 2216 1072 2232 1088
rect 2328 1072 2344 1088
rect 2456 1072 2472 1088
rect 2520 1072 2536 1088
rect 2632 1072 2648 1088
rect 2696 1072 2712 1088
rect 2808 1072 2824 1088
rect 2872 1072 2888 1088
rect 2904 1072 2920 1088
rect 3032 1072 3048 1088
rect 3064 1072 3080 1088
rect 3096 1072 3112 1088
rect 3144 1072 3160 1088
rect 1256 1052 1272 1068
rect 1592 1052 1608 1068
rect 1688 1052 1704 1068
rect 1848 1052 1864 1068
rect 1912 1052 1928 1068
rect 2328 1052 2344 1068
rect 2440 1052 2456 1068
rect 2584 1052 2600 1068
rect 2792 1052 2808 1068
rect 2872 1052 2888 1068
rect 2968 1052 2984 1068
rect 3192 1052 3208 1068
rect 376 1032 392 1048
rect 840 1032 856 1048
rect 888 1032 904 1048
rect 1224 1032 1240 1048
rect 1432 1032 1448 1048
rect 1672 1032 1688 1048
rect 1704 1032 1720 1048
rect 1832 1032 1848 1048
rect 1880 1032 1896 1048
rect 1928 1032 1944 1048
rect 2504 1032 2520 1048
rect 2600 1032 2616 1048
rect 2744 1032 2760 1048
rect 2776 1032 2792 1048
rect 2888 1032 2904 1048
rect 3016 1032 3032 1048
rect 3080 1032 3096 1048
rect 2077 1002 2113 1018
rect 216 972 232 988
rect 472 972 488 988
rect 616 972 632 988
rect 712 972 728 988
rect 872 972 888 988
rect 1000 972 1016 988
rect 1784 972 1800 988
rect 2392 972 2408 988
rect 2472 972 2488 988
rect 2696 972 2712 988
rect 344 952 360 968
rect 408 952 424 968
rect 488 952 504 968
rect 520 952 536 968
rect 568 952 584 968
rect 600 952 616 968
rect 888 952 920 968
rect 1368 952 1384 968
rect 1416 952 1432 968
rect 24 932 40 948
rect 232 932 264 948
rect 312 932 328 948
rect 360 932 376 948
rect 424 932 440 948
rect 584 932 600 948
rect 632 932 648 948
rect 696 932 712 948
rect 760 932 776 948
rect 792 932 808 948
rect 824 932 840 948
rect 856 932 872 948
rect 936 932 952 948
rect 1176 932 1192 948
rect 1208 932 1240 948
rect 1288 932 1304 948
rect 1400 932 1416 948
rect 1432 932 1464 948
rect 1544 952 1560 968
rect 1576 952 1592 968
rect 1768 952 1784 968
rect 2136 952 2168 968
rect 2344 952 2360 968
rect 2408 952 2424 968
rect 2536 952 2552 968
rect 2664 952 2680 968
rect 1624 932 1640 948
rect 1688 932 1704 948
rect 1800 932 1816 948
rect 1832 932 1848 948
rect 1896 932 1912 948
rect 1992 932 2008 948
rect 2040 932 2056 948
rect 2104 932 2120 948
rect 2344 932 2360 948
rect 2424 944 2440 948
rect 2424 932 2456 944
rect 2504 932 2520 948
rect 2616 932 2632 948
rect 2744 932 2760 948
rect 2792 932 2808 948
rect 2920 932 2952 948
rect 3000 932 3016 948
rect 3048 932 3080 948
rect 3192 932 3208 948
rect 2440 928 2456 932
rect 8 912 40 928
rect 72 912 104 928
rect 120 912 136 928
rect 168 912 184 928
rect 232 912 248 928
rect 312 912 328 928
rect 440 912 456 928
rect 488 912 504 928
rect 536 912 552 928
rect 648 912 664 928
rect 744 912 760 928
rect 824 912 856 928
rect 920 912 936 928
rect 952 912 968 928
rect 984 912 1000 928
rect 1032 912 1064 928
rect 1096 912 1128 928
rect 1160 912 1176 928
rect 1240 912 1256 928
rect 200 892 216 908
rect 296 892 312 908
rect 408 892 424 908
rect 472 892 488 908
rect 664 892 680 908
rect 696 892 728 908
rect 776 892 792 908
rect 1252 892 1268 908
rect 1304 912 1320 928
rect 1416 912 1432 928
rect 1480 912 1496 928
rect 1576 912 1592 928
rect 1720 912 1736 928
rect 1816 912 1832 928
rect 1848 912 1864 928
rect 1912 912 1928 928
rect 1336 892 1352 908
rect 1656 892 1672 908
rect 1704 892 1720 908
rect 1848 892 1864 908
rect 1880 892 1896 908
rect 2088 912 2104 928
rect 2200 912 2216 928
rect 2248 912 2264 928
rect 2280 912 2296 928
rect 2312 912 2328 928
rect 2360 912 2376 928
rect 2488 912 2504 928
rect 2568 912 2584 928
rect 2616 912 2632 928
rect 2728 912 2744 928
rect 2776 912 2792 928
rect 2824 912 2840 928
rect 2904 912 2920 928
rect 2952 912 2968 928
rect 2984 912 3016 928
rect 3032 912 3048 928
rect 3096 912 3112 928
rect 3144 912 3160 928
rect 1960 892 1976 908
rect 2008 892 2024 908
rect 2152 892 2168 908
rect 2184 892 2200 908
rect 2248 892 2264 908
rect 2536 892 2568 908
rect 2600 892 2616 908
rect 2744 892 2760 908
rect 2808 892 2824 908
rect 2872 892 2888 908
rect 1736 872 1752 888
rect 2216 872 2232 888
rect 2584 872 2600 888
rect 2840 872 2856 888
rect 152 832 168 848
rect 1192 832 1208 848
rect 1528 832 1544 848
rect 1592 832 1608 848
rect 1720 832 1736 848
rect 1912 832 1928 848
rect 2024 832 2040 848
rect 2168 832 2184 848
rect 2200 832 2216 848
rect 2664 832 2680 848
rect 2856 832 2872 848
rect 2904 832 2920 848
rect 3128 832 3144 848
rect 1037 802 1073 818
rect 40 772 56 788
rect 600 772 616 788
rect 824 772 840 788
rect 1208 772 1224 788
rect 1720 772 1736 788
rect 2296 772 2312 788
rect 2728 772 2744 788
rect 2936 772 2952 788
rect 3192 752 3208 768
rect 680 732 696 748
rect 1592 732 1608 748
rect 1992 732 2008 748
rect 2456 732 2472 748
rect 3128 732 3144 748
rect 264 712 296 728
rect 372 712 388 728
rect 392 712 408 728
rect 504 712 520 728
rect 568 712 584 728
rect 632 712 664 728
rect 1000 712 1016 728
rect 1128 712 1160 728
rect 1224 712 1240 728
rect 1272 712 1288 728
rect 1400 712 1416 728
rect 8 692 24 708
rect 88 692 104 708
rect 216 692 232 708
rect 312 692 328 708
rect 424 692 440 708
rect 488 692 520 708
rect 584 692 616 708
rect 664 692 680 708
rect 872 692 888 708
rect 920 692 968 708
rect 1032 692 1048 708
rect 72 672 88 688
rect 136 672 152 688
rect 216 672 232 688
rect 328 672 360 688
rect 408 672 424 688
rect 472 672 488 688
rect 520 672 536 688
rect 584 672 600 688
rect 712 672 728 688
rect 808 672 824 688
rect 856 672 872 688
rect 1048 672 1064 688
rect 1096 672 1112 688
rect 1176 672 1192 688
rect 1352 692 1368 708
rect 1416 692 1432 708
rect 1560 712 1576 728
rect 1624 712 1640 728
rect 1704 712 1720 728
rect 2024 712 2040 728
rect 2136 712 2152 728
rect 2216 712 2248 728
rect 2328 712 2344 728
rect 1496 692 1512 708
rect 1528 692 1544 708
rect 1608 692 1624 708
rect 1640 692 1656 708
rect 1912 692 1928 708
rect 2008 692 2024 708
rect 2040 692 2056 708
rect 2088 692 2104 708
rect 2184 692 2200 708
rect 2296 692 2312 708
rect 2344 692 2360 708
rect 2408 692 2424 708
rect 2584 692 2600 708
rect 2760 692 2776 708
rect 2824 692 2840 708
rect 2888 692 2920 708
rect 3016 692 3032 708
rect 3096 692 3112 708
rect 3144 692 3160 708
rect 1880 688 1896 692
rect 1240 672 1256 688
rect 1304 672 1320 688
rect 1336 672 1368 688
rect 1416 672 1432 688
rect 1496 672 1512 688
rect 1656 672 1672 688
rect 1736 672 1752 688
rect 1784 672 1800 688
rect 1880 676 1912 688
rect 1896 672 1912 676
rect 1928 672 1944 688
rect 120 652 136 668
rect 200 652 216 668
rect 840 652 856 668
rect 968 652 984 668
rect 1288 652 1304 668
rect 1464 652 1480 668
rect 1688 652 1704 668
rect 1752 652 1768 668
rect 2072 652 2088 668
rect 2168 672 2184 688
rect 2264 672 2296 688
rect 2360 672 2376 688
rect 2392 672 2408 688
rect 2424 672 2440 688
rect 2520 672 2536 688
rect 2600 672 2616 688
rect 2712 672 2728 688
rect 2776 672 2792 688
rect 3000 672 3016 688
rect 3000 652 3032 668
rect 456 632 472 648
rect 568 632 584 648
rect 680 632 696 648
rect 776 632 792 648
rect 1128 632 1144 648
rect 1256 632 1272 648
rect 1432 632 1448 648
rect 1480 632 1496 648
rect 1560 632 1576 648
rect 1608 632 1624 648
rect 1672 632 1688 648
rect 1832 632 1848 648
rect 1944 632 1960 648
rect 2056 632 2072 648
rect 2216 632 2232 648
rect 2248 632 2264 648
rect 2360 632 2376 648
rect 2552 632 2568 648
rect 2664 632 2680 648
rect 2856 632 2872 648
rect 2077 602 2113 618
rect 200 572 216 588
rect 520 572 536 588
rect 584 572 600 588
rect 648 572 664 588
rect 824 572 840 588
rect 1368 572 1384 588
rect 1688 572 1704 588
rect 1736 572 1752 588
rect 1960 572 1976 588
rect 2168 572 2184 588
rect 2264 572 2280 588
rect 2392 572 2408 588
rect 184 552 200 568
rect 840 552 856 568
rect 1160 552 1176 568
rect 1256 552 1272 568
rect 1400 552 1416 568
rect 1464 552 1480 568
rect 1816 552 1832 568
rect 1848 552 1864 568
rect 2040 552 2056 568
rect 2184 552 2200 568
rect 2248 552 2264 568
rect 2920 552 2936 568
rect 56 532 72 548
rect 24 512 40 528
rect 136 532 152 548
rect 408 532 424 548
rect 472 532 488 548
rect 600 532 616 548
rect 776 532 792 548
rect 808 532 824 548
rect 952 532 968 548
rect 120 512 136 528
rect 184 512 200 528
rect 232 512 248 528
rect 296 512 312 528
rect 376 512 392 528
rect 456 512 472 528
rect 488 512 504 528
rect 536 512 568 528
rect 616 512 632 528
rect 792 512 808 528
rect 872 512 888 528
rect 920 512 936 528
rect 1176 532 1192 548
rect 1240 532 1256 548
rect 1384 532 1400 548
rect 1432 532 1448 548
rect 1576 532 1592 548
rect 1848 532 1864 548
rect 2152 532 2168 548
rect 2200 532 2216 548
rect 2344 532 2360 548
rect 2408 532 2424 548
rect 2520 532 2552 548
rect 2584 532 2600 548
rect 2616 532 2632 548
rect 2712 532 2744 548
rect 2824 532 2840 548
rect 1016 512 1048 528
rect 1064 512 1080 528
rect 1192 512 1208 528
rect 1224 512 1240 528
rect 1272 512 1288 528
rect 1320 512 1336 528
rect 1480 512 1512 528
rect 1544 512 1560 528
rect 1592 512 1608 528
rect 1640 512 1672 528
rect 1784 512 1800 528
rect 1880 512 1896 528
rect 1928 512 1944 528
rect 2024 512 2040 528
rect 2296 512 2312 528
rect 2360 512 2376 528
rect 2424 512 2440 528
rect 2472 512 2520 528
rect 2536 512 2552 528
rect 2568 512 2584 528
rect 2600 512 2616 528
rect 2872 532 2888 548
rect 2920 532 2936 548
rect 3080 532 3096 548
rect 3112 532 3128 548
rect 3192 532 3208 548
rect 2888 512 2904 528
rect 2984 512 3000 528
rect 3032 512 3048 528
rect 3064 512 3080 528
rect 3128 512 3160 528
rect 8 492 24 508
rect 168 492 184 508
rect 216 492 232 508
rect 296 492 312 508
rect 392 492 408 508
rect 568 492 584 508
rect 856 492 872 508
rect 920 492 936 508
rect 1000 492 1016 508
rect 1096 492 1112 508
rect 1336 492 1352 508
rect 1400 492 1416 508
rect 1464 492 1480 508
rect 1672 492 1688 508
rect 1944 492 1960 508
rect 2120 492 2136 508
rect 2216 492 2248 508
rect 2280 492 2296 508
rect 2392 492 2408 508
rect 2472 492 2488 508
rect 2872 492 2888 508
rect 2920 492 2936 508
rect 3048 492 3064 508
rect 3080 492 3096 508
rect 232 472 264 488
rect 312 472 328 488
rect 360 472 376 488
rect 888 472 904 488
rect 1304 472 1320 488
rect 1624 472 1640 488
rect 1912 472 1928 488
rect 2312 472 2328 488
rect 2648 472 2664 488
rect 3016 472 3032 488
rect 296 452 312 468
rect 872 452 888 468
rect 88 432 104 448
rect 264 432 280 448
rect 376 432 392 448
rect 712 432 728 448
rect 1224 432 1240 448
rect 1320 432 1336 448
rect 1864 432 1880 448
rect 1928 432 1944 448
rect 2328 432 2344 448
rect 3000 432 3016 448
rect 1037 402 1073 418
rect 488 372 504 388
rect 728 372 744 388
rect 792 372 808 388
rect 1000 372 1016 388
rect 1288 372 1304 388
rect 1352 372 1368 388
rect 2408 372 2424 388
rect 3128 372 3144 388
rect 664 352 680 368
rect 1992 352 2008 368
rect 472 332 488 348
rect 552 332 568 348
rect 648 332 664 348
rect 712 332 728 348
rect 776 332 792 348
rect 1016 332 1032 348
rect 1160 332 1176 348
rect 1272 332 1288 348
rect 1336 332 1352 348
rect 1816 332 1832 348
rect 1848 332 1864 348
rect 2168 332 2184 348
rect 24 292 40 308
rect 56 292 72 308
rect 104 292 120 308
rect 152 312 168 328
rect 248 312 264 328
rect 408 312 424 328
rect 504 312 520 328
rect 616 312 632 328
rect 680 312 696 328
rect 744 312 760 328
rect 808 312 840 328
rect 936 312 952 328
rect 984 312 1000 328
rect 1112 312 1144 328
rect 1304 312 1320 328
rect 1368 312 1384 328
rect 1432 312 1448 328
rect 1496 312 1512 328
rect 1544 312 1560 328
rect 1656 312 1688 328
rect 1880 312 1896 328
rect 1944 312 1960 328
rect 2104 312 2120 328
rect 2200 312 2216 328
rect 2232 312 2248 328
rect 2264 312 2280 328
rect 2312 312 2328 328
rect 2344 312 2360 328
rect 2376 312 2392 328
rect 2456 312 2472 328
rect 2488 312 2520 328
rect 216 292 232 308
rect 280 292 296 308
rect 8 272 24 288
rect 72 286 104 288
rect 56 272 104 286
rect 184 272 216 288
rect 248 272 280 288
rect 344 292 360 308
rect 376 292 392 308
rect 488 292 504 308
rect 520 292 536 308
rect 664 292 680 308
rect 728 292 744 308
rect 792 292 808 308
rect 1000 292 1016 308
rect 1144 292 1160 308
rect 1224 292 1240 308
rect 1288 292 1304 308
rect 1352 292 1368 308
rect 1400 292 1416 308
rect 1464 292 1480 308
rect 1576 292 1608 308
rect 1624 292 1640 308
rect 1672 292 1688 308
rect 1768 292 1784 308
rect 1816 292 1848 308
rect 2008 292 2024 308
rect 2184 292 2200 308
rect 2232 292 2248 308
rect 2344 292 2360 308
rect 2408 292 2424 308
rect 2760 292 2776 308
rect 2872 292 2888 308
rect 2904 292 2920 308
rect 2968 292 2984 308
rect 3000 292 3016 308
rect 3064 292 3080 308
rect 56 270 72 272
rect 376 270 392 286
rect 440 272 456 288
rect 568 272 584 288
rect 856 272 872 288
rect 888 272 904 288
rect 968 272 984 288
rect 1080 272 1096 288
rect 1176 272 1192 288
rect 1240 272 1256 288
rect 1384 272 1400 288
rect 1448 272 1464 288
rect 1512 272 1528 288
rect 1608 272 1624 288
rect 1688 272 1704 288
rect 1720 272 1736 288
rect 1832 272 1848 288
rect 1896 272 1912 288
rect 1976 272 1992 288
rect 2136 272 2152 288
rect 2216 272 2232 288
rect 2280 272 2296 288
rect 2328 272 2344 288
rect 2392 272 2408 288
rect 2456 272 2472 288
rect 2488 272 2504 288
rect 2552 272 2568 288
rect 2584 272 2600 288
rect 2712 272 2728 288
rect 2744 272 2760 288
rect 2888 272 2904 288
rect 2920 272 2936 288
rect 2952 272 2968 288
rect 3048 272 3064 288
rect 3112 272 3128 288
rect 136 252 152 268
rect 824 252 840 268
rect 920 252 936 268
rect 1432 252 1448 268
rect 1496 252 1512 268
rect 1560 252 1576 268
rect 1736 252 1752 268
rect 1784 252 1800 268
rect 2008 252 2024 268
rect 2056 252 2088 268
rect 2488 252 2504 268
rect 2584 252 2600 268
rect 2728 252 2744 268
rect 168 232 184 248
rect 600 232 616 248
rect 904 232 920 248
rect 952 232 968 248
rect 1112 232 1128 248
rect 1192 232 1208 248
rect 1544 232 1560 248
rect 1912 232 1928 248
rect 1944 232 1960 248
rect 2040 232 2056 248
rect 2152 232 2168 248
rect 2296 232 2312 248
rect 2632 232 2648 248
rect 2792 232 2808 248
rect 2840 232 2856 248
rect 2936 232 2952 248
rect 3032 232 3048 248
rect 3096 232 3112 248
rect 2077 202 2113 218
rect 56 172 72 188
rect 408 172 424 188
rect 504 172 520 188
rect 552 172 568 188
rect 1528 172 1544 188
rect 1576 172 1592 188
rect 1928 172 1944 188
rect 2248 172 2264 188
rect 2952 172 2968 188
rect 232 152 248 168
rect 536 152 552 168
rect 1032 152 1048 168
rect 1176 152 1192 168
rect 1304 152 1320 168
rect 1368 152 1384 168
rect 1608 152 1624 168
rect 1640 152 1656 168
rect 1704 152 1736 168
rect 1768 152 1784 168
rect 1800 152 1816 168
rect 2024 152 2040 168
rect 2296 152 2312 168
rect 2408 152 2424 168
rect 2488 152 2504 168
rect 2952 152 2968 168
rect 8 132 24 148
rect 104 132 120 148
rect 152 132 168 148
rect 312 132 328 148
rect 488 132 504 148
rect 840 132 856 148
rect 936 132 952 148
rect 1000 132 1016 148
rect 1064 132 1080 148
rect 1256 132 1288 148
rect 1384 144 1400 148
rect 1384 132 1416 144
rect 1496 132 1528 148
rect 1608 132 1624 148
rect 1656 132 1688 148
rect 1736 132 1752 148
rect 1864 132 1896 148
rect 2120 132 2136 148
rect 2184 132 2200 148
rect 2296 132 2312 148
rect 2472 132 2488 148
rect 2600 132 2616 148
rect 2984 132 3000 148
rect 3192 132 3208 148
rect 1400 128 1416 132
rect 88 112 104 128
rect 120 112 136 128
rect 200 112 216 128
rect 264 112 280 128
rect 328 112 344 128
rect 376 112 392 128
rect 456 112 472 128
rect 584 112 600 128
rect 664 112 680 128
rect 728 112 744 128
rect 792 112 824 128
rect 888 112 904 128
rect 952 112 968 128
rect 984 112 1000 128
rect 1112 112 1128 128
rect 1144 112 1160 128
rect 184 92 200 108
rect 248 92 264 108
rect 344 92 376 108
rect 424 92 440 108
rect 472 92 488 108
rect 520 92 536 108
rect 616 92 632 108
rect 680 92 696 108
rect 744 92 760 108
rect 888 92 904 108
rect 968 92 984 108
rect 1128 92 1144 108
rect 1224 112 1240 128
rect 1256 112 1272 128
rect 1336 112 1352 128
rect 1448 112 1464 128
rect 1480 112 1496 128
rect 1688 112 1704 128
rect 1752 112 1768 128
rect 1800 112 1816 128
rect 1848 112 1864 128
rect 1896 112 1912 128
rect 1944 112 1960 128
rect 1992 112 2008 128
rect 2024 112 2040 128
rect 2136 112 2152 128
rect 2408 112 2424 128
rect 2440 112 2456 128
rect 2536 112 2552 128
rect 2584 112 2600 128
rect 2616 112 2632 128
rect 2664 112 2680 128
rect 2712 112 2728 128
rect 2776 112 2792 128
rect 2808 112 2824 128
rect 2856 112 2872 128
rect 2936 112 2952 128
rect 3032 112 3064 128
rect 3096 112 3112 128
rect 3144 112 3160 128
rect 1224 92 1240 108
rect 1304 92 1336 108
rect 1448 92 1464 108
rect 1480 92 1496 108
rect 1544 92 1576 108
rect 1816 92 1832 108
rect 2008 92 2024 108
rect 2148 92 2164 108
rect 2168 92 2184 108
rect 2424 92 2440 108
rect 2552 92 2568 108
rect 2584 92 2600 108
rect 2760 92 2776 108
rect 216 72 232 88
rect 280 72 296 88
rect 392 72 408 88
rect 440 72 456 88
rect 648 72 664 88
rect 712 72 728 88
rect 776 72 792 88
rect 872 72 888 88
rect 936 72 952 88
rect 1096 72 1112 88
rect 1352 72 1368 88
rect 1800 72 1816 88
rect 2392 72 2408 88
rect 2792 72 2808 88
rect 264 52 280 68
rect 664 52 680 68
rect 728 52 744 68
rect 792 52 808 68
rect 888 52 904 68
rect 1112 52 1128 68
rect 584 32 600 48
rect 1976 32 1992 48
rect 2104 32 2120 48
rect 2360 32 2376 48
rect 2504 32 2520 48
rect 2648 32 2664 48
rect 2696 32 2712 48
rect 2744 32 2760 48
rect 2824 32 2840 48
rect 3000 32 3016 48
rect 3080 32 3096 48
rect 3128 32 3144 48
rect 1037 2 1073 18
<< metal2 >>
rect 93 2128 99 2263
rect 13 1908 19 2112
rect 13 1568 19 1712
rect 13 1508 19 1552
rect 13 1328 19 1452
rect 13 1048 19 1312
rect 29 1188 35 1892
rect 61 1748 67 2112
rect 93 2108 99 2112
rect 141 2088 147 2112
rect 157 1928 163 2132
rect 189 2128 195 2172
rect 237 2128 243 2263
rect 285 2128 291 2263
rect 349 2128 355 2132
rect 365 2128 371 2152
rect 381 2128 387 2132
rect 477 2128 483 2132
rect 541 2128 547 2152
rect 669 2128 675 2263
rect 701 2148 707 2152
rect 717 2128 723 2263
rect 781 2148 787 2152
rect 749 2128 755 2132
rect 189 2088 195 2112
rect 157 1908 163 1912
rect 189 1908 195 1912
rect 77 1888 83 1892
rect 93 1748 99 1892
rect 173 1888 179 1892
rect 157 1868 163 1872
rect 237 1848 243 1892
rect 221 1808 227 1832
rect 77 1728 83 1732
rect 189 1728 195 1732
rect 77 1508 83 1712
rect 93 1688 99 1712
rect 141 1708 147 1712
rect 173 1668 179 1672
rect 93 1508 99 1572
rect 173 1548 179 1652
rect 141 1508 147 1532
rect 45 1448 51 1472
rect 45 1328 51 1432
rect 77 1368 83 1372
rect 125 1368 131 1432
rect 141 1408 147 1492
rect 173 1463 179 1532
rect 221 1468 227 1492
rect 237 1488 243 1712
rect 253 1708 259 2112
rect 285 1888 291 2112
rect 333 2108 339 2112
rect 397 1908 403 2052
rect 525 2048 531 2112
rect 669 2068 675 2112
rect 733 2068 739 2112
rect 413 1988 419 2032
rect 509 1948 515 2032
rect 557 1928 563 1952
rect 573 1908 579 2032
rect 733 2028 739 2052
rect 333 1888 339 1892
rect 349 1888 355 1892
rect 269 1768 275 1872
rect 269 1728 275 1752
rect 317 1748 323 1752
rect 349 1728 355 1752
rect 365 1588 371 1712
rect 381 1508 387 1532
rect 397 1528 403 1892
rect 413 1728 419 1892
rect 525 1888 531 1892
rect 429 1848 435 1852
rect 573 1788 579 1892
rect 429 1728 435 1732
rect 445 1728 451 1752
rect 477 1728 483 1732
rect 637 1728 643 1892
rect 653 1768 659 1892
rect 733 1868 739 1912
rect 781 1908 787 2012
rect 797 1968 803 2132
rect 861 2128 867 2263
rect 1101 2228 1107 2263
rect 1064 2157 1107 2163
rect 893 2128 899 2152
rect 925 2128 931 2152
rect 1005 2148 1011 2152
rect 1101 2148 1107 2157
rect 1085 2128 1091 2132
rect 1149 2128 1155 2152
rect 813 1968 819 2112
rect 861 2048 867 2112
rect 877 2068 883 2112
rect 925 2028 931 2112
rect 941 2108 947 2112
rect 957 2008 963 2032
rect 797 1888 803 1952
rect 877 1888 883 1912
rect 669 1788 675 1812
rect 813 1768 819 1832
rect 509 1568 515 1712
rect 541 1708 547 1712
rect 445 1508 451 1552
rect 285 1488 291 1492
rect 157 1457 179 1463
rect 77 1328 83 1352
rect 45 968 51 1312
rect 141 1308 147 1332
rect 61 1288 67 1292
rect 93 1108 99 1112
rect 13 928 19 952
rect 29 908 35 912
rect 45 788 51 912
rect 13 708 19 772
rect 61 548 67 972
rect 77 928 83 1032
rect 109 988 115 1232
rect 93 928 99 952
rect 93 708 99 852
rect 93 608 99 692
rect 13 328 19 492
rect 29 308 35 512
rect 61 308 67 312
rect 93 308 99 432
rect 109 308 115 952
rect 125 928 131 1192
rect 141 1108 147 1132
rect 125 908 131 912
rect 141 768 147 1072
rect 157 923 163 1457
rect 173 1348 179 1432
rect 221 1328 227 1392
rect 269 1328 275 1372
rect 173 968 179 1232
rect 253 1168 259 1232
rect 285 1208 291 1472
rect 333 1448 339 1492
rect 333 1388 339 1432
rect 301 1328 307 1352
rect 365 1348 371 1492
rect 429 1468 435 1472
rect 413 1348 419 1432
rect 365 1328 371 1332
rect 493 1328 499 1512
rect 525 1468 531 1492
rect 541 1488 547 1692
rect 589 1668 595 1712
rect 637 1648 643 1712
rect 557 1588 563 1632
rect 653 1628 659 1752
rect 701 1728 707 1752
rect 685 1703 691 1712
rect 685 1697 696 1703
rect 605 1508 611 1612
rect 701 1588 707 1692
rect 717 1588 723 1732
rect 765 1728 771 1732
rect 845 1648 851 1692
rect 685 1508 691 1532
rect 733 1508 739 1572
rect 765 1508 771 1552
rect 781 1548 787 1632
rect 845 1508 851 1632
rect 541 1328 547 1372
rect 557 1328 563 1492
rect 573 1448 579 1492
rect 573 1428 579 1432
rect 605 1368 611 1472
rect 621 1348 627 1472
rect 637 1348 643 1432
rect 333 1128 339 1312
rect 413 1188 419 1232
rect 205 1088 211 1092
rect 221 988 227 1112
rect 349 1108 355 1132
rect 413 1108 419 1152
rect 157 917 168 923
rect 157 868 163 917
rect 157 808 163 832
rect 141 688 147 752
rect 189 568 195 932
rect 205 908 211 952
rect 237 948 243 1092
rect 269 1088 275 1092
rect 237 928 243 932
rect 301 928 307 1092
rect 317 1048 323 1092
rect 477 1068 483 1072
rect 349 968 355 1012
rect 381 988 387 1032
rect 493 1028 499 1072
rect 509 1068 515 1232
rect 541 1108 547 1152
rect 605 1128 611 1312
rect 605 1108 611 1112
rect 621 1108 627 1332
rect 653 1128 659 1452
rect 685 1448 691 1492
rect 749 1388 755 1492
rect 861 1488 867 1712
rect 893 1648 899 1852
rect 909 1848 915 1892
rect 957 1888 963 1972
rect 989 1968 995 2092
rect 1021 2048 1027 2112
rect 1069 2108 1075 2112
rect 1085 2068 1091 2112
rect 1229 2108 1235 2263
rect 1309 2148 1315 2152
rect 1517 2148 1523 2263
rect 1645 2148 1651 2152
rect 1501 2137 1512 2143
rect 1293 2108 1299 2112
rect 1021 1928 1027 1992
rect 1064 1937 1107 1943
rect 1101 1923 1107 1937
rect 1101 1917 1112 1923
rect 989 1897 1043 1903
rect 989 1883 995 1897
rect 1037 1888 1043 1897
rect 1053 1888 1059 1912
rect 1085 1908 1091 1912
rect 973 1877 995 1883
rect 973 1863 979 1877
rect 968 1857 979 1863
rect 925 1748 931 1832
rect 909 1708 915 1712
rect 909 1648 915 1692
rect 861 1408 867 1452
rect 749 1328 755 1372
rect 829 1328 835 1392
rect 861 1328 867 1372
rect 877 1328 883 1512
rect 957 1508 963 1752
rect 989 1748 995 1752
rect 973 1708 979 1732
rect 989 1668 995 1692
rect 1005 1488 1011 1792
rect 1021 1748 1027 1872
rect 1133 1868 1139 1912
rect 1165 1908 1171 1952
rect 1181 1908 1187 1932
rect 1101 1788 1107 1812
rect 1037 1748 1043 1752
rect 1149 1748 1155 1792
rect 1181 1748 1187 1872
rect 1021 1708 1027 1712
rect 1085 1708 1091 1732
rect 1021 1508 1027 1512
rect 701 1168 707 1312
rect 893 1288 899 1432
rect 1021 1348 1027 1492
rect 1069 1488 1075 1532
rect 1128 1517 1139 1523
rect 1037 1328 1043 1392
rect 1101 1328 1107 1452
rect 1133 1388 1139 1517
rect 1165 1508 1171 1712
rect 1165 1483 1171 1492
rect 1197 1488 1203 2092
rect 1213 1883 1219 2072
rect 1309 1968 1315 2112
rect 1373 2088 1379 2132
rect 1389 2128 1395 2132
rect 1245 1888 1251 1892
rect 1213 1877 1224 1883
rect 1229 1788 1235 1832
rect 1213 1748 1219 1752
rect 1245 1728 1251 1752
rect 1261 1748 1267 1952
rect 1277 1848 1283 1932
rect 1309 1928 1315 1952
rect 1293 1908 1299 1912
rect 1309 1897 1320 1903
rect 1309 1883 1315 1897
rect 1341 1888 1347 1912
rect 1389 1908 1395 1912
rect 1421 1908 1427 1912
rect 1304 1877 1315 1883
rect 1373 1848 1379 1852
rect 1277 1828 1283 1832
rect 1357 1748 1363 1752
rect 1437 1748 1443 1872
rect 1469 1808 1475 1892
rect 1485 1888 1491 1912
rect 1501 1868 1507 2137
rect 1597 2128 1603 2132
rect 1805 2128 1811 2263
rect 1965 2208 1971 2263
rect 1917 2128 1923 2152
rect 1517 1888 1523 1892
rect 1517 1848 1523 1852
rect 1501 1808 1507 1832
rect 1373 1728 1379 1732
rect 1437 1728 1443 1732
rect 1213 1688 1219 1712
rect 1309 1688 1315 1692
rect 1341 1628 1347 1632
rect 1389 1588 1395 1712
rect 1453 1688 1459 1712
rect 1501 1708 1507 1712
rect 1485 1588 1491 1632
rect 1389 1568 1395 1572
rect 1165 1477 1187 1483
rect 1165 1328 1171 1392
rect 1181 1368 1187 1477
rect 1197 1408 1203 1452
rect 1213 1348 1219 1532
rect 1277 1488 1283 1552
rect 1373 1488 1379 1492
rect 973 1308 979 1312
rect 1149 1308 1155 1312
rect 893 1263 899 1272
rect 877 1257 899 1263
rect 477 988 483 992
rect 221 723 227 912
rect 205 717 227 723
rect 205 688 211 717
rect 237 708 243 912
rect 317 908 323 912
rect 301 748 307 892
rect 285 728 291 732
rect 317 723 323 892
rect 301 717 323 723
rect 205 668 211 672
rect 221 643 227 672
rect 205 637 227 643
rect 205 588 211 637
rect 141 548 147 552
rect 125 528 131 532
rect 93 288 99 292
rect 13 248 19 272
rect 77 268 83 272
rect 61 188 67 232
rect 13 128 19 132
rect 93 128 99 212
rect 125 128 131 512
rect 157 308 163 312
rect 173 308 179 492
rect 189 288 195 372
rect 221 328 227 492
rect 237 303 243 472
rect 269 428 275 432
rect 285 308 291 652
rect 301 528 307 717
rect 349 688 355 792
rect 381 728 387 932
rect 445 928 451 952
rect 477 928 483 932
rect 413 908 419 912
rect 477 908 483 912
rect 493 908 499 912
rect 397 728 403 732
rect 413 688 419 752
rect 429 708 435 712
rect 477 688 483 752
rect 509 728 515 1012
rect 541 928 547 1092
rect 589 1088 595 1092
rect 653 1088 659 1112
rect 765 1108 771 1172
rect 797 1108 803 1232
rect 813 1108 819 1112
rect 845 1108 851 1152
rect 877 1088 883 1257
rect 893 1188 899 1232
rect 941 1108 947 1252
rect 989 1108 995 1232
rect 1117 1128 1123 1232
rect 1117 1108 1123 1112
rect 909 1088 915 1092
rect 621 988 627 1012
rect 541 788 547 912
rect 589 868 595 932
rect 509 708 515 712
rect 525 688 531 752
rect 589 708 595 852
rect 637 848 643 932
rect 669 908 675 1032
rect 717 988 723 1052
rect 765 1048 771 1072
rect 701 948 707 972
rect 765 948 771 1032
rect 845 1008 851 1032
rect 797 948 803 952
rect 829 948 835 972
rect 861 963 867 1052
rect 877 988 883 992
rect 893 968 899 1032
rect 909 968 915 992
rect 925 988 931 1092
rect 941 1008 947 1092
rect 845 957 867 963
rect 717 908 723 932
rect 845 928 851 957
rect 941 948 947 952
rect 605 788 611 832
rect 669 748 675 892
rect 685 748 691 812
rect 749 768 755 912
rect 829 788 835 912
rect 333 668 339 672
rect 301 468 307 472
rect 232 297 243 303
rect 205 288 211 292
rect 253 288 259 292
rect 173 128 179 232
rect 253 108 259 192
rect 269 148 275 272
rect 285 268 291 292
rect 317 188 323 472
rect 349 323 355 672
rect 461 528 467 632
rect 477 548 483 632
rect 525 588 531 612
rect 589 588 595 652
rect 493 528 499 552
rect 605 548 611 692
rect 637 668 643 712
rect 813 688 819 772
rect 829 748 835 772
rect 845 708 851 912
rect 861 848 867 932
rect 957 928 963 1092
rect 925 908 931 912
rect 925 708 931 712
rect 941 708 947 712
rect 957 708 963 712
rect 973 683 979 992
rect 989 928 995 1092
rect 1005 1028 1011 1072
rect 1005 988 1011 1012
rect 1053 988 1059 1092
rect 957 677 979 683
rect 717 648 723 672
rect 381 348 387 432
rect 333 317 355 323
rect 333 143 339 317
rect 328 137 339 143
rect 317 128 323 132
rect 349 108 355 132
rect 365 108 371 312
rect 381 308 387 312
rect 397 308 403 492
rect 493 388 499 472
rect 413 328 419 332
rect 509 328 515 392
rect 525 308 531 532
rect 605 528 611 532
rect 621 528 627 532
rect 541 508 547 512
rect 504 297 515 303
rect 397 208 403 292
rect 493 288 499 292
rect 413 188 419 192
rect 509 188 515 297
rect 573 288 579 492
rect 653 348 659 372
rect 621 328 627 332
rect 685 328 691 632
rect 717 556 723 632
rect 781 568 787 632
rect 829 588 835 632
rect 861 563 867 672
rect 856 557 867 563
rect 717 408 723 432
rect 717 348 723 352
rect 749 328 755 492
rect 797 468 803 512
rect 813 488 819 532
rect 781 348 787 372
rect 829 328 835 332
rect 397 88 403 92
rect 445 88 451 172
rect 541 168 547 252
rect 557 188 563 252
rect 493 148 499 152
rect 525 108 531 132
rect 541 88 547 152
rect 589 128 595 132
rect 605 103 611 232
rect 669 128 675 292
rect 685 188 691 312
rect 733 268 739 292
rect 749 248 755 312
rect 621 108 627 112
rect 669 108 675 112
rect 685 108 691 172
rect 749 108 755 232
rect 797 208 803 292
rect 813 208 819 312
rect 813 128 819 192
rect 845 168 851 552
rect 957 548 963 677
rect 861 488 867 492
rect 893 468 899 472
rect 893 288 899 352
rect 925 348 931 492
rect 989 363 995 912
rect 1005 728 1011 932
rect 1053 868 1059 912
rect 1069 908 1075 1092
rect 1149 1068 1155 1172
rect 1181 1108 1187 1232
rect 1197 1108 1203 1332
rect 1229 1328 1235 1332
rect 1261 1328 1267 1472
rect 1389 1468 1395 1552
rect 1453 1508 1459 1532
rect 1485 1528 1491 1572
rect 1293 1288 1299 1292
rect 1101 928 1107 972
rect 1117 928 1123 952
rect 1181 948 1187 952
rect 1197 943 1203 1092
rect 1213 1088 1219 1092
rect 1229 988 1235 1032
rect 1197 937 1208 943
rect 1037 728 1043 752
rect 1037 708 1043 712
rect 1053 628 1059 672
rect 1037 528 1043 572
rect 1069 528 1075 732
rect 1101 688 1107 852
rect 1133 728 1139 832
rect 1005 468 1011 492
rect 1005 388 1011 452
rect 989 357 1011 363
rect 941 328 947 332
rect 989 308 995 312
rect 1005 308 1011 357
rect 845 148 851 152
rect 861 128 867 272
rect 1005 268 1011 292
rect 925 248 931 252
rect 909 228 915 232
rect 605 97 616 103
rect 877 88 883 172
rect 941 128 947 132
rect 957 128 963 232
rect 973 108 979 232
rect 1021 188 1027 332
rect 1117 328 1123 332
rect 1133 328 1139 632
rect 1149 628 1155 712
rect 1165 568 1171 912
rect 1229 908 1235 932
rect 1245 928 1251 1132
rect 1277 1083 1283 1232
rect 1293 1088 1299 1112
rect 1309 1108 1315 1172
rect 1325 1128 1331 1212
rect 1341 1188 1347 1432
rect 1373 1168 1379 1352
rect 1405 1328 1411 1332
rect 1421 1328 1427 1392
rect 1453 1288 1459 1492
rect 1485 1368 1491 1492
rect 1517 1488 1523 1512
rect 1533 1508 1539 2112
rect 1565 1708 1571 2032
rect 1613 1948 1619 2112
rect 1661 2108 1667 2112
rect 1693 2108 1699 2112
rect 1709 2088 1715 2112
rect 1725 2088 1731 2092
rect 1629 1908 1635 2072
rect 1645 1908 1651 1912
rect 1661 1888 1667 1972
rect 1709 1928 1715 2032
rect 1773 1928 1779 2032
rect 1805 1908 1811 2112
rect 1837 1908 1843 1912
rect 1736 1897 1747 1903
rect 1693 1868 1699 1872
rect 1709 1868 1715 1872
rect 1629 1728 1635 1812
rect 1533 1488 1539 1492
rect 1517 1328 1523 1332
rect 1549 1328 1555 1592
rect 1565 1368 1571 1432
rect 1581 1423 1587 1632
rect 1597 1488 1603 1552
rect 1581 1417 1603 1423
rect 1581 1328 1587 1392
rect 1373 1108 1379 1152
rect 1272 1077 1283 1083
rect 1261 888 1267 892
rect 1197 728 1203 832
rect 1213 788 1219 812
rect 1277 748 1283 1077
rect 1373 1008 1379 1092
rect 1293 948 1299 952
rect 1229 728 1235 732
rect 1197 688 1203 712
rect 1245 688 1251 692
rect 1245 563 1251 672
rect 1261 608 1267 632
rect 1277 588 1283 712
rect 1293 668 1299 932
rect 1309 788 1315 912
rect 1389 908 1395 1232
rect 1469 1228 1475 1232
rect 1405 1048 1411 1092
rect 1421 968 1427 1132
rect 1453 1108 1459 1112
rect 1469 1108 1475 1192
rect 1485 1148 1491 1292
rect 1501 1108 1507 1132
rect 1453 1068 1459 1092
rect 1485 1088 1491 1092
rect 1341 888 1347 892
rect 1405 888 1411 932
rect 1437 928 1443 932
rect 1453 928 1459 932
rect 1421 908 1427 912
rect 1357 708 1363 732
rect 1405 708 1411 712
rect 1421 708 1427 852
rect 1357 648 1363 672
rect 1245 557 1256 563
rect 1165 363 1171 552
rect 1181 528 1187 532
rect 1325 528 1331 592
rect 1373 588 1379 612
rect 1389 548 1395 592
rect 1197 488 1203 512
rect 1293 477 1304 483
rect 1197 468 1203 472
rect 1293 388 1299 477
rect 1325 403 1331 432
rect 1341 428 1347 492
rect 1325 397 1347 403
rect 1149 357 1171 363
rect 1133 308 1139 312
rect 1149 308 1155 357
rect 1085 268 1091 272
rect 1101 88 1107 172
rect 1117 148 1123 232
rect 1133 108 1139 292
rect 1149 288 1155 292
rect 1149 128 1155 212
rect 1165 188 1171 332
rect 1277 288 1283 332
rect 1325 328 1331 372
rect 1341 363 1347 397
rect 1357 388 1363 492
rect 1405 428 1411 472
rect 1421 468 1427 672
rect 1437 608 1443 632
rect 1453 543 1459 772
rect 1469 668 1475 892
rect 1485 808 1491 912
rect 1501 688 1507 692
rect 1469 568 1475 652
rect 1485 608 1491 632
rect 1501 588 1507 672
rect 1448 537 1459 543
rect 1485 528 1491 572
rect 1517 548 1523 1312
rect 1565 1308 1571 1312
rect 1597 1308 1603 1417
rect 1613 1408 1619 1492
rect 1613 1328 1619 1332
rect 1629 1328 1635 1632
rect 1645 1508 1651 1512
rect 1661 1463 1667 1852
rect 1693 1848 1699 1852
rect 1677 1828 1683 1832
rect 1741 1788 1747 1897
rect 1821 1868 1827 1872
rect 1757 1808 1763 1832
rect 1677 1728 1683 1772
rect 1757 1648 1763 1712
rect 1773 1683 1779 1732
rect 1789 1728 1795 1832
rect 1805 1728 1811 1832
rect 1853 1788 1859 1872
rect 1821 1708 1827 1772
rect 1901 1768 1907 1832
rect 1837 1728 1843 1752
rect 1869 1728 1875 1732
rect 1773 1677 1784 1683
rect 1885 1648 1891 1712
rect 1917 1648 1923 2112
rect 1933 2088 1939 2092
rect 1949 2088 1955 2112
rect 1933 1868 1939 2072
rect 1965 1968 1971 2072
rect 1981 1988 1987 2072
rect 1997 1908 2003 2192
rect 2045 2128 2051 2132
rect 2109 2108 2115 2132
rect 2173 2068 2179 2132
rect 2189 2108 2195 2112
rect 2045 1908 2051 1912
rect 2061 1908 2067 2032
rect 1949 1848 1955 1852
rect 1965 1788 1971 1892
rect 1997 1888 2003 1892
rect 1965 1728 1971 1772
rect 1677 1508 1683 1612
rect 1693 1528 1699 1532
rect 1661 1457 1683 1463
rect 1661 1348 1667 1412
rect 1677 1328 1683 1457
rect 1629 1268 1635 1272
rect 1533 1128 1539 1212
rect 1613 1168 1619 1232
rect 1629 1208 1635 1212
rect 1533 1108 1539 1112
rect 1565 1028 1571 1092
rect 1549 968 1555 992
rect 1581 968 1587 1152
rect 1629 1108 1635 1192
rect 1677 1188 1683 1312
rect 1613 1088 1619 1092
rect 1645 948 1651 1092
rect 1661 1088 1667 1092
rect 1693 1068 1699 1432
rect 1709 1368 1715 1632
rect 1773 1628 1779 1632
rect 1773 1528 1779 1552
rect 1725 1368 1731 1412
rect 1741 1403 1747 1432
rect 1789 1408 1795 1432
rect 1741 1397 1763 1403
rect 1709 1108 1715 1112
rect 1661 968 1667 972
rect 1629 928 1635 932
rect 1645 928 1651 932
rect 1581 888 1587 912
rect 1661 908 1667 952
rect 1533 768 1539 832
rect 1597 788 1603 832
rect 1597 748 1603 752
rect 1565 728 1571 732
rect 1629 708 1635 712
rect 1645 708 1651 712
rect 1613 688 1619 692
rect 1661 668 1667 672
rect 1677 668 1683 1032
rect 1709 1028 1715 1032
rect 1709 908 1715 952
rect 1725 908 1731 912
rect 1741 888 1747 1252
rect 1757 1188 1763 1397
rect 1821 1368 1827 1632
rect 1901 1568 1907 1632
rect 1981 1603 1987 1832
rect 2061 1808 2067 1872
rect 2157 1868 2163 1932
rect 2221 1908 2227 1932
rect 2237 1908 2243 2032
rect 2253 1892 2259 2263
rect 2301 2188 2307 2263
rect 2333 2257 2355 2263
rect 2269 2148 2275 2172
rect 2333 2148 2339 2172
rect 2349 2128 2355 2257
rect 2381 2243 2387 2263
rect 2365 2237 2387 2243
rect 2333 1988 2339 2092
rect 2061 1788 2067 1792
rect 2045 1768 2051 1772
rect 2029 1708 2035 1732
rect 2125 1728 2131 1832
rect 2173 1763 2179 1852
rect 2168 1757 2179 1763
rect 2189 1708 2195 1832
rect 2237 1748 2243 1872
rect 1997 1628 2003 1692
rect 2029 1688 2035 1692
rect 2237 1668 2243 1732
rect 2253 1728 2259 1876
rect 2285 1748 2291 1832
rect 2301 1728 2307 1912
rect 2349 1908 2355 2012
rect 2365 2003 2371 2237
rect 2397 2148 2403 2152
rect 2509 2148 2515 2152
rect 2541 2148 2547 2263
rect 2861 2148 2867 2263
rect 2909 2228 2915 2263
rect 2413 2108 2419 2112
rect 2541 2108 2547 2132
rect 2589 2128 2595 2132
rect 2685 2128 2691 2132
rect 2669 2108 2675 2112
rect 2381 2028 2387 2032
rect 2365 1997 2387 2003
rect 2381 1908 2387 1997
rect 2333 1768 2339 1872
rect 2349 1828 2355 1872
rect 2365 1868 2371 1872
rect 2317 1703 2323 1752
rect 2349 1748 2355 1772
rect 2381 1723 2387 1892
rect 2413 1808 2419 2032
rect 2461 1948 2467 2092
rect 2557 2088 2563 2092
rect 2749 2088 2755 2132
rect 2765 2088 2771 2112
rect 2781 2108 2787 2132
rect 2829 2128 2835 2132
rect 2493 1968 2499 2032
rect 2509 1888 2515 1912
rect 2376 1717 2387 1723
rect 2413 1708 2419 1712
rect 2429 1708 2435 1832
rect 2477 1748 2483 1812
rect 2445 1728 2451 1732
rect 2493 1708 2499 1712
rect 2312 1697 2323 1703
rect 2397 1688 2403 1692
rect 1965 1597 1987 1603
rect 1965 1508 1971 1597
rect 1981 1508 1987 1572
rect 1965 1488 1971 1492
rect 2013 1468 2019 1632
rect 2029 1508 2035 1552
rect 1933 1448 1939 1452
rect 1837 1348 1843 1352
rect 1869 1288 1875 1432
rect 1885 1348 1891 1432
rect 1997 1348 2003 1432
rect 2013 1368 2019 1452
rect 2029 1388 2035 1472
rect 2061 1408 2067 1632
rect 2093 1468 2099 1632
rect 2205 1528 2211 1532
rect 2237 1508 2243 1612
rect 2221 1468 2227 1492
rect 2093 1448 2099 1452
rect 2221 1448 2227 1452
rect 2061 1368 2067 1372
rect 1773 1268 1779 1272
rect 1789 1168 1795 1232
rect 1869 1168 1875 1232
rect 1757 1088 1763 1092
rect 1757 948 1763 1072
rect 1789 1068 1795 1112
rect 1853 1068 1859 1152
rect 1885 1148 1891 1312
rect 2013 1288 2019 1312
rect 1869 1108 1875 1112
rect 1901 1088 1907 1212
rect 1981 1088 1987 1092
rect 1917 1068 1923 1072
rect 1837 1028 1843 1032
rect 1885 1008 1891 1032
rect 1773 968 1779 992
rect 1789 988 1795 992
rect 1837 948 1843 952
rect 1725 808 1731 832
rect 1693 668 1699 792
rect 1549 508 1555 512
rect 1565 468 1571 632
rect 1613 568 1619 632
rect 1581 528 1587 532
rect 1677 528 1683 632
rect 1693 588 1699 632
rect 1709 628 1715 712
rect 1741 688 1747 812
rect 1757 708 1763 912
rect 1741 648 1747 672
rect 1757 668 1763 692
rect 1789 688 1795 712
rect 1741 588 1747 632
rect 1597 508 1603 512
rect 1629 488 1635 492
rect 1341 357 1363 363
rect 1197 128 1203 232
rect 1309 168 1315 292
rect 1325 188 1331 312
rect 1357 308 1363 357
rect 1373 328 1379 352
rect 1405 308 1411 412
rect 1437 328 1443 352
rect 1501 328 1507 352
rect 1517 288 1523 452
rect 1565 323 1571 452
rect 1560 317 1571 323
rect 1597 308 1603 432
rect 1645 328 1651 512
rect 1661 428 1667 512
rect 1805 508 1811 932
rect 1853 928 1859 932
rect 1917 928 1923 932
rect 1821 828 1827 912
rect 1885 848 1891 892
rect 1917 728 1923 832
rect 1933 703 1939 1032
rect 1965 908 1971 992
rect 1997 948 2003 1072
rect 2013 923 2019 1252
rect 2045 1168 2051 1352
rect 2093 1308 2099 1332
rect 2109 1228 2115 1312
rect 2141 1308 2147 1392
rect 2173 1388 2179 1432
rect 2237 1368 2243 1472
rect 2253 1408 2259 1512
rect 2189 1348 2195 1352
rect 2253 1348 2259 1352
rect 2269 1323 2275 1632
rect 2317 1488 2323 1572
rect 2285 1328 2291 1452
rect 2301 1368 2307 1472
rect 2365 1468 2371 1632
rect 2381 1508 2387 1572
rect 2413 1488 2419 1512
rect 2429 1488 2435 1692
rect 2509 1548 2515 1832
rect 2525 1768 2531 1872
rect 2525 1728 2531 1752
rect 2525 1708 2531 1712
rect 2573 1708 2579 1892
rect 2621 1888 2627 2032
rect 2637 1908 2643 1932
rect 2685 1888 2691 2032
rect 2733 1908 2739 2032
rect 2781 1988 2787 2052
rect 2749 1908 2755 1912
rect 2781 1908 2787 1952
rect 2813 1948 2819 2032
rect 2605 1748 2611 1752
rect 2621 1728 2627 1732
rect 2573 1508 2579 1692
rect 2413 1468 2419 1472
rect 2365 1328 2371 1432
rect 2253 1317 2275 1323
rect 2045 948 2051 1092
rect 2061 1088 2067 1212
rect 2141 1188 2147 1272
rect 2237 1248 2243 1312
rect 2125 1128 2131 1132
rect 2157 1128 2163 1212
rect 2253 1123 2259 1317
rect 2269 1288 2275 1292
rect 2301 1268 2307 1272
rect 2253 1117 2264 1123
rect 2301 1108 2307 1192
rect 2317 1128 2323 1232
rect 2173 1088 2179 1092
rect 2333 1088 2339 1292
rect 2141 968 2147 992
rect 1997 917 2019 923
rect 1933 697 1955 703
rect 1677 448 1683 492
rect 1661 388 1667 412
rect 1661 328 1667 332
rect 1677 328 1683 332
rect 1773 308 1779 492
rect 1821 488 1827 552
rect 1725 268 1731 272
rect 1533 188 1539 232
rect 1261 128 1267 132
rect 269 68 275 72
rect 669 68 675 72
rect 733 68 739 72
rect 893 68 899 72
rect 1117 68 1123 72
rect 1277 48 1283 132
rect 1325 128 1331 172
rect 1501 148 1507 172
rect 1517 148 1523 152
rect 1341 128 1347 132
rect 1325 108 1331 112
rect 1389 88 1395 132
rect 1549 108 1555 232
rect 1565 208 1571 252
rect 1581 188 1587 212
rect 1613 168 1619 172
rect 1613 148 1619 152
rect 1677 108 1683 132
rect 1693 128 1699 232
rect 1741 208 1747 252
rect 1789 208 1795 252
rect 1805 168 1811 432
rect 1837 348 1843 632
rect 1885 628 1891 676
rect 1917 608 1923 692
rect 1949 663 1955 697
rect 1965 688 1971 792
rect 1997 748 2003 917
rect 2109 908 2115 932
rect 2205 928 2211 1012
rect 2013 888 2019 892
rect 2221 868 2227 872
rect 2029 728 2035 832
rect 2013 688 2019 692
rect 1933 657 1955 663
rect 1853 568 1859 572
rect 1853 548 1859 552
rect 1869 368 1875 432
rect 1821 323 1827 332
rect 1885 328 1891 352
rect 1821 317 1843 323
rect 1837 308 1843 317
rect 1821 228 1827 292
rect 1901 288 1907 592
rect 1933 528 1939 657
rect 1949 608 1955 632
rect 1965 588 1971 672
rect 2077 668 2083 812
rect 2093 708 2099 732
rect 2173 688 2179 832
rect 2189 708 2195 732
rect 2205 688 2211 832
rect 2253 828 2259 892
rect 2221 708 2227 712
rect 2269 688 2275 952
rect 2285 928 2291 972
rect 2317 928 2323 932
rect 2301 788 2307 832
rect 2333 743 2339 1052
rect 2349 1028 2355 1312
rect 2381 1288 2387 1452
rect 2397 1348 2403 1432
rect 2397 988 2403 1312
rect 2429 1188 2435 1412
rect 2461 1348 2467 1432
rect 2525 1428 2531 1472
rect 2557 1408 2563 1432
rect 2493 1348 2499 1352
rect 2525 1328 2531 1372
rect 2557 1348 2563 1392
rect 2461 1308 2467 1312
rect 2557 1308 2563 1312
rect 2461 1288 2467 1292
rect 2413 1068 2419 1092
rect 2445 1068 2451 1092
rect 2413 968 2419 1012
rect 2509 988 2515 1032
rect 2445 944 2451 952
rect 2349 808 2355 932
rect 2365 908 2371 912
rect 2413 768 2419 812
rect 2509 808 2515 932
rect 2333 737 2355 743
rect 2301 708 2307 712
rect 2349 708 2355 737
rect 1917 448 1923 472
rect 1981 468 1987 552
rect 2045 488 2051 552
rect 2061 483 2067 632
rect 2125 608 2131 672
rect 2365 668 2371 672
rect 2189 568 2195 572
rect 2157 528 2163 532
rect 2189 528 2195 552
rect 2205 548 2211 632
rect 2221 528 2227 632
rect 2253 608 2259 632
rect 2269 588 2275 632
rect 2365 608 2371 632
rect 2061 477 2083 483
rect 1837 268 1843 272
rect 1917 228 1923 232
rect 1821 208 1827 212
rect 1933 203 1939 432
rect 1949 328 1955 352
rect 1981 288 1987 452
rect 2013 268 2019 292
rect 1933 197 1955 203
rect 1773 148 1779 152
rect 1741 128 1747 132
rect 1805 128 1811 132
rect 1821 108 1827 172
rect 1869 148 1875 172
rect 1885 148 1891 152
rect 1933 148 1939 172
rect 1949 128 1955 197
rect 1565 68 1571 92
rect 1901 28 1907 112
rect 1965 28 1971 232
rect 2029 168 2035 352
rect 2061 328 2067 452
rect 2061 268 2067 312
rect 2077 308 2083 477
rect 2109 328 2115 472
rect 2125 428 2131 492
rect 2237 448 2243 492
rect 2253 468 2259 552
rect 2285 508 2291 592
rect 2141 288 2147 412
rect 2173 348 2179 372
rect 2317 328 2323 472
rect 2333 368 2339 432
rect 2237 248 2243 292
rect 2045 188 2051 232
rect 2029 128 2035 152
rect 2125 148 2131 152
rect 2157 123 2163 232
rect 2253 188 2259 272
rect 2333 268 2339 272
rect 2301 188 2307 232
rect 2152 117 2163 123
rect 2173 108 2179 172
rect 2285 157 2296 163
rect 2252 150 2260 152
rect 2285 108 2291 157
rect 2317 143 2323 192
rect 2349 168 2355 292
rect 2312 137 2323 143
rect 2365 68 2371 512
rect 2381 468 2387 712
rect 2397 688 2403 732
rect 2413 708 2419 752
rect 2429 688 2435 772
rect 2525 728 2531 1072
rect 2541 968 2547 972
rect 2557 908 2563 1132
rect 2573 1108 2579 1492
rect 2589 1388 2595 1712
rect 2669 1703 2675 1832
rect 2685 1768 2691 1872
rect 2701 1848 2707 1892
rect 2733 1748 2739 1832
rect 2797 1788 2803 1872
rect 2829 1768 2835 1852
rect 2733 1728 2739 1732
rect 2845 1728 2851 2032
rect 2877 1908 2883 2212
rect 3037 2168 3043 2263
rect 3085 2188 3091 2263
rect 3053 2157 3064 2163
rect 2909 2128 2915 2132
rect 2925 2088 2931 2132
rect 2973 2088 2979 2112
rect 2989 2088 2995 2132
rect 3037 2128 3043 2152
rect 3053 2128 3059 2157
rect 2973 2028 2979 2032
rect 2861 1868 2867 1892
rect 2877 1788 2883 1852
rect 2909 1728 2915 2012
rect 2989 1908 2995 1912
rect 3005 1908 3011 1912
rect 3037 1908 3043 1912
rect 2909 1708 2915 1712
rect 2669 1697 2680 1703
rect 2797 1688 2803 1692
rect 2669 1568 2675 1632
rect 2605 1428 2611 1472
rect 2589 1308 2595 1332
rect 2589 1068 2595 1272
rect 2605 1128 2611 1332
rect 2605 928 2611 1032
rect 2621 948 2627 1532
rect 2637 1528 2643 1532
rect 2637 1117 2648 1123
rect 2637 1108 2643 1117
rect 2637 1008 2643 1072
rect 2669 968 2675 1432
rect 2701 1163 2707 1552
rect 2749 1468 2755 1632
rect 2797 1548 2803 1572
rect 2781 1468 2787 1472
rect 2733 1368 2739 1432
rect 2781 1388 2787 1452
rect 2797 1328 2803 1512
rect 2813 1508 2819 1632
rect 2925 1588 2931 1892
rect 2941 1868 2947 1872
rect 2957 1848 2963 1892
rect 3053 1888 3059 1952
rect 2957 1748 2963 1832
rect 2957 1728 2963 1732
rect 2877 1528 2883 1532
rect 2957 1528 2963 1712
rect 2989 1708 2995 1712
rect 2989 1568 2995 1632
rect 2909 1508 2915 1512
rect 2717 1248 2723 1292
rect 2685 1157 2707 1163
rect 2685 1128 2691 1157
rect 2717 1143 2723 1232
rect 2749 1148 2755 1232
rect 2701 1137 2723 1143
rect 2701 1088 2707 1137
rect 2797 1128 2803 1312
rect 2717 1108 2723 1112
rect 2701 988 2707 1052
rect 2717 968 2723 1092
rect 2765 1088 2771 1092
rect 2797 1068 2803 1112
rect 2813 1048 2819 1072
rect 2749 963 2755 1032
rect 2749 957 2771 963
rect 2765 923 2771 957
rect 2781 943 2787 1032
rect 2781 937 2792 943
rect 2829 928 2835 932
rect 2765 917 2776 923
rect 2589 708 2595 712
rect 2525 688 2531 692
rect 2605 688 2611 852
rect 2621 848 2627 912
rect 2813 908 2819 912
rect 2733 897 2744 903
rect 2669 728 2675 832
rect 2733 788 2739 897
rect 2845 903 2851 1312
rect 2861 1128 2867 1472
rect 2877 1428 2883 1432
rect 2877 1348 2883 1412
rect 2973 1348 2979 1492
rect 3005 1488 3011 1852
rect 3037 1708 3043 1712
rect 3053 1608 3059 1872
rect 3069 1848 3075 1912
rect 3117 1868 3123 1872
rect 3085 1748 3091 1852
rect 3101 1748 3107 1752
rect 3133 1743 3139 1832
rect 3149 1768 3155 2032
rect 3165 1908 3171 1912
rect 3181 1888 3187 1952
rect 3133 1737 3155 1743
rect 3117 1488 3123 1712
rect 3021 1448 3027 1472
rect 2909 1088 2915 1132
rect 2941 1123 2947 1232
rect 2925 1117 2947 1123
rect 2925 1108 2931 1117
rect 2829 897 2851 903
rect 2733 768 2739 772
rect 2829 708 2835 897
rect 2893 903 2899 1032
rect 2909 928 2915 1072
rect 2925 948 2931 1092
rect 2941 1088 2947 1092
rect 3037 1088 3043 1232
rect 3053 1088 3059 1092
rect 3085 1083 3091 1432
rect 3133 1408 3139 1492
rect 3149 1356 3155 1737
rect 3181 1283 3187 1712
rect 3165 1277 3187 1283
rect 3117 1088 3123 1112
rect 3149 1088 3155 1232
rect 3165 1188 3171 1277
rect 3080 1077 3091 1083
rect 2973 1068 2979 1072
rect 2941 908 2947 932
rect 2957 928 2963 952
rect 2888 897 2899 903
rect 2861 748 2867 832
rect 2909 728 2915 832
rect 2973 788 2979 1052
rect 3005 948 3011 952
rect 3005 908 3011 912
rect 2765 688 2771 692
rect 2781 688 2787 692
rect 2909 688 2915 692
rect 2557 648 2563 672
rect 2541 548 2547 632
rect 2557 548 2563 632
rect 2669 588 2675 632
rect 2717 548 2723 672
rect 2733 548 2739 612
rect 2861 548 2867 632
rect 2877 548 2883 572
rect 2909 548 2915 672
rect 2493 508 2499 512
rect 2541 508 2547 512
rect 2477 468 2483 492
rect 2381 328 2387 452
rect 2397 288 2403 392
rect 2413 388 2419 412
rect 2472 317 2483 323
rect 2477 283 2483 317
rect 2493 308 2499 312
rect 2557 288 2563 532
rect 2573 308 2579 512
rect 2589 508 2595 532
rect 2621 528 2627 532
rect 2605 488 2611 512
rect 2653 488 2659 492
rect 2477 277 2488 283
rect 2493 168 2499 172
rect 2573 148 2579 292
rect 2589 268 2595 272
rect 2605 188 2611 392
rect 2717 288 2723 532
rect 2925 508 2931 532
rect 2877 488 2883 492
rect 2765 308 2771 312
rect 2877 308 2883 352
rect 2749 288 2755 292
rect 2893 288 2899 292
rect 2925 288 2931 352
rect 2973 308 2979 712
rect 3005 688 3011 732
rect 3021 708 3027 1032
rect 3069 948 3075 1012
rect 3085 968 3091 1032
rect 3101 948 3107 1072
rect 3101 928 3107 932
rect 3197 928 3203 932
rect 2989 528 2995 532
rect 2989 388 2995 512
rect 3021 488 3027 652
rect 3037 528 3043 912
rect 3133 768 3139 832
rect 3133 728 3139 732
rect 3149 708 3155 732
rect 3117 548 3123 552
rect 3085 528 3091 532
rect 3133 528 3139 532
rect 3197 528 3203 532
rect 3005 323 3011 432
rect 3069 348 3075 512
rect 2989 317 3011 323
rect 2605 148 2611 172
rect 2477 128 2483 132
rect 2541 128 2547 132
rect 2621 128 2627 132
rect 2637 128 2643 232
rect 2669 128 2675 232
rect 2717 208 2723 272
rect 2733 248 2739 252
rect 2781 128 2787 132
rect 2717 108 2723 112
rect 2397 88 2403 92
rect 2429 88 2435 92
rect 2557 88 2563 92
rect 2797 88 2803 232
rect 2845 123 2851 232
rect 2941 148 2947 232
rect 2989 148 2995 317
rect 3053 288 3059 332
rect 3069 308 3075 312
rect 3117 288 3123 392
rect 3037 128 3043 232
rect 3053 128 3059 172
rect 3101 128 3107 232
rect 3149 128 3155 132
rect 3197 128 3203 132
rect 2845 117 2856 123
rect 1981 28 1987 32
rect 2109 28 2115 32
rect 1965 -43 1971 12
rect 2045 -43 2051 12
rect 2173 -43 2179 12
rect 2365 -43 2371 32
rect 2429 -43 2435 12
rect 2477 -43 2483 52
rect 2509 -43 2515 32
rect 2653 -43 2659 32
rect 2701 -43 2707 32
rect 2749 -43 2755 32
rect 2829 -43 2835 32
rect 3005 -43 3011 32
rect 3085 -43 3091 32
rect 3133 -43 3139 32
<< m3contact >>
rect 40 2152 56 2168
rect 184 2172 200 2188
rect 56 2112 72 2128
rect 24 1892 40 1908
rect 8 1552 24 1568
rect 8 1492 24 1508
rect 8 1452 24 1468
rect 8 1312 24 1328
rect 88 2092 104 2108
rect 136 2072 152 2088
rect 248 2132 264 2148
rect 360 2152 376 2168
rect 536 2152 552 2168
rect 376 2132 392 2148
rect 472 2132 488 2148
rect 696 2132 712 2148
rect 776 2152 792 2168
rect 744 2132 760 2148
rect 776 2132 792 2148
rect 168 2112 184 2128
rect 264 2112 280 2128
rect 344 2112 360 2128
rect 424 2112 440 2128
rect 568 2112 584 2128
rect 712 2112 728 2128
rect 184 2072 200 2088
rect 152 1912 168 1928
rect 184 1912 200 1928
rect 72 1872 88 1888
rect 168 1872 184 1888
rect 152 1852 168 1868
rect 232 1832 248 1848
rect 216 1792 232 1808
rect 216 1772 232 1788
rect 88 1732 104 1748
rect 184 1732 200 1748
rect 72 1712 88 1728
rect 152 1712 168 1728
rect 232 1712 248 1728
rect 136 1692 152 1708
rect 88 1672 104 1688
rect 168 1672 184 1688
rect 168 1652 184 1668
rect 88 1572 104 1588
rect 136 1532 152 1548
rect 72 1492 88 1508
rect 40 1472 56 1488
rect 72 1372 88 1388
rect 200 1472 216 1488
rect 264 1892 280 1908
rect 328 2092 344 2108
rect 392 2052 408 2068
rect 600 2072 616 2088
rect 760 2092 776 2108
rect 664 2052 680 2068
rect 728 2052 744 2068
rect 520 2032 536 2048
rect 568 2032 584 2048
rect 408 1972 424 1988
rect 552 1952 568 1968
rect 504 1932 520 1948
rect 728 2012 744 2028
rect 776 2012 792 2028
rect 696 1912 708 1928
rect 708 1912 712 1928
rect 328 1892 344 1908
rect 472 1892 488 1908
rect 520 1892 536 1908
rect 648 1892 664 1908
rect 680 1892 696 1908
rect 264 1872 296 1888
rect 344 1872 360 1888
rect 376 1832 392 1848
rect 264 1752 280 1768
rect 344 1752 360 1768
rect 312 1732 328 1748
rect 280 1712 296 1728
rect 328 1712 344 1728
rect 360 1712 376 1728
rect 248 1692 264 1708
rect 376 1532 392 1548
rect 504 1872 520 1888
rect 424 1832 440 1848
rect 616 1832 632 1848
rect 440 1752 456 1768
rect 424 1732 440 1748
rect 664 1872 680 1888
rect 1096 2212 1112 2228
rect 888 2152 904 2168
rect 1000 2152 1016 2168
rect 1144 2152 1160 2168
rect 1176 2152 1192 2168
rect 1080 2132 1096 2148
rect 1192 2132 1208 2148
rect 808 2112 824 2128
rect 920 2112 936 2128
rect 872 2052 888 2068
rect 856 2032 872 2048
rect 936 2092 952 2108
rect 920 2012 936 2028
rect 952 1992 968 2008
rect 952 1972 968 1988
rect 792 1952 824 1968
rect 872 1912 888 1928
rect 840 1892 856 1908
rect 760 1872 776 1888
rect 728 1852 744 1868
rect 888 1852 904 1868
rect 664 1812 680 1828
rect 648 1752 664 1768
rect 696 1752 712 1768
rect 808 1752 824 1768
rect 408 1712 424 1728
rect 472 1712 488 1728
rect 600 1712 616 1728
rect 408 1672 424 1688
rect 536 1692 552 1708
rect 440 1552 456 1568
rect 504 1552 520 1568
rect 392 1512 408 1528
rect 488 1512 504 1528
rect 296 1492 312 1508
rect 360 1492 376 1508
rect 280 1472 296 1488
rect 136 1392 152 1408
rect 72 1352 88 1368
rect 120 1352 136 1368
rect 136 1332 152 1348
rect 40 1312 56 1328
rect 88 1312 104 1328
rect 8 1032 24 1048
rect 56 1292 72 1308
rect 56 1132 72 1148
rect 88 1112 104 1128
rect 56 1072 72 1088
rect 72 1032 88 1048
rect 56 972 72 988
rect 8 952 24 968
rect 40 952 56 968
rect 24 932 40 948
rect 40 912 56 928
rect 24 892 40 908
rect 8 772 24 788
rect 8 692 24 708
rect 120 1192 136 1208
rect 104 972 120 988
rect 88 952 120 968
rect 88 852 104 868
rect 72 672 88 688
rect 88 592 104 608
rect 8 312 24 328
rect 56 312 72 328
rect 136 1132 152 1148
rect 136 1072 152 1088
rect 120 892 136 908
rect 216 1452 232 1468
rect 216 1392 232 1408
rect 168 1332 184 1348
rect 184 1332 200 1348
rect 264 1372 280 1388
rect 168 1312 184 1328
rect 328 1432 344 1448
rect 328 1372 344 1388
rect 424 1472 440 1488
rect 408 1332 424 1348
rect 504 1492 520 1508
rect 584 1652 600 1668
rect 552 1632 568 1648
rect 632 1632 648 1648
rect 744 1732 760 1748
rect 792 1732 808 1748
rect 872 1732 888 1748
rect 696 1692 712 1708
rect 600 1612 616 1628
rect 648 1612 664 1628
rect 760 1712 776 1728
rect 808 1712 824 1728
rect 856 1712 872 1728
rect 808 1652 824 1668
rect 840 1632 856 1648
rect 712 1572 744 1588
rect 680 1532 696 1548
rect 760 1552 776 1568
rect 776 1532 792 1548
rect 552 1492 568 1508
rect 664 1492 680 1508
rect 744 1492 760 1508
rect 536 1472 552 1488
rect 520 1452 536 1468
rect 536 1372 552 1388
rect 616 1472 632 1488
rect 568 1432 584 1448
rect 568 1412 584 1428
rect 600 1352 616 1368
rect 648 1452 664 1468
rect 296 1312 312 1328
rect 392 1312 408 1328
rect 456 1312 472 1328
rect 600 1312 616 1328
rect 280 1192 296 1208
rect 248 1152 264 1168
rect 568 1292 584 1308
rect 408 1172 424 1188
rect 408 1152 424 1168
rect 344 1132 360 1148
rect 248 1112 264 1128
rect 200 1092 216 1108
rect 440 1132 456 1148
rect 232 1092 248 1108
rect 248 1092 264 1108
rect 264 1092 280 1108
rect 312 1092 328 1108
rect 168 952 184 968
rect 200 952 216 968
rect 184 932 200 948
rect 152 852 168 868
rect 152 792 168 808
rect 136 752 152 768
rect 136 672 152 688
rect 120 652 136 668
rect 280 1072 296 1088
rect 248 932 264 948
rect 472 1072 488 1088
rect 312 1032 328 1048
rect 344 1012 360 1028
rect 536 1152 552 1168
rect 600 1112 616 1128
rect 680 1432 696 1448
rect 1064 2092 1080 2108
rect 1304 2152 1320 2168
rect 1352 2134 1368 2148
rect 1352 2132 1368 2134
rect 1256 2112 1272 2128
rect 1288 2112 1320 2128
rect 1352 2112 1368 2128
rect 1224 2092 1240 2108
rect 1080 2052 1096 2068
rect 1016 2032 1032 2048
rect 1016 1992 1032 2008
rect 1037 2002 1073 2018
rect 984 1952 1000 1968
rect 1160 1952 1176 1968
rect 1080 1912 1096 1928
rect 1128 1912 1144 1928
rect 968 1892 984 1908
rect 920 1872 936 1888
rect 1016 1872 1032 1888
rect 1032 1872 1048 1888
rect 904 1832 936 1848
rect 1000 1792 1016 1808
rect 952 1752 968 1768
rect 984 1752 1000 1768
rect 904 1732 920 1748
rect 904 1692 920 1708
rect 888 1632 920 1648
rect 936 1632 952 1648
rect 872 1512 888 1528
rect 856 1472 872 1488
rect 824 1392 840 1408
rect 856 1392 872 1408
rect 744 1372 760 1388
rect 728 1352 744 1368
rect 664 1332 680 1348
rect 856 1372 872 1388
rect 968 1732 984 1748
rect 984 1652 1000 1668
rect 984 1492 1000 1508
rect 1176 1932 1192 1948
rect 1112 1832 1128 1848
rect 1096 1812 1112 1828
rect 1144 1792 1160 1808
rect 1032 1752 1048 1768
rect 1016 1732 1032 1748
rect 1112 1732 1128 1748
rect 1176 1732 1192 1748
rect 1112 1712 1128 1728
rect 1160 1712 1176 1728
rect 1016 1692 1032 1708
rect 1144 1692 1160 1708
rect 1037 1602 1073 1618
rect 1064 1532 1080 1548
rect 1016 1512 1032 1528
rect 968 1472 984 1488
rect 680 1312 696 1328
rect 776 1312 792 1328
rect 664 1232 680 1248
rect 1080 1492 1096 1508
rect 1112 1492 1128 1508
rect 1096 1472 1112 1488
rect 1096 1452 1112 1468
rect 1032 1392 1048 1408
rect 1016 1332 1032 1348
rect 1176 1492 1192 1508
rect 1208 2072 1224 2088
rect 1224 1972 1240 1988
rect 1384 2112 1400 2128
rect 1432 2112 1448 2128
rect 1368 2072 1384 2088
rect 1256 1952 1272 1968
rect 1304 1952 1320 1968
rect 1240 1892 1256 1908
rect 1240 1872 1256 1888
rect 1224 1832 1240 1848
rect 1208 1752 1224 1768
rect 1288 1912 1304 1928
rect 1336 1912 1368 1928
rect 1384 1912 1400 1928
rect 1416 1912 1432 1928
rect 1480 1912 1496 1928
rect 1288 1892 1304 1908
rect 1448 1892 1464 1908
rect 1400 1872 1416 1888
rect 1272 1832 1288 1848
rect 1368 1832 1384 1848
rect 1272 1812 1288 1828
rect 1352 1752 1368 1768
rect 1640 2132 1656 2148
rect 1960 2192 1976 2208
rect 1992 2192 2008 2208
rect 2077 2202 2113 2218
rect 1528 2112 1544 2128
rect 1592 2112 1608 2128
rect 1672 2112 1688 2128
rect 1688 2112 1704 2128
rect 1864 2112 1880 2128
rect 1912 2112 1928 2128
rect 1512 1892 1528 1908
rect 1496 1852 1512 1868
rect 1512 1832 1528 1848
rect 1464 1792 1480 1808
rect 1496 1792 1512 1808
rect 1432 1732 1448 1748
rect 1240 1712 1256 1728
rect 1304 1712 1320 1728
rect 1336 1712 1352 1728
rect 1368 1712 1384 1728
rect 1496 1712 1512 1728
rect 1272 1692 1288 1708
rect 1208 1672 1224 1688
rect 1304 1672 1320 1688
rect 1336 1612 1352 1628
rect 1496 1692 1512 1708
rect 1448 1672 1464 1688
rect 1384 1572 1400 1588
rect 1480 1572 1496 1588
rect 1272 1552 1288 1568
rect 1384 1552 1400 1568
rect 1208 1532 1224 1548
rect 1144 1452 1160 1468
rect 1160 1392 1176 1408
rect 1128 1372 1144 1388
rect 1192 1472 1208 1488
rect 1192 1392 1208 1408
rect 1192 1372 1208 1388
rect 1176 1352 1192 1368
rect 1256 1492 1272 1508
rect 1320 1492 1336 1508
rect 1368 1472 1384 1488
rect 1240 1352 1256 1368
rect 1192 1332 1208 1348
rect 1224 1332 1240 1348
rect 952 1312 968 1328
rect 1016 1312 1032 1328
rect 1096 1312 1112 1328
rect 968 1292 984 1308
rect 1144 1292 1160 1308
rect 888 1272 904 1288
rect 760 1172 776 1188
rect 696 1152 712 1168
rect 648 1112 664 1128
rect 584 1092 600 1108
rect 616 1092 632 1108
rect 520 1072 536 1088
rect 504 1052 520 1068
rect 488 1012 520 1028
rect 472 992 488 1008
rect 376 972 392 988
rect 408 952 424 968
rect 440 952 456 968
rect 488 952 504 968
rect 312 932 328 948
rect 360 932 376 948
rect 376 932 392 948
rect 424 932 440 948
rect 216 912 232 928
rect 296 912 312 928
rect 312 892 328 908
rect 280 732 312 748
rect 264 712 280 728
rect 344 792 360 808
rect 232 692 248 708
rect 200 672 216 688
rect 280 652 296 668
rect 136 552 152 568
rect 184 552 200 568
rect 120 532 136 548
rect 184 512 200 528
rect 232 512 248 528
rect 88 292 104 308
rect 56 286 72 288
rect 56 272 72 286
rect 72 252 88 268
rect 8 232 24 248
rect 56 232 72 248
rect 88 212 104 228
rect 104 132 120 148
rect 184 372 200 388
rect 152 292 184 308
rect 248 472 264 488
rect 216 312 232 328
rect 200 292 216 308
rect 264 412 280 428
rect 248 312 264 328
rect 312 692 328 708
rect 472 932 488 948
rect 408 912 424 928
rect 472 912 488 928
rect 488 892 504 908
rect 408 752 424 768
rect 472 752 488 768
rect 392 732 408 748
rect 424 712 440 728
rect 520 952 536 968
rect 840 1152 856 1168
rect 808 1112 824 1128
rect 696 1092 728 1108
rect 792 1092 808 1108
rect 936 1252 952 1268
rect 888 1172 904 1188
rect 1176 1232 1192 1248
rect 1037 1202 1073 1218
rect 1144 1172 1160 1188
rect 1112 1112 1128 1128
rect 952 1092 968 1108
rect 792 1072 808 1088
rect 904 1072 920 1088
rect 648 1052 664 1068
rect 680 1052 696 1068
rect 712 1052 728 1068
rect 664 1032 680 1048
rect 616 1012 632 1028
rect 568 952 584 968
rect 584 952 600 968
rect 584 852 600 868
rect 536 772 552 788
rect 520 752 536 768
rect 504 712 520 728
rect 488 692 504 708
rect 568 712 584 728
rect 648 912 664 928
rect 856 1052 872 1068
rect 872 1052 888 1068
rect 760 1032 776 1048
rect 696 972 712 988
rect 840 992 856 1008
rect 824 972 840 988
rect 792 952 808 968
rect 872 992 888 1008
rect 904 992 920 1008
rect 936 992 952 1008
rect 920 972 936 988
rect 712 932 728 948
rect 936 952 952 968
rect 696 892 712 908
rect 600 832 616 848
rect 632 832 648 848
rect 680 812 696 828
rect 776 892 792 908
rect 808 772 824 788
rect 744 752 760 768
rect 664 732 680 748
rect 664 712 680 728
rect 568 672 584 688
rect 328 652 344 668
rect 296 492 312 508
rect 296 472 312 488
rect 312 472 328 488
rect 248 292 264 308
rect 136 252 152 268
rect 152 132 168 148
rect 248 192 264 208
rect 232 152 248 168
rect 8 112 24 128
rect 168 112 184 128
rect 200 112 216 128
rect 280 252 296 268
rect 584 652 600 668
rect 472 632 488 648
rect 568 632 584 648
rect 408 532 424 548
rect 520 612 536 628
rect 488 552 504 568
rect 664 692 680 708
rect 824 732 840 748
rect 968 992 984 1008
rect 952 912 968 928
rect 920 892 936 908
rect 856 832 872 848
rect 920 712 968 728
rect 840 692 856 708
rect 872 692 888 708
rect 1000 1072 1016 1088
rect 1032 1072 1048 1088
rect 1000 1012 1016 1028
rect 1048 972 1064 988
rect 1000 932 1016 948
rect 632 652 648 668
rect 824 652 840 668
rect 712 632 728 648
rect 824 632 840 648
rect 648 572 664 588
rect 520 532 536 548
rect 616 532 632 548
rect 392 512 408 528
rect 392 492 408 508
rect 360 472 376 488
rect 376 332 392 348
rect 312 172 328 188
rect 264 132 280 148
rect 360 312 392 328
rect 344 292 360 308
rect 344 132 360 148
rect 264 112 280 128
rect 312 112 328 128
rect 328 112 344 128
rect 488 472 504 488
rect 504 392 520 408
rect 408 332 424 348
rect 472 332 488 348
rect 504 312 520 328
rect 536 512 568 528
rect 600 512 616 528
rect 536 492 552 508
rect 568 492 584 508
rect 552 332 568 348
rect 392 292 408 308
rect 376 286 392 288
rect 376 272 392 286
rect 440 272 456 288
rect 488 272 504 288
rect 392 192 424 208
rect 648 372 664 388
rect 664 352 680 368
rect 616 332 632 348
rect 776 552 792 568
rect 792 532 808 548
rect 744 492 760 508
rect 712 392 728 408
rect 728 372 744 388
rect 712 352 728 368
rect 808 472 824 488
rect 792 452 808 468
rect 776 372 792 388
rect 792 372 808 388
rect 824 332 840 348
rect 664 292 680 308
rect 536 252 568 268
rect 440 172 456 188
rect 376 112 392 128
rect 184 92 200 108
rect 360 92 376 108
rect 392 92 408 108
rect 424 92 440 108
rect 488 152 504 168
rect 520 132 536 148
rect 456 112 472 128
rect 472 92 488 108
rect 584 132 600 148
rect 728 252 744 268
rect 744 232 760 248
rect 680 172 696 188
rect 616 112 632 128
rect 728 112 744 128
rect 824 252 840 268
rect 792 192 824 208
rect 968 652 984 668
rect 872 512 888 528
rect 920 512 936 528
rect 856 492 872 508
rect 856 472 872 488
rect 872 452 888 468
rect 888 452 904 468
rect 888 352 904 368
rect 1016 912 1032 928
rect 1128 1072 1144 1088
rect 1448 1532 1464 1548
rect 1496 1532 1512 1548
rect 1464 1512 1480 1528
rect 1480 1512 1496 1528
rect 1512 1512 1528 1528
rect 1480 1492 1496 1508
rect 1320 1452 1336 1468
rect 1432 1452 1448 1468
rect 1304 1372 1320 1388
rect 1256 1312 1272 1328
rect 1288 1272 1304 1288
rect 1240 1132 1256 1148
rect 1192 1092 1208 1108
rect 1208 1092 1224 1108
rect 1144 1052 1160 1068
rect 1176 1052 1192 1068
rect 1096 972 1112 988
rect 1112 952 1128 968
rect 1176 952 1192 968
rect 1224 972 1240 988
rect 1160 912 1176 928
rect 1064 892 1080 908
rect 1048 852 1064 868
rect 1096 852 1112 868
rect 1037 802 1073 818
rect 1032 752 1048 768
rect 1064 732 1080 748
rect 1032 712 1048 728
rect 1048 612 1064 628
rect 1032 572 1048 588
rect 1128 832 1144 848
rect 1016 512 1032 528
rect 1096 492 1112 508
rect 1000 452 1016 468
rect 1037 402 1073 418
rect 920 332 952 348
rect 1112 332 1128 348
rect 984 292 1000 308
rect 856 272 872 288
rect 968 272 984 288
rect 840 152 856 168
rect 1000 252 1016 268
rect 920 232 936 248
rect 968 232 984 248
rect 904 212 920 228
rect 872 172 888 188
rect 776 112 792 128
rect 856 112 872 128
rect 664 92 680 108
rect 888 112 904 128
rect 936 112 952 128
rect 1144 612 1160 628
rect 1256 1092 1272 1108
rect 1320 1212 1336 1228
rect 1304 1172 1320 1188
rect 1288 1112 1304 1128
rect 1416 1392 1432 1408
rect 1368 1352 1384 1368
rect 1352 1312 1368 1328
rect 1336 1172 1352 1188
rect 1400 1332 1416 1348
rect 1544 1712 1560 1728
rect 1656 2092 1672 2108
rect 1720 2092 1736 2108
rect 1624 2072 1640 2088
rect 1704 2072 1720 2088
rect 1608 1932 1624 1948
rect 1656 1972 1672 1988
rect 1640 1912 1656 1928
rect 1592 1892 1608 1908
rect 1704 1912 1720 1928
rect 1768 1912 1784 1928
rect 1896 2092 1912 2108
rect 1848 2072 1864 2088
rect 1832 1912 1848 1928
rect 1592 1872 1608 1888
rect 1688 1872 1704 1888
rect 1592 1852 1608 1868
rect 1656 1852 1672 1868
rect 1704 1852 1720 1868
rect 1624 1812 1640 1828
rect 1560 1692 1576 1708
rect 1640 1692 1656 1708
rect 1560 1672 1576 1688
rect 1544 1592 1560 1608
rect 1528 1472 1544 1488
rect 1480 1352 1496 1368
rect 1512 1332 1528 1348
rect 1592 1552 1608 1568
rect 1576 1392 1592 1408
rect 1560 1352 1576 1368
rect 1464 1312 1480 1328
rect 1544 1312 1560 1328
rect 1368 1152 1384 1168
rect 1256 1052 1272 1068
rect 1224 892 1240 908
rect 1256 872 1272 888
rect 1208 812 1224 828
rect 1336 1072 1352 1088
rect 1368 992 1384 1008
rect 1288 952 1304 968
rect 1368 952 1384 968
rect 1224 732 1240 748
rect 1272 732 1288 748
rect 1192 712 1208 728
rect 1240 692 1256 708
rect 1176 672 1192 688
rect 1192 672 1208 688
rect 1256 592 1272 608
rect 1304 912 1320 928
rect 1464 1212 1480 1228
rect 1464 1192 1480 1208
rect 1416 1132 1432 1148
rect 1400 1032 1416 1048
rect 1448 1112 1464 1128
rect 1480 1132 1512 1148
rect 1480 1092 1496 1108
rect 1448 1052 1464 1068
rect 1432 1032 1448 1048
rect 1384 892 1400 908
rect 1432 912 1464 928
rect 1416 892 1432 908
rect 1464 892 1480 908
rect 1336 872 1352 888
rect 1400 872 1416 888
rect 1416 852 1432 868
rect 1304 772 1320 788
rect 1352 732 1368 748
rect 1448 772 1464 788
rect 1400 692 1416 708
rect 1304 672 1320 688
rect 1336 672 1352 688
rect 1352 632 1368 648
rect 1368 612 1384 628
rect 1320 592 1336 608
rect 1272 572 1288 588
rect 1240 532 1256 548
rect 1384 592 1400 608
rect 1400 552 1416 568
rect 1176 512 1192 528
rect 1224 512 1240 528
rect 1272 512 1288 528
rect 1352 492 1368 508
rect 1400 492 1416 508
rect 1192 472 1208 488
rect 1192 452 1208 468
rect 1224 432 1240 448
rect 1336 412 1352 428
rect 1320 372 1336 388
rect 1128 292 1144 308
rect 1080 252 1096 268
rect 1016 172 1032 188
rect 1096 172 1112 188
rect 1032 152 1048 168
rect 984 132 1000 148
rect 1064 132 1080 148
rect 984 112 1000 128
rect 888 92 904 108
rect 1112 132 1128 148
rect 1112 112 1128 128
rect 1144 272 1160 288
rect 1144 212 1160 228
rect 1208 292 1224 308
rect 1400 472 1416 488
rect 1432 592 1448 608
rect 1480 792 1496 808
rect 1480 592 1496 608
rect 1480 572 1512 588
rect 1608 1392 1624 1408
rect 1608 1332 1624 1348
rect 1640 1492 1656 1508
rect 1688 1832 1704 1848
rect 1672 1812 1688 1828
rect 1800 1892 1816 1908
rect 1864 1892 1880 1908
rect 1768 1872 1784 1888
rect 1816 1852 1832 1868
rect 1800 1832 1816 1848
rect 1752 1792 1768 1808
rect 1672 1772 1688 1788
rect 1720 1752 1736 1768
rect 1768 1732 1784 1748
rect 1688 1672 1704 1688
rect 1816 1772 1832 1788
rect 1784 1712 1800 1728
rect 1832 1752 1848 1768
rect 1896 1752 1912 1768
rect 1864 1732 1880 1748
rect 1832 1712 1848 1728
rect 1928 2072 1960 2088
rect 1976 2072 1992 2088
rect 1960 1952 1976 1968
rect 2024 2152 2040 2168
rect 2104 2152 2120 2168
rect 2040 2132 2056 2148
rect 2104 2132 2120 2148
rect 2056 2112 2072 2128
rect 2184 2092 2200 2108
rect 2168 2052 2184 2068
rect 2040 1912 2056 1928
rect 2152 1932 2168 1948
rect 2216 1932 2232 1948
rect 2136 1912 2152 1928
rect 1960 1892 1976 1908
rect 1992 1892 2008 1908
rect 2056 1892 2072 1908
rect 1944 1852 1960 1868
rect 1944 1832 1960 1848
rect 2008 1872 2024 1888
rect 1960 1772 1976 1788
rect 1928 1732 1944 1748
rect 1928 1692 1944 1708
rect 1960 1692 1976 1708
rect 1752 1632 1768 1648
rect 1816 1632 1832 1648
rect 1880 1632 1896 1648
rect 1912 1632 1928 1648
rect 1672 1612 1688 1628
rect 1688 1512 1704 1528
rect 1656 1412 1672 1428
rect 1624 1312 1640 1328
rect 1560 1292 1576 1308
rect 1528 1252 1544 1268
rect 1624 1252 1640 1268
rect 1528 1212 1544 1228
rect 1624 1212 1640 1228
rect 1624 1192 1640 1208
rect 1576 1152 1592 1168
rect 1608 1152 1624 1168
rect 1528 1092 1544 1108
rect 1544 1072 1560 1088
rect 1560 1012 1576 1028
rect 1544 992 1560 1008
rect 1672 1172 1688 1188
rect 1656 1092 1672 1108
rect 1608 1072 1624 1088
rect 1592 1052 1608 1068
rect 1768 1612 1784 1628
rect 1768 1552 1784 1568
rect 1736 1512 1752 1528
rect 1784 1492 1800 1508
rect 1752 1472 1768 1488
rect 1800 1472 1816 1488
rect 1720 1412 1736 1428
rect 1736 1372 1752 1388
rect 1704 1352 1720 1368
rect 1704 1332 1720 1348
rect 1720 1292 1736 1308
rect 1736 1252 1752 1268
rect 1704 1092 1720 1108
rect 1656 972 1672 988
rect 1656 952 1672 968
rect 1640 932 1656 948
rect 1624 912 1656 928
rect 1576 872 1592 888
rect 1592 772 1608 788
rect 1528 752 1544 768
rect 1592 752 1608 768
rect 1560 732 1576 748
rect 1640 712 1656 728
rect 1528 692 1544 708
rect 1624 692 1640 708
rect 1608 672 1624 688
rect 1704 1012 1720 1028
rect 1704 952 1720 968
rect 1688 932 1704 948
rect 1720 892 1736 908
rect 1784 1392 1800 1408
rect 2232 1892 2248 1908
rect 2264 2172 2280 2188
rect 2296 2172 2312 2188
rect 2328 2172 2344 2188
rect 2296 2132 2312 2148
rect 2280 2112 2296 2128
rect 2344 2112 2360 2128
rect 2344 2012 2360 2028
rect 2200 1872 2216 1888
rect 2104 1852 2136 1868
rect 2168 1852 2184 1868
rect 2120 1832 2136 1848
rect 2056 1792 2072 1808
rect 2077 1802 2113 1818
rect 2040 1772 2072 1788
rect 2168 1732 2184 1748
rect 2152 1712 2168 1728
rect 2024 1692 2040 1708
rect 2184 1692 2200 1708
rect 2024 1672 2040 1688
rect 2280 1732 2296 1748
rect 2392 2152 2408 2168
rect 2504 2152 2520 2168
rect 2552 2152 2568 2168
rect 2872 2212 2888 2228
rect 2904 2212 2920 2228
rect 2520 2132 2536 2148
rect 2680 2132 2696 2148
rect 2744 2132 2760 2148
rect 2776 2132 2792 2148
rect 2824 2132 2840 2148
rect 2856 2132 2872 2148
rect 2584 2112 2600 2128
rect 2616 2112 2632 2128
rect 2664 2112 2680 2128
rect 2408 2092 2424 2108
rect 2536 2092 2552 2108
rect 2600 2092 2616 2108
rect 2376 2012 2392 2028
rect 2328 1872 2344 1888
rect 2312 1772 2328 1788
rect 2360 1852 2376 1868
rect 2344 1812 2360 1828
rect 2344 1772 2360 1788
rect 2312 1752 2328 1768
rect 2296 1712 2312 1728
rect 2760 2112 2776 2128
rect 2808 2092 2824 2108
rect 2552 2072 2568 2088
rect 2632 2072 2648 2088
rect 2696 2072 2712 2088
rect 2776 2052 2792 2068
rect 2488 1952 2504 1968
rect 2456 1932 2472 1948
rect 2504 1912 2520 1928
rect 2472 1892 2488 1908
rect 2568 1892 2584 1908
rect 2600 1892 2616 1908
rect 2488 1852 2504 1868
rect 2408 1792 2424 1808
rect 2408 1752 2424 1768
rect 2408 1712 2424 1728
rect 2472 1812 2488 1828
rect 2440 1732 2456 1748
rect 2472 1732 2488 1748
rect 2424 1692 2440 1708
rect 2488 1692 2504 1708
rect 2392 1672 2408 1688
rect 2232 1652 2248 1668
rect 2008 1632 2024 1648
rect 1992 1612 2008 1628
rect 1896 1552 1912 1568
rect 1976 1572 1992 1588
rect 1944 1492 1960 1508
rect 1912 1472 1928 1488
rect 1960 1472 1976 1488
rect 2024 1552 2040 1568
rect 1880 1432 1896 1448
rect 1928 1432 1944 1448
rect 1832 1352 1848 1368
rect 1784 1312 1800 1328
rect 1800 1292 1816 1308
rect 2232 1612 2248 1628
rect 2200 1532 2216 1548
rect 2152 1512 2168 1528
rect 2184 1512 2200 1528
rect 2248 1512 2264 1528
rect 2104 1472 2120 1488
rect 2216 1452 2232 1468
rect 2088 1432 2104 1448
rect 2216 1432 2232 1448
rect 2056 1392 2072 1408
rect 2077 1402 2113 1418
rect 2136 1392 2152 1408
rect 2056 1372 2072 1388
rect 2008 1352 2024 1368
rect 1880 1332 1896 1348
rect 1944 1332 1960 1348
rect 1992 1332 2008 1348
rect 1880 1312 1896 1328
rect 1960 1312 1976 1328
rect 1992 1312 2008 1328
rect 1864 1272 1880 1288
rect 1768 1252 1784 1268
rect 1752 1172 1768 1188
rect 1784 1152 1800 1168
rect 1848 1152 1880 1168
rect 1752 1092 1768 1108
rect 1800 1072 1816 1088
rect 1896 1292 1912 1308
rect 1928 1292 1944 1308
rect 2008 1272 2024 1288
rect 2008 1252 2024 1268
rect 1896 1212 1912 1228
rect 1880 1132 1896 1148
rect 1864 1092 1880 1108
rect 1976 1092 1992 1108
rect 1912 1072 1944 1088
rect 1992 1072 2008 1088
rect 1784 1052 1800 1068
rect 1832 1012 1848 1028
rect 1768 992 1800 1008
rect 1880 992 1896 1008
rect 1832 952 1848 968
rect 1752 932 1768 948
rect 1848 932 1864 948
rect 1880 932 1896 948
rect 1912 932 1928 948
rect 1752 912 1768 928
rect 1736 812 1752 828
rect 1688 792 1704 808
rect 1720 792 1736 808
rect 1720 772 1736 788
rect 1656 652 1688 668
rect 1688 632 1704 648
rect 1512 532 1528 548
rect 1496 512 1512 528
rect 1464 492 1480 508
rect 1544 492 1560 508
rect 1608 552 1624 568
rect 1784 712 1800 728
rect 1752 692 1768 708
rect 1736 632 1752 648
rect 1704 612 1720 628
rect 1576 512 1592 528
rect 1640 512 1656 528
rect 1672 512 1688 528
rect 1784 512 1800 528
rect 1592 492 1608 508
rect 1624 492 1640 508
rect 1416 452 1432 468
rect 1512 452 1528 468
rect 1560 452 1576 468
rect 1400 412 1416 428
rect 1336 332 1352 348
rect 1304 312 1320 328
rect 1320 312 1336 328
rect 1288 292 1304 308
rect 1304 292 1320 308
rect 1176 272 1192 288
rect 1240 272 1256 288
rect 1272 272 1288 288
rect 1160 172 1176 188
rect 1176 152 1192 168
rect 1368 352 1384 368
rect 1432 352 1448 368
rect 1496 352 1512 368
rect 1400 292 1416 308
rect 1464 292 1480 308
rect 1592 432 1608 448
rect 1848 892 1864 908
rect 1880 832 1896 848
rect 1816 812 1832 828
rect 1912 712 1928 728
rect 1960 992 1976 1008
rect 1992 932 2008 948
rect 2088 1292 2104 1308
rect 2168 1372 2184 1388
rect 2248 1392 2264 1408
rect 2184 1352 2200 1368
rect 2232 1352 2264 1368
rect 2200 1332 2216 1348
rect 2168 1312 2184 1328
rect 2312 1572 2328 1588
rect 2280 1492 2296 1508
rect 2328 1476 2344 1488
rect 2328 1472 2344 1476
rect 2280 1452 2296 1468
rect 2376 1572 2392 1588
rect 2408 1512 2424 1528
rect 2488 1672 2504 1688
rect 2520 1752 2536 1768
rect 2536 1732 2552 1748
rect 2520 1712 2536 1728
rect 2632 1932 2648 1948
rect 2840 2032 2856 2048
rect 2776 1952 2792 1968
rect 2808 1932 2824 1948
rect 2824 1912 2840 1928
rect 2696 1892 2712 1908
rect 2728 1892 2760 1908
rect 2616 1872 2632 1888
rect 2600 1752 2616 1768
rect 2616 1732 2632 1748
rect 2584 1712 2600 1728
rect 2568 1692 2584 1708
rect 2504 1532 2520 1548
rect 2568 1492 2584 1508
rect 2408 1472 2424 1488
rect 2360 1452 2392 1468
rect 2296 1352 2312 1368
rect 2136 1292 2152 1308
rect 2200 1292 2216 1308
rect 2136 1272 2152 1288
rect 2120 1232 2136 1248
rect 2056 1212 2072 1228
rect 2104 1212 2120 1228
rect 2040 1152 2056 1168
rect 2024 1112 2040 1128
rect 2040 1092 2056 1108
rect 2232 1232 2248 1248
rect 2152 1212 2168 1228
rect 2120 1112 2136 1128
rect 2328 1292 2344 1308
rect 2264 1272 2280 1288
rect 2296 1272 2312 1288
rect 2296 1252 2312 1268
rect 2296 1192 2312 1208
rect 2312 1112 2328 1128
rect 2136 1092 2152 1108
rect 2168 1092 2184 1108
rect 2232 1092 2248 1108
rect 2216 1072 2232 1088
rect 2077 1002 2113 1018
rect 2200 1012 2216 1028
rect 2136 992 2152 1008
rect 2152 952 2168 968
rect 1960 792 1976 808
rect 1768 492 1784 508
rect 1800 492 1816 508
rect 1672 432 1688 448
rect 1656 412 1672 428
rect 1656 372 1672 388
rect 1656 332 1688 348
rect 1640 312 1656 328
rect 1816 472 1832 488
rect 1800 432 1816 448
rect 1576 292 1592 308
rect 1624 292 1640 308
rect 1672 292 1688 308
rect 1368 272 1384 288
rect 1432 272 1448 288
rect 1608 272 1624 288
rect 1688 272 1704 288
rect 1432 252 1448 268
rect 1496 252 1512 268
rect 1720 252 1736 268
rect 1528 232 1544 248
rect 1320 172 1336 188
rect 1496 172 1512 188
rect 1304 152 1320 168
rect 1192 112 1208 128
rect 1224 112 1240 128
rect 1256 112 1272 128
rect 1224 92 1240 108
rect 216 72 232 88
rect 264 72 280 88
rect 280 72 296 88
rect 440 72 456 88
rect 536 72 552 88
rect 648 72 664 88
rect 664 72 680 88
rect 712 72 728 88
rect 728 72 744 88
rect 776 72 792 88
rect 888 72 904 88
rect 936 72 952 88
rect 1112 72 1128 88
rect 792 52 808 68
rect 1368 152 1384 168
rect 1512 152 1528 168
rect 1336 132 1352 148
rect 1400 144 1416 148
rect 1400 132 1416 144
rect 1320 112 1336 128
rect 1304 92 1320 108
rect 1448 112 1464 128
rect 1480 112 1496 128
rect 1688 232 1704 248
rect 1576 212 1592 228
rect 1560 192 1576 208
rect 1608 172 1624 188
rect 1640 152 1656 168
rect 1656 132 1672 148
rect 1736 192 1752 208
rect 1784 192 1800 208
rect 1896 672 1912 688
rect 1880 612 1896 628
rect 1928 672 1944 688
rect 2088 912 2104 928
rect 2280 972 2296 988
rect 2264 952 2280 968
rect 2248 912 2264 928
rect 2104 892 2120 908
rect 2152 892 2168 908
rect 2184 892 2200 908
rect 2008 872 2024 888
rect 2216 852 2232 868
rect 2072 812 2088 828
rect 2040 692 2056 708
rect 1960 672 1976 688
rect 2008 672 2024 688
rect 1896 592 1928 608
rect 1848 572 1864 588
rect 1880 512 1896 528
rect 1864 352 1896 368
rect 1832 332 1848 348
rect 1848 332 1864 348
rect 1944 592 1960 608
rect 2088 732 2104 748
rect 2136 712 2152 728
rect 2184 732 2200 748
rect 2248 812 2264 828
rect 2232 712 2248 728
rect 2216 692 2232 708
rect 2312 932 2328 948
rect 2312 912 2328 928
rect 2296 832 2312 848
rect 2424 1412 2440 1428
rect 2408 1332 2424 1348
rect 2376 1272 2392 1288
rect 2344 1012 2360 1028
rect 2408 1252 2424 1268
rect 2520 1412 2536 1428
rect 2552 1392 2568 1408
rect 2520 1372 2536 1388
rect 2488 1352 2504 1368
rect 2488 1332 2504 1348
rect 2536 1332 2552 1348
rect 2552 1332 2568 1348
rect 2456 1292 2472 1308
rect 2552 1292 2568 1308
rect 2456 1272 2472 1288
rect 2552 1132 2568 1148
rect 2504 1112 2520 1128
rect 2440 1092 2456 1108
rect 2472 1092 2488 1108
rect 2456 1072 2472 1088
rect 2408 1052 2424 1068
rect 2408 1012 2424 1028
rect 2472 972 2488 988
rect 2504 972 2520 988
rect 2344 952 2360 968
rect 2440 952 2456 968
rect 2424 932 2440 948
rect 2472 912 2488 928
rect 2360 892 2376 908
rect 2408 812 2424 828
rect 2344 792 2360 808
rect 2504 792 2520 808
rect 2424 772 2440 788
rect 2408 752 2424 768
rect 2296 712 2312 728
rect 2328 712 2344 728
rect 2392 732 2408 748
rect 2376 712 2392 728
rect 2120 672 2136 688
rect 2200 672 2216 688
rect 2280 672 2296 688
rect 1976 552 1992 568
rect 1944 492 1960 508
rect 2024 512 2040 528
rect 2040 472 2056 488
rect 2077 602 2113 618
rect 2360 652 2376 668
rect 2200 632 2216 648
rect 2264 632 2280 648
rect 2120 592 2136 608
rect 2168 572 2184 588
rect 2184 572 2200 588
rect 2248 592 2264 608
rect 2280 592 2296 608
rect 2360 592 2376 608
rect 2152 512 2168 528
rect 2184 512 2200 528
rect 2216 512 2232 528
rect 2216 492 2232 508
rect 1976 452 1992 468
rect 2056 452 2072 468
rect 1912 432 1928 448
rect 1832 252 1848 268
rect 1816 212 1832 228
rect 1912 212 1928 228
rect 1816 192 1832 208
rect 1944 352 1960 368
rect 1992 352 2008 368
rect 2024 352 2040 368
rect 2008 252 2024 268
rect 1944 232 1960 248
rect 1960 232 1976 248
rect 1816 172 1832 188
rect 1864 172 1880 188
rect 1704 152 1736 168
rect 1768 132 1784 148
rect 1800 132 1816 148
rect 1736 112 1752 128
rect 1768 112 1784 128
rect 1880 152 1896 168
rect 1928 132 1944 148
rect 1832 112 1848 128
rect 1944 112 1960 128
rect 1448 92 1464 108
rect 1480 92 1496 108
rect 1672 92 1688 108
rect 1352 72 1368 88
rect 1384 72 1400 88
rect 1800 72 1816 88
rect 1560 52 1576 68
rect 584 32 600 48
rect 1272 32 1288 48
rect 2056 312 2072 328
rect 2104 472 2120 488
rect 2344 532 2360 548
rect 2296 512 2312 528
rect 2360 512 2376 528
rect 2312 472 2328 488
rect 2248 452 2264 468
rect 2232 432 2248 448
rect 2120 412 2152 428
rect 2072 292 2088 308
rect 2168 372 2184 388
rect 2328 352 2344 368
rect 2200 312 2216 328
rect 2232 312 2248 328
rect 2264 312 2280 328
rect 2344 312 2360 328
rect 2184 292 2200 308
rect 2216 272 2232 288
rect 2072 252 2088 268
rect 2248 272 2264 288
rect 2280 272 2296 288
rect 2232 232 2248 248
rect 2077 202 2113 218
rect 2040 172 2056 188
rect 2120 152 2136 168
rect 1992 112 2008 128
rect 2328 252 2344 268
rect 2312 192 2328 208
rect 2168 172 2184 188
rect 2296 172 2312 188
rect 2248 152 2264 168
rect 2184 132 2200 148
rect 2344 152 2360 168
rect 2008 92 2024 108
rect 2152 92 2164 108
rect 2164 92 2168 108
rect 2280 92 2296 108
rect 2456 732 2472 748
rect 2536 972 2552 988
rect 2696 1832 2712 1848
rect 2824 1852 2840 1868
rect 2728 1732 2744 1748
rect 2760 1732 2776 1748
rect 2856 1912 2872 1928
rect 2904 2132 2936 2148
rect 2984 2132 3000 2148
rect 2888 2092 2904 2108
rect 2952 2092 2968 2108
rect 3112 2132 3128 2148
rect 3032 2112 3048 2128
rect 3112 2112 3128 2128
rect 2904 2072 2920 2088
rect 2968 2072 2984 2088
rect 2984 2072 3000 2088
rect 3016 2072 3032 2088
rect 2904 2032 2920 2048
rect 2904 2012 2920 2028
rect 2968 2012 2984 2028
rect 2888 1912 2904 1928
rect 2872 1872 2888 1888
rect 2856 1852 2888 1868
rect 3048 1952 3064 1968
rect 2920 1912 2936 1928
rect 2952 1912 2968 1928
rect 3032 1912 3048 1928
rect 2952 1892 2968 1908
rect 2984 1892 3016 1908
rect 2840 1712 2856 1728
rect 2904 1692 2920 1708
rect 2648 1672 2664 1688
rect 2696 1672 2712 1688
rect 2792 1672 2808 1688
rect 2664 1552 2680 1568
rect 2696 1552 2712 1568
rect 2616 1532 2648 1548
rect 2600 1492 2616 1508
rect 2600 1412 2616 1428
rect 2584 1372 2600 1388
rect 2584 1332 2600 1348
rect 2584 1272 2600 1288
rect 2600 1112 2616 1128
rect 2584 1052 2600 1068
rect 2648 1472 2664 1488
rect 2680 1472 2696 1488
rect 2648 1452 2664 1468
rect 2632 1332 2648 1348
rect 2632 1312 2648 1328
rect 2648 1092 2664 1108
rect 2632 992 2648 1008
rect 2680 1312 2696 1328
rect 2712 1512 2728 1528
rect 2792 1572 2808 1588
rect 2792 1532 2808 1548
rect 2792 1512 2808 1528
rect 2760 1492 2776 1508
rect 2744 1452 2760 1468
rect 2728 1432 2744 1448
rect 2744 1352 2760 1368
rect 2936 1852 2952 1868
rect 3000 1872 3016 1888
rect 3000 1852 3016 1868
rect 2952 1832 2968 1848
rect 2984 1732 3000 1748
rect 2952 1712 2968 1728
rect 2920 1572 2936 1588
rect 2872 1532 2888 1548
rect 2984 1692 3000 1708
rect 2984 1552 3000 1568
rect 2984 1532 3000 1548
rect 2904 1512 2920 1528
rect 2808 1492 2824 1508
rect 2840 1492 2856 1508
rect 2904 1492 2920 1508
rect 2952 1492 2968 1508
rect 2968 1492 2984 1508
rect 2984 1492 3000 1508
rect 2824 1472 2840 1488
rect 2888 1472 2904 1488
rect 2824 1332 2840 1348
rect 2840 1312 2856 1328
rect 2712 1292 2728 1308
rect 2744 1132 2760 1148
rect 2712 1112 2728 1128
rect 2792 1112 2808 1128
rect 2696 1072 2712 1088
rect 2696 1052 2712 1068
rect 2760 1072 2776 1088
rect 2824 1092 2840 1108
rect 2808 1032 2824 1048
rect 2712 952 2728 968
rect 2744 932 2760 948
rect 2568 912 2584 928
rect 2600 912 2616 928
rect 2728 912 2744 928
rect 2824 932 2840 948
rect 2808 912 2824 928
rect 2536 892 2552 908
rect 2600 892 2616 908
rect 2568 872 2584 888
rect 2600 852 2616 868
rect 2520 712 2536 728
rect 2584 712 2600 728
rect 2520 692 2536 708
rect 2616 832 2632 848
rect 2872 1432 2888 1448
rect 2872 1412 2888 1428
rect 3032 1712 3048 1728
rect 3080 1892 3096 1908
rect 3080 1852 3096 1868
rect 3112 1852 3128 1868
rect 3064 1832 3080 1848
rect 3096 1732 3112 1748
rect 3176 1952 3192 1968
rect 3160 1912 3176 1928
rect 3144 1752 3160 1768
rect 3064 1712 3080 1728
rect 3112 1712 3128 1728
rect 3128 1712 3144 1728
rect 3048 1592 3064 1608
rect 3016 1432 3032 1448
rect 2872 1332 2888 1348
rect 2952 1332 2968 1348
rect 3064 1332 3080 1348
rect 2904 1312 2920 1328
rect 2904 1132 2920 1148
rect 2968 1092 2984 1108
rect 2872 1072 2888 1088
rect 2888 1052 2904 1068
rect 2728 752 2744 768
rect 2664 712 2680 728
rect 2936 1072 2952 1088
rect 2968 1072 2984 1088
rect 3048 1072 3064 1088
rect 3128 1392 3144 1408
rect 3192 1552 3208 1568
rect 3112 1072 3128 1088
rect 2952 952 2968 968
rect 2936 892 2952 908
rect 2840 872 2856 888
rect 2856 732 2872 748
rect 3000 952 3016 968
rect 2984 912 3000 928
rect 3000 892 3016 908
rect 2936 772 2952 788
rect 2968 772 2984 788
rect 3000 732 3016 748
rect 2904 712 2920 728
rect 2968 712 2984 728
rect 2776 692 2792 708
rect 2824 692 2840 708
rect 2888 692 2904 708
rect 2552 672 2568 688
rect 2760 672 2776 688
rect 2904 672 2920 688
rect 2536 632 2552 648
rect 2392 572 2408 588
rect 2664 572 2680 588
rect 2728 612 2744 628
rect 2872 572 2888 588
rect 2920 552 2936 568
rect 2408 532 2424 548
rect 2520 532 2536 548
rect 2552 532 2568 548
rect 2712 532 2728 548
rect 2824 532 2840 548
rect 2856 532 2872 548
rect 2904 532 2920 548
rect 2424 512 2440 528
rect 2472 512 2488 528
rect 2504 512 2520 528
rect 2392 492 2408 508
rect 2488 492 2504 508
rect 2536 492 2552 508
rect 2376 452 2392 468
rect 2472 452 2488 468
rect 2408 412 2424 428
rect 2392 392 2408 408
rect 2376 312 2392 328
rect 2408 292 2424 308
rect 2392 272 2408 288
rect 2456 272 2472 288
rect 2504 312 2520 328
rect 2488 292 2504 308
rect 2616 512 2632 528
rect 2584 492 2600 508
rect 2648 492 2664 508
rect 2600 472 2616 488
rect 2600 392 2616 408
rect 2568 292 2584 308
rect 2552 272 2568 288
rect 2488 252 2504 268
rect 2488 172 2504 188
rect 2408 152 2424 168
rect 2584 252 2600 268
rect 2888 512 2904 528
rect 2872 492 2888 508
rect 2920 492 2936 508
rect 2872 472 2888 488
rect 2872 352 2888 368
rect 2920 352 2936 368
rect 2760 312 2776 328
rect 2744 292 2760 308
rect 2888 292 2904 308
rect 3064 1012 3080 1028
rect 3080 952 3096 968
rect 3192 1052 3208 1068
rect 3048 932 3064 948
rect 3096 932 3112 948
rect 3144 912 3160 928
rect 3192 912 3208 928
rect 3016 692 3032 708
rect 2984 652 3000 668
rect 2984 532 3000 548
rect 3128 752 3144 768
rect 3192 752 3208 768
rect 3144 732 3160 748
rect 3128 712 3144 728
rect 3096 692 3112 708
rect 3112 552 3128 568
rect 3128 532 3144 548
rect 3080 512 3096 528
rect 3144 512 3160 528
rect 3192 512 3208 528
rect 3048 492 3064 508
rect 2984 372 3000 388
rect 3080 492 3096 508
rect 3112 392 3128 408
rect 3048 332 3080 348
rect 2968 292 2984 308
rect 2952 272 2968 288
rect 2664 232 2680 248
rect 2600 172 2616 188
rect 2536 132 2552 148
rect 2568 132 2584 148
rect 2616 132 2632 148
rect 2728 232 2744 248
rect 2712 192 2728 208
rect 2776 132 2792 148
rect 2408 112 2424 128
rect 2440 112 2456 128
rect 2472 112 2488 128
rect 2584 112 2600 128
rect 2632 112 2648 128
rect 2392 92 2408 108
rect 2584 92 2600 108
rect 2712 92 2728 108
rect 2744 92 2760 108
rect 2808 112 2824 128
rect 2952 172 2968 188
rect 2952 152 2968 168
rect 3000 292 3016 308
rect 3064 312 3080 328
rect 3128 372 3144 388
rect 2936 132 2952 148
rect 3048 172 3064 188
rect 3144 132 3160 148
rect 2936 112 2952 128
rect 3192 112 3208 128
rect 2424 72 2440 88
rect 2552 72 2568 88
rect 2360 52 2376 68
rect 2472 52 2488 68
rect 1037 2 1073 18
rect 1896 12 1912 28
rect 1960 12 1992 28
rect 2040 12 2056 28
rect 2104 12 2120 28
rect 2168 12 2184 28
rect 2424 12 2440 28
<< metal3 >>
rect 1976 2197 1992 2203
rect 2888 2217 2904 2223
rect 200 2177 2264 2183
rect 2280 2177 2296 2183
rect 2312 2177 2328 2183
rect 56 2157 360 2163
rect 376 2157 536 2163
rect 552 2157 776 2163
rect 904 2157 1000 2163
rect 1069 2157 1144 2163
rect 264 2137 376 2143
rect 392 2137 472 2143
rect 712 2137 744 2143
rect 1069 2143 1075 2157
rect 1192 2157 1304 2163
rect 2040 2157 2104 2163
rect 2408 2157 2504 2163
rect 2520 2157 2552 2163
rect 792 2137 1075 2143
rect 1096 2137 1192 2143
rect 1368 2137 1624 2143
rect 1656 2137 2040 2143
rect 2120 2137 2296 2143
rect 2536 2137 2680 2143
rect 2696 2137 2744 2143
rect 2792 2137 2824 2143
rect 2840 2137 2856 2143
rect 2872 2137 2904 2143
rect 2936 2137 2984 2143
rect 72 2117 168 2123
rect 184 2117 264 2123
rect 360 2117 424 2123
rect 440 2117 568 2123
rect 728 2117 808 2123
rect 936 2117 1240 2123
rect 1320 2117 1352 2123
rect 1368 2117 1384 2123
rect 1448 2117 1528 2123
rect 1608 2117 1672 2123
rect 1880 2117 1891 2123
rect 1928 2117 2056 2123
rect 2296 2117 2344 2123
rect 2600 2117 2616 2123
rect 2632 2117 2664 2123
rect 2680 2117 2760 2123
rect 2776 2117 3032 2123
rect 3080 2117 3112 2123
rect 104 2097 328 2103
rect 344 2097 440 2103
rect 776 2097 936 2103
rect 1080 2097 1096 2103
rect 1240 2097 1256 2103
rect 1672 2097 1720 2103
rect 1912 2097 2184 2103
rect 2424 2097 2536 2103
rect 2552 2097 2600 2103
rect 2616 2097 2808 2103
rect 2824 2097 2888 2103
rect 2904 2097 2952 2103
rect 152 2077 184 2083
rect 616 2077 1208 2083
rect 1224 2077 1368 2083
rect 1640 2077 1704 2083
rect 1720 2077 1848 2083
rect 1864 2077 1928 2083
rect 1960 2077 1976 2083
rect 2568 2077 2632 2083
rect 2648 2077 2696 2083
rect 2712 2077 2904 2083
rect 2920 2077 2968 2083
rect 3000 2077 3016 2083
rect 408 2057 664 2063
rect 744 2057 872 2063
rect 888 2057 1080 2063
rect 2184 2057 2776 2063
rect 536 2037 568 2043
rect 872 2037 1000 2043
rect 2856 2037 2904 2043
rect 792 2017 920 2023
rect 968 1997 1016 2003
rect 2360 2017 2376 2023
rect 2920 2017 2968 2023
rect 424 1977 952 1983
rect 1240 1977 1656 1983
rect 568 1957 792 1963
rect 1000 1957 1160 1963
rect 1176 1957 1256 1963
rect 1272 1957 1304 1963
rect 1976 1957 2488 1963
rect 2504 1957 2776 1963
rect 3064 1957 3176 1963
rect 3192 1957 3251 1963
rect 520 1937 1176 1943
rect 1192 1937 1608 1943
rect 2168 1937 2216 1943
rect 2232 1937 2456 1943
rect 2472 1937 2632 1943
rect 2648 1937 2808 1943
rect 168 1917 184 1923
rect 712 1917 856 1923
rect 888 1917 1080 1923
rect 1096 1917 1128 1923
rect 1144 1917 1288 1923
rect 1432 1917 1480 1923
rect 1656 1917 1704 1923
rect 2056 1917 2136 1923
rect 2520 1917 2824 1923
rect 2872 1917 2888 1923
rect 2936 1917 2952 1923
rect 3048 1917 3160 1923
rect 3176 1917 3251 1923
rect 40 1897 264 1903
rect 344 1897 472 1903
rect 488 1897 520 1903
rect 536 1897 648 1903
rect 696 1897 840 1903
rect 984 1897 1128 1903
rect 1144 1897 1240 1903
rect 1304 1897 1448 1903
rect 1464 1897 1512 1903
rect 1608 1897 1800 1903
rect 1816 1897 1864 1903
rect 1976 1897 1992 1903
rect 2072 1897 2136 1903
rect 2184 1897 2232 1903
rect 2488 1897 2499 1903
rect 2584 1897 2600 1903
rect 2712 1897 2728 1903
rect 2760 1897 2899 1903
rect 88 1877 168 1883
rect 184 1877 264 1883
rect 296 1877 344 1883
rect 520 1877 664 1883
rect 776 1877 920 1883
rect 936 1877 1016 1883
rect 1048 1877 1224 1883
rect 1256 1877 1400 1883
rect 1416 1877 1592 1883
rect 1704 1877 1768 1883
rect 1784 1877 2008 1883
rect 2216 1877 2328 1883
rect 2344 1877 2616 1883
rect 2776 1877 2872 1883
rect 2893 1883 2899 1897
rect 2968 1897 2984 1903
rect 3016 1897 3080 1903
rect 2893 1877 3000 1883
rect 168 1857 728 1863
rect 744 1857 872 1863
rect 904 1857 1496 1863
rect 1512 1857 1592 1863
rect 1608 1857 1656 1863
rect 1832 1857 1896 1863
rect 1960 1857 2104 1863
rect 2136 1857 2168 1863
rect 2840 1857 2856 1863
rect 2888 1857 2936 1863
rect 2952 1857 3000 1863
rect 3016 1857 3080 1863
rect 3096 1857 3112 1863
rect 248 1837 376 1843
rect 392 1837 424 1843
rect 632 1837 904 1843
rect 1128 1837 1208 1843
rect 1240 1837 1272 1843
rect 1384 1837 1512 1843
rect 1528 1837 1688 1843
rect 1816 1837 1944 1843
rect 2136 1837 2696 1843
rect 2968 1837 3064 1843
rect 680 1817 1080 1823
rect 1112 1817 1267 1823
rect 232 1797 1000 1803
rect 1016 1797 1144 1803
rect 1261 1803 1267 1817
rect 1288 1817 1624 1823
rect 1688 1817 2040 1823
rect 1261 1797 1464 1803
rect 1512 1797 1624 1803
rect 1768 1797 1832 1803
rect 1853 1797 2056 1803
rect 232 1777 1075 1783
rect 280 1757 344 1763
rect 360 1757 440 1763
rect 664 1757 696 1763
rect 824 1757 952 1763
rect 1069 1763 1075 1777
rect 1096 1777 1656 1783
rect 1853 1783 1859 1797
rect 2360 1817 2472 1823
rect 2200 1797 2408 1803
rect 1832 1777 1859 1783
rect 1976 1777 2040 1783
rect 2072 1777 2312 1783
rect 1069 1757 1208 1763
rect 1224 1757 1336 1763
rect 1368 1757 1496 1763
rect 1512 1757 1720 1763
rect 1736 1757 1832 1763
rect 1912 1757 1976 1763
rect 1992 1757 2051 1763
rect 104 1737 184 1743
rect 328 1737 408 1743
rect 440 1737 744 1743
rect 760 1737 792 1743
rect 920 1737 968 1743
rect 989 1737 995 1752
rect 1032 1737 1112 1743
rect 1128 1737 1176 1743
rect 1448 1737 1768 1743
rect 1885 1743 1891 1752
rect 1880 1737 1891 1743
rect 2045 1743 2051 1757
rect 2328 1757 2408 1763
rect 2536 1757 2600 1763
rect 2045 1737 2168 1743
rect 2296 1737 2424 1743
rect 2488 1737 2536 1743
rect 2552 1737 2616 1743
rect 2744 1737 2760 1743
rect 3000 1737 3096 1743
rect 1373 1728 1379 1732
rect 88 1717 152 1723
rect 248 1717 280 1723
rect 344 1717 360 1723
rect 424 1717 472 1723
rect 488 1717 600 1723
rect 616 1717 728 1723
rect 744 1717 760 1723
rect 824 1717 856 1723
rect 1176 1717 1240 1723
rect 1320 1717 1336 1723
rect 1512 1717 1544 1723
rect 1848 1717 2152 1723
rect 2312 1717 2408 1723
rect 2424 1717 2520 1723
rect 2600 1717 2840 1723
rect 2968 1717 3032 1723
rect 3080 1717 3112 1723
rect 152 1697 248 1703
rect 552 1697 584 1703
rect 712 1697 856 1703
rect 920 1697 1016 1703
rect 1160 1697 1267 1703
rect 104 1677 168 1683
rect 424 1677 840 1683
rect 872 1677 1208 1683
rect 1261 1683 1267 1697
rect 1288 1697 1496 1703
rect 1576 1697 1640 1703
rect 1944 1697 1960 1703
rect 2040 1697 2184 1703
rect 2440 1697 2488 1703
rect 2584 1697 2904 1703
rect 3000 1697 3016 1703
rect 1261 1677 1304 1683
rect 1352 1677 1448 1683
rect 1576 1677 1688 1683
rect 1704 1677 2024 1683
rect 2408 1677 2488 1683
rect 2664 1677 2696 1683
rect 2712 1677 2792 1683
rect 184 1657 584 1663
rect 824 1657 984 1663
rect 1096 1657 2232 1663
rect 568 1637 632 1643
rect 856 1637 888 1643
rect 952 1637 1752 1643
rect 1768 1637 1816 1643
rect 1896 1637 1912 1643
rect 1928 1637 2008 1643
rect 616 1617 648 1623
rect 1352 1617 1656 1623
rect 1688 1617 1768 1623
rect 2008 1617 2232 1623
rect 1560 1597 3048 1603
rect -51 1577 88 1583
rect 104 1577 712 1583
rect 744 1577 1384 1583
rect 1496 1577 1976 1583
rect 2328 1577 2376 1583
rect 2808 1577 2920 1583
rect 24 1557 88 1563
rect 104 1557 440 1563
rect 456 1557 504 1563
rect 520 1557 760 1563
rect 1144 1557 1272 1563
rect 1400 1557 1592 1563
rect 1672 1557 1768 1563
rect 2040 1557 2664 1563
rect 2712 1557 2984 1563
rect 3208 1557 3251 1563
rect -51 1537 136 1543
rect 152 1537 376 1543
rect 392 1537 680 1543
rect 792 1537 1064 1543
rect 1080 1537 1208 1543
rect 1224 1537 1448 1543
rect 1512 1537 1672 1543
rect 1720 1537 2200 1543
rect 2520 1537 2616 1543
rect 2648 1537 2792 1543
rect 2888 1537 2984 1543
rect 1693 1528 1699 1532
rect 408 1517 488 1523
rect 504 1517 872 1523
rect 888 1517 984 1523
rect 1069 1517 1464 1523
rect -51 1497 8 1503
rect 88 1497 296 1503
rect 376 1497 504 1503
rect 520 1497 552 1503
rect 568 1497 664 1503
rect 680 1497 744 1503
rect 1069 1503 1075 1517
rect 1496 1517 1512 1523
rect 1725 1517 1736 1523
rect 2200 1517 2248 1523
rect 2424 1517 2712 1523
rect 2728 1517 2792 1523
rect 2920 1517 3251 1523
rect 1000 1497 1075 1503
rect 1096 1497 1112 1503
rect 1192 1497 1256 1503
rect 1336 1497 1464 1503
rect 1656 1497 1704 1503
rect 1800 1497 1816 1503
rect 1960 1497 2280 1503
rect 2584 1497 2600 1503
rect 2776 1497 2808 1503
rect 2856 1497 2904 1503
rect 56 1477 200 1483
rect 296 1477 424 1483
rect 440 1477 536 1483
rect 632 1477 856 1483
rect 984 1477 1096 1483
rect 1384 1477 1528 1483
rect 1768 1477 1784 1483
rect 1928 1477 1960 1483
rect 2120 1477 2131 1483
rect 2168 1477 2328 1483
rect 2344 1477 2408 1483
rect 2664 1477 2680 1483
rect 2840 1477 2888 1483
rect 24 1457 216 1463
rect 232 1457 520 1463
rect 536 1457 632 1463
rect 1112 1457 1144 1463
rect 1309 1457 1320 1463
rect 1448 1457 2216 1463
rect 2296 1457 2360 1463
rect 2392 1457 2648 1463
rect 2664 1457 2744 1463
rect 2760 1457 2872 1463
rect 344 1437 568 1443
rect 696 1437 1880 1443
rect 2104 1437 2120 1443
rect 2232 1437 2728 1443
rect 2888 1437 3016 1443
rect 1933 1428 1939 1432
rect 584 1417 1656 1423
rect 1672 1417 1720 1423
rect 152 1397 216 1403
rect 605 1397 824 1403
rect 88 1377 264 1383
rect 280 1377 328 1383
rect 360 1377 536 1383
rect 605 1383 611 1397
rect 872 1397 1032 1403
rect 1048 1397 1160 1403
rect 1176 1397 1192 1403
rect 1208 1397 1416 1403
rect 1432 1397 1576 1403
rect 1592 1397 1608 1403
rect 1800 1397 2024 1403
rect 2440 1417 2504 1423
rect 2536 1417 2600 1423
rect 2616 1417 2872 1423
rect 2152 1397 2248 1403
rect 2264 1397 2552 1403
rect 2792 1397 3000 1403
rect 3016 1397 3128 1403
rect 552 1377 611 1383
rect 760 1377 856 1383
rect 1144 1377 1192 1383
rect 1320 1377 1496 1383
rect 1752 1377 2056 1383
rect 2184 1377 2504 1383
rect 2536 1377 2552 1383
rect 2568 1377 2584 1383
rect -51 1357 72 1363
rect 136 1357 600 1363
rect 744 1357 1176 1363
rect 1256 1357 1368 1363
rect 1384 1357 1480 1363
rect 1848 1357 2008 1363
rect 2200 1357 2232 1363
rect 2264 1357 2296 1363
rect 2312 1357 2488 1363
rect 2840 1357 3251 1363
rect 152 1337 168 1343
rect 200 1337 408 1343
rect 424 1337 552 1343
rect 680 1337 1016 1343
rect 1032 1337 1192 1343
rect 1240 1337 1256 1343
rect 1272 1337 1400 1343
rect 1416 1337 1512 1343
rect 1624 1337 1704 1343
rect 1896 1337 1944 1343
rect 2024 1337 2200 1343
rect 2232 1337 2408 1343
rect 2504 1337 2536 1343
rect 2568 1337 2584 1343
rect 2840 1337 2872 1343
rect 2968 1337 3064 1343
rect -51 1317 8 1323
rect 56 1317 88 1323
rect 104 1317 168 1323
rect 200 1317 296 1323
rect 312 1317 392 1323
rect 445 1317 456 1323
rect 616 1317 680 1323
rect 712 1317 776 1323
rect 824 1317 952 1323
rect 968 1317 1016 1323
rect 1032 1317 1080 1323
rect 1112 1317 1251 1323
rect 72 1297 488 1303
rect 504 1297 568 1303
rect 984 1297 1000 1303
rect 1016 1297 1144 1303
rect 1245 1303 1251 1317
rect 1272 1317 1352 1323
rect 1368 1317 1464 1323
rect 1480 1317 1544 1323
rect 1640 1317 1784 1323
rect 1896 1317 1960 1323
rect 2008 1317 2168 1323
rect 2184 1317 2248 1323
rect 2648 1317 2680 1323
rect 2696 1317 2824 1323
rect 2856 1317 2904 1323
rect 2920 1317 3251 1323
rect 1245 1297 1560 1303
rect 1576 1297 1704 1303
rect 1816 1297 1896 1303
rect 1944 1297 2088 1303
rect 2152 1297 2200 1303
rect 2344 1297 2456 1303
rect 2568 1297 2712 1303
rect 904 1277 1288 1283
rect 1304 1277 1368 1283
rect 1880 1277 1928 1283
rect 1944 1277 2008 1283
rect 2152 1277 2264 1283
rect 2312 1277 2376 1283
rect 2472 1277 2584 1283
rect 952 1257 1480 1263
rect 1496 1257 1528 1263
rect 1640 1257 1688 1263
rect 1704 1257 1736 1263
rect 1752 1257 1768 1263
rect 1784 1257 2008 1263
rect 2024 1257 2296 1263
rect 2424 1257 2776 1263
rect 680 1237 1171 1243
rect 1165 1223 1171 1237
rect 2136 1237 2232 1243
rect 2248 1237 2344 1243
rect 136 1197 280 1203
rect 1165 1217 1320 1223
rect 1480 1217 1528 1223
rect 1640 1217 1896 1223
rect 1912 1217 2056 1223
rect 2072 1217 2104 1223
rect 2120 1217 2152 1223
rect 1480 1197 1576 1203
rect 1592 1197 1624 1203
rect 2056 1197 2296 1203
rect 392 1177 408 1183
rect 776 1177 888 1183
rect 904 1177 1080 1183
rect 1160 1177 1304 1183
rect 1320 1177 1336 1183
rect 1448 1177 1672 1183
rect 1768 1177 2392 1183
rect 264 1157 312 1163
rect 424 1157 536 1163
rect 552 1157 696 1163
rect 856 1157 920 1163
rect 936 1157 1368 1163
rect 1592 1157 1608 1163
rect 1800 1157 1848 1163
rect 1880 1157 1896 1163
rect 72 1137 136 1143
rect 152 1137 344 1143
rect 456 1137 1240 1143
rect 1256 1137 1416 1143
rect 1432 1137 1480 1143
rect 1512 1137 1880 1143
rect 2040 1137 2552 1143
rect 2760 1137 2904 1143
rect 264 1117 600 1123
rect 664 1117 808 1123
rect 1128 1117 1144 1123
rect 1224 1117 1288 1123
rect 1464 1117 2024 1123
rect 2040 1117 2120 1123
rect 2328 1117 2408 1123
rect 2520 1117 2600 1123
rect 2728 1117 2792 1123
rect 1213 1108 1219 1112
rect 216 1097 232 1103
rect 280 1097 312 1103
rect 600 1097 616 1103
rect 632 1097 696 1103
rect 728 1097 792 1103
rect 808 1097 840 1103
rect 968 1097 1192 1103
rect 1272 1097 1288 1103
rect 1624 1097 1656 1103
rect 2056 1097 2120 1103
rect 2152 1097 2168 1103
rect 2248 1097 2440 1103
rect 2456 1097 2472 1103
rect 2488 1097 2648 1103
rect 2664 1097 2824 1103
rect 1757 1088 1763 1092
rect 1981 1088 1987 1092
rect 152 1077 280 1083
rect 296 1077 472 1083
rect 536 1077 680 1083
rect 696 1077 792 1083
rect 920 1077 1000 1083
rect 1048 1077 1064 1083
rect 1144 1077 1331 1083
rect 696 1057 712 1063
rect 888 1057 1144 1063
rect 1192 1057 1256 1063
rect 1325 1063 1331 1077
rect 1352 1077 1528 1083
rect 1560 1077 1608 1083
rect 1624 1077 1736 1083
rect 2040 1077 2216 1083
rect 2248 1077 2456 1083
rect 2712 1077 2760 1083
rect 2888 1077 2936 1083
rect 2984 1077 3048 1083
rect 3064 1077 3112 1083
rect 1325 1057 1448 1063
rect 1608 1057 1784 1063
rect 1800 1057 2408 1063
rect 2600 1057 2696 1063
rect 3032 1057 3192 1063
rect 3208 1057 3251 1063
rect 24 1037 72 1043
rect 328 1037 664 1043
rect 776 1037 1400 1043
rect 1448 1037 2808 1043
rect 88 1017 344 1023
rect 360 1017 488 1023
rect 632 1017 984 1023
rect 1016 1017 1560 1023
rect 1656 1017 1704 1023
rect 1848 1017 1880 1023
rect 488 997 824 1003
rect 952 997 968 1003
rect 1384 997 1544 1003
rect 1560 997 1592 1003
rect 1640 997 1768 1003
rect 1800 997 1864 1003
rect 1896 997 1960 1003
rect 1976 997 2008 1003
rect 2216 1017 2344 1023
rect 2520 1017 3064 1023
rect 2237 997 2632 1003
rect 72 977 104 983
rect 392 977 696 983
rect 712 977 824 983
rect 840 977 920 983
rect 936 977 1048 983
rect 1064 977 1096 983
rect 2237 983 2243 997
rect 1672 977 2243 983
rect 2296 977 2472 983
rect 2520 977 2536 983
rect -51 957 8 963
rect 56 957 88 963
rect 120 957 168 963
rect 184 957 200 963
rect 456 957 488 963
rect 536 957 568 963
rect 600 957 611 963
rect 808 957 936 963
rect 952 957 1064 963
rect 1128 957 1144 963
rect 1192 957 1288 963
rect 1384 957 1656 963
rect 1816 957 1832 963
rect 1848 957 2152 963
rect 2280 957 2344 963
rect 2360 957 2440 963
rect 2456 957 2712 963
rect 2968 957 3000 963
rect 3016 957 3080 963
rect 40 937 184 943
rect 200 937 248 943
rect 328 937 360 943
rect 392 937 424 943
rect 488 937 712 943
rect 728 937 1000 943
rect 1016 937 1640 943
rect 1704 937 1752 943
rect 1768 937 1848 943
rect 1928 937 1992 943
rect 2328 937 2424 943
rect 2760 937 2824 943
rect 3064 937 3096 943
rect -51 917 8 923
rect 56 917 72 923
rect 152 917 216 923
rect 232 917 296 923
rect 424 917 472 923
rect 664 917 952 923
rect 1032 917 1043 923
rect 1096 917 1160 923
rect 1320 917 1432 923
rect 1656 917 1752 923
rect 1768 917 2056 923
rect 2072 917 2088 923
rect 2136 917 2248 923
rect 2296 917 2312 923
rect 2584 917 2600 923
rect 3000 917 3144 923
rect 3208 917 3251 923
rect 317 908 323 912
rect 493 908 499 912
rect 2365 908 2371 912
rect 40 897 120 903
rect 712 897 776 903
rect 936 897 1048 903
rect 1080 897 1224 903
rect 1240 897 1384 903
rect 1400 897 1416 903
rect 1432 897 1464 903
rect 1736 897 1848 903
rect 1880 897 2104 903
rect 2168 897 2184 903
rect 2552 897 2584 903
rect 2616 897 2936 903
rect 2952 897 3000 903
rect 1272 877 1336 883
rect 1416 877 1576 883
rect 1592 877 2008 883
rect 2584 877 2595 883
rect 2616 877 2840 883
rect 24 857 88 863
rect 104 857 152 863
rect 600 857 1048 863
rect 1064 857 1096 863
rect 1432 857 2216 863
rect 2360 857 2600 863
rect 616 837 632 843
rect 648 837 856 843
rect 1144 837 1304 843
rect 1725 837 1864 843
rect 168 797 344 803
rect 1725 823 1731 837
rect 1896 837 2296 843
rect 2392 837 2616 843
rect 1224 817 1731 823
rect 1752 817 1816 823
rect 2088 817 2248 823
rect 2264 817 2408 823
rect 1144 797 1480 803
rect 1704 797 1720 803
rect 1976 797 2344 803
rect 2360 797 2504 803
rect 24 777 536 783
rect 824 777 1304 783
rect 1464 777 1592 783
rect 1736 777 2408 783
rect 2952 777 2968 783
rect 152 757 408 763
rect 424 757 472 763
rect 488 757 520 763
rect 760 757 1032 763
rect 1544 757 1592 763
rect 2424 757 2728 763
rect 3208 757 3251 763
rect 312 737 392 743
rect 408 737 600 743
rect 840 737 1064 743
rect 1288 737 1352 743
rect 1608 737 2088 743
rect 2104 737 2184 743
rect 2408 737 2456 743
rect 2872 737 3000 743
rect 3016 737 3144 743
rect 1229 728 1235 732
rect 280 717 408 723
rect 440 717 504 723
rect 584 717 648 723
rect 1048 717 1192 723
rect 1800 717 1912 723
rect 2152 717 2232 723
rect 2248 717 2296 723
rect 2344 717 2376 723
rect 2392 717 2520 723
rect 2568 717 2584 723
rect 2680 717 2728 723
rect 2920 717 2968 723
rect 3144 717 3251 723
rect 925 708 931 712
rect -51 697 8 703
rect 248 697 312 703
rect 504 697 664 703
rect 792 697 840 703
rect 941 703 947 712
rect 1405 708 1411 712
rect 941 697 952 703
rect 1160 697 1240 703
rect 1496 697 1528 703
rect 1640 697 1752 703
rect 2008 697 2040 703
rect 2072 697 2216 703
rect 2232 697 2520 703
rect 2536 697 2776 703
rect 2840 697 2888 703
rect 3032 697 3096 703
rect 88 677 136 683
rect 216 677 536 683
rect 616 677 1128 683
rect 1144 677 1176 683
rect 1208 677 1304 683
rect 1352 677 1608 683
rect 1944 677 1960 683
rect 2024 677 2120 683
rect 2152 677 2200 683
rect 2296 677 2552 683
rect 2776 677 2904 683
rect 136 657 280 663
rect 296 657 328 663
rect 600 657 632 663
rect 984 657 1656 663
rect 1725 657 2360 663
rect 488 637 568 643
rect 584 637 712 643
rect 840 637 1352 643
rect 1725 643 1731 657
rect 1704 637 1731 643
rect 1752 637 2200 643
rect 2280 637 2360 643
rect 2408 637 2536 643
rect 536 617 1048 623
rect 1064 617 1144 623
rect 1384 617 1704 623
rect 104 597 1096 603
rect 1240 597 1256 603
rect 1336 597 1384 603
rect 1400 597 1432 603
rect 1496 597 1896 603
rect 1960 597 2056 603
rect 2264 617 2728 623
rect 2136 597 2211 603
rect 664 577 1032 583
rect 1048 577 1272 583
rect 1288 577 1480 583
rect 1864 577 2168 583
rect 2205 583 2211 597
rect 2264 597 2280 603
rect 2376 597 2536 603
rect 2205 577 2392 583
rect 2680 577 2872 583
rect 152 557 184 563
rect 792 557 808 563
rect 1416 557 1592 563
rect 1624 557 1960 563
rect 1992 557 2488 563
rect 2936 557 3064 563
rect 3080 557 3112 563
rect 136 537 408 543
rect 424 537 520 543
rect 536 537 616 543
rect 808 537 1240 543
rect 1528 537 2344 543
rect 2360 537 2408 543
rect 2536 537 2552 543
rect 2728 537 2824 543
rect 2840 537 2856 543
rect 2920 537 2984 543
rect 200 517 232 523
rect 408 517 536 523
rect 568 517 600 523
rect 888 517 920 523
rect 1032 517 1176 523
rect 1208 517 1224 523
rect 1288 517 1496 523
rect 1592 517 1640 523
rect 1800 517 1880 523
rect 1896 517 1928 523
rect 1944 517 2024 523
rect 2168 517 2184 523
rect 2232 517 2296 523
rect 2376 517 2424 523
rect 2488 517 2504 523
rect 2520 517 2616 523
rect 2904 517 3064 523
rect 3208 517 3251 523
rect 312 497 392 503
rect 552 497 568 503
rect 760 497 808 503
rect 824 497 856 503
rect 1112 497 1336 503
rect 1368 497 1400 503
rect 1480 497 1544 503
rect 1640 497 1768 503
rect 1784 497 1800 503
rect 1960 497 2120 503
rect 2232 497 2376 503
rect 2408 497 2488 503
rect 2600 497 2648 503
rect 2888 497 2920 503
rect 3064 497 3080 503
rect 264 477 296 483
rect 328 477 360 483
rect 504 477 808 483
rect 872 477 1192 483
rect 1416 477 1816 483
rect 1832 477 2040 483
rect 2056 477 2104 483
rect 2328 477 2600 483
rect 2616 477 2872 483
rect 808 457 872 463
rect 904 457 1000 463
rect 1208 457 1416 463
rect 1432 457 1512 463
rect 1576 457 1976 463
rect 2072 457 2248 463
rect 2392 457 2472 463
rect 1240 437 1592 443
rect 1608 437 1672 443
rect 1816 437 1912 443
rect 2072 437 2232 443
rect 280 417 792 423
rect 520 397 712 403
rect 1352 417 1400 423
rect 1672 417 2120 423
rect 2168 417 2408 423
rect 1112 397 2392 403
rect 2616 397 2872 403
rect 2888 397 3112 403
rect 200 377 648 383
rect 744 377 776 383
rect 808 377 1304 383
rect 1336 377 1656 383
rect 1976 377 2168 383
rect 3000 377 3128 383
rect 680 357 712 363
rect 728 357 888 363
rect 1384 357 1400 363
rect 1416 357 1432 363
rect 1448 357 1496 363
rect 1512 357 1608 363
rect 1624 357 1864 363
rect 1960 357 1992 363
rect 2040 357 2136 363
rect 2344 357 2872 363
rect 2888 357 2920 363
rect 392 337 408 343
rect 424 337 472 343
rect 568 337 616 343
rect 632 337 824 343
rect 840 337 920 343
rect 952 337 1112 343
rect 1320 337 1336 343
rect 1816 337 1832 343
rect 1864 337 3048 343
rect 24 317 56 323
rect 72 317 216 323
rect 232 317 248 323
rect 264 317 360 323
rect 392 317 504 323
rect 520 317 1304 323
rect 1656 317 2056 323
rect 2216 317 2232 323
rect 2280 317 2344 323
rect 2392 317 2504 323
rect 2552 317 2760 323
rect 3069 308 3075 312
rect 104 297 152 303
rect 184 297 200 303
rect 264 297 344 303
rect 408 297 664 303
rect 680 297 984 303
rect 1000 297 1128 303
rect 1240 297 1288 303
rect 1320 297 1400 303
rect 1416 297 1464 303
rect 1592 297 1624 303
rect 1688 297 2040 303
rect 2088 297 2184 303
rect 2440 297 2488 303
rect 2584 297 2744 303
rect 2904 297 2915 303
rect 2984 297 3000 303
rect 72 277 360 283
rect 392 277 424 283
rect 456 277 488 283
rect 984 277 1144 283
rect 1192 277 1240 283
rect 1256 277 1272 283
rect 1448 277 1459 283
rect 1485 277 1608 283
rect 88 257 136 263
rect 296 257 536 263
rect 568 257 584 263
rect 744 257 824 263
rect 1016 257 1080 263
rect 1485 263 1491 277
rect 1704 277 1864 283
rect 1896 277 2216 283
rect 2264 277 2280 283
rect 2408 277 2456 283
rect 2477 277 2552 283
rect 1448 257 1491 263
rect 1512 257 1720 263
rect 2024 257 2072 263
rect 2477 263 2483 277
rect 2616 277 2952 283
rect 2344 257 2483 263
rect 2504 257 2584 263
rect 2733 248 2739 252
rect 24 237 56 243
rect 760 237 920 243
rect 936 237 968 243
rect 1544 237 1683 243
rect 104 217 488 223
rect 920 217 1144 223
rect 1592 217 1656 223
rect 1677 223 1683 237
rect 1704 237 1944 243
rect 1976 237 2232 243
rect 2680 237 2728 243
rect 1677 217 1816 223
rect 1848 217 1912 223
rect 264 197 392 203
rect 424 197 792 203
rect 824 197 1560 203
rect 1576 197 1736 203
rect 1752 197 1784 203
rect 1832 197 2056 203
rect 2328 197 2712 203
rect 328 177 440 183
rect 456 177 680 183
rect 696 177 872 183
rect 888 177 1016 183
rect 1032 177 1096 183
rect 1112 177 1160 183
rect 1336 177 1496 183
rect 1624 177 1816 183
rect 1880 177 2040 183
rect 2184 177 2296 183
rect 2504 177 2600 183
rect 2968 177 3048 183
rect 1613 168 1619 172
rect 248 157 472 163
rect 856 157 1032 163
rect 1048 157 1176 163
rect 1192 157 1304 163
rect 1384 157 1512 163
rect 1656 157 1704 163
rect 1736 157 1864 163
rect 2264 157 2344 163
rect 2424 157 2952 163
rect 1885 148 1891 152
rect 120 137 152 143
rect 168 137 264 143
rect 280 137 344 143
rect 360 137 520 143
rect 536 137 584 143
rect 1080 137 1096 143
rect 1128 137 1336 143
rect 1352 137 1400 143
rect 1672 137 1768 143
rect 1944 137 2184 143
rect 2584 137 2616 143
rect 2792 137 2936 143
rect 1805 128 1811 132
rect 3149 128 3155 132
rect -51 117 8 123
rect 184 117 200 123
rect 280 117 312 123
rect 344 117 376 123
rect 472 117 488 123
rect 632 117 728 123
rect 872 117 888 123
rect 952 117 984 123
rect 1032 117 1112 123
rect 1208 117 1224 123
rect 1272 117 1320 123
rect 1464 117 1480 123
rect 1757 117 1768 123
rect 1960 117 1992 123
rect 2424 117 2440 123
rect 2488 117 2584 123
rect 2600 117 2632 123
rect 2824 117 2936 123
rect 3208 117 3251 123
rect 200 97 360 103
rect 408 97 424 103
rect 488 97 664 103
rect 680 97 888 103
rect 1240 97 1288 103
rect 1320 97 1448 103
rect 1496 97 1672 103
rect 2024 97 2136 103
rect 2168 97 2280 103
rect 2296 97 2392 103
rect 2600 97 2712 103
rect 2760 97 2771 103
rect 232 77 264 83
rect 296 77 440 83
rect 552 77 648 83
rect 680 77 712 83
rect 744 77 776 83
rect 904 77 936 83
rect 1128 77 1352 83
rect 1368 77 1384 83
rect 1816 77 2424 83
rect 2440 77 2552 83
rect 808 57 1560 63
rect 2376 57 2472 63
rect 600 37 1272 43
rect 1912 17 1960 23
rect 1992 17 2040 23
rect 2120 17 2168 23
<< m4contact >>
rect 1096 2212 1112 2228
rect 2078 2202 2106 2218
rect 1624 2132 1640 2148
rect 3096 2132 3112 2148
rect 1240 2112 1256 2128
rect 1864 2112 1880 2128
rect 3064 2112 3080 2128
rect 440 2092 456 2108
rect 1096 2092 1112 2108
rect 1256 2092 1272 2108
rect 1656 2092 1672 2108
rect 184 2072 200 2088
rect 1000 2032 1016 2048
rect 728 2012 744 2028
rect 1038 2002 1066 2018
rect 2376 2012 2392 2028
rect 808 1952 824 1968
rect 856 1912 872 1928
rect 1336 1912 1352 1928
rect 1368 1912 1384 1928
rect 1384 1912 1400 1928
rect 1752 1912 1768 1928
rect 1816 1912 1832 1928
rect 664 1892 680 1908
rect 1128 1892 1144 1908
rect 2136 1892 2152 1908
rect 2168 1892 2184 1908
rect 2472 1892 2488 1908
rect 344 1872 360 1888
rect 1224 1872 1240 1888
rect 2760 1872 2776 1888
rect 872 1852 888 1868
rect 1688 1852 1704 1868
rect 1896 1852 1912 1868
rect 2344 1852 2360 1868
rect 2504 1852 2520 1868
rect 1208 1832 1224 1848
rect 1080 1812 1096 1828
rect 2040 1812 2056 1828
rect 1624 1792 1640 1808
rect 1832 1792 1848 1808
rect 984 1752 1000 1768
rect 1016 1752 1032 1768
rect 1080 1772 1096 1788
rect 1656 1772 1672 1788
rect 2078 1802 2106 1818
rect 2184 1792 2200 1808
rect 2344 1772 2360 1788
rect 1336 1752 1352 1768
rect 1496 1752 1512 1768
rect 1880 1752 1896 1768
rect 1976 1752 1992 1768
rect 408 1732 424 1748
rect 856 1732 872 1748
rect 1016 1732 1032 1748
rect 1368 1732 1384 1748
rect 1944 1732 1960 1748
rect 3144 1752 3160 1768
rect 2424 1732 2440 1748
rect 2968 1732 2984 1748
rect 728 1712 744 1728
rect 1128 1712 1144 1728
rect 1240 1712 1256 1728
rect 1784 1712 1800 1728
rect 136 1692 152 1708
rect 584 1692 600 1708
rect 856 1692 872 1708
rect 840 1672 872 1688
rect 1272 1692 1288 1708
rect 3016 1692 3032 1708
rect 1336 1672 1352 1688
rect 1080 1652 1096 1668
rect 1038 1602 1066 1618
rect 1656 1612 1672 1628
rect 2376 1572 2392 1588
rect 88 1552 104 1568
rect 1128 1552 1144 1568
rect 1656 1552 1672 1568
rect 1912 1552 1928 1568
rect 1672 1532 1720 1548
rect 984 1512 1000 1528
rect 1016 1512 1032 1528
rect 1736 1512 1752 1528
rect 2168 1512 2184 1528
rect 1464 1492 1480 1508
rect 1496 1492 1512 1508
rect 1704 1492 1720 1508
rect 1816 1492 1832 1508
rect 2280 1492 2296 1508
rect 1192 1472 1208 1488
rect 1784 1472 1800 1488
rect 2104 1472 2120 1488
rect 2152 1472 2168 1488
rect 2808 1472 2824 1488
rect 632 1452 648 1468
rect 664 1452 680 1468
rect 1096 1452 1112 1468
rect 1320 1452 1336 1468
rect 2872 1452 2888 1468
rect 2120 1432 2136 1448
rect 1928 1412 1944 1428
rect 344 1372 360 1388
rect 840 1392 856 1408
rect 2024 1392 2040 1408
rect 2056 1392 2072 1408
rect 2078 1402 2106 1418
rect 2504 1412 2520 1428
rect 2776 1392 2792 1408
rect 3000 1392 3016 1408
rect 1496 1372 1512 1388
rect 2504 1372 2520 1388
rect 2552 1372 2568 1388
rect 1576 1352 1592 1368
rect 1720 1352 1736 1368
rect 2760 1352 2776 1368
rect 2824 1352 2840 1368
rect 552 1332 568 1348
rect 1256 1332 1272 1348
rect 1992 1332 2008 1348
rect 2008 1332 2024 1348
rect 2216 1332 2232 1348
rect 2648 1332 2664 1348
rect 184 1312 200 1328
rect 456 1312 472 1328
rect 696 1312 712 1328
rect 808 1312 824 1328
rect 1080 1312 1096 1328
rect 488 1292 504 1308
rect 1000 1292 1016 1308
rect 2248 1312 2264 1328
rect 2824 1312 2840 1328
rect 1704 1292 1720 1308
rect 1736 1292 1752 1308
rect 1368 1272 1384 1288
rect 1928 1272 1944 1288
rect 1480 1252 1496 1268
rect 1688 1252 1704 1268
rect 2776 1252 2792 1268
rect 1192 1232 1208 1248
rect 2344 1232 2360 1248
rect 1038 1202 1066 1218
rect 1576 1192 1592 1208
rect 2040 1192 2056 1208
rect 376 1172 392 1188
rect 1080 1172 1096 1188
rect 1432 1172 1448 1188
rect 2392 1172 2408 1188
rect 312 1152 328 1168
rect 920 1152 936 1168
rect 1896 1152 1912 1168
rect 2040 1152 2056 1168
rect 2024 1132 2040 1148
rect 88 1112 104 1128
rect 1144 1112 1160 1128
rect 1208 1112 1224 1128
rect 2408 1112 2424 1128
rect 840 1092 856 1108
rect 1288 1092 1304 1108
rect 1480 1092 1496 1108
rect 1544 1092 1560 1108
rect 1608 1092 1624 1108
rect 1688 1092 1704 1108
rect 1848 1092 1864 1108
rect 2120 1092 2136 1108
rect 2984 1092 3000 1108
rect 72 1072 88 1088
rect 680 1072 696 1088
rect 1064 1072 1080 1088
rect 504 1052 520 1068
rect 664 1052 680 1068
rect 1528 1072 1544 1088
rect 1736 1072 1768 1088
rect 1816 1072 1832 1088
rect 1912 1072 1928 1088
rect 1944 1072 1960 1088
rect 1976 1072 1992 1088
rect 2024 1072 2040 1088
rect 2232 1072 2248 1088
rect 2872 1052 2888 1068
rect 3016 1052 3032 1068
rect 72 1012 88 1028
rect 984 1012 1000 1028
rect 1640 1012 1656 1028
rect 1880 1012 1896 1028
rect 824 992 840 1008
rect 856 992 872 1008
rect 872 992 888 1008
rect 888 992 904 1008
rect 1592 992 1608 1008
rect 1624 992 1640 1008
rect 1864 992 1880 1008
rect 2008 992 2024 1008
rect 2078 1002 2106 1018
rect 2408 1012 2424 1028
rect 2504 1012 2520 1028
rect 2136 992 2152 1008
rect 1224 972 1240 988
rect 424 952 440 968
rect 584 952 600 968
rect 1064 952 1080 968
rect 1144 952 1160 968
rect 1720 952 1736 968
rect 1800 952 1816 968
rect 1896 932 1912 948
rect 8 912 24 928
rect 72 912 88 928
rect 136 912 152 928
rect 312 912 328 928
rect 488 912 504 928
rect 1016 912 1032 928
rect 1080 912 1096 928
rect 1432 912 1448 928
rect 1464 912 1480 928
rect 1624 912 1640 928
rect 2056 912 2072 928
rect 2120 912 2136 928
rect 2280 912 2296 928
rect 2360 912 2376 928
rect 2488 912 2504 928
rect 2744 912 2760 928
rect 2792 912 2808 928
rect 1048 892 1064 908
rect 1864 892 1880 908
rect 2584 892 2600 908
rect 2568 872 2584 888
rect 2600 872 2616 888
rect 8 852 24 868
rect 2344 852 2360 868
rect 1304 832 1320 848
rect 680 812 696 828
rect 1038 802 1066 818
rect 1864 832 1880 848
rect 2376 832 2392 848
rect 1128 792 1144 808
rect 2408 772 2424 788
rect 2424 772 2440 788
rect 3128 752 3144 768
rect 600 732 616 748
rect 664 732 680 748
rect 1544 732 1560 748
rect 1592 732 1608 748
rect 408 712 424 728
rect 648 712 664 728
rect 968 712 984 728
rect 1224 712 1240 728
rect 1400 712 1416 728
rect 1640 712 1656 728
rect 2552 712 2568 728
rect 2728 712 2744 728
rect 776 692 792 708
rect 856 692 872 708
rect 920 692 936 708
rect 952 692 968 708
rect 1144 692 1160 708
rect 1480 692 1496 708
rect 1992 692 2008 708
rect 2056 692 2072 708
rect 536 672 552 688
rect 584 672 616 688
rect 1128 672 1144 688
rect 1912 672 1928 688
rect 2136 672 2152 688
rect 2744 672 2760 688
rect 840 652 856 668
rect 1672 652 1688 668
rect 3000 652 3016 668
rect 2360 632 2376 648
rect 2392 632 2408 648
rect 1896 612 1912 628
rect 1096 592 1112 608
rect 1224 592 1240 608
rect 2056 592 2072 608
rect 2078 602 2106 618
rect 2248 612 2264 628
rect 2184 572 2200 588
rect 2536 592 2552 608
rect 504 552 520 568
rect 808 552 824 568
rect 1592 552 1608 568
rect 1960 552 1976 568
rect 2488 552 2504 568
rect 3064 552 3080 568
rect 776 532 792 548
rect 3112 532 3128 548
rect 376 512 392 528
rect 1192 512 1208 528
rect 1656 512 1672 528
rect 1928 512 1944 528
rect 3064 512 3080 528
rect 3128 512 3144 528
rect 808 492 824 508
rect 1336 492 1352 508
rect 1576 492 1592 508
rect 2120 492 2136 508
rect 2376 492 2392 508
rect 2520 492 2536 508
rect 2040 472 2056 488
rect 2056 432 2072 448
rect 792 412 808 428
rect 1038 402 1066 418
rect 2152 412 2168 428
rect 1096 392 1112 408
rect 2872 392 2888 408
rect 664 372 680 388
rect 1304 372 1320 388
rect 1960 372 1976 388
rect 1400 352 1416 368
rect 1608 352 1624 368
rect 1880 352 1896 368
rect 2136 352 2152 368
rect 1304 332 1320 348
rect 1656 332 1688 348
rect 1800 332 1816 348
rect 2536 312 2552 328
rect 1224 292 1240 308
rect 2040 292 2056 308
rect 2424 292 2440 308
rect 2888 292 2904 308
rect 3064 292 3080 308
rect 360 272 376 288
rect 424 272 440 288
rect 840 272 856 288
rect 1384 272 1400 288
rect 1432 272 1448 288
rect 584 252 600 268
rect 1864 272 1896 288
rect 1816 252 1832 268
rect 2600 272 2616 288
rect 2728 252 2744 268
rect 488 212 504 228
rect 1656 212 1672 228
rect 1832 212 1848 228
rect 2056 192 2072 208
rect 2078 202 2106 218
rect 472 152 488 168
rect 504 152 520 168
rect 1608 152 1624 168
rect 1864 152 1880 168
rect 2104 152 2120 168
rect 1000 132 1016 148
rect 1096 132 1112 148
rect 1880 132 1896 148
rect 2536 132 2552 148
rect 488 112 504 128
rect 792 112 808 128
rect 1016 112 1032 128
rect 1720 112 1736 128
rect 1768 112 1784 128
rect 1800 112 1816 128
rect 1848 112 1864 128
rect 3144 112 3160 128
rect 1288 92 1304 108
rect 2136 92 2152 108
rect 2744 92 2760 108
rect 1038 2 1066 18
rect 2424 12 2440 28
<< metal4 >>
rect 1101 2108 1107 2212
rect 2106 2206 2112 2214
rect 1629 2124 1635 2132
rect 1628 2116 1636 2124
rect 1884 2123 1892 2124
rect 1880 2117 1892 2123
rect 1884 2116 1892 2117
rect 93 1128 99 1552
rect 77 1028 83 1072
rect 77 928 83 1012
rect 141 928 147 1692
rect 189 1328 195 2072
rect 349 1388 355 1872
rect 412 1756 420 1764
rect 413 1748 419 1756
rect 445 1324 451 2092
rect 588 1716 596 1724
rect 589 1708 595 1716
rect 669 1468 675 1892
rect 733 1728 739 2012
rect 556 1436 564 1444
rect 557 1348 563 1436
rect 444 1323 452 1324
rect 444 1317 456 1323
rect 444 1316 452 1317
rect 317 928 323 1152
rect 13 868 19 912
rect 381 528 387 1172
rect 493 928 499 1292
rect 509 924 515 1052
rect 637 964 643 1452
rect 813 1328 819 1952
rect 876 1876 884 1884
rect 877 1868 883 1876
rect 1005 1844 1011 2032
rect 1066 2006 1072 2014
rect 1004 1836 1012 1844
rect 989 1744 995 1752
rect 988 1736 996 1744
rect 861 1708 867 1732
rect 844 1696 852 1704
rect 845 1688 851 1696
rect 861 1688 867 1692
rect 988 1656 996 1664
rect 989 1528 995 1656
rect 845 1384 851 1392
rect 844 1376 852 1384
rect 1005 1308 1011 1836
rect 1085 1788 1091 1812
rect 1036 1763 1044 1764
rect 1032 1757 1044 1763
rect 1036 1756 1044 1757
rect 1021 1528 1027 1732
rect 1066 1606 1072 1614
rect 1085 1328 1091 1652
rect 1101 1468 1107 2092
rect 1228 1896 1236 1904
rect 1133 1728 1139 1892
rect 1229 1888 1235 1896
rect 1212 1856 1220 1864
rect 1213 1848 1219 1856
rect 1245 1728 1251 2112
rect 1133 1568 1139 1712
rect 1066 1206 1072 1214
rect 669 1044 675 1052
rect 668 1036 676 1044
rect 604 963 612 964
rect 600 957 612 963
rect 604 956 612 957
rect 636 956 644 964
rect 508 916 516 924
rect 429 264 435 272
rect 428 256 436 264
rect 493 228 499 912
rect 509 568 515 916
rect 685 828 691 1072
rect 605 688 611 732
rect 653 704 659 712
rect 652 696 660 704
rect 493 128 499 212
rect 509 168 515 552
rect 541 184 547 672
rect 589 268 595 672
rect 669 388 675 732
rect 781 548 787 692
rect 845 668 851 1092
rect 908 1003 916 1004
rect 904 997 916 1003
rect 908 996 916 997
rect 861 708 867 992
rect 877 944 883 992
rect 876 936 884 944
rect 925 708 931 1152
rect 1068 1096 1076 1104
rect 1069 1088 1075 1096
rect 988 1056 996 1064
rect 989 1028 995 1056
rect 1069 924 1075 952
rect 1085 928 1091 1172
rect 1036 923 1044 924
rect 1032 917 1044 923
rect 1036 916 1044 917
rect 1068 916 1076 924
rect 956 723 964 724
rect 956 717 968 723
rect 956 716 964 717
rect 940 703 948 704
rect 940 697 952 703
rect 940 696 948 697
rect 813 508 819 552
rect 540 176 548 184
rect 797 128 803 412
rect 845 288 851 652
rect 1004 156 1012 164
rect 1005 148 1011 156
rect 1021 128 1027 912
rect 1066 806 1072 814
rect 1133 808 1139 1552
rect 1197 1248 1203 1472
rect 1261 1348 1267 2092
rect 1341 1904 1347 1912
rect 1373 1904 1379 1912
rect 1340 1896 1348 1904
rect 1372 1896 1380 1904
rect 1389 1884 1395 1912
rect 1388 1876 1396 1884
rect 1292 1703 1300 1704
rect 1288 1697 1300 1703
rect 1292 1696 1300 1697
rect 1341 1688 1347 1752
rect 1308 1463 1316 1464
rect 1308 1457 1320 1463
rect 1308 1456 1316 1457
rect 1149 968 1155 1112
rect 1133 688 1139 792
rect 1149 708 1155 952
rect 1066 406 1072 414
rect 1101 408 1107 592
rect 1197 528 1203 1232
rect 1213 1104 1219 1112
rect 1212 1096 1220 1104
rect 1229 728 1235 972
rect 1309 848 1315 1456
rect 1373 1288 1379 1732
rect 1501 1508 1507 1752
rect 1500 1476 1508 1484
rect 1501 1388 1507 1476
rect 1437 928 1443 1172
rect 1485 1108 1491 1252
rect 1581 1208 1587 1352
rect 1452 923 1460 924
rect 1452 917 1464 923
rect 1452 916 1460 917
rect 1229 308 1235 592
rect 1309 348 1315 372
rect 1405 368 1411 712
rect 1485 708 1491 1092
rect 1549 748 1555 1092
rect 1613 1084 1619 1092
rect 1612 1076 1620 1084
rect 1629 1008 1635 1792
rect 1661 1788 1667 2092
rect 1836 1923 1844 1924
rect 1832 1917 1844 1923
rect 1836 1916 1844 1917
rect 1708 1863 1716 1864
rect 1704 1857 1716 1863
rect 1708 1856 1716 1857
rect 1661 1568 1667 1612
rect 1677 1524 1683 1532
rect 1676 1516 1684 1524
rect 1693 1268 1699 1532
rect 1709 1508 1715 1532
rect 1724 1523 1732 1524
rect 1724 1517 1736 1523
rect 1724 1516 1732 1517
rect 1708 1116 1716 1124
rect 1709 1104 1715 1116
rect 1708 1103 1716 1104
rect 1704 1097 1716 1103
rect 1708 1096 1716 1097
rect 1597 748 1603 992
rect 1629 904 1635 912
rect 1628 896 1636 904
rect 1645 728 1651 1012
rect 1725 968 1731 1352
rect 1740 1336 1748 1344
rect 1741 1308 1747 1336
rect 1740 1096 1748 1104
rect 1741 1088 1747 1096
rect 1757 1088 1763 1912
rect 1789 1488 1795 1712
rect 1804 1503 1812 1504
rect 1804 1497 1816 1503
rect 1804 1496 1812 1497
rect 1821 1064 1827 1072
rect 1820 1056 1828 1064
rect 1837 924 1843 1792
rect 1885 1744 1891 1752
rect 1884 1736 1892 1744
rect 1901 1364 1907 1852
rect 1949 1724 1955 1732
rect 1948 1716 1956 1724
rect 1900 1356 1908 1364
rect 1868 1103 1876 1104
rect 1864 1097 1876 1103
rect 1868 1096 1876 1097
rect 1868 1056 1876 1064
rect 1869 1008 1875 1056
rect 1836 916 1844 924
rect 1869 848 1875 892
rect 1597 544 1603 552
rect 1596 536 1604 544
rect 1596 503 1604 504
rect 1592 497 1604 503
rect 1596 496 1604 497
rect 1452 283 1460 284
rect 1448 277 1460 283
rect 1452 276 1460 277
rect 1389 264 1395 272
rect 1388 256 1396 264
rect 1613 168 1619 352
rect 1661 348 1667 512
rect 1677 348 1683 652
rect 1885 368 1891 1012
rect 1901 963 1907 1152
rect 1917 1088 1923 1552
rect 1932 1436 1940 1444
rect 1933 1428 1939 1436
rect 1901 957 1923 963
rect 1917 688 1923 957
rect 1901 584 1907 612
rect 1900 576 1908 584
rect 1933 528 1939 1272
rect 1981 1088 1987 1752
rect 1949 1044 1955 1072
rect 1948 1036 1956 1044
rect 1997 708 2003 1332
rect 2029 1148 2035 1392
rect 2045 1208 2051 1812
rect 2106 1806 2112 1814
rect 2124 1483 2132 1484
rect 2120 1477 2132 1483
rect 2124 1476 2132 1477
rect 2106 1406 2112 1414
rect 2028 1116 2036 1124
rect 2029 1088 2035 1116
rect 2012 1076 2020 1084
rect 2013 1008 2019 1076
rect 1965 388 1971 552
rect 2045 488 2051 1152
rect 2061 928 2067 1392
rect 2125 1108 2131 1432
rect 2106 1006 2112 1014
rect 2141 1008 2147 1892
rect 2173 1528 2179 1892
rect 2349 1844 2355 1852
rect 2348 1836 2356 1844
rect 2157 1464 2163 1472
rect 2156 1456 2164 1464
rect 2106 606 2112 614
rect 2061 504 2067 592
rect 2125 508 2131 912
rect 2060 496 2068 504
rect 1660 256 1668 264
rect 1661 228 1667 256
rect 1805 128 1811 332
rect 1836 263 1844 264
rect 1832 257 1844 263
rect 1836 256 1844 257
rect 1292 116 1300 124
rect 1293 108 1299 116
rect 1740 123 1748 124
rect 1736 117 1748 123
rect 1740 116 1748 117
rect 1756 123 1764 124
rect 1756 117 1768 123
rect 1756 116 1764 117
rect 1837 124 1843 212
rect 1885 184 1891 272
rect 2061 208 2067 432
rect 2141 368 2147 672
rect 2189 588 2195 1792
rect 2349 1788 2355 1836
rect 2381 1588 2387 2012
rect 2492 1903 2500 1904
rect 2488 1897 2500 1903
rect 2492 1896 2500 1897
rect 2220 1356 2228 1364
rect 2221 1348 2227 1356
rect 2253 628 2259 1312
rect 2285 928 2291 1492
rect 2349 868 2355 1232
rect 2365 648 2371 912
rect 2156 576 2164 584
rect 2157 428 2163 576
rect 2381 508 2387 832
rect 2397 648 2403 1172
rect 2413 1028 2419 1112
rect 2412 876 2420 884
rect 2413 788 2419 876
rect 2429 788 2435 1732
rect 2509 1428 2515 1852
rect 2765 1384 2771 1872
rect 2973 1664 2979 1732
rect 2972 1656 2980 1664
rect 2764 1376 2772 1384
rect 2509 1028 2515 1372
rect 2493 568 2499 912
rect 2557 728 2563 1372
rect 2765 1368 2771 1376
rect 2653 1304 2659 1332
rect 2652 1296 2660 1304
rect 2781 1268 2787 1392
rect 2813 1324 2819 1472
rect 2829 1328 2835 1352
rect 2812 1316 2820 1324
rect 2877 1068 2883 1452
rect 2989 1064 2995 1092
rect 2988 1056 2996 1064
rect 2812 923 2820 924
rect 2808 917 2820 923
rect 2812 916 2820 917
rect 2600 897 2611 903
rect 2605 888 2611 897
rect 2588 883 2596 884
rect 2584 877 2596 883
rect 2588 876 2596 877
rect 2541 328 2547 592
rect 2106 206 2112 214
rect 1884 176 1892 184
rect 1885 148 1891 176
rect 2124 163 2132 164
rect 2120 157 2132 163
rect 2124 156 2132 157
rect 1852 136 1860 144
rect 1853 128 1859 136
rect 1836 116 1844 124
rect 2429 28 2435 292
rect 2541 148 2547 312
rect 2733 268 2739 712
rect 2749 688 2755 912
rect 2877 408 2883 1052
rect 3005 668 3011 1392
rect 3021 1068 3027 1692
rect 3069 568 3075 2112
rect 3101 544 3107 2132
rect 3100 536 3108 544
rect 3133 528 3139 752
rect 3069 308 3075 512
rect 2908 303 2916 304
rect 2904 297 2916 303
rect 2908 296 2916 297
rect 3149 128 3155 1752
rect 2764 103 2772 104
rect 2760 97 2772 103
rect 2764 96 2772 97
rect 1066 6 1072 14
use BUFX4  BUFX4_27
timestamp 1515334672
transform 1 0 8 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_41
timestamp 1515334672
transform 1 0 72 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_38
timestamp 1515334672
transform 1 0 168 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_43
timestamp 1515334672
transform 1 0 264 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_44
timestamp 1515334672
transform 1 0 360 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_39
timestamp 1515334672
transform -1 0 552 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_48
timestamp 1515334672
transform 1 0 552 0 -1 2210
box 0 0 96 200
use MUX2X1  MUX2X1_47
timestamp 1515334672
transform -1 0 744 0 -1 2210
box 0 0 96 200
use NOR2X1  NOR2X1_41
timestamp 1515334672
transform -1 0 792 0 -1 2210
box 0 0 48 200
use MUX2X1  MUX2X1_49
timestamp 1515334672
transform -1 0 888 0 -1 2210
box 0 0 96 200
use NOR2X1  NOR2X1_40
timestamp 1515334672
transform -1 0 936 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_86
timestamp 1515334672
transform 1 0 936 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_50
timestamp 1515334672
transform -1 0 1096 0 -1 2210
box 0 0 96 200
use FILL  FILL_10_0_0
timestamp 1515334672
transform 1 0 1096 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_0_1
timestamp 1515334672
transform 1 0 1112 0 -1 2210
box 0 0 16 200
use OAI21X1  OAI21X1_97
timestamp 1515334672
transform 1 0 1128 0 -1 2210
box 0 0 64 200
use NAND2X1  NAND2X1_64
timestamp 1515334672
transform 1 0 1192 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_98
timestamp 1515334672
transform 1 0 1240 0 -1 2210
box 0 0 64 200
use OAI22X1  OAI22X1_5
timestamp 1515334672
transform 1 0 1304 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_6
timestamp 1515334672
transform -1 0 1448 0 -1 2210
box 0 0 64 200
use INVX8  INVX8_2
timestamp 1515334672
transform -1 0 1528 0 -1 2210
box 0 0 80 200
use BUFX4  BUFX4_7
timestamp 1515334672
transform 1 0 1528 0 -1 2210
box 0 0 64 200
use MUX2X1  MUX2X1_40
timestamp 1515334672
transform -1 0 1688 0 -1 2210
box 0 0 96 200
use NAND3X1  NAND3X1_49
timestamp 1515334672
transform 1 0 1688 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_12
timestamp 1515334672
transform -1 0 1816 0 -1 2210
box 0 0 64 200
use BUFX4  BUFX4_11
timestamp 1515334672
transform 1 0 1816 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_45
timestamp 1515334672
transform -1 0 1928 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_54
timestamp 1515334672
transform 1 0 1928 0 -1 2210
box 0 0 64 200
use NOR2X1  NOR2X1_44
timestamp 1515334672
transform 1 0 1992 0 -1 2210
box 0 0 48 200
use OAI21X1  OAI21X1_63
timestamp 1515334672
transform 1 0 2040 0 -1 2210
box 0 0 64 200
use FILL  FILL_10_1_0
timestamp 1515334672
transform 1 0 2104 0 -1 2210
box 0 0 16 200
use FILL  FILL_10_1_1
timestamp 1515334672
transform 1 0 2120 0 -1 2210
box 0 0 16 200
use NOR3X1  NOR3X1_7
timestamp 1515334672
transform 1 0 2136 0 -1 2210
box 0 0 128 200
use OAI21X1  OAI21X1_62
timestamp 1515334672
transform 1 0 2264 0 -1 2210
box 0 0 64 200
use AND2X2  AND2X2_18
timestamp 1515334672
transform 1 0 2328 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_8
timestamp 1515334672
transform 1 0 2392 0 -1 2210
box 0 0 64 200
use OAI21X1  OAI21X1_69
timestamp 1515334672
transform -1 0 2520 0 -1 2210
box 0 0 64 200
use INVX2  INVX2_3
timestamp 1515334672
transform -1 0 2552 0 -1 2210
box 0 0 32 200
use NAND2X1  NAND2X1_5
timestamp 1515334672
transform -1 0 2600 0 -1 2210
box 0 0 48 200
use NAND3X1  NAND3X1_2
timestamp 1515334672
transform 1 0 2600 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_3
timestamp 1515334672
transform 1 0 2664 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_4
timestamp 1515334672
transform -1 0 2792 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_1
timestamp 1515334672
transform 1 0 2792 0 -1 2210
box 0 0 64 200
use INVX2  INVX2_2
timestamp 1515334672
transform 1 0 2856 0 -1 2210
box 0 0 32 200
use NAND3X1  NAND3X1_6
timestamp 1515334672
transform 1 0 2888 0 -1 2210
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1515334672
transform 1 0 2952 0 -1 2210
box 0 0 64 200
use INVX1  INVX1_3
timestamp 1515334672
transform -1 0 3048 0 -1 2210
box 0 0 32 200
use BUFX2  BUFX2_17
timestamp 1515334672
transform 1 0 3048 0 -1 2210
box 0 0 48 200
use AND2X2  AND2X2_10
timestamp 1515334672
transform 1 0 3096 0 -1 2210
box 0 0 64 200
use FILL  FILL_11_1
timestamp 1515334672
transform -1 0 3176 0 -1 2210
box 0 0 16 200
use FILL  FILL_11_2
timestamp 1515334672
transform -1 0 3192 0 -1 2210
box 0 0 16 200
use BUFX4  BUFX4_26
timestamp 1515334672
transform 1 0 8 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_42
timestamp 1515334672
transform 1 0 72 0 1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_46
timestamp 1515334672
transform 1 0 168 0 1 1810
box 0 0 96 200
use BUFX4  BUFX4_24
timestamp 1515334672
transform 1 0 264 0 1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_45
timestamp 1515334672
transform -1 0 424 0 1 1810
box 0 0 96 200
use INVX1  INVX1_29
timestamp 1515334672
transform 1 0 424 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_81
timestamp 1515334672
transform 1 0 456 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_58
timestamp 1515334672
transform 1 0 520 0 1 1810
box 0 0 48 200
use MUX2X1  MUX2X1_34
timestamp 1515334672
transform -1 0 664 0 1 1810
box 0 0 96 200
use OAI21X1  OAI21X1_82
timestamp 1515334672
transform 1 0 664 0 1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_59
timestamp 1515334672
transform -1 0 776 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_33
timestamp 1515334672
transform 1 0 776 0 1 1810
box 0 0 64 200
use OR2X2  OR2X2_2
timestamp 1515334672
transform -1 0 904 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_4
timestamp 1515334672
transform 1 0 904 0 1 1810
box 0 0 80 200
use NAND2X1  NAND2X1_61
timestamp 1515334672
transform -1 0 1032 0 1 1810
box 0 0 48 200
use FILL  FILL_9_0_0
timestamp 1515334672
transform 1 0 1032 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1515334672
transform 1 0 1048 0 1 1810
box 0 0 16 200
use OAI21X1  OAI21X1_87
timestamp 1515334672
transform 1 0 1064 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_7
timestamp 1515334672
transform 1 0 1128 0 1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_6
timestamp 1515334672
transform 1 0 1176 0 1 1810
box 0 0 80 200
use NAND3X1  NAND3X1_47
timestamp 1515334672
transform -1 0 1320 0 1 1810
box 0 0 64 200
use AOI21X1  AOI21X1_26
timestamp 1515334672
transform 1 0 1320 0 1 1810
box 0 0 64 200
use AOI22X1  AOI22X1_2
timestamp 1515334672
transform -1 0 1464 0 1 1810
box 0 0 80 200
use AOI21X1  AOI21X1_24
timestamp 1515334672
transform 1 0 1464 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_9
timestamp 1515334672
transform -1 0 1592 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_4
timestamp 1515334672
transform 1 0 1592 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_29
timestamp 1515334672
transform 1 0 1640 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_88
timestamp 1515334672
transform 1 0 1704 0 1 1810
box 0 0 64 200
use INVX2  INVX2_8
timestamp 1515334672
transform 1 0 1768 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_83
timestamp 1515334672
transform -1 0 1864 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_10
timestamp 1515334672
transform 1 0 1864 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_8
timestamp 1515334672
transform 1 0 1928 0 1 1810
box 0 0 48 200
use INVX2  INVX2_5
timestamp 1515334672
transform -1 0 2008 0 1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_68
timestamp 1515334672
transform -1 0 2072 0 1 1810
box 0 0 64 200
use FILL  FILL_9_1_0
timestamp 1515334672
transform 1 0 2072 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1515334672
transform 1 0 2088 0 1 1810
box 0 0 16 200
use INVX1  INVX1_15
timestamp 1515334672
transform 1 0 2104 0 1 1810
box 0 0 32 200
use INVX1  INVX1_24
timestamp 1515334672
transform -1 0 2168 0 1 1810
box 0 0 32 200
use AOI21X1  AOI21X1_6
timestamp 1515334672
transform -1 0 2232 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_22
timestamp 1515334672
transform 1 0 2232 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_61
timestamp 1515334672
transform -1 0 2360 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_23
timestamp 1515334672
transform 1 0 2360 0 1 1810
box 0 0 64 200
use NOR3X1  NOR3X1_4
timestamp 1515334672
transform -1 0 2552 0 1 1810
box 0 0 128 200
use BUFX4  BUFX4_39
timestamp 1515334672
transform -1 0 2616 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_1
timestamp 1515334672
transform 1 0 2616 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_2
timestamp 1515334672
transform 1 0 2680 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_101
timestamp 1515334672
transform -1 0 2808 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_72
timestamp 1515334672
transform 1 0 2808 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_71
timestamp 1515334672
transform 1 0 2872 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_70
timestamp 1515334672
transform 1 0 2936 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_100
timestamp 1515334672
transform -1 0 3064 0 1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_99
timestamp 1515334672
transform -1 0 3128 0 1 1810
box 0 0 64 200
use AND2X2  AND2X2_27
timestamp 1515334672
transform -1 0 3192 0 1 1810
box 0 0 64 200
use BUFX4  BUFX4_17
timestamp 1515334672
transform 1 0 8 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_35
timestamp 1515334672
transform -1 0 168 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_36
timestamp 1515334672
transform -1 0 264 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_32
timestamp 1515334672
transform -1 0 360 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_26
timestamp 1515334672
transform -1 0 456 0 -1 1810
box 0 0 96 200
use BUFX4  BUFX4_16
timestamp 1515334672
transform -1 0 520 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_33
timestamp 1515334672
transform -1 0 616 0 -1 1810
box 0 0 96 200
use MUX2X1  MUX2X1_30
timestamp 1515334672
transform -1 0 712 0 -1 1810
box 0 0 96 200
use NAND2X1  NAND2X1_26
timestamp 1515334672
transform 1 0 712 0 -1 1810
box 0 0 48 200
use INVX2  INVX2_1
timestamp 1515334672
transform 1 0 760 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_43
timestamp 1515334672
transform 1 0 792 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_52
timestamp 1515334672
transform 1 0 856 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_53
timestamp 1515334672
transform 1 0 920 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_44
timestamp 1515334672
transform -1 0 1048 0 -1 1810
box 0 0 64 200
use FILL  FILL_8_0_0
timestamp 1515334672
transform -1 0 1064 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1515334672
transform -1 0 1080 0 -1 1810
box 0 0 16 200
use NAND2X1  NAND2X1_48
timestamp 1515334672
transform -1 0 1128 0 -1 1810
box 0 0 48 200
use AOI22X1  AOI22X1_5
timestamp 1515334672
transform -1 0 1208 0 -1 1810
box 0 0 80 200
use NOR2X1  NOR2X1_11
timestamp 1515334672
transform -1 0 1256 0 -1 1810
box 0 0 48 200
use NAND2X1  NAND2X1_54
timestamp 1515334672
transform 1 0 1256 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_74
timestamp 1515334672
transform -1 0 1368 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_6
timestamp 1515334672
transform 1 0 1368 0 -1 1810
box 0 0 64 200
use MUX2X1  MUX2X1_37
timestamp 1515334672
transform -1 0 1528 0 -1 1810
box 0 0 96 200
use NAND3X1  NAND3X1_30
timestamp 1515334672
transform 1 0 1528 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_19
timestamp 1515334672
transform -1 0 1656 0 -1 1810
box 0 0 64 200
use NAND3X1  NAND3X1_34
timestamp 1515334672
transform 1 0 1656 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_39
timestamp 1515334672
transform 1 0 1720 0 -1 1810
box 0 0 48 200
use NAND3X1  NAND3X1_8
timestamp 1515334672
transform -1 0 1832 0 -1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_38
timestamp 1515334672
transform 1 0 1832 0 -1 1810
box 0 0 48 200
use OAI21X1  OAI21X1_45
timestamp 1515334672
transform 1 0 1880 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_42
timestamp 1515334672
transform 1 0 1944 0 -1 1810
box 0 0 64 200
use INVX2  INVX2_7
timestamp 1515334672
transform -1 0 2040 0 -1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_6
timestamp 1515334672
transform 1 0 2040 0 -1 1810
box 0 0 48 200
use FILL  FILL_8_1_0
timestamp 1515334672
transform -1 0 2104 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1515334672
transform -1 0 2120 0 -1 1810
box 0 0 16 200
use NOR2X1  NOR2X1_32
timestamp 1515334672
transform -1 0 2168 0 -1 1810
box 0 0 48 200
use INVX8  INVX8_1
timestamp 1515334672
transform 1 0 2168 0 -1 1810
box 0 0 80 200
use OAI21X1  OAI21X1_79
timestamp 1515334672
transform 1 0 2248 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_12
timestamp 1515334672
transform -1 0 2344 0 -1 1810
box 0 0 32 200
use OAI21X1  OAI21X1_85
timestamp 1515334672
transform 1 0 2344 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_78
timestamp 1515334672
transform -1 0 2472 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_84
timestamp 1515334672
transform 1 0 2472 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_22
timestamp 1515334672
transform -1 0 2600 0 -1 1810
box 0 0 64 200
use AND2X2  AND2X2_3
timestamp 1515334672
transform 1 0 2600 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_32
timestamp 1515334672
transform -1 0 2696 0 -1 1810
box 0 0 32 200
use NAND3X1  NAND3X1_7
timestamp 1515334672
transform 1 0 2696 0 -1 1810
box 0 0 64 200
use NAND2X1  NAND2X1_50
timestamp 1515334672
transform 1 0 2760 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_26
timestamp 1515334672
transform -1 0 2840 0 -1 1810
box 0 0 32 200
use BUFX4  BUFX4_21
timestamp 1515334672
transform 1 0 2840 0 -1 1810
box 0 0 64 200
use BUFX4  BUFX4_38
timestamp 1515334672
transform 1 0 2904 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_76
timestamp 1515334672
transform 1 0 2968 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_75
timestamp 1515334672
transform -1 0 3096 0 -1 1810
box 0 0 64 200
use INVX1  INVX1_27
timestamp 1515334672
transform 1 0 3096 0 -1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_36
timestamp 1515334672
transform 1 0 3128 0 -1 1810
box 0 0 48 200
use FILL  FILL_9_1
timestamp 1515334672
transform -1 0 3192 0 -1 1810
box 0 0 16 200
use BUFX4  BUFX4_18
timestamp 1515334672
transform 1 0 8 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_10
timestamp 1515334672
transform 1 0 72 0 1 1410
box 0 0 96 200
use NAND2X1  NAND2X1_2
timestamp 1515334672
transform -1 0 216 0 1 1410
box 0 0 48 200
use MUX2X1  MUX2X1_31
timestamp 1515334672
transform -1 0 312 0 1 1410
box 0 0 96 200
use MUX2X1  MUX2X1_25
timestamp 1515334672
transform 1 0 312 0 1 1410
box 0 0 96 200
use INVX1  INVX1_9
timestamp 1515334672
transform -1 0 440 0 1 1410
box 0 0 32 200
use BUFX4  BUFX4_13
timestamp 1515334672
transform 1 0 440 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_29
timestamp 1515334672
transform 1 0 504 0 1 1410
box 0 0 96 200
use AOI21X1  AOI21X1_3
timestamp 1515334672
transform 1 0 600 0 1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_22
timestamp 1515334672
transform 1 0 664 0 1 1410
box 0 0 96 200
use BUFX4  BUFX4_14
timestamp 1515334672
transform 1 0 760 0 1 1410
box 0 0 64 200
use NOR3X1  NOR3X1_1
timestamp 1515334672
transform 1 0 824 0 1 1410
box 0 0 128 200
use AOI22X1  AOI22X1_9
timestamp 1515334672
transform 1 0 952 0 1 1410
box 0 0 80 200
use FILL  FILL_7_0_0
timestamp 1515334672
transform 1 0 1032 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1515334672
transform 1 0 1048 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_93
timestamp 1515334672
transform 1 0 1064 0 1 1410
box 0 0 64 200
use INVX1  INVX1_31
timestamp 1515334672
transform -1 0 1160 0 1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_3
timestamp 1515334672
transform -1 0 1208 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_28
timestamp 1515334672
transform -1 0 1256 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_2
timestamp 1515334672
transform 1 0 1256 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_5
timestamp 1515334672
transform -1 0 1384 0 1 1410
box 0 0 64 200
use INVX1  INVX1_1
timestamp 1515334672
transform 1 0 1384 0 1 1410
box 0 0 32 200
use NOR2X1  NOR2X1_1
timestamp 1515334672
transform 1 0 1416 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_94
timestamp 1515334672
transform -1 0 1528 0 1 1410
box 0 0 64 200
use BUFX4  BUFX4_8
timestamp 1515334672
transform 1 0 1528 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_13
timestamp 1515334672
transform 1 0 1592 0 1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1515334672
transform 1 0 1656 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_62
timestamp 1515334672
transform -1 0 1768 0 1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_55
timestamp 1515334672
transform -1 0 1816 0 1 1410
box 0 0 48 200
use XNOR2X1  XNOR2X1_2
timestamp 1515334672
transform 1 0 1816 0 1 1410
box 0 0 112 200
use NOR2X1  NOR2X1_22
timestamp 1515334672
transform 1 0 1928 0 1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_28
timestamp 1515334672
transform -1 0 2024 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_35
timestamp 1515334672
transform 1 0 2024 0 1 1410
box 0 0 64 200
use FILL  FILL_7_1_0
timestamp 1515334672
transform 1 0 2088 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1515334672
transform 1 0 2104 0 1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_102
timestamp 1515334672
transform 1 0 2120 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_12
timestamp 1515334672
transform -1 0 2248 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_41
timestamp 1515334672
transform -1 0 2312 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_19
timestamp 1515334672
transform 1 0 2312 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_31
timestamp 1515334672
transform -1 0 2424 0 1 1410
box 0 0 48 200
use XNOR2X1  XNOR2X1_10
timestamp 1515334672
transform 1 0 2424 0 1 1410
box 0 0 112 200
use BUFX4  BUFX4_36
timestamp 1515334672
transform -1 0 2600 0 1 1410
box 0 0 64 200
use NAND2X1  NAND2X1_51
timestamp 1515334672
transform 1 0 2600 0 1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_27
timestamp 1515334672
transform -1 0 2712 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_73
timestamp 1515334672
transform -1 0 2776 0 1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_35
timestamp 1515334672
transform 1 0 2776 0 1 1410
box 0 0 48 200
use OAI21X1  OAI21X1_66
timestamp 1515334672
transform 1 0 2824 0 1 1410
box 0 0 64 200
use AND2X2  AND2X2_20
timestamp 1515334672
transform 1 0 2888 0 1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_65
timestamp 1515334672
transform -1 0 3016 0 1 1410
box 0 0 64 200
use XNOR2X1  XNOR2X1_8
timestamp 1515334672
transform -1 0 3128 0 1 1410
box 0 0 112 200
use BUFX2  BUFX2_13
timestamp 1515334672
transform 1 0 3128 0 1 1410
box 0 0 48 200
use FILL  FILL_8_1
timestamp 1515334672
transform 1 0 3176 0 1 1410
box 0 0 16 200
use MUX2X1  MUX2X1_9
timestamp 1515334672
transform -1 0 104 0 -1 1410
box 0 0 96 200
use INVX1  INVX1_8
timestamp 1515334672
transform -1 0 136 0 -1 1410
box 0 0 32 200
use OAI21X1  OAI21X1_5
timestamp 1515334672
transform -1 0 200 0 -1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_18
timestamp 1515334672
transform 1 0 200 0 -1 1410
box 0 0 96 200
use INVX1  INVX1_10
timestamp 1515334672
transform 1 0 296 0 -1 1410
box 0 0 32 200
use NAND2X1  NAND2X1_3
timestamp 1515334672
transform -1 0 376 0 -1 1410
box 0 0 48 200
use MUX2X1  MUX2X1_19
timestamp 1515334672
transform 1 0 376 0 -1 1410
box 0 0 96 200
use MUX2X1  MUX2X1_15
timestamp 1515334672
transform -1 0 568 0 -1 1410
box 0 0 96 200
use NAND2X1  NAND2X1_6
timestamp 1515334672
transform -1 0 616 0 -1 1410
box 0 0 48 200
use AOI22X1  AOI22X1_1
timestamp 1515334672
transform 1 0 616 0 -1 1410
box 0 0 80 200
use BUFX4  BUFX4_40
timestamp 1515334672
transform 1 0 696 0 -1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_5
timestamp 1515334672
transform 1 0 760 0 -1 1410
box 0 0 96 200
use MUX2X1  MUX2X1_6
timestamp 1515334672
transform 1 0 856 0 -1 1410
box 0 0 96 200
use MUX2X1  MUX2X1_16
timestamp 1515334672
transform -1 0 1048 0 -1 1410
box 0 0 96 200
use FILL  FILL_6_0_0
timestamp 1515334672
transform -1 0 1064 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1515334672
transform -1 0 1080 0 -1 1410
box 0 0 16 200
use MUX2X1  MUX2X1_3
timestamp 1515334672
transform -1 0 1176 0 -1 1410
box 0 0 96 200
use AOI21X1  AOI21X1_32
timestamp 1515334672
transform -1 0 1240 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_30
timestamp 1515334672
transform 1 0 1240 0 -1 1410
box 0 0 48 200
use NAND2X1  NAND2X1_45
timestamp 1515334672
transform -1 0 1336 0 -1 1410
box 0 0 48 200
use MUX2X1  MUX2X1_2
timestamp 1515334672
transform -1 0 1432 0 -1 1410
box 0 0 96 200
use NAND3X1  NAND3X1_10
timestamp 1515334672
transform -1 0 1496 0 -1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_14
timestamp 1515334672
transform -1 0 1592 0 -1 1410
box 0 0 96 200
use NAND3X1  NAND3X1_31
timestamp 1515334672
transform 1 0 1592 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_30
timestamp 1515334672
transform 1 0 1656 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_16
timestamp 1515334672
transform 1 0 1720 0 -1 1410
box 0 0 32 200
use NAND3X1  NAND3X1_20
timestamp 1515334672
transform -1 0 1816 0 -1 1410
box 0 0 64 200
use OR2X2  OR2X2_3
timestamp 1515334672
transform 1 0 1816 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_22
timestamp 1515334672
transform 1 0 1880 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_8
timestamp 1515334672
transform 1 0 1944 0 -1 1410
box 0 0 64 200
use NOR2X1  NOR2X1_43
timestamp 1515334672
transform -1 0 2056 0 -1 1410
box 0 0 48 200
use NOR2X1  NOR2X1_12
timestamp 1515334672
transform 1 0 2056 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_1_0
timestamp 1515334672
transform -1 0 2120 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1515334672
transform -1 0 2136 0 -1 1410
box 0 0 16 200
use OAI21X1  OAI21X1_21
timestamp 1515334672
transform -1 0 2200 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_29
timestamp 1515334672
transform -1 0 2264 0 -1 1410
box 0 0 64 200
use NAND3X1  NAND3X1_51
timestamp 1515334672
transform 1 0 2264 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_64
timestamp 1515334672
transform -1 0 2392 0 -1 1410
box 0 0 64 200
use AOI22X1  AOI22X1_8
timestamp 1515334672
transform -1 0 2472 0 -1 1410
box 0 0 80 200
use BUFX4  BUFX4_19
timestamp 1515334672
transform -1 0 2536 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_89
timestamp 1515334672
transform 1 0 2536 0 -1 1410
box 0 0 64 200
use OAI21X1  OAI21X1_90
timestamp 1515334672
transform -1 0 2664 0 -1 1410
box 0 0 64 200
use AND2X2  AND2X2_24
timestamp 1515334672
transform 1 0 2664 0 -1 1410
box 0 0 64 200
use INVX1  INVX1_2
timestamp 1515334672
transform 1 0 2728 0 -1 1410
box 0 0 32 200
use INVX1  INVX1_25
timestamp 1515334672
transform 1 0 2760 0 -1 1410
box 0 0 32 200
use INVX4  INVX4_1
timestamp 1515334672
transform -1 0 2840 0 -1 1410
box 0 0 48 200
use BUFX4  BUFX4_35
timestamp 1515334672
transform 1 0 2840 0 -1 1410
box 0 0 64 200
use BUFX4  BUFX4_34
timestamp 1515334672
transform 1 0 2904 0 -1 1410
box 0 0 64 200
use XNOR2X1  XNOR2X1_7
timestamp 1515334672
transform 1 0 2968 0 -1 1410
box 0 0 112 200
use XNOR2X1  XNOR2X1_12
timestamp 1515334672
transform -1 0 3192 0 -1 1410
box 0 0 112 200
use INVX8  INVX8_3
timestamp 1515334672
transform -1 0 88 0 1 1010
box 0 0 80 200
use BUFX4  BUFX4_15
timestamp 1515334672
transform 1 0 88 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_23
timestamp 1515334672
transform 1 0 152 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_10
timestamp 1515334672
transform -1 0 280 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_6
timestamp 1515334672
transform 1 0 280 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_25
timestamp 1515334672
transform 1 0 344 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_41
timestamp 1515334672
transform 1 0 408 0 1 1010
box 0 0 64 200
use OR2X2  OR2X2_1
timestamp 1515334672
transform 1 0 472 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_44
timestamp 1515334672
transform 1 0 536 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_20
timestamp 1515334672
transform -1 0 648 0 1 1010
box 0 0 48 200
use NOR2X1  NOR2X1_21
timestamp 1515334672
transform -1 0 696 0 1 1010
box 0 0 48 200
use MUX2X1  MUX2X1_12
timestamp 1515334672
transform 1 0 696 0 1 1010
box 0 0 96 200
use OAI22X1  OAI22X1_1
timestamp 1515334672
transform 1 0 792 0 1 1010
box 0 0 80 200
use NOR2X1  NOR2X1_24
timestamp 1515334672
transform 1 0 872 0 1 1010
box 0 0 48 200
use MUX2X1  MUX2X1_27
timestamp 1515334672
transform 1 0 920 0 1 1010
box 0 0 96 200
use FILL  FILL_5_0_0
timestamp 1515334672
transform 1 0 1016 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1515334672
transform 1 0 1032 0 1 1010
box 0 0 16 200
use MUX2X1  MUX2X1_11
timestamp 1515334672
transform 1 0 1048 0 1 1010
box 0 0 96 200
use NOR2X1  NOR2X1_16
timestamp 1515334672
transform 1 0 1144 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_22
timestamp 1515334672
transform 1 0 1192 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_10
timestamp 1515334672
transform -1 0 1320 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_11
timestamp 1515334672
transform -1 0 1384 0 1 1010
box 0 0 64 200
use MUX2X1  MUX2X1_13
timestamp 1515334672
transform -1 0 1480 0 1 1010
box 0 0 96 200
use OAI21X1  OAI21X1_17
timestamp 1515334672
transform 1 0 1480 0 1 1010
box 0 0 64 200
use MUX2X1  MUX2X1_21
timestamp 1515334672
transform -1 0 1640 0 1 1010
box 0 0 96 200
use AOI21X1  AOI21X1_4
timestamp 1515334672
transform 1 0 1640 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_33
timestamp 1515334672
transform -1 0 1752 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_16
timestamp 1515334672
transform 1 0 1752 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_7
timestamp 1515334672
transform 1 0 1800 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_40
timestamp 1515334672
transform -1 0 1912 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_14
timestamp 1515334672
transform -1 0 1976 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_38
timestamp 1515334672
transform 1 0 1976 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_37
timestamp 1515334672
transform -1 0 2072 0 1 1010
box 0 0 48 200
use FILL  FILL_5_1_0
timestamp 1515334672
transform -1 0 2088 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1515334672
transform -1 0 2104 0 1 1010
box 0 0 16 200
use NAND3X1  NAND3X1_50
timestamp 1515334672
transform -1 0 2168 0 1 1010
box 0 0 64 200
use INVX4  INVX4_2
timestamp 1515334672
transform 1 0 2168 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_80
timestamp 1515334672
transform 1 0 2216 0 1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_5
timestamp 1515334672
transform 1 0 2280 0 1 1010
box 0 0 128 200
use NOR2X1  NOR2X1_34
timestamp 1515334672
transform -1 0 2456 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_91
timestamp 1515334672
transform 1 0 2456 0 1 1010
box 0 0 64 200
use BUFX4  BUFX4_37
timestamp 1515334672
transform -1 0 2584 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_37
timestamp 1515334672
transform 1 0 2584 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_77
timestamp 1515334672
transform 1 0 2632 0 1 1010
box 0 0 64 200
use AND2X2  AND2X2_25
timestamp 1515334672
transform 1 0 2696 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_42
timestamp 1515334672
transform -1 0 2808 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_67
timestamp 1515334672
transform 1 0 2808 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_1
timestamp 1515334672
transform -1 0 2936 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_33
timestamp 1515334672
transform -1 0 2984 0 1 1010
box 0 0 48 200
use AOI22X1  AOI22X1_3
timestamp 1515334672
transform -1 0 3064 0 1 1010
box 0 0 80 200
use NAND2X1  NAND2X1_56
timestamp 1515334672
transform 1 0 3064 0 1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_65
timestamp 1515334672
transform -1 0 3160 0 1 1010
box 0 0 48 200
use INVX1  INVX1_28
timestamp 1515334672
transform -1 0 3192 0 1 1010
box 0 0 32 200
use MUX2X1  MUX2X1_17
timestamp 1515334672
transform -1 0 104 0 -1 1010
box 0 0 96 200
use MUX2X1  MUX2X1_23
timestamp 1515334672
transform 1 0 104 0 -1 1010
box 0 0 96 200
use NAND2X1  NAND2X1_7
timestamp 1515334672
transform -1 0 248 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_19
timestamp 1515334672
transform 1 0 248 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_10
timestamp 1515334672
transform -1 0 360 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_20
timestamp 1515334672
transform 1 0 360 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_28
timestamp 1515334672
transform 1 0 424 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_14
timestamp 1515334672
transform -1 0 536 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_42
timestamp 1515334672
transform 1 0 536 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_5
timestamp 1515334672
transform -1 0 664 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_25
timestamp 1515334672
transform -1 0 712 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_40
timestamp 1515334672
transform -1 0 776 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1515334672
transform -1 0 840 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_17
timestamp 1515334672
transform 1 0 840 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_8
timestamp 1515334672
transform -1 0 968 0 -1 1010
box 0 0 64 200
use MUX2X1  MUX2X1_20
timestamp 1515334672
transform -1 0 1064 0 -1 1010
box 0 0 96 200
use FILL  FILL_4_0_0
timestamp 1515334672
transform 1 0 1064 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1515334672
transform 1 0 1080 0 -1 1010
box 0 0 16 200
use MUX2X1  MUX2X1_24
timestamp 1515334672
transform 1 0 1096 0 -1 1010
box 0 0 96 200
use INVX2  INVX2_6
timestamp 1515334672
transform -1 0 1224 0 -1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_24
timestamp 1515334672
transform 1 0 1224 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_25
timestamp 1515334672
transform 1 0 1288 0 -1 1010
box 0 0 64 200
use NOR3X1  NOR3X1_2
timestamp 1515334672
transform -1 0 1480 0 -1 1010
box 0 0 128 200
use AOI21X1  AOI21X1_20
timestamp 1515334672
transform 1 0 1480 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_27
timestamp 1515334672
transform 1 0 1544 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_9
timestamp 1515334672
transform -1 0 1656 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_24
timestamp 1515334672
transform -1 0 1704 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_35
timestamp 1515334672
transform 1 0 1704 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_25
timestamp 1515334672
transform -1 0 1832 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_36
timestamp 1515334672
transform 1 0 1832 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_49
timestamp 1515334672
transform 1 0 1896 0 -1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_41
timestamp 1515334672
transform -1 0 2008 0 -1 1010
box 0 0 48 200
use NAND2X1  NAND2X1_63
timestamp 1515334672
transform -1 0 2056 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_1_0
timestamp 1515334672
transform 1 0 2056 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1515334672
transform 1 0 2072 0 -1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_23
timestamp 1515334672
transform 1 0 2088 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_18
timestamp 1515334672
transform 1 0 2152 0 -1 1010
box 0 0 32 200
use NAND3X1  NAND3X1_46
timestamp 1515334672
transform 1 0 2184 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_46
timestamp 1515334672
transform -1 0 2312 0 -1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_23
timestamp 1515334672
transform -1 0 2360 0 -1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_30
timestamp 1515334672
transform 1 0 2360 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_13
timestamp 1515334672
transform 1 0 2424 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_31
timestamp 1515334672
transform 1 0 2488 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_48
timestamp 1515334672
transform 1 0 2552 0 -1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_28
timestamp 1515334672
transform 1 0 2616 0 -1 1010
box 0 0 64 200
use BUFX4  BUFX4_29
timestamp 1515334672
transform -1 0 2744 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_92
timestamp 1515334672
transform -1 0 2808 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_52
timestamp 1515334672
transform 1 0 2808 0 -1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_1
timestamp 1515334672
transform -1 0 2936 0 -1 1010
box 0 0 64 200
use AND2X2  AND2X2_21
timestamp 1515334672
transform 1 0 2936 0 -1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_13
timestamp 1515334672
transform 1 0 3000 0 -1 1010
box 0 0 80 200
use AND2X2  AND2X2_28
timestamp 1515334672
transform 1 0 3080 0 -1 1010
box 0 0 64 200
use BUFX2  BUFX2_11
timestamp 1515334672
transform 1 0 3144 0 -1 1010
box 0 0 48 200
use BUFX4  BUFX4_43
timestamp 1515334672
transform 1 0 8 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_16
timestamp 1515334672
transform 1 0 72 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_13
timestamp 1515334672
transform 1 0 136 0 1 610
box 0 0 48 200
use INVX1  INVX1_13
timestamp 1515334672
transform -1 0 216 0 1 610
box 0 0 32 200
use AOI21X1  AOI21X1_11
timestamp 1515334672
transform 1 0 216 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_33
timestamp 1515334672
transform -1 0 344 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_27
timestamp 1515334672
transform 1 0 344 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_4
timestamp 1515334672
transform 1 0 408 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_9
timestamp 1515334672
transform 1 0 472 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_2
timestamp 1515334672
transform 1 0 520 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_18
timestamp 1515334672
transform 1 0 584 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_11
timestamp 1515334672
transform 1 0 648 0 1 610
box 0 0 64 200
use XNOR2X1  XNOR2X1_3
timestamp 1515334672
transform 1 0 712 0 1 610
box 0 0 112 200
use INVX1  INVX1_6
timestamp 1515334672
transform -1 0 856 0 1 610
box 0 0 32 200
use MUX2X1  MUX2X1_1
timestamp 1515334672
transform -1 0 952 0 1 610
box 0 0 96 200
use NOR2X1  NOR2X1_17
timestamp 1515334672
transform -1 0 1000 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_34
timestamp 1515334672
transform -1 0 1064 0 1 610
box 0 0 64 200
use FILL  FILL_3_0_0
timestamp 1515334672
transform 1 0 1064 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1515334672
transform 1 0 1080 0 1 610
box 0 0 16 200
use NAND2X1  NAND2X1_1
timestamp 1515334672
transform 1 0 1096 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_46
timestamp 1515334672
transform -1 0 1192 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_47
timestamp 1515334672
transform 1 0 1192 0 1 610
box 0 0 48 200
use NAND2X1  NAND2X1_21
timestamp 1515334672
transform 1 0 1240 0 1 610
box 0 0 48 200
use OR2X2  OR2X2_4
timestamp 1515334672
transform 1 0 1288 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_60
timestamp 1515334672
transform 1 0 1352 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_20
timestamp 1515334672
transform 1 0 1416 0 1 610
box 0 0 48 200
use NOR2X1  NOR2X1_13
timestamp 1515334672
transform 1 0 1464 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_15
timestamp 1515334672
transform 1 0 1512 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_42
timestamp 1515334672
transform -1 0 1640 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_12
timestamp 1515334672
transform 1 0 1640 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_53
timestamp 1515334672
transform -1 0 1752 0 1 610
box 0 0 48 200
use INVX1  INVX1_21
timestamp 1515334672
transform 1 0 1752 0 1 610
box 0 0 32 200
use OAI21X1  OAI21X1_54
timestamp 1515334672
transform 1 0 1784 0 1 610
box 0 0 64 200
use AND2X2  AND2X2_15
timestamp 1515334672
transform -1 0 1912 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_34
timestamp 1515334672
transform 1 0 1912 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_53
timestamp 1515334672
transform -1 0 2040 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_29
timestamp 1515334672
transform -1 0 2088 0 1 610
box 0 0 48 200
use FILL  FILL_3_1_0
timestamp 1515334672
transform -1 0 2104 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1515334672
transform -1 0 2120 0 1 610
box 0 0 16 200
use NOR2X1  NOR2X1_18
timestamp 1515334672
transform -1 0 2168 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_38
timestamp 1515334672
transform 1 0 2168 0 1 610
box 0 0 64 200
use NAND2X1  NAND2X1_34
timestamp 1515334672
transform -1 0 2280 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_35
timestamp 1515334672
transform 1 0 2280 0 1 610
box 0 0 64 200
use AOI22X1  AOI22X1_7
timestamp 1515334672
transform -1 0 2424 0 1 610
box 0 0 80 200
use XNOR2X1  XNOR2X1_9
timestamp 1515334672
transform 1 0 2424 0 1 610
box 0 0 112 200
use BUFX4  BUFX4_20
timestamp 1515334672
transform -1 0 2600 0 1 610
box 0 0 64 200
use XNOR2X1  XNOR2X1_5
timestamp 1515334672
transform 1 0 2600 0 1 610
box 0 0 112 200
use BUFX4  BUFX4_30
timestamp 1515334672
transform -1 0 2776 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_33
timestamp 1515334672
transform -1 0 2840 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_32
timestamp 1515334672
transform -1 0 2904 0 1 610
box 0 0 64 200
use BUFX4  BUFX4_31
timestamp 1515334672
transform 1 0 2904 0 1 610
box 0 0 64 200
use NOR3X1  NOR3X1_9
timestamp 1515334672
transform 1 0 2968 0 1 610
box 0 0 128 200
use BUFX2  BUFX2_9
timestamp 1515334672
transform 1 0 3096 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_14
timestamp 1515334672
transform 1 0 3144 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_4
timestamp 1515334672
transform -1 0 72 0 -1 610
box 0 0 64 200
use BUFX4  BUFX4_3
timestamp 1515334672
transform -1 0 136 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_12
timestamp 1515334672
transform 1 0 136 0 -1 610
box 0 0 48 200
use INVX1  INVX1_17
timestamp 1515334672
transform 1 0 184 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_15
timestamp 1515334672
transform 1 0 216 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_14
timestamp 1515334672
transform 1 0 280 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_33
timestamp 1515334672
transform -1 0 408 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_3
timestamp 1515334672
transform -1 0 472 0 -1 610
box 0 0 64 200
use MUX2X1  MUX2X1_28
timestamp 1515334672
transform -1 0 568 0 -1 610
box 0 0 96 200
use NAND2X1  NAND2X1_17
timestamp 1515334672
transform -1 0 616 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_4
timestamp 1515334672
transform 1 0 616 0 -1 610
box 0 0 64 200
use XNOR2X1  XNOR2X1_1
timestamp 1515334672
transform 1 0 680 0 -1 610
box 0 0 112 200
use AOI21X1  AOI21X1_21
timestamp 1515334672
transform 1 0 792 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_44
timestamp 1515334672
transform 1 0 856 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_29
timestamp 1515334672
transform -1 0 968 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_30
timestamp 1515334672
transform 1 0 968 0 -1 610
box 0 0 48 200
use FILL  FILL_2_0_0
timestamp 1515334672
transform 1 0 1016 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1515334672
transform 1 0 1032 0 -1 610
box 0 0 16 200
use MUX2X1  MUX2X1_7
timestamp 1515334672
transform 1 0 1048 0 -1 610
box 0 0 96 200
use INVX1  INVX1_7
timestamp 1515334672
transform -1 0 1176 0 -1 610
box 0 0 32 200
use OAI22X1  OAI22X1_3
timestamp 1515334672
transform -1 0 1256 0 -1 610
box 0 0 80 200
use INVX1  INVX1_5
timestamp 1515334672
transform 1 0 1256 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_23
timestamp 1515334672
transform -1 0 1352 0 -1 610
box 0 0 64 200
use NAND2X1  NAND2X1_52
timestamp 1515334672
transform -1 0 1400 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_27
timestamp 1515334672
transform -1 0 1448 0 -1 610
box 0 0 48 200
use INVX1  INVX1_4
timestamp 1515334672
transform -1 0 1480 0 -1 610
box 0 0 32 200
use MUX2X1  MUX2X1_4
timestamp 1515334672
transform 1 0 1480 0 -1 610
box 0 0 96 200
use MUX2X1  MUX2X1_8
timestamp 1515334672
transform -1 0 1672 0 -1 610
box 0 0 96 200
use NAND2X1  NAND2X1_57
timestamp 1515334672
transform -1 0 1720 0 -1 610
box 0 0 48 200
use NOR3X1  NOR3X1_3
timestamp 1515334672
transform -1 0 1848 0 -1 610
box 0 0 128 200
use NOR2X1  NOR2X1_5
timestamp 1515334672
transform 1 0 1848 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_41
timestamp 1515334672
transform -1 0 1960 0 -1 610
box 0 0 64 200
use NOR3X1  NOR3X1_6
timestamp 1515334672
transform -1 0 2088 0 -1 610
box 0 0 128 200
use FILL  FILL_2_1_0
timestamp 1515334672
transform -1 0 2104 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1515334672
transform -1 0 2120 0 -1 610
box 0 0 16 200
use NAND2X1  NAND2X1_60
timestamp 1515334672
transform -1 0 2168 0 -1 610
box 0 0 48 200
use INVX1  INVX1_11
timestamp 1515334672
transform -1 0 2200 0 -1 610
box 0 0 32 200
use NAND2X1  NAND2X1_49
timestamp 1515334672
transform 1 0 2200 0 -1 610
box 0 0 48 200
use INVX1  INVX1_30
timestamp 1515334672
transform 1 0 2248 0 -1 610
box 0 0 32 200
use NAND3X1  NAND3X1_36
timestamp 1515334672
transform 1 0 2280 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_96
timestamp 1515334672
transform 1 0 2344 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_26
timestamp 1515334672
transform 1 0 2408 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_95
timestamp 1515334672
transform -1 0 2536 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_10
timestamp 1515334672
transform -1 0 2616 0 -1 610
box 0 0 80 200
use XNOR2X1  XNOR2X1_11
timestamp 1515334672
transform 1 0 2616 0 -1 610
box 0 0 112 200
use XNOR2X1  XNOR2X1_4
timestamp 1515334672
transform 1 0 2728 0 -1 610
box 0 0 112 200
use NAND2X1  NAND2X1_18
timestamp 1515334672
transform 1 0 2840 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_19
timestamp 1515334672
transform 1 0 2888 0 -1 610
box 0 0 48 200
use BUFX4  BUFX4_28
timestamp 1515334672
transform -1 0 3000 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_57
timestamp 1515334672
transform -1 0 3064 0 -1 610
box 0 0 64 200
use AOI22X1  AOI22X1_12
timestamp 1515334672
transform -1 0 3144 0 -1 610
box 0 0 80 200
use BUFX2  BUFX2_16
timestamp 1515334672
transform 1 0 3144 0 -1 610
box 0 0 48 200
use OAI22X1  OAI22X1_2
timestamp 1515334672
transform 1 0 8 0 1 210
box 0 0 80 200
use OAI21X1  OAI21X1_7
timestamp 1515334672
transform 1 0 88 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_4
timestamp 1515334672
transform -1 0 200 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_31
timestamp 1515334672
transform 1 0 200 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_11
timestamp 1515334672
transform 1 0 264 0 1 210
box 0 0 64 200
use OAI22X1  OAI22X1_4
timestamp 1515334672
transform 1 0 328 0 1 210
box 0 0 80 200
use NAND2X1  NAND2X1_32
timestamp 1515334672
transform -1 0 456 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_45
timestamp 1515334672
transform -1 0 520 0 1 210
box 0 0 64 200
use BUFX4  BUFX4_2
timestamp 1515334672
transform 1 0 520 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_14
timestamp 1515334672
transform 1 0 584 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_26
timestamp 1515334672
transform -1 0 696 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_27
timestamp 1515334672
transform -1 0 760 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_28
timestamp 1515334672
transform -1 0 824 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_23
timestamp 1515334672
transform -1 0 872 0 1 210
box 0 0 48 200
use AOI21X1  AOI21X1_18
timestamp 1515334672
transform 1 0 872 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_36
timestamp 1515334672
transform -1 0 984 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_32
timestamp 1515334672
transform 1 0 984 0 1 210
box 0 0 64 200
use FILL  FILL_1_0_0
timestamp 1515334672
transform 1 0 1048 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1515334672
transform 1 0 1064 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_10
timestamp 1515334672
transform 1 0 1080 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_21
timestamp 1515334672
transform 1 0 1128 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_16
timestamp 1515334672
transform -1 0 1256 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_22
timestamp 1515334672
transform -1 0 1320 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_29
timestamp 1515334672
transform -1 0 1384 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_32
timestamp 1515334672
transform 1 0 1384 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1515334672
transform 1 0 1448 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_8
timestamp 1515334672
transform 1 0 1512 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_15
timestamp 1515334672
transform 1 0 1560 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_37
timestamp 1515334672
transform 1 0 1608 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_14
timestamp 1515334672
transform -1 0 1736 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_2
timestamp 1515334672
transform 1 0 1736 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_9
timestamp 1515334672
transform 1 0 1784 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_23
timestamp 1515334672
transform 1 0 1832 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_43
timestamp 1515334672
transform 1 0 1896 0 1 210
box 0 0 48 200
use NAND2X1  NAND2X1_39
timestamp 1515334672
transform -1 0 1992 0 1 210
box 0 0 48 200
use INVX1  INVX1_20
timestamp 1515334672
transform -1 0 2024 0 1 210
box 0 0 32 200
use NOR2X1  NOR2X1_19
timestamp 1515334672
transform -1 0 2072 0 1 210
box 0 0 48 200
use FILL  FILL_1_1_0
timestamp 1515334672
transform -1 0 2088 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1515334672
transform -1 0 2104 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_35
timestamp 1515334672
transform -1 0 2152 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_43
timestamp 1515334672
transform -1 0 2216 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_58
timestamp 1515334672
transform 1 0 2216 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_44
timestamp 1515334672
transform 1 0 2280 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_57
timestamp 1515334672
transform 1 0 2328 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_51
timestamp 1515334672
transform 1 0 2392 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_42
timestamp 1515334672
transform 1 0 2456 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_50
timestamp 1515334672
transform -1 0 2568 0 1 210
box 0 0 64 200
use INVX1  INVX1_22
timestamp 1515334672
transform -1 0 2600 0 1 210
box 0 0 32 200
use XOR2X1  XOR2X1_1
timestamp 1515334672
transform 1 0 2600 0 1 210
box 0 0 112 200
use NOR3X1  NOR3X1_8
timestamp 1515334672
transform 1 0 2712 0 1 210
box 0 0 128 200
use AND2X2  AND2X2_12
timestamp 1515334672
transform -1 0 2904 0 1 210
box 0 0 64 200
use AOI22X1  AOI22X1_11
timestamp 1515334672
transform 1 0 2904 0 1 210
box 0 0 80 200
use AND2X2  AND2X2_7
timestamp 1515334672
transform 1 0 2984 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_9
timestamp 1515334672
transform 1 0 3048 0 1 210
box 0 0 64 200
use INVX8  INVX8_4
timestamp 1515334672
transform 1 0 3112 0 1 210
box 0 0 80 200
use BUFX2  BUFX2_19
timestamp 1515334672
transform -1 0 56 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_5
timestamp 1515334672
transform -1 0 120 0 -1 210
box 0 0 64 200
use BUFX4  BUFX4_1
timestamp 1515334672
transform 1 0 120 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_38
timestamp 1515334672
transform 1 0 184 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_37
timestamp 1515334672
transform 1 0 248 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_22
timestamp 1515334672
transform 1 0 312 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_25
timestamp 1515334672
transform 1 0 360 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_24
timestamp 1515334672
transform -1 0 488 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_31
timestamp 1515334672
transform 1 0 488 0 -1 210
box 0 0 48 200
use INVX1  INVX1_14
timestamp 1515334672
transform 1 0 536 0 -1 210
box 0 0 32 200
use OAI21X1  OAI21X1_47
timestamp 1515334672
transform 1 0 568 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_16
timestamp 1515334672
transform -1 0 696 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_17
timestamp 1515334672
transform -1 0 760 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_18
timestamp 1515334672
transform -1 0 824 0 -1 210
box 0 0 64 200
use INVX2  INVX2_4
timestamp 1515334672
transform -1 0 856 0 -1 210
box 0 0 32 200
use NAND3X1  NAND3X1_39
timestamp 1515334672
transform -1 0 920 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_40
timestamp 1515334672
transform -1 0 984 0 -1 210
box 0 0 64 200
use AOI21X1  AOI21X1_13
timestamp 1515334672
transform 1 0 984 0 -1 210
box 0 0 64 200
use FILL  FILL_0_0_0
timestamp 1515334672
transform -1 0 1064 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1515334672
transform -1 0 1080 0 -1 210
box 0 0 16 200
use NAND3X1  NAND3X1_12
timestamp 1515334672
transform -1 0 1144 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_26
timestamp 1515334672
transform -1 0 1192 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_56
timestamp 1515334672
transform -1 0 1256 0 -1 210
box 0 0 64 200
use AOI21X1  AOI21X1_15
timestamp 1515334672
transform 1 0 1256 0 -1 210
box 0 0 64 200
use NAND3X1  NAND3X1_13
timestamp 1515334672
transform 1 0 1320 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_14
timestamp 1515334672
transform 1 0 1384 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_48
timestamp 1515334672
transform -1 0 1512 0 -1 210
box 0 0 64 200
use NAND2X1  NAND2X1_11
timestamp 1515334672
transform 1 0 1512 0 -1 210
box 0 0 48 200
use NAND2X1  NAND2X1_15
timestamp 1515334672
transform -1 0 1608 0 -1 210
box 0 0 48 200
use INVX1  INVX1_19
timestamp 1515334672
transform 1 0 1608 0 -1 210
box 0 0 32 200
use AOI21X1  AOI21X1_16
timestamp 1515334672
transform -1 0 1704 0 -1 210
box 0 0 64 200
use AOI21X1  AOI21X1_19
timestamp 1515334672
transform -1 0 1768 0 -1 210
box 0 0 64 200
use NOR2X1  NOR2X1_25
timestamp 1515334672
transform 1 0 1768 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_39
timestamp 1515334672
transform -1 0 1880 0 -1 210
box 0 0 64 200
use AND2X2  AND2X2_17
timestamp 1515334672
transform 1 0 1880 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_5
timestamp 1515334672
transform 1 0 1944 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_46
timestamp 1515334672
transform -1 0 2040 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_8
timestamp 1515334672
transform 1 0 2040 0 -1 210
box 0 0 48 200
use FILL  FILL_0_1_0
timestamp 1515334672
transform 1 0 2088 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1515334672
transform 1 0 2104 0 -1 210
box 0 0 16 200
use OAI21X1  OAI21X1_59
timestamp 1515334672
transform 1 0 2120 0 -1 210
box 0 0 64 200
use XNOR2X1  XNOR2X1_6
timestamp 1515334672
transform 1 0 2184 0 -1 210
box 0 0 112 200
use INVX1  INVX1_23
timestamp 1515334672
transform 1 0 2296 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_7
timestamp 1515334672
transform 1 0 2328 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_56
timestamp 1515334672
transform -1 0 2440 0 -1 210
box 0 0 64 200
use OR2X2  OR2X2_5
timestamp 1515334672
transform -1 0 2504 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_12
timestamp 1515334672
transform -1 0 2552 0 -1 210
box 0 0 48 200
use OAI21X1  OAI21X1_55
timestamp 1515334672
transform -1 0 2616 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_15
timestamp 1515334672
transform 1 0 2616 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_10
timestamp 1515334672
transform 1 0 2664 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_6
timestamp 1515334672
transform 1 0 2712 0 -1 210
box 0 0 48 200
use NAND3X1  NAND3X1_55
timestamp 1515334672
transform 1 0 2760 0 -1 210
box 0 0 64 200
use BUFX2  BUFX2_4
timestamp 1515334672
transform -1 0 2872 0 -1 210
box 0 0 48 200
use NOR3X1  NOR3X1_10
timestamp 1515334672
transform -1 0 3000 0 -1 210
box 0 0 128 200
use BUFX2  BUFX2_1
timestamp 1515334672
transform -1 0 3048 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_18
timestamp 1515334672
transform 1 0 3048 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_2
timestamp 1515334672
transform 1 0 3096 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_3
timestamp 1515334672
transform 1 0 3144 0 -1 210
box 0 0 48 200
<< labels >>
flabel space 1268 42 1276 136 6 FreeSans 48 0 0 0 vdd
port 0 nsew
flabel space 2308 42 2316 136 6 FreeSans 48 0 0 0 gnd
port 1 nsew
flabel metal3 -48 1580 -48 1580 7 FreeSans 48 0 0 0 ULA_A<0>
port 2 nsew
flabel metal3 -48 1540 -48 1540 7 FreeSans 48 0 0 0 ULA_A<1>
port 3 nsew
flabel metal3 -48 1360 -48 1360 7 FreeSans 48 0 0 0 ULA_A<2>
port 4 nsew
flabel metal3 -48 1320 -48 1320 7 FreeSans 48 0 0 0 ULA_A<3>
port 5 nsew
flabel metal3 -48 960 -48 960 7 FreeSans 48 0 0 0 ULA_A<4>
port 6 nsew
flabel metal3 -48 920 -48 920 7 FreeSans 48 0 0 0 ULA_A<5>
port 7 nsew
flabel metal2 240 2260 240 2260 3 FreeSans 48 90 0 0 ULA_A<6>
port 8 nsew
flabel metal2 2304 2260 2304 2260 3 FreeSans 48 90 0 0 ULA_A<7>
port 9 nsew
flabel metal2 96 2260 96 2260 3 FreeSans 48 90 0 0 ULA_A<8>
port 10 nsew
flabel metal2 288 2260 288 2260 3 FreeSans 48 90 0 0 ULA_A<9>
port 11 nsew
flabel metal2 672 2260 672 2260 3 FreeSans 48 90 0 0 ULA_A<10>
port 12 nsew
flabel metal2 720 2260 720 2260 3 FreeSans 48 90 0 0 ULA_A<11>
port 13 nsew
flabel metal2 864 2260 864 2260 3 FreeSans 48 90 0 0 ULA_A<12>
port 14 nsew
flabel metal2 1104 2260 1104 2260 3 FreeSans 48 90 0 0 ULA_A<13>
port 15 nsew
flabel metal2 1232 2260 1232 2260 3 FreeSans 48 90 0 0 ULA_A<14>
port 16 nsew
flabel metal3 3248 1960 3248 1960 3 FreeSans 48 0 0 0 ULA_A<15>
port 17 nsew
flabel metal3 -48 1500 -48 1500 7 FreeSans 48 0 0 0 ULA_B<0>
port 18 nsew
flabel metal3 -48 700 -48 700 7 FreeSans 48 0 0 0 ULA_B<1>
port 19 nsew
flabel metal2 1520 2260 1520 2260 3 FreeSans 48 90 0 0 ULA_B<2>
port 20 nsew
flabel metal2 1808 2260 1808 2260 3 FreeSans 48 90 0 0 ULA_B<3>
port 21 nsew
flabel metal2 1968 2260 1968 2260 3 FreeSans 48 90 0 0 ULA_B<4>
port 22 nsew
flabel metal2 2432 -40 2432 -40 7 FreeSans 48 270 0 0 ULA_B<5>
port 23 nsew
flabel metal2 1968 -40 1968 -40 7 FreeSans 48 270 0 0 ULA_B<6>
port 24 nsew
flabel metal2 2336 2260 2336 2260 3 FreeSans 48 90 0 0 ULA_B<7>
port 25 nsew
flabel metal3 3248 1520 3248 1520 3 FreeSans 48 0 0 0 ULA_B<8>
port 26 nsew
flabel metal2 2912 2260 2912 2260 3 FreeSans 48 90 0 0 ULA_B<9>
port 27 nsew
flabel metal3 3248 1060 3248 1060 3 FreeSans 48 0 0 0 ULA_B<10>
port 28 nsew
flabel metal2 2256 2260 2256 2260 3 FreeSans 48 90 0 0 ULA_B<11>
port 29 nsew
flabel metal2 2384 2260 2384 2260 3 FreeSans 48 90 0 0 ULA_B<12>
port 30 nsew
flabel metal3 3248 1360 3248 1360 3 FreeSans 48 0 0 0 ULA_B<13>
port 31 nsew
flabel metal2 2480 -40 2480 -40 7 FreeSans 48 270 0 0 ULA_B<14>
port 32 nsew
flabel metal3 3248 1920 3248 1920 3 FreeSans 48 0 0 0 ULA_B<15>
port 33 nsew
flabel metal3 3248 1320 3248 1320 3 FreeSans 48 0 0 0 ULA_ctrl<0>
port 34 nsew
flabel metal2 2864 2260 2864 2260 3 FreeSans 48 90 0 0 ULA_ctrl<1>
port 35 nsew
flabel metal2 2544 2260 2544 2260 3 FreeSans 48 90 0 0 ULA_ctrl<2>
port 36 nsew
flabel metal2 3040 2260 3040 2260 3 FreeSans 48 90 0 0 ULA_ctrl<3>
port 37 nsew
flabel metal2 3008 -40 3008 -40 7 FreeSans 48 270 0 0 ULA_OUT<0>
port 38 nsew
flabel metal2 3136 -40 3136 -40 7 FreeSans 48 270 0 0 ULA_OUT<1>
port 39 nsew
flabel metal3 3248 120 3248 120 3 FreeSans 48 0 0 0 ULA_OUT<2>
port 40 nsew
flabel metal2 2832 -40 2832 -40 7 FreeSans 48 270 0 0 ULA_OUT<3>
port 41 nsew
flabel metal2 2048 -40 2048 -40 7 FreeSans 48 270 0 0 ULA_OUT<4>
port 42 nsew
flabel metal2 2752 -40 2752 -40 7 FreeSans 48 270 0 0 ULA_OUT<5>
port 43 nsew
flabel metal2 2368 -40 2368 -40 7 FreeSans 48 270 0 0 ULA_OUT<6>
port 44 nsew
flabel metal2 2176 -40 2176 -40 7 FreeSans 48 270 0 0 ULA_OUT<7>
port 45 nsew
flabel metal3 3248 720 3248 720 3 FreeSans 48 0 0 0 ULA_OUT<8>
port 46 nsew
flabel metal2 2704 -40 2704 -40 7 FreeSans 48 270 0 0 ULA_OUT<9>
port 47 nsew
flabel metal3 3248 920 3248 920 3 FreeSans 48 0 0 0 ULA_OUT<10>
port 48 nsew
flabel metal2 2512 -40 2512 -40 7 FreeSans 48 270 0 0 ULA_OUT<11>
port 49 nsew
flabel metal3 3248 1560 3248 1560 3 FreeSans 48 0 0 0 ULA_OUT<12>
port 50 nsew
flabel metal3 3248 760 3248 760 3 FreeSans 48 0 0 0 ULA_OUT<13>
port 51 nsew
flabel metal2 2656 -40 2656 -40 7 FreeSans 48 270 0 0 ULA_OUT<14>
port 52 nsew
flabel metal3 3248 520 3248 520 3 FreeSans 48 0 0 0 ULA_OUT<15>
port 53 nsew
flabel metal2 3088 2260 3088 2260 3 FreeSans 48 90 0 0 ULA_flags<0>
port 54 nsew
flabel metal2 3088 -40 3088 -40 7 FreeSans 48 270 0 0 ULA_flags<1>
port 55 nsew
flabel metal3 -48 120 -48 120 7 FreeSans 48 0 0 0 ULA_flags<2>
port 56 nsew
<< end >>
